module configurable_sync_fifo (almost_empty,
    almost_full,
    clk,
    empty,
    full,
    rd_en,
    rst_n,
    wr_en,
    data_in,
    data_out,
    fill_level);
 output almost_empty;
 output almost_full;
 input clk;
 output empty;
 output full;
 input rd_en;
 input rst_n;
 input wr_en;
 input [7:0] data_in;
 output [7:0] data_out;
 output [4:0] fill_level;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire \memory[0][0] ;
 wire \memory[0][1] ;
 wire \memory[0][2] ;
 wire \memory[0][3] ;
 wire \memory[0][4] ;
 wire \memory[0][5] ;
 wire \memory[0][6] ;
 wire \memory[0][7] ;
 wire \memory[10][0] ;
 wire \memory[10][1] ;
 wire \memory[10][2] ;
 wire \memory[10][3] ;
 wire \memory[10][4] ;
 wire \memory[10][5] ;
 wire \memory[10][6] ;
 wire \memory[10][7] ;
 wire \memory[11][0] ;
 wire \memory[11][1] ;
 wire \memory[11][2] ;
 wire \memory[11][3] ;
 wire \memory[11][4] ;
 wire \memory[11][5] ;
 wire \memory[11][6] ;
 wire \memory[11][7] ;
 wire \memory[12][0] ;
 wire \memory[12][1] ;
 wire \memory[12][2] ;
 wire \memory[12][3] ;
 wire \memory[12][4] ;
 wire \memory[12][5] ;
 wire \memory[12][6] ;
 wire \memory[12][7] ;
 wire \memory[13][0] ;
 wire \memory[13][1] ;
 wire \memory[13][2] ;
 wire \memory[13][3] ;
 wire \memory[13][4] ;
 wire \memory[13][5] ;
 wire \memory[13][6] ;
 wire \memory[13][7] ;
 wire \memory[14][0] ;
 wire \memory[14][1] ;
 wire \memory[14][2] ;
 wire \memory[14][3] ;
 wire \memory[14][4] ;
 wire \memory[14][5] ;
 wire \memory[14][6] ;
 wire \memory[14][7] ;
 wire \memory[15][0] ;
 wire \memory[15][1] ;
 wire \memory[15][2] ;
 wire \memory[15][3] ;
 wire \memory[15][4] ;
 wire \memory[15][5] ;
 wire \memory[15][6] ;
 wire \memory[15][7] ;
 wire \memory[1][0] ;
 wire \memory[1][1] ;
 wire \memory[1][2] ;
 wire \memory[1][3] ;
 wire \memory[1][4] ;
 wire \memory[1][5] ;
 wire \memory[1][6] ;
 wire \memory[1][7] ;
 wire \memory[2][0] ;
 wire \memory[2][1] ;
 wire \memory[2][2] ;
 wire \memory[2][3] ;
 wire \memory[2][4] ;
 wire \memory[2][5] ;
 wire \memory[2][6] ;
 wire \memory[2][7] ;
 wire \memory[3][0] ;
 wire \memory[3][1] ;
 wire \memory[3][2] ;
 wire \memory[3][3] ;
 wire \memory[3][4] ;
 wire \memory[3][5] ;
 wire \memory[3][6] ;
 wire \memory[3][7] ;
 wire \memory[4][0] ;
 wire \memory[4][1] ;
 wire \memory[4][2] ;
 wire \memory[4][3] ;
 wire \memory[4][4] ;
 wire \memory[4][5] ;
 wire \memory[4][6] ;
 wire \memory[4][7] ;
 wire \memory[5][0] ;
 wire \memory[5][1] ;
 wire \memory[5][2] ;
 wire \memory[5][3] ;
 wire \memory[5][4] ;
 wire \memory[5][5] ;
 wire \memory[5][6] ;
 wire \memory[5][7] ;
 wire \memory[6][0] ;
 wire \memory[6][1] ;
 wire \memory[6][2] ;
 wire \memory[6][3] ;
 wire \memory[6][4] ;
 wire \memory[6][5] ;
 wire \memory[6][6] ;
 wire \memory[6][7] ;
 wire \memory[7][0] ;
 wire \memory[7][1] ;
 wire \memory[7][2] ;
 wire \memory[7][3] ;
 wire \memory[7][4] ;
 wire \memory[7][5] ;
 wire \memory[7][6] ;
 wire \memory[7][7] ;
 wire \memory[8][0] ;
 wire \memory[8][1] ;
 wire \memory[8][2] ;
 wire \memory[8][3] ;
 wire \memory[8][4] ;
 wire \memory[8][5] ;
 wire \memory[8][6] ;
 wire \memory[8][7] ;
 wire \memory[9][0] ;
 wire \memory[9][1] ;
 wire \memory[9][2] ;
 wire \memory[9][3] ;
 wire \memory[9][4] ;
 wire \memory[9][5] ;
 wire \memory[9][6] ;
 wire \memory[9][7] ;
 wire \rd_ptr[0] ;
 wire \rd_ptr[1] ;
 wire \rd_ptr[2] ;
 wire \rd_ptr[3] ;
 wire \wr_ptr[0] ;
 wire \wr_ptr[1] ;
 wire \wr_ptr[2] ;
 wire \wr_ptr[3] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net30;
 wire net31;
 wire net32;
 wire net33;

 sky130_fd_sc_hd__inv_1 _275_ (.A(net28),
    .Y(_038_));
 sky130_fd_sc_hd__or4_1 _276_ (.A(net25),
    .B(net24),
    .C(net27),
    .D(net26),
    .X(_039_));
 sky130_fd_sc_hd__nor2_1 _277_ (.A(_038_),
    .B(_039_),
    .Y(net29));
 sky130_fd_sc_hd__nor2b_1 _278_ (.A(net29),
    .B_N(net12),
    .Y(_040_));
 sky130_fd_sc_hd__clkbuf_4 _279_ (.A(_040_),
    .X(_243_));
 sky130_fd_sc_hd__nor2_1 _280_ (.A(net28),
    .B(_039_),
    .Y(net23));
 sky130_fd_sc_hd__nand3_4 _281_ (.A(net11),
    .B(_252_),
    .C(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__buf_6 _282_ (.A(\wr_ptr[2] ),
    .X(_042_));
 sky130_fd_sc_hd__buf_6 _283_ (.A(\wr_ptr[3] ),
    .X(_043_));
 sky130_fd_sc_hd__nand2_8 _284_ (.A(_042_),
    .B(_043_),
    .Y(_044_));
 sky130_fd_sc_hd__nor2_8 _285_ (.A(_041_),
    .B(_044_),
    .Y(_002_));
 sky130_fd_sc_hd__nand3_4 _286_ (.A(net11),
    .B(_254_),
    .C(_243_),
    .Y(_045_));
 sky130_fd_sc_hd__nand2b_4 _287_ (.A_N(_042_),
    .B(_043_),
    .Y(_046_));
 sky130_fd_sc_hd__nor2_4 _288_ (.A(_045_),
    .B(_046_),
    .Y(_004_));
 sky130_fd_sc_hd__inv_1 _289_ (.A(net24),
    .Y(_016_));
 sky130_fd_sc_hd__nand3_4 _290_ (.A(net11),
    .B(_248_),
    .C(_243_),
    .Y(_047_));
 sky130_fd_sc_hd__nor3_4 _291_ (.A(_042_),
    .B(_043_),
    .C(_047_),
    .Y(_015_));
 sky130_fd_sc_hd__nor3_4 _292_ (.A(_042_),
    .B(_043_),
    .C(_041_),
    .Y(_014_));
 sky130_fd_sc_hd__nand3_4 _293_ (.A(net11),
    .B(_250_),
    .C(_243_),
    .Y(_048_));
 sky130_fd_sc_hd__nor3_4 _294_ (.A(_042_),
    .B(_043_),
    .C(_048_),
    .Y(_013_));
 sky130_fd_sc_hd__nor3_4 _295_ (.A(_042_),
    .B(_043_),
    .C(_045_),
    .Y(_012_));
 sky130_fd_sc_hd__nand2b_4 _296_ (.A_N(_043_),
    .B(_042_),
    .Y(_049_));
 sky130_fd_sc_hd__nor2_4 _297_ (.A(_047_),
    .B(_049_),
    .Y(_011_));
 sky130_fd_sc_hd__nor2_8 _298_ (.A(_041_),
    .B(_049_),
    .Y(_010_));
 sky130_fd_sc_hd__nor2_8 _299_ (.A(_048_),
    .B(_049_),
    .Y(_009_));
 sky130_fd_sc_hd__nor2_4 _300_ (.A(_045_),
    .B(_049_),
    .Y(_008_));
 sky130_fd_sc_hd__nor2_4 _301_ (.A(_046_),
    .B(_047_),
    .Y(_007_));
 sky130_fd_sc_hd__nor2_8 _302_ (.A(_041_),
    .B(_046_),
    .Y(_006_));
 sky130_fd_sc_hd__nor2_8 _303_ (.A(_044_),
    .B(_045_),
    .Y(_000_));
 sky130_fd_sc_hd__nor2_4 _304_ (.A(_044_),
    .B(_047_),
    .Y(_003_));
 sky130_fd_sc_hd__nor2_8 _305_ (.A(_046_),
    .B(_048_),
    .Y(_005_));
 sky130_fd_sc_hd__nor2_4 _306_ (.A(_044_),
    .B(_048_),
    .Y(_001_));
 sky130_fd_sc_hd__inv_1 _307_ (.A(net25),
    .Y(_239_));
 sky130_fd_sc_hd__inv_1 _308_ (.A(\wr_ptr[0] ),
    .Y(_246_));
 sky130_fd_sc_hd__inv_1 _309_ (.A(\rd_ptr[0] ),
    .Y(_256_));
 sky130_fd_sc_hd__o21a_2 _310_ (.A1(net28),
    .A2(_039_),
    .B1(net10),
    .X(_050_));
 sky130_fd_sc_hd__inv_2 _311_ (.A(_050_),
    .Y(_051_));
 sky130_fd_sc_hd__buf_6 _312_ (.A(_051_),
    .X(_244_));
 sky130_fd_sc_hd__inv_1 _313_ (.A(\wr_ptr[1] ),
    .Y(_247_));
 sky130_fd_sc_hd__inv_1 _314_ (.A(\rd_ptr[1] ),
    .Y(_257_));
 sky130_fd_sc_hd__inv_1 _315_ (.A(_240_),
    .Y(_266_));
 sky130_fd_sc_hd__buf_2 _316_ (.A(_050_),
    .X(_052_));
 sky130_fd_sc_hd__buf_4 _317_ (.A(_262_),
    .X(_053_));
 sky130_fd_sc_hd__buf_4 _318_ (.A(_053_),
    .X(_054_));
 sky130_fd_sc_hd__inv_1 _319_ (.A(\memory[1][0] ),
    .Y(_055_));
 sky130_fd_sc_hd__clkbuf_2 _320_ (.A(\rd_ptr[3] ),
    .X(_056_));
 sky130_fd_sc_hd__or2_2 _321_ (.A(\rd_ptr[2] ),
    .B(_056_),
    .X(_057_));
 sky130_fd_sc_hd__clkbuf_4 _322_ (.A(\rd_ptr[2] ),
    .X(_058_));
 sky130_fd_sc_hd__buf_4 _323_ (.A(_056_),
    .X(_059_));
 sky130_fd_sc_hd__buf_4 _324_ (.A(_059_),
    .X(_060_));
 sky130_fd_sc_hd__nand3_1 _325_ (.A(_058_),
    .B(_060_),
    .C(\memory[13][0] ),
    .Y(_061_));
 sky130_fd_sc_hd__o21ai_0 _326_ (.A1(_055_),
    .A2(_057_),
    .B1(_061_),
    .Y(_062_));
 sky130_fd_sc_hd__o21ai_1 _327_ (.A1(_058_),
    .A2(_059_),
    .B1(_258_),
    .Y(_063_));
 sky130_fd_sc_hd__nor3_1 _328_ (.A(_264_),
    .B(_260_),
    .C(_262_),
    .Y(_064_));
 sky130_fd_sc_hd__and2_0 _329_ (.A(_063_),
    .B(_064_),
    .X(_065_));
 sky130_fd_sc_hd__nand2b_2 _330_ (.A_N(\rd_ptr[2] ),
    .B(_056_),
    .Y(_066_));
 sky130_fd_sc_hd__buf_4 _331_ (.A(_258_),
    .X(_067_));
 sky130_fd_sc_hd__clkbuf_4 _332_ (.A(_053_),
    .X(_068_));
 sky130_fd_sc_hd__a22oi_1 _333_ (.A1(\memory[8][0] ),
    .A2(_067_),
    .B1(_068_),
    .B2(\memory[9][0] ),
    .Y(_069_));
 sky130_fd_sc_hd__nand2_2 _334_ (.A(_058_),
    .B(_264_),
    .Y(_070_));
 sky130_fd_sc_hd__mux2i_2 _335_ (.A0(\memory[7][0] ),
    .A1(\memory[15][0] ),
    .S(_059_),
    .Y(_071_));
 sky130_fd_sc_hd__clkbuf_4 _336_ (.A(_058_),
    .X(_072_));
 sky130_fd_sc_hd__buf_4 _337_ (.A(_258_),
    .X(_073_));
 sky130_fd_sc_hd__mux2_1 _338_ (.A0(\memory[4][0] ),
    .A1(\memory[12][0] ),
    .S(_059_),
    .X(_074_));
 sky130_fd_sc_hd__nand3_1 _339_ (.A(_072_),
    .B(_073_),
    .C(_074_),
    .Y(_075_));
 sky130_fd_sc_hd__o221ai_2 _340_ (.A1(_066_),
    .A2(_069_),
    .B1(_070_),
    .B2(_071_),
    .C1(_075_),
    .Y(_076_));
 sky130_fd_sc_hd__a211oi_1 _341_ (.A1(_054_),
    .A2(_062_),
    .B1(_065_),
    .C1(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__buf_4 _342_ (.A(_059_),
    .X(_078_));
 sky130_fd_sc_hd__clkbuf_4 _343_ (.A(_260_),
    .X(_079_));
 sky130_fd_sc_hd__clkbuf_4 _344_ (.A(_079_),
    .X(_080_));
 sky130_fd_sc_hd__a22oi_2 _345_ (.A1(\memory[6][0] ),
    .A2(_080_),
    .B1(_068_),
    .B2(\memory[5][0] ),
    .Y(_081_));
 sky130_fd_sc_hd__nand3_1 _346_ (.A(_078_),
    .B(\memory[14][0] ),
    .C(_080_),
    .Y(_082_));
 sky130_fd_sc_hd__clkbuf_4 _347_ (.A(_058_),
    .X(_083_));
 sky130_fd_sc_hd__o211ai_2 _348_ (.A1(_078_),
    .A2(_081_),
    .B1(_082_),
    .C1(_083_),
    .Y(_084_));
 sky130_fd_sc_hd__clkbuf_4 _349_ (.A(_264_),
    .X(_085_));
 sky130_fd_sc_hd__clkbuf_4 _350_ (.A(_085_),
    .X(_086_));
 sky130_fd_sc_hd__buf_4 _351_ (.A(_260_),
    .X(_087_));
 sky130_fd_sc_hd__a221o_1 _352_ (.A1(_086_),
    .A2(\memory[3][0] ),
    .B1(\memory[2][0] ),
    .B2(_087_),
    .C1(_057_),
    .X(_088_));
 sky130_fd_sc_hd__a221o_1 _353_ (.A1(_086_),
    .A2(\memory[11][0] ),
    .B1(\memory[10][0] ),
    .B2(_087_),
    .C1(_066_),
    .X(_089_));
 sky130_fd_sc_hd__nand3_1 _354_ (.A(_084_),
    .B(_088_),
    .C(_089_),
    .Y(_090_));
 sky130_fd_sc_hd__nand2_2 _355_ (.A(_063_),
    .B(_064_),
    .Y(_091_));
 sky130_fd_sc_hd__or3_1 _356_ (.A(\memory[0][0] ),
    .B(_051_),
    .C(_091_),
    .X(_092_));
 sky130_fd_sc_hd__o21ai_0 _357_ (.A1(net15),
    .A2(_050_),
    .B1(_092_),
    .Y(_093_));
 sky130_fd_sc_hd__a31oi_1 _358_ (.A1(_052_),
    .A2(_077_),
    .A3(_090_),
    .B1(_093_),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _359_ (.A(_059_),
    .Y(_094_));
 sky130_fd_sc_hd__a22oi_1 _360_ (.A1(\memory[12][1] ),
    .A2(_073_),
    .B1(_080_),
    .B2(\memory[14][1] ),
    .Y(_095_));
 sky130_fd_sc_hd__mux2i_1 _361_ (.A0(\memory[7][1] ),
    .A1(\memory[15][1] ),
    .S(_060_),
    .Y(_096_));
 sky130_fd_sc_hd__inv_1 _362_ (.A(_086_),
    .Y(_097_));
 sky130_fd_sc_hd__o22ai_1 _363_ (.A1(_094_),
    .A2(_095_),
    .B1(_096_),
    .B2(_097_),
    .Y(_098_));
 sky130_fd_sc_hd__a221oi_1 _364_ (.A1(\memory[10][1] ),
    .A2(_087_),
    .B1(_068_),
    .B2(\memory[9][1] ),
    .C1(_094_),
    .Y(_099_));
 sky130_fd_sc_hd__a21oi_1 _365_ (.A1(_086_),
    .A2(\memory[3][1] ),
    .B1(_078_),
    .Y(_100_));
 sky130_fd_sc_hd__nor3_1 _366_ (.A(_083_),
    .B(_099_),
    .C(_100_),
    .Y(_101_));
 sky130_fd_sc_hd__a21oi_1 _367_ (.A1(_083_),
    .A2(_098_),
    .B1(_101_),
    .Y(_102_));
 sky130_fd_sc_hd__a22oi_1 _368_ (.A1(\memory[4][1] ),
    .A2(_258_),
    .B1(_053_),
    .B2(\memory[5][1] ),
    .Y(_103_));
 sky130_fd_sc_hd__nand2_1 _369_ (.A(\memory[6][1] ),
    .B(_087_),
    .Y(_104_));
 sky130_fd_sc_hd__a21oi_1 _370_ (.A1(\memory[1][1] ),
    .A2(_068_),
    .B1(_058_),
    .Y(_105_));
 sky130_fd_sc_hd__a311oi_2 _371_ (.A1(_058_),
    .A2(_103_),
    .A3(_104_),
    .B1(_060_),
    .C1(_105_),
    .Y(_106_));
 sky130_fd_sc_hd__nand2_2 _372_ (.A(_058_),
    .B(_059_),
    .Y(_107_));
 sky130_fd_sc_hd__nand2_1 _373_ (.A(\memory[13][1] ),
    .B(_054_),
    .Y(_108_));
 sky130_fd_sc_hd__nand2_1 _374_ (.A(\memory[2][1] ),
    .B(_080_),
    .Y(_109_));
 sky130_fd_sc_hd__o22ai_1 _375_ (.A1(_107_),
    .A2(_108_),
    .B1(_109_),
    .B2(_057_),
    .Y(_110_));
 sky130_fd_sc_hd__a22oi_1 _376_ (.A1(_086_),
    .A2(\memory[11][1] ),
    .B1(\memory[8][1] ),
    .B2(_073_),
    .Y(_111_));
 sky130_fd_sc_hd__o21ai_0 _377_ (.A1(_066_),
    .A2(_111_),
    .B1(_091_),
    .Y(_112_));
 sky130_fd_sc_hd__nor4_1 _378_ (.A(_244_),
    .B(_106_),
    .C(_110_),
    .D(_112_),
    .Y(_113_));
 sky130_fd_sc_hd__or3_1 _379_ (.A(\memory[0][1] ),
    .B(_244_),
    .C(_091_),
    .X(_114_));
 sky130_fd_sc_hd__o21ai_0 _380_ (.A1(net16),
    .A2(_052_),
    .B1(_114_),
    .Y(_115_));
 sky130_fd_sc_hd__a21oi_1 _381_ (.A1(_102_),
    .A2(_113_),
    .B1(_115_),
    .Y(_023_));
 sky130_fd_sc_hd__nand2_2 _382_ (.A(_050_),
    .B(_091_),
    .Y(_116_));
 sky130_fd_sc_hd__nor2b_1 _383_ (.A(_058_),
    .B_N(_085_),
    .Y(_117_));
 sky130_fd_sc_hd__a32oi_1 _384_ (.A1(_072_),
    .A2(\memory[5][2] ),
    .A3(_054_),
    .B1(_117_),
    .B2(\memory[3][2] ),
    .Y(_118_));
 sky130_fd_sc_hd__mux2i_2 _385_ (.A0(\memory[7][2] ),
    .A1(\memory[15][2] ),
    .S(_060_),
    .Y(_119_));
 sky130_fd_sc_hd__o22ai_1 _386_ (.A1(_078_),
    .A2(_118_),
    .B1(_119_),
    .B2(_070_),
    .Y(_120_));
 sky130_fd_sc_hd__nor2_1 _387_ (.A(_116_),
    .B(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__a22oi_1 _388_ (.A1(\memory[12][2] ),
    .A2(_073_),
    .B1(_080_),
    .B2(\memory[14][2] ),
    .Y(_122_));
 sky130_fd_sc_hd__nand2_1 _389_ (.A(\memory[13][2] ),
    .B(_054_),
    .Y(_123_));
 sky130_fd_sc_hd__a221oi_1 _390_ (.A1(\memory[4][2] ),
    .A2(_067_),
    .B1(_080_),
    .B2(\memory[6][2] ),
    .C1(_060_),
    .Y(_124_));
 sky130_fd_sc_hd__a31oi_1 _391_ (.A1(_078_),
    .A2(_122_),
    .A3(_123_),
    .B1(_124_),
    .Y(_125_));
 sky130_fd_sc_hd__a22oi_1 _392_ (.A1(_086_),
    .A2(\memory[11][2] ),
    .B1(\memory[8][2] ),
    .B2(_073_),
    .Y(_126_));
 sky130_fd_sc_hd__a22oi_1 _393_ (.A1(\memory[10][2] ),
    .A2(_087_),
    .B1(_068_),
    .B2(\memory[9][2] ),
    .Y(_127_));
 sky130_fd_sc_hd__a221oi_1 _394_ (.A1(\memory[2][2] ),
    .A2(_087_),
    .B1(_053_),
    .B2(\memory[1][2] ),
    .C1(_060_),
    .Y(_128_));
 sky130_fd_sc_hd__a311oi_1 _395_ (.A1(_078_),
    .A2(_126_),
    .A3(_127_),
    .B1(_128_),
    .C1(_083_),
    .Y(_129_));
 sky130_fd_sc_hd__a21oi_1 _396_ (.A1(_083_),
    .A2(_125_),
    .B1(_129_),
    .Y(_130_));
 sky130_fd_sc_hd__or3_1 _397_ (.A(\memory[0][2] ),
    .B(_244_),
    .C(_091_),
    .X(_131_));
 sky130_fd_sc_hd__o21ai_0 _398_ (.A1(net17),
    .A2(_052_),
    .B1(_131_),
    .Y(_132_));
 sky130_fd_sc_hd__a21oi_1 _399_ (.A1(_121_),
    .A2(_130_),
    .B1(_132_),
    .Y(_024_));
 sky130_fd_sc_hd__a222oi_1 _400_ (.A1(\memory[14][3] ),
    .A2(_079_),
    .B1(_053_),
    .B2(\memory[13][3] ),
    .C1(\memory[12][3] ),
    .C2(_067_),
    .Y(_133_));
 sky130_fd_sc_hd__nand3_1 _401_ (.A(_094_),
    .B(\memory[4][3] ),
    .C(_073_),
    .Y(_134_));
 sky130_fd_sc_hd__o21ai_1 _402_ (.A1(_094_),
    .A2(_133_),
    .B1(_134_),
    .Y(_135_));
 sky130_fd_sc_hd__a222oi_1 _403_ (.A1(_264_),
    .A2(\memory[3][3] ),
    .B1(\memory[2][3] ),
    .B2(_260_),
    .C1(_262_),
    .C2(\memory[1][3] ),
    .Y(_136_));
 sky130_fd_sc_hd__mux2i_1 _404_ (.A0(\memory[7][3] ),
    .A1(\memory[15][3] ),
    .S(_056_),
    .Y(_137_));
 sky130_fd_sc_hd__o22ai_1 _405_ (.A1(_057_),
    .A2(_136_),
    .B1(_137_),
    .B2(_070_),
    .Y(_138_));
 sky130_fd_sc_hd__a22oi_1 _406_ (.A1(\memory[6][3] ),
    .A2(_260_),
    .B1(_262_),
    .B2(\memory[5][3] ),
    .Y(_139_));
 sky130_fd_sc_hd__nand2b_4 _407_ (.A_N(_056_),
    .B(\rd_ptr[2] ),
    .Y(_140_));
 sky130_fd_sc_hd__nor2_1 _408_ (.A(_139_),
    .B(_140_),
    .Y(_141_));
 sky130_fd_sc_hd__a22oi_1 _409_ (.A1(\memory[10][3] ),
    .A2(_079_),
    .B1(_053_),
    .B2(\memory[9][3] ),
    .Y(_142_));
 sky130_fd_sc_hd__a22oi_1 _410_ (.A1(_085_),
    .A2(\memory[11][3] ),
    .B1(\memory[8][3] ),
    .B2(_258_),
    .Y(_143_));
 sky130_fd_sc_hd__a21oi_1 _411_ (.A1(_142_),
    .A2(_143_),
    .B1(_066_),
    .Y(_144_));
 sky130_fd_sc_hd__or3_1 _412_ (.A(_138_),
    .B(_141_),
    .C(_144_),
    .X(_145_));
 sky130_fd_sc_hd__a21oi_1 _413_ (.A1(_083_),
    .A2(_135_),
    .B1(_145_),
    .Y(_146_));
 sky130_fd_sc_hd__nor2_1 _414_ (.A(net18),
    .B(_052_),
    .Y(_147_));
 sky130_fd_sc_hd__a21oi_1 _415_ (.A1(\memory[0][3] ),
    .A2(_065_),
    .B1(_244_),
    .Y(_148_));
 sky130_fd_sc_hd__o22ai_1 _416_ (.A1(_116_),
    .A2(_146_),
    .B1(_147_),
    .B2(_148_),
    .Y(_025_));
 sky130_fd_sc_hd__a222oi_1 _417_ (.A1(\memory[14][4] ),
    .A2(_079_),
    .B1(_053_),
    .B2(\memory[13][4] ),
    .C1(\memory[12][4] ),
    .C2(_067_),
    .Y(_149_));
 sky130_fd_sc_hd__nand3_1 _418_ (.A(_094_),
    .B(\memory[4][4] ),
    .C(_073_),
    .Y(_150_));
 sky130_fd_sc_hd__o21ai_1 _419_ (.A1(_094_),
    .A2(_149_),
    .B1(_150_),
    .Y(_151_));
 sky130_fd_sc_hd__a222oi_1 _420_ (.A1(_264_),
    .A2(\memory[3][4] ),
    .B1(\memory[2][4] ),
    .B2(_260_),
    .C1(_262_),
    .C2(\memory[1][4] ),
    .Y(_152_));
 sky130_fd_sc_hd__mux2i_1 _421_ (.A0(\memory[7][4] ),
    .A1(\memory[15][4] ),
    .S(_056_),
    .Y(_153_));
 sky130_fd_sc_hd__o22ai_1 _422_ (.A1(_057_),
    .A2(_152_),
    .B1(_153_),
    .B2(_070_),
    .Y(_154_));
 sky130_fd_sc_hd__a22oi_1 _423_ (.A1(\memory[6][4] ),
    .A2(_079_),
    .B1(_053_),
    .B2(\memory[5][4] ),
    .Y(_155_));
 sky130_fd_sc_hd__nor2_1 _424_ (.A(_140_),
    .B(_155_),
    .Y(_156_));
 sky130_fd_sc_hd__a22oi_1 _425_ (.A1(\memory[10][4] ),
    .A2(_079_),
    .B1(_053_),
    .B2(\memory[9][4] ),
    .Y(_157_));
 sky130_fd_sc_hd__a22oi_2 _426_ (.A1(_264_),
    .A2(\memory[11][4] ),
    .B1(\memory[8][4] ),
    .B2(_258_),
    .Y(_158_));
 sky130_fd_sc_hd__a21oi_1 _427_ (.A1(_157_),
    .A2(_158_),
    .B1(_066_),
    .Y(_159_));
 sky130_fd_sc_hd__or3_1 _428_ (.A(_154_),
    .B(_156_),
    .C(_159_),
    .X(_160_));
 sky130_fd_sc_hd__a21oi_1 _429_ (.A1(_083_),
    .A2(_151_),
    .B1(_160_),
    .Y(_161_));
 sky130_fd_sc_hd__nor2_1 _430_ (.A(net19),
    .B(_052_),
    .Y(_162_));
 sky130_fd_sc_hd__a21oi_1 _431_ (.A1(\memory[0][4] ),
    .A2(_065_),
    .B1(_244_),
    .Y(_163_));
 sky130_fd_sc_hd__o22ai_1 _432_ (.A1(_116_),
    .A2(_161_),
    .B1(_162_),
    .B2(_163_),
    .Y(_026_));
 sky130_fd_sc_hd__nor2_1 _433_ (.A(_072_),
    .B(_094_),
    .Y(_164_));
 sky130_fd_sc_hd__a22oi_1 _434_ (.A1(_085_),
    .A2(\memory[11][5] ),
    .B1(\memory[10][5] ),
    .B2(_079_),
    .Y(_165_));
 sky130_fd_sc_hd__nand2_1 _435_ (.A(\memory[8][5] ),
    .B(_067_),
    .Y(_166_));
 sky130_fd_sc_hd__a21oi_1 _436_ (.A1(_086_),
    .A2(\memory[3][5] ),
    .B1(_059_),
    .Y(_167_));
 sky130_fd_sc_hd__a311oi_1 _437_ (.A1(_060_),
    .A2(_165_),
    .A3(_166_),
    .B1(_167_),
    .C1(_072_),
    .Y(_168_));
 sky130_fd_sc_hd__a222oi_1 _438_ (.A1(_085_),
    .A2(\memory[7][5] ),
    .B1(\memory[6][5] ),
    .B2(_087_),
    .C1(_068_),
    .C2(\memory[5][5] ),
    .Y(_169_));
 sky130_fd_sc_hd__a22o_1 _439_ (.A1(_085_),
    .A2(\memory[15][5] ),
    .B1(\memory[14][5] ),
    .B2(_079_),
    .X(_170_));
 sky130_fd_sc_hd__a221oi_1 _440_ (.A1(\memory[12][5] ),
    .A2(_067_),
    .B1(_068_),
    .B2(\memory[13][5] ),
    .C1(_170_),
    .Y(_171_));
 sky130_fd_sc_hd__o22ai_2 _441_ (.A1(_140_),
    .A2(_169_),
    .B1(_171_),
    .B2(_107_),
    .Y(_172_));
 sky130_fd_sc_hd__a311oi_2 _442_ (.A1(\memory[9][5] ),
    .A2(_054_),
    .A3(_164_),
    .B1(_168_),
    .C1(_172_),
    .Y(_173_));
 sky130_fd_sc_hd__a22oi_1 _443_ (.A1(\memory[2][5] ),
    .A2(_080_),
    .B1(_054_),
    .B2(\memory[1][5] ),
    .Y(_174_));
 sky130_fd_sc_hd__nand3_1 _444_ (.A(_072_),
    .B(\memory[4][5] ),
    .C(_073_),
    .Y(_175_));
 sky130_fd_sc_hd__o21ai_0 _445_ (.A1(_072_),
    .A2(_174_),
    .B1(_175_),
    .Y(_176_));
 sky130_fd_sc_hd__a21oi_1 _446_ (.A1(_094_),
    .A2(_176_),
    .B1(_116_),
    .Y(_177_));
 sky130_fd_sc_hd__or3_1 _447_ (.A(\memory[0][5] ),
    .B(_244_),
    .C(_091_),
    .X(_178_));
 sky130_fd_sc_hd__o21ai_0 _448_ (.A1(net20),
    .A2(_052_),
    .B1(_178_),
    .Y(_179_));
 sky130_fd_sc_hd__a21oi_1 _449_ (.A1(_173_),
    .A2(_177_),
    .B1(_179_),
    .Y(_027_));
 sky130_fd_sc_hd__a32oi_1 _450_ (.A1(_058_),
    .A2(\memory[5][6] ),
    .A3(_054_),
    .B1(_117_),
    .B2(\memory[3][6] ),
    .Y(_180_));
 sky130_fd_sc_hd__mux2i_2 _451_ (.A0(\memory[7][6] ),
    .A1(\memory[15][6] ),
    .S(_060_),
    .Y(_181_));
 sky130_fd_sc_hd__o22ai_1 _452_ (.A1(_078_),
    .A2(_180_),
    .B1(_181_),
    .B2(_070_),
    .Y(_182_));
 sky130_fd_sc_hd__nor2_1 _453_ (.A(_116_),
    .B(_182_),
    .Y(_183_));
 sky130_fd_sc_hd__a22oi_1 _454_ (.A1(\memory[12][6] ),
    .A2(_073_),
    .B1(_080_),
    .B2(\memory[14][6] ),
    .Y(_184_));
 sky130_fd_sc_hd__nand2_1 _455_ (.A(\memory[13][6] ),
    .B(_054_),
    .Y(_185_));
 sky130_fd_sc_hd__a221oi_1 _456_ (.A1(\memory[4][6] ),
    .A2(_067_),
    .B1(_080_),
    .B2(\memory[6][6] ),
    .C1(_060_),
    .Y(_186_));
 sky130_fd_sc_hd__a31oi_2 _457_ (.A1(_078_),
    .A2(_184_),
    .A3(_185_),
    .B1(_186_),
    .Y(_187_));
 sky130_fd_sc_hd__a22oi_1 _458_ (.A1(_086_),
    .A2(\memory[11][6] ),
    .B1(\memory[8][6] ),
    .B2(_067_),
    .Y(_188_));
 sky130_fd_sc_hd__a22oi_2 _459_ (.A1(\memory[10][6] ),
    .A2(_087_),
    .B1(_068_),
    .B2(\memory[9][6] ),
    .Y(_189_));
 sky130_fd_sc_hd__a221oi_1 _460_ (.A1(\memory[2][6] ),
    .A2(_087_),
    .B1(_053_),
    .B2(\memory[1][6] ),
    .C1(_059_),
    .Y(_190_));
 sky130_fd_sc_hd__a311oi_2 _461_ (.A1(_078_),
    .A2(_188_),
    .A3(_189_),
    .B1(_190_),
    .C1(_072_),
    .Y(_191_));
 sky130_fd_sc_hd__a21oi_1 _462_ (.A1(_083_),
    .A2(_187_),
    .B1(_191_),
    .Y(_192_));
 sky130_fd_sc_hd__or3_1 _463_ (.A(\memory[0][6] ),
    .B(_244_),
    .C(_091_),
    .X(_193_));
 sky130_fd_sc_hd__o21ai_0 _464_ (.A1(net21),
    .A2(_050_),
    .B1(_193_),
    .Y(_194_));
 sky130_fd_sc_hd__a21oi_1 _465_ (.A1(_183_),
    .A2(_192_),
    .B1(_194_),
    .Y(_028_));
 sky130_fd_sc_hd__a22oi_2 _466_ (.A1(_085_),
    .A2(\memory[11][7] ),
    .B1(\memory[10][7] ),
    .B2(_079_),
    .Y(_195_));
 sky130_fd_sc_hd__nand2_1 _467_ (.A(\memory[8][7] ),
    .B(_067_),
    .Y(_196_));
 sky130_fd_sc_hd__a21oi_1 _468_ (.A1(_085_),
    .A2(\memory[3][7] ),
    .B1(_059_),
    .Y(_197_));
 sky130_fd_sc_hd__a311oi_2 _469_ (.A1(_060_),
    .A2(_195_),
    .A3(_196_),
    .B1(_197_),
    .C1(_072_),
    .Y(_198_));
 sky130_fd_sc_hd__a222oi_1 _470_ (.A1(_085_),
    .A2(\memory[7][7] ),
    .B1(\memory[6][7] ),
    .B2(_087_),
    .C1(_068_),
    .C2(\memory[5][7] ),
    .Y(_199_));
 sky130_fd_sc_hd__a22o_1 _471_ (.A1(_085_),
    .A2(\memory[15][7] ),
    .B1(\memory[14][7] ),
    .B2(_079_),
    .X(_200_));
 sky130_fd_sc_hd__a221oi_2 _472_ (.A1(\memory[12][7] ),
    .A2(_067_),
    .B1(_068_),
    .B2(\memory[13][7] ),
    .C1(_200_),
    .Y(_201_));
 sky130_fd_sc_hd__o22ai_4 _473_ (.A1(_140_),
    .A2(_199_),
    .B1(_201_),
    .B2(_107_),
    .Y(_202_));
 sky130_fd_sc_hd__a311oi_4 _474_ (.A1(\memory[9][7] ),
    .A2(_054_),
    .A3(_164_),
    .B1(_198_),
    .C1(_202_),
    .Y(_203_));
 sky130_fd_sc_hd__a22oi_1 _475_ (.A1(\memory[2][7] ),
    .A2(_080_),
    .B1(_054_),
    .B2(\memory[1][7] ),
    .Y(_204_));
 sky130_fd_sc_hd__nand3_1 _476_ (.A(_072_),
    .B(\memory[4][7] ),
    .C(_073_),
    .Y(_205_));
 sky130_fd_sc_hd__o21ai_0 _477_ (.A1(_072_),
    .A2(_204_),
    .B1(_205_),
    .Y(_206_));
 sky130_fd_sc_hd__a21oi_1 _478_ (.A1(_094_),
    .A2(_206_),
    .B1(_116_),
    .Y(_207_));
 sky130_fd_sc_hd__or3_1 _479_ (.A(\memory[0][7] ),
    .B(_244_),
    .C(_091_),
    .X(_208_));
 sky130_fd_sc_hd__o21ai_0 _480_ (.A1(net22),
    .A2(_050_),
    .B1(_208_),
    .Y(_209_));
 sky130_fd_sc_hd__a21oi_1 _481_ (.A1(_203_),
    .A2(_207_),
    .B1(_209_),
    .Y(_029_));
 sky130_fd_sc_hd__o211ai_1 _482_ (.A1(_097_),
    .A2(_107_),
    .B1(_052_),
    .C1(_256_),
    .Y(_210_));
 sky130_fd_sc_hd__o21ai_0 _483_ (.A1(_256_),
    .A2(_052_),
    .B1(_210_),
    .Y(_030_));
 sky130_fd_sc_hd__nand2_1 _484_ (.A(_259_),
    .B(_052_),
    .Y(_211_));
 sky130_fd_sc_hd__o21ai_0 _485_ (.A1(_257_),
    .A2(_052_),
    .B1(_211_),
    .Y(_031_));
 sky130_fd_sc_hd__nand2_1 _486_ (.A(_086_),
    .B(_050_),
    .Y(_212_));
 sky130_fd_sc_hd__xnor2_1 _487_ (.A(_083_),
    .B(_212_),
    .Y(_032_));
 sky130_fd_sc_hd__a21oi_1 _488_ (.A1(\rd_ptr[0] ),
    .A2(\rd_ptr[1] ),
    .B1(_086_),
    .Y(_213_));
 sky130_fd_sc_hd__nand2_1 _489_ (.A(_083_),
    .B(_050_),
    .Y(_214_));
 sky130_fd_sc_hd__o21ai_0 _490_ (.A1(_213_),
    .A2(_214_),
    .B1(_078_),
    .Y(_215_));
 sky130_fd_sc_hd__o41ai_1 _491_ (.A1(_256_),
    .A2(_257_),
    .A3(_244_),
    .A4(_140_),
    .B1(_215_),
    .Y(_033_));
 sky130_fd_sc_hd__nand3_1 _492_ (.A(_042_),
    .B(_043_),
    .C(_254_),
    .Y(_216_));
 sky130_fd_sc_hd__nand3_1 _493_ (.A(_246_),
    .B(_243_),
    .C(_216_),
    .Y(_217_));
 sky130_fd_sc_hd__o21ai_0 _494_ (.A1(_246_),
    .A2(_243_),
    .B1(_217_),
    .Y(_034_));
 sky130_fd_sc_hd__nand2_1 _495_ (.A(_249_),
    .B(_243_),
    .Y(_218_));
 sky130_fd_sc_hd__o21ai_0 _496_ (.A1(_247_),
    .A2(_243_),
    .B1(_218_),
    .Y(_035_));
 sky130_fd_sc_hd__nand2_1 _497_ (.A(_254_),
    .B(_243_),
    .Y(_219_));
 sky130_fd_sc_hd__xnor2_1 _498_ (.A(_042_),
    .B(_219_),
    .Y(_036_));
 sky130_fd_sc_hd__a21o_1 _499_ (.A1(\wr_ptr[0] ),
    .A2(\wr_ptr[1] ),
    .B1(_254_),
    .X(_220_));
 sky130_fd_sc_hd__nand3_1 _500_ (.A(_042_),
    .B(_040_),
    .C(_220_),
    .Y(_221_));
 sky130_fd_sc_hd__nor3_1 _501_ (.A(_246_),
    .B(_247_),
    .C(_049_),
    .Y(_222_));
 sky130_fd_sc_hd__a22o_1 _502_ (.A1(_043_),
    .A2(_221_),
    .B1(_222_),
    .B2(_243_),
    .X(_037_));
 sky130_fd_sc_hd__clkbuf_2 _503_ (.A(_245_),
    .X(_223_));
 sky130_fd_sc_hd__xnor2_1 _504_ (.A(net24),
    .B(_223_),
    .Y(_017_));
 sky130_fd_sc_hd__mux2i_1 _505_ (.A0(_242_),
    .A1(_239_),
    .S(_223_),
    .Y(_018_));
 sky130_fd_sc_hd__xor2_1 _506_ (.A(_270_),
    .B(_241_),
    .X(_224_));
 sky130_fd_sc_hd__nand2_1 _507_ (.A(net26),
    .B(_223_),
    .Y(_225_));
 sky130_fd_sc_hd__o21ai_0 _508_ (.A1(_223_),
    .A2(_224_),
    .B1(_225_),
    .Y(_019_));
 sky130_fd_sc_hd__nand3_1 _509_ (.A(net24),
    .B(_268_),
    .C(_274_),
    .Y(_226_));
 sky130_fd_sc_hd__a21oi_1 _510_ (.A1(_270_),
    .A2(_267_),
    .B1(_269_),
    .Y(_227_));
 sky130_fd_sc_hd__nand2_1 _511_ (.A(_226_),
    .B(_227_),
    .Y(_228_));
 sky130_fd_sc_hd__xnor2_1 _512_ (.A(_272_),
    .B(_228_),
    .Y(_229_));
 sky130_fd_sc_hd__nand2_1 _513_ (.A(net27),
    .B(_223_),
    .Y(_230_));
 sky130_fd_sc_hd__o21ai_0 _514_ (.A1(_223_),
    .A2(_229_),
    .B1(_230_),
    .Y(_020_));
 sky130_fd_sc_hd__nor2_1 _515_ (.A(_266_),
    .B(_223_),
    .Y(_231_));
 sky130_fd_sc_hd__nor2_1 _516_ (.A(_240_),
    .B(_223_),
    .Y(_232_));
 sky130_fd_sc_hd__inv_1 _517_ (.A(_241_),
    .Y(_233_));
 sky130_fd_sc_hd__a21o_1 _518_ (.A1(_233_),
    .A2(_274_),
    .B1(_269_),
    .X(_234_));
 sky130_fd_sc_hd__a21oi_1 _519_ (.A1(_272_),
    .A2(_234_),
    .B1(_271_),
    .Y(_235_));
 sky130_fd_sc_hd__mux2i_1 _520_ (.A0(_231_),
    .A1(_232_),
    .S(_235_),
    .Y(_236_));
 sky130_fd_sc_hd__xnor2_1 _521_ (.A(net28),
    .B(_236_),
    .Y(_021_));
 sky130_fd_sc_hd__o21a_1 _522_ (.A1(net25),
    .A2(net24),
    .B1(net26),
    .X(_237_));
 sky130_fd_sc_hd__nor3_1 _523_ (.A(net27),
    .B(net28),
    .C(_237_),
    .Y(net13));
 sky130_fd_sc_hd__nand2_1 _524_ (.A(net27),
    .B(net26),
    .Y(_238_));
 sky130_fd_sc_hd__nand2_1 _525_ (.A(_038_),
    .B(_238_),
    .Y(net14));
 sky130_fd_sc_hd__fa_1 _526_ (.A(_016_),
    .B(_239_),
    .CIN(_240_),
    .COUT(_241_),
    .SUM(_242_));
 sky130_fd_sc_hd__ha_1 _527_ (.A(_243_),
    .B(_244_),
    .COUT(_240_),
    .SUM(_245_));
 sky130_fd_sc_hd__ha_1 _528_ (.A(_246_),
    .B(_247_),
    .COUT(_248_),
    .SUM(_249_));
 sky130_fd_sc_hd__ha_1 _529_ (.A(_246_),
    .B(\wr_ptr[1] ),
    .COUT(_250_),
    .SUM(_251_));
 sky130_fd_sc_hd__ha_1 _530_ (.A(\wr_ptr[0] ),
    .B(_247_),
    .COUT(_252_),
    .SUM(_253_));
 sky130_fd_sc_hd__ha_1 _531_ (.A(\wr_ptr[0] ),
    .B(\wr_ptr[1] ),
    .COUT(_254_),
    .SUM(_255_));
 sky130_fd_sc_hd__ha_2 _532_ (.A(_256_),
    .B(_257_),
    .COUT(_258_),
    .SUM(_259_));
 sky130_fd_sc_hd__ha_2 _533_ (.A(_256_),
    .B(\rd_ptr[1] ),
    .COUT(_260_),
    .SUM(_261_));
 sky130_fd_sc_hd__ha_1 _534_ (.A(\rd_ptr[0] ),
    .B(_257_),
    .COUT(_262_),
    .SUM(_263_));
 sky130_fd_sc_hd__ha_2 _535_ (.A(\rd_ptr[0] ),
    .B(\rd_ptr[1] ),
    .COUT(_264_),
    .SUM(_265_));
 sky130_fd_sc_hd__ha_1 _536_ (.A(net25),
    .B(_266_),
    .COUT(_267_),
    .SUM(_268_));
 sky130_fd_sc_hd__ha_1 _537_ (.A(net26),
    .B(_266_),
    .COUT(_269_),
    .SUM(_270_));
 sky130_fd_sc_hd__ha_1 _538_ (.A(net27),
    .B(_266_),
    .COUT(_271_),
    .SUM(_272_));
 sky130_fd_sc_hd__ha_1 _539_ (.A(net26),
    .B(_266_),
    .COUT(_273_),
    .SUM(_274_));
 sky130_fd_sc_hd__dfrtp_2 \count[0]$_DFFE_PN0P_  (.D(_017_),
    .Q(net24),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \count[1]$_DFFE_PN0P_  (.D(_018_),
    .Q(net25),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \count[2]$_DFFE_PN0P_  (.D(_019_),
    .Q(net26),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \count[3]$_DFFE_PN0P_  (.D(_020_),
    .Q(net27),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \count[4]$_DFFE_PN0P_  (.D(_021_),
    .Q(net28),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out[0]$_DFFE_PN0P_  (.D(_022_),
    .Q(net15),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out[1]$_DFFE_PN0P_  (.D(_023_),
    .Q(net16),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out[2]$_DFFE_PN0P_  (.D(_024_),
    .Q(net17),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out[3]$_DFFE_PN0P_  (.D(_025_),
    .Q(net18),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out[4]$_DFFE_PN0P_  (.D(_026_),
    .Q(net19),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out[5]$_DFFE_PN0P_  (.D(_027_),
    .Q(net20),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out[6]$_DFFE_PN0P_  (.D(_028_),
    .Q(net21),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \data_out[7]$_DFFE_PN0P_  (.D(_029_),
    .Q(net22),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[0][0]$_DFFE_PP_  (.D(net2),
    .DE(_015_),
    .Q(\memory[0][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[0][1]$_DFFE_PP_  (.D(net3),
    .DE(_015_),
    .Q(\memory[0][1] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[0][2]$_DFFE_PP_  (.D(net4),
    .DE(_015_),
    .Q(\memory[0][2] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[0][3]$_DFFE_PP_  (.D(net5),
    .DE(_015_),
    .Q(\memory[0][3] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[0][4]$_DFFE_PP_  (.D(net6),
    .DE(_015_),
    .Q(\memory[0][4] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[0][5]$_DFFE_PP_  (.D(net7),
    .DE(_015_),
    .Q(\memory[0][5] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[0][6]$_DFFE_PP_  (.D(net8),
    .DE(_015_),
    .Q(\memory[0][6] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[0][7]$_DFFE_PP_  (.D(net9),
    .DE(_015_),
    .Q(\memory[0][7] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[10][0]$_DFFE_PP_  (.D(net2),
    .DE(_005_),
    .Q(\memory[10][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[10][1]$_DFFE_PP_  (.D(net3),
    .DE(_005_),
    .Q(\memory[10][1] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[10][2]$_DFFE_PP_  (.D(net4),
    .DE(_005_),
    .Q(\memory[10][2] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[10][3]$_DFFE_PP_  (.D(net5),
    .DE(_005_),
    .Q(\memory[10][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[10][4]$_DFFE_PP_  (.D(net6),
    .DE(_005_),
    .Q(\memory[10][4] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[10][5]$_DFFE_PP_  (.D(net7),
    .DE(_005_),
    .Q(\memory[10][5] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[10][6]$_DFFE_PP_  (.D(net8),
    .DE(_005_),
    .Q(\memory[10][6] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[10][7]$_DFFE_PP_  (.D(net9),
    .DE(_005_),
    .Q(\memory[10][7] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[11][0]$_DFFE_PP_  (.D(net2),
    .DE(_004_),
    .Q(\memory[11][0] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[11][1]$_DFFE_PP_  (.D(net3),
    .DE(_004_),
    .Q(\memory[11][1] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[11][2]$_DFFE_PP_  (.D(net4),
    .DE(_004_),
    .Q(\memory[11][2] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[11][3]$_DFFE_PP_  (.D(net5),
    .DE(_004_),
    .Q(\memory[11][3] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[11][4]$_DFFE_PP_  (.D(net6),
    .DE(_004_),
    .Q(\memory[11][4] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[11][5]$_DFFE_PP_  (.D(net7),
    .DE(_004_),
    .Q(\memory[11][5] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[11][6]$_DFFE_PP_  (.D(net8),
    .DE(_004_),
    .Q(\memory[11][6] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[11][7]$_DFFE_PP_  (.D(net9),
    .DE(_004_),
    .Q(\memory[11][7] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[12][0]$_DFFE_PP_  (.D(net2),
    .DE(_003_),
    .Q(\memory[12][0] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[12][1]$_DFFE_PP_  (.D(net3),
    .DE(_003_),
    .Q(\memory[12][1] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[12][2]$_DFFE_PP_  (.D(net4),
    .DE(_003_),
    .Q(\memory[12][2] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[12][3]$_DFFE_PP_  (.D(net5),
    .DE(_003_),
    .Q(\memory[12][3] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[12][4]$_DFFE_PP_  (.D(net6),
    .DE(_003_),
    .Q(\memory[12][4] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[12][5]$_DFFE_PP_  (.D(net7),
    .DE(_003_),
    .Q(\memory[12][5] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[12][6]$_DFFE_PP_  (.D(net8),
    .DE(_003_),
    .Q(\memory[12][6] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[12][7]$_DFFE_PP_  (.D(net9),
    .DE(_003_),
    .Q(\memory[12][7] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[13][0]$_DFFE_PP_  (.D(net2),
    .DE(_002_),
    .Q(\memory[13][0] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[13][1]$_DFFE_PP_  (.D(net3),
    .DE(_002_),
    .Q(\memory[13][1] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[13][2]$_DFFE_PP_  (.D(net4),
    .DE(_002_),
    .Q(\memory[13][2] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[13][3]$_DFFE_PP_  (.D(net5),
    .DE(_002_),
    .Q(\memory[13][3] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[13][4]$_DFFE_PP_  (.D(net6),
    .DE(_002_),
    .Q(\memory[13][4] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[13][5]$_DFFE_PP_  (.D(net7),
    .DE(_002_),
    .Q(\memory[13][5] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[13][6]$_DFFE_PP_  (.D(net8),
    .DE(_002_),
    .Q(\memory[13][6] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[13][7]$_DFFE_PP_  (.D(net9),
    .DE(_002_),
    .Q(\memory[13][7] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[14][0]$_DFFE_PP_  (.D(net2),
    .DE(_001_),
    .Q(\memory[14][0] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[14][1]$_DFFE_PP_  (.D(net3),
    .DE(_001_),
    .Q(\memory[14][1] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[14][2]$_DFFE_PP_  (.D(net4),
    .DE(_001_),
    .Q(\memory[14][2] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[14][3]$_DFFE_PP_  (.D(net5),
    .DE(_001_),
    .Q(\memory[14][3] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[14][4]$_DFFE_PP_  (.D(net6),
    .DE(_001_),
    .Q(\memory[14][4] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[14][5]$_DFFE_PP_  (.D(net7),
    .DE(_001_),
    .Q(\memory[14][5] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[14][6]$_DFFE_PP_  (.D(net8),
    .DE(_001_),
    .Q(\memory[14][6] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[14][7]$_DFFE_PP_  (.D(net9),
    .DE(_001_),
    .Q(\memory[14][7] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[15][0]$_DFFE_PP_  (.D(net2),
    .DE(_000_),
    .Q(\memory[15][0] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[15][1]$_DFFE_PP_  (.D(net3),
    .DE(_000_),
    .Q(\memory[15][1] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[15][2]$_DFFE_PP_  (.D(net4),
    .DE(_000_),
    .Q(\memory[15][2] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[15][3]$_DFFE_PP_  (.D(net5),
    .DE(_000_),
    .Q(\memory[15][3] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[15][4]$_DFFE_PP_  (.D(net6),
    .DE(_000_),
    .Q(\memory[15][4] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[15][5]$_DFFE_PP_  (.D(net7),
    .DE(_000_),
    .Q(\memory[15][5] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[15][6]$_DFFE_PP_  (.D(net8),
    .DE(_000_),
    .Q(\memory[15][6] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[15][7]$_DFFE_PP_  (.D(net9),
    .DE(_000_),
    .Q(\memory[15][7] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[1][0]$_DFFE_PP_  (.D(net2),
    .DE(_014_),
    .Q(\memory[1][0] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[1][1]$_DFFE_PP_  (.D(net3),
    .DE(_014_),
    .Q(\memory[1][1] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[1][2]$_DFFE_PP_  (.D(net4),
    .DE(_014_),
    .Q(\memory[1][2] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[1][3]$_DFFE_PP_  (.D(net5),
    .DE(_014_),
    .Q(\memory[1][3] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[1][4]$_DFFE_PP_  (.D(net6),
    .DE(_014_),
    .Q(\memory[1][4] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[1][5]$_DFFE_PP_  (.D(net7),
    .DE(_014_),
    .Q(\memory[1][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[1][6]$_DFFE_PP_  (.D(net8),
    .DE(_014_),
    .Q(\memory[1][6] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[1][7]$_DFFE_PP_  (.D(net9),
    .DE(_014_),
    .Q(\memory[1][7] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[2][0]$_DFFE_PP_  (.D(net2),
    .DE(_013_),
    .Q(\memory[2][0] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[2][1]$_DFFE_PP_  (.D(net3),
    .DE(_013_),
    .Q(\memory[2][1] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[2][2]$_DFFE_PP_  (.D(net4),
    .DE(_013_),
    .Q(\memory[2][2] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[2][3]$_DFFE_PP_  (.D(net5),
    .DE(_013_),
    .Q(\memory[2][3] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[2][4]$_DFFE_PP_  (.D(net6),
    .DE(_013_),
    .Q(\memory[2][4] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[2][5]$_DFFE_PP_  (.D(net7),
    .DE(_013_),
    .Q(\memory[2][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[2][6]$_DFFE_PP_  (.D(net8),
    .DE(_013_),
    .Q(\memory[2][6] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[2][7]$_DFFE_PP_  (.D(net9),
    .DE(_013_),
    .Q(\memory[2][7] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[3][0]$_DFFE_PP_  (.D(net2),
    .DE(_012_),
    .Q(\memory[3][0] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[3][1]$_DFFE_PP_  (.D(net3),
    .DE(_012_),
    .Q(\memory[3][1] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[3][2]$_DFFE_PP_  (.D(net4),
    .DE(_012_),
    .Q(\memory[3][2] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[3][3]$_DFFE_PP_  (.D(net5),
    .DE(_012_),
    .Q(\memory[3][3] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[3][4]$_DFFE_PP_  (.D(net6),
    .DE(_012_),
    .Q(\memory[3][4] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[3][5]$_DFFE_PP_  (.D(net7),
    .DE(_012_),
    .Q(\memory[3][5] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[3][6]$_DFFE_PP_  (.D(net8),
    .DE(_012_),
    .Q(\memory[3][6] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[3][7]$_DFFE_PP_  (.D(net9),
    .DE(_012_),
    .Q(\memory[3][7] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[4][0]$_DFFE_PP_  (.D(net2),
    .DE(_011_),
    .Q(\memory[4][0] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[4][1]$_DFFE_PP_  (.D(net3),
    .DE(_011_),
    .Q(\memory[4][1] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[4][2]$_DFFE_PP_  (.D(net4),
    .DE(_011_),
    .Q(\memory[4][2] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[4][3]$_DFFE_PP_  (.D(net5),
    .DE(_011_),
    .Q(\memory[4][3] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[4][4]$_DFFE_PP_  (.D(net6),
    .DE(_011_),
    .Q(\memory[4][4] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[4][5]$_DFFE_PP_  (.D(net7),
    .DE(_011_),
    .Q(\memory[4][5] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[4][6]$_DFFE_PP_  (.D(net8),
    .DE(_011_),
    .Q(\memory[4][6] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[4][7]$_DFFE_PP_  (.D(net9),
    .DE(_011_),
    .Q(\memory[4][7] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[5][0]$_DFFE_PP_  (.D(net2),
    .DE(_010_),
    .Q(\memory[5][0] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[5][1]$_DFFE_PP_  (.D(net3),
    .DE(_010_),
    .Q(\memory[5][1] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[5][2]$_DFFE_PP_  (.D(net4),
    .DE(_010_),
    .Q(\memory[5][2] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[5][3]$_DFFE_PP_  (.D(net5),
    .DE(_010_),
    .Q(\memory[5][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[5][4]$_DFFE_PP_  (.D(net6),
    .DE(_010_),
    .Q(\memory[5][4] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[5][5]$_DFFE_PP_  (.D(net7),
    .DE(_010_),
    .Q(\memory[5][5] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[5][6]$_DFFE_PP_  (.D(net8),
    .DE(_010_),
    .Q(\memory[5][6] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[5][7]$_DFFE_PP_  (.D(net9),
    .DE(_010_),
    .Q(\memory[5][7] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[6][0]$_DFFE_PP_  (.D(net2),
    .DE(_009_),
    .Q(\memory[6][0] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[6][1]$_DFFE_PP_  (.D(net3),
    .DE(_009_),
    .Q(\memory[6][1] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[6][2]$_DFFE_PP_  (.D(net4),
    .DE(_009_),
    .Q(\memory[6][2] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[6][3]$_DFFE_PP_  (.D(net5),
    .DE(_009_),
    .Q(\memory[6][3] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[6][4]$_DFFE_PP_  (.D(net6),
    .DE(_009_),
    .Q(\memory[6][4] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[6][5]$_DFFE_PP_  (.D(net7),
    .DE(_009_),
    .Q(\memory[6][5] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[6][6]$_DFFE_PP_  (.D(net8),
    .DE(_009_),
    .Q(\memory[6][6] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[6][7]$_DFFE_PP_  (.D(net9),
    .DE(_009_),
    .Q(\memory[6][7] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[7][0]$_DFFE_PP_  (.D(net2),
    .DE(_008_),
    .Q(\memory[7][0] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[7][1]$_DFFE_PP_  (.D(net3),
    .DE(_008_),
    .Q(\memory[7][1] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[7][2]$_DFFE_PP_  (.D(net4),
    .DE(_008_),
    .Q(\memory[7][2] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[7][3]$_DFFE_PP_  (.D(net5),
    .DE(_008_),
    .Q(\memory[7][3] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[7][4]$_DFFE_PP_  (.D(net6),
    .DE(_008_),
    .Q(\memory[7][4] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[7][5]$_DFFE_PP_  (.D(net7),
    .DE(_008_),
    .Q(\memory[7][5] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[7][6]$_DFFE_PP_  (.D(net8),
    .DE(_008_),
    .Q(\memory[7][6] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[7][7]$_DFFE_PP_  (.D(net9),
    .DE(_008_),
    .Q(\memory[7][7] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[8][0]$_DFFE_PP_  (.D(net2),
    .DE(_007_),
    .Q(\memory[8][0] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[8][1]$_DFFE_PP_  (.D(net3),
    .DE(_007_),
    .Q(\memory[8][1] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[8][2]$_DFFE_PP_  (.D(net4),
    .DE(_007_),
    .Q(\memory[8][2] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[8][3]$_DFFE_PP_  (.D(net5),
    .DE(_007_),
    .Q(\memory[8][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[8][4]$_DFFE_PP_  (.D(net6),
    .DE(_007_),
    .Q(\memory[8][4] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[8][5]$_DFFE_PP_  (.D(net7),
    .DE(_007_),
    .Q(\memory[8][5] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[8][6]$_DFFE_PP_  (.D(net8),
    .DE(_007_),
    .Q(\memory[8][6] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[8][7]$_DFFE_PP_  (.D(net9),
    .DE(_007_),
    .Q(\memory[8][7] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[9][0]$_DFFE_PP_  (.D(net2),
    .DE(_006_),
    .Q(\memory[9][0] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[9][1]$_DFFE_PP_  (.D(net3),
    .DE(_006_),
    .Q(\memory[9][1] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[9][2]$_DFFE_PP_  (.D(net4),
    .DE(_006_),
    .Q(\memory[9][2] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[9][3]$_DFFE_PP_  (.D(net5),
    .DE(_006_),
    .Q(\memory[9][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[9][4]$_DFFE_PP_  (.D(net6),
    .DE(_006_),
    .Q(\memory[9][4] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[9][5]$_DFFE_PP_  (.D(net7),
    .DE(_006_),
    .Q(\memory[9][5] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[9][6]$_DFFE_PP_  (.D(net8),
    .DE(_006_),
    .Q(\memory[9][6] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \memory[9][7]$_DFFE_PP_  (.D(net9),
    .DE(_006_),
    .Q(\memory[9][7] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[0]$_DFFE_PN0P_  (.D(_030_),
    .Q(\rd_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[1]$_DFFE_PN0P_  (.D(_031_),
    .Q(\rd_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \rd_ptr[2]$_DFFE_PN0P_  (.D(_032_),
    .Q(\rd_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[3]$_DFFE_PN0P_  (.D(_033_),
    .Q(\rd_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[0]$_DFFE_PN0P_  (.D(_034_),
    .Q(\wr_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[1]$_DFFE_PN0P_  (.D(_035_),
    .Q(\wr_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[2]$_DFFE_PN0P_  (.D(_036_),
    .Q(\wr_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[3]$_DFFE_PN0P_  (.D(_037_),
    .Q(\wr_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__buf_8 hold1 (.A(net11),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_135 ();
 sky130_fd_sc_hd__buf_4 input1 (.A(net33),
    .X(net2));
 sky130_fd_sc_hd__buf_4 input2 (.A(data_in[1]),
    .X(net3));
 sky130_fd_sc_hd__buf_4 input3 (.A(data_in[2]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input4 (.A(data_in[3]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input5 (.A(data_in[4]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_8 input6 (.A(net32),
    .X(net7));
 sky130_fd_sc_hd__buf_6 input7 (.A(net31),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input8 (.A(data_in[7]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(rd_en),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(net30),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(wr_en),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 output12 (.A(net13),
    .X(almost_empty));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net14),
    .X(almost_full));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net15),
    .X(data_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net16),
    .X(data_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net17),
    .X(data_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net18),
    .X(data_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net19),
    .X(data_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net20),
    .X(data_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net21),
    .X(data_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net22),
    .X(data_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net23),
    .X(empty));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net24),
    .X(fill_level[0]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net25),
    .X(fill_level[1]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net26),
    .X(fill_level[2]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net27),
    .X(fill_level[3]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net28),
    .X(fill_level[4]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net29),
    .X(full));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload0 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload1 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__inv_6 clkload2 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload3 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload4 (.A(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload5 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload6 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload7 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__inv_6 clkload8 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload9 (.A(clknet_4_10_0_clk));
 sky130_fd_sc_hd__inv_6 clkload10 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__inv_8 clkload11 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__inv_6 clkload12 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__inv_8 clkload13 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload14 (.A(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net30));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(data_in[6]),
    .X(net31));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(data_in[5]),
    .X(net32));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(data_in[0]),
    .X(net33));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_76 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_87 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_126 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_182 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_102 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_219 ();
endmodule
