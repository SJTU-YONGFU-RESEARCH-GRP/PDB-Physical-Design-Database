module arbiter_rr (active,
    clk,
    rst_n,
    grant,
    request);
 output active;
 input clk;
 input rst_n;
 output [3:0] grant;
 input [3:0] request;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire \priority_ptr[0] ;
 wire \priority_ptr[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 INV_X1 _082_ (.A(net5),
    .ZN(_006_));
 NOR4_X4 _083_ (.A1(net1),
    .A2(net2),
    .A3(net3),
    .A4(net4),
    .ZN(_007_));
 OR2_X1 _084_ (.A1(_006_),
    .A2(_007_),
    .ZN(_008_));
 BUF_X2 _085_ (.A(\priority_ptr[1] ),
    .Z(_009_));
 MUX2_X1 _086_ (.A(net2),
    .B(net4),
    .S(_009_),
    .Z(_010_));
 MUX2_X1 _087_ (.A(net1),
    .B(net3),
    .S(_009_),
    .Z(_011_));
 BUF_X2 _088_ (.A(\priority_ptr[0] ),
    .Z(_012_));
 INV_X1 _089_ (.A(_012_),
    .ZN(_013_));
 MUX2_X1 _090_ (.A(_010_),
    .B(_011_),
    .S(_013_),
    .Z(_014_));
 BUF_X4 _091_ (.A(_014_),
    .Z(_015_));
 BUF_X4 _092_ (.A(_067_),
    .Z(_016_));
 MUX2_X1 _093_ (.A(net4),
    .B(net2),
    .S(_016_),
    .Z(_017_));
 MUX2_X1 _094_ (.A(net3),
    .B(net1),
    .S(_016_),
    .Z(_018_));
 MUX2_X1 _095_ (.A(_017_),
    .B(_018_),
    .S(_012_),
    .Z(_019_));
 BUF_X8 _096_ (.A(_019_),
    .Z(_020_));
 MUX2_X1 _097_ (.A(net3),
    .B(net1),
    .S(_009_),
    .Z(_021_));
 NOR2_X1 _098_ (.A1(_012_),
    .A2(_021_),
    .ZN(_022_));
 MUX2_X1 _099_ (.A(net4),
    .B(net2),
    .S(_009_),
    .Z(_023_));
 NOR2_X1 _100_ (.A1(_013_),
    .A2(_023_),
    .ZN(_024_));
 NOR3_X2 _101_ (.A1(_022_),
    .A2(_024_),
    .A3(_020_),
    .ZN(_025_));
 AOI22_X1 _102_ (.A1(_076_),
    .A2(_020_),
    .B1(_025_),
    .B2(_072_),
    .ZN(_026_));
 OR2_X1 _103_ (.A1(_015_),
    .A2(_026_),
    .ZN(_027_));
 MUX2_X1 _104_ (.A(_021_),
    .B(_023_),
    .S(_012_),
    .Z(_028_));
 MUX2_X1 _105_ (.A(net2),
    .B(net4),
    .S(_016_),
    .Z(_029_));
 NOR2_X1 _106_ (.A1(_012_),
    .A2(_029_),
    .ZN(_030_));
 MUX2_X1 _107_ (.A(net1),
    .B(net3),
    .S(_016_),
    .Z(_031_));
 NOR2_X1 _108_ (.A1(_013_),
    .A2(_031_),
    .ZN(_032_));
 NOR3_X1 _109_ (.A1(_028_),
    .A2(_030_),
    .A3(_032_),
    .ZN(_033_));
 NOR2_X1 _110_ (.A1(_015_),
    .A2(_020_),
    .ZN(_034_));
 AND2_X1 _111_ (.A1(_033_),
    .A2(_034_),
    .ZN(_035_));
 AOI22_X1 _112_ (.A1(_066_),
    .A2(_015_),
    .B1(_035_),
    .B2(_080_),
    .ZN(_036_));
 AOI21_X1 _113_ (.A(_008_),
    .B1(_027_),
    .B2(_036_),
    .ZN(_000_));
 AOI22_X1 _114_ (.A1(_072_),
    .A2(_020_),
    .B1(_025_),
    .B2(_080_),
    .ZN(_037_));
 OR2_X1 _115_ (.A1(_015_),
    .A2(_037_),
    .ZN(_038_));
 AOI22_X1 _116_ (.A1(_074_),
    .A2(_015_),
    .B1(_035_),
    .B2(_068_),
    .ZN(_039_));
 AOI21_X1 _117_ (.A(_008_),
    .B1(_038_),
    .B2(_039_),
    .ZN(_001_));
 AOI22_X1 _118_ (.A1(_080_),
    .A2(_020_),
    .B1(_025_),
    .B2(_068_),
    .ZN(_040_));
 OR2_X1 _119_ (.A1(_015_),
    .A2(_040_),
    .ZN(_041_));
 AOI22_X1 _120_ (.A1(_070_),
    .A2(_015_),
    .B1(_035_),
    .B2(_076_),
    .ZN(_042_));
 AOI21_X1 _121_ (.A(_008_),
    .B1(_041_),
    .B2(_042_),
    .ZN(_002_));
 AOI22_X1 _122_ (.A1(_068_),
    .A2(_020_),
    .B1(_025_),
    .B2(_076_),
    .ZN(_043_));
 OR2_X1 _123_ (.A1(_015_),
    .A2(_043_),
    .ZN(_044_));
 AOI22_X1 _124_ (.A1(_078_),
    .A2(_015_),
    .B1(_035_),
    .B2(_072_),
    .ZN(_045_));
 AOI21_X1 _125_ (.A(_008_),
    .B1(_044_),
    .B2(_045_),
    .ZN(_003_));
 NOR2_X1 _126_ (.A1(_007_),
    .A2(_020_),
    .ZN(_046_));
 INV_X1 _127_ (.A(_064_),
    .ZN(_047_));
 NOR4_X1 _128_ (.A1(_047_),
    .A2(_022_),
    .A3(_024_),
    .A4(_015_),
    .ZN(_048_));
 NOR3_X1 _129_ (.A1(_012_),
    .A2(_021_),
    .A3(_029_),
    .ZN(_049_));
 OAI21_X1 _130_ (.A(_046_),
    .B1(_048_),
    .B2(_049_),
    .ZN(_050_));
 OR2_X1 _131_ (.A1(_012_),
    .A2(_011_),
    .ZN(_051_));
 OAI21_X1 _132_ (.A(_051_),
    .B1(_007_),
    .B2(_013_),
    .ZN(_052_));
 NOR2_X1 _133_ (.A1(_013_),
    .A2(_010_),
    .ZN(_053_));
 OAI21_X1 _134_ (.A(_053_),
    .B1(_020_),
    .B2(_033_),
    .ZN(_054_));
 NAND4_X1 _135_ (.A1(net5),
    .A2(_050_),
    .A3(_052_),
    .A4(_054_),
    .ZN(_004_));
 AOI21_X1 _136_ (.A(_006_),
    .B1(_007_),
    .B2(_009_),
    .ZN(_055_));
 OR3_X1 _137_ (.A1(_047_),
    .A2(_030_),
    .A3(_032_),
    .ZN(_056_));
 NOR2_X1 _138_ (.A1(_028_),
    .A2(_020_),
    .ZN(_057_));
 AOI221_X2 _139_ (.A(_014_),
    .B1(_056_),
    .B2(_057_),
    .C1(_020_),
    .C2(_064_),
    .ZN(_058_));
 XOR2_X1 _140_ (.A(_016_),
    .B(_058_),
    .Z(_059_));
 OAI21_X1 _141_ (.A(_055_),
    .B1(_059_),
    .B2(_007_),
    .ZN(_005_));
 OR4_X1 _142_ (.A1(net8),
    .A2(net7),
    .A3(net10),
    .A4(net9),
    .ZN(net6));
 HA_X1 _143_ (.A(_064_),
    .B(_065_),
    .CO(_066_),
    .S(_067_));
 HA_X1 _144_ (.A(_064_),
    .B(_065_),
    .CO(_068_),
    .S(_069_));
 HA_X1 _145_ (.A(_064_),
    .B(\priority_ptr[1] ),
    .CO(_070_),
    .S(_071_));
 HA_X1 _146_ (.A(_064_),
    .B(\priority_ptr[1] ),
    .CO(_072_),
    .S(_073_));
 HA_X1 _147_ (.A(\priority_ptr[0] ),
    .B(_065_),
    .CO(_074_),
    .S(_075_));
 HA_X1 _148_ (.A(\priority_ptr[0] ),
    .B(_065_),
    .CO(_076_),
    .S(_077_));
 HA_X1 _149_ (.A(\priority_ptr[0] ),
    .B(\priority_ptr[1] ),
    .CO(_078_),
    .S(_079_));
 HA_X1 _150_ (.A(\priority_ptr[0] ),
    .B(\priority_ptr[1] ),
    .CO(_080_),
    .S(_081_));
 DFF_X1 \grant[0]$_SDFF_PN0_  (.D(_000_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net7),
    .QN(_063_));
 DFF_X1 \grant[1]$_SDFF_PN0_  (.D(_001_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net8),
    .QN(_062_));
 DFF_X1 \grant[2]$_SDFF_PN0_  (.D(_002_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net9),
    .QN(_061_));
 DFF_X1 \grant[3]$_SDFF_PN0_  (.D(_003_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net10),
    .QN(_060_));
 DFF_X2 \priority_ptr[0]$_SDFFE_PN1P_  (.D(_004_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\priority_ptr[0] ),
    .QN(_064_));
 DFF_X2 \priority_ptr[1]$_SDFFE_PN1P_  (.D(_005_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\priority_ptr[1] ),
    .QN(_065_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_49 ();
 CLKBUF_X2 input1 (.A(request[0]),
    .Z(net1));
 CLKBUF_X2 input2 (.A(request[1]),
    .Z(net2));
 CLKBUF_X2 input3 (.A(request[2]),
    .Z(net3));
 CLKBUF_X2 input4 (.A(request[3]),
    .Z(net4));
 BUF_X1 input5 (.A(rst_n),
    .Z(net5));
 BUF_X1 output6 (.A(net6),
    .Z(active));
 BUF_X1 output7 (.A(net7),
    .Z(grant[0]));
 BUF_X1 output8 (.A(net8),
    .Z(grant[1]));
 BUF_X1 output9 (.A(net9),
    .Z(grant[2]));
 BUF_X1 output10 (.A(net10),
    .Z(grant[3]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 CLKBUF_X1 clkload0 (.A(clknet_1_0__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X16 FILLER_0_33 ();
 FILLCELL_X8 FILLER_0_49 ();
 FILLCELL_X4 FILLER_0_57 ();
 FILLCELL_X1 FILLER_0_61 ();
 FILLCELL_X16 FILLER_0_78 ();
 FILLCELL_X1 FILLER_0_94 ();
 FILLCELL_X32 FILLER_0_98 ();
 FILLCELL_X32 FILLER_0_130 ();
 FILLCELL_X16 FILLER_0_162 ();
 FILLCELL_X8 FILLER_0_178 ();
 FILLCELL_X2 FILLER_0_186 ();
 FILLCELL_X1 FILLER_0_188 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X4 FILLER_1_65 ();
 FILLCELL_X2 FILLER_1_69 ();
 FILLCELL_X32 FILLER_1_106 ();
 FILLCELL_X32 FILLER_1_138 ();
 FILLCELL_X16 FILLER_1_170 ();
 FILLCELL_X2 FILLER_1_186 ();
 FILLCELL_X1 FILLER_1_188 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X4 FILLER_2_65 ();
 FILLCELL_X4 FILLER_2_110 ();
 FILLCELL_X1 FILLER_2_117 ();
 FILLCELL_X1 FILLER_2_121 ();
 FILLCELL_X32 FILLER_2_127 ();
 FILLCELL_X16 FILLER_2_159 ();
 FILLCELL_X8 FILLER_2_175 ();
 FILLCELL_X4 FILLER_2_183 ();
 FILLCELL_X2 FILLER_2_187 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X4 FILLER_3_65 ();
 FILLCELL_X2 FILLER_3_90 ();
 FILLCELL_X1 FILLER_3_92 ();
 FILLCELL_X1 FILLER_3_116 ();
 FILLCELL_X4 FILLER_3_140 ();
 FILLCELL_X2 FILLER_3_144 ();
 FILLCELL_X32 FILLER_3_153 ();
 FILLCELL_X4 FILLER_3_185 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X2 FILLER_4_105 ();
 FILLCELL_X2 FILLER_4_110 ();
 FILLCELL_X1 FILLER_4_112 ();
 FILLCELL_X2 FILLER_4_117 ();
 FILLCELL_X1 FILLER_4_119 ();
 FILLCELL_X32 FILLER_4_143 ();
 FILLCELL_X8 FILLER_4_175 ();
 FILLCELL_X4 FILLER_4_183 ();
 FILLCELL_X2 FILLER_4_187 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_104 ();
 FILLCELL_X32 FILLER_5_136 ();
 FILLCELL_X16 FILLER_5_168 ();
 FILLCELL_X4 FILLER_5_184 ();
 FILLCELL_X1 FILLER_5_188 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X16 FILLER_6_65 ();
 FILLCELL_X8 FILLER_6_81 ();
 FILLCELL_X4 FILLER_6_89 ();
 FILLCELL_X32 FILLER_6_107 ();
 FILLCELL_X32 FILLER_6_139 ();
 FILLCELL_X16 FILLER_6_171 ();
 FILLCELL_X2 FILLER_6_187 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X16 FILLER_7_65 ();
 FILLCELL_X8 FILLER_7_81 ();
 FILLCELL_X4 FILLER_7_89 ();
 FILLCELL_X8 FILLER_7_101 ();
 FILLCELL_X1 FILLER_7_109 ();
 FILLCELL_X16 FILLER_7_114 ();
 FILLCELL_X4 FILLER_7_130 ();
 FILLCELL_X4 FILLER_7_144 ();
 FILLCELL_X1 FILLER_7_148 ();
 FILLCELL_X16 FILLER_7_169 ();
 FILLCELL_X4 FILLER_7_185 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X2 FILLER_8_97 ();
 FILLCELL_X8 FILLER_8_116 ();
 FILLCELL_X1 FILLER_8_124 ();
 FILLCELL_X16 FILLER_8_171 ();
 FILLCELL_X2 FILLER_8_187 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X16 FILLER_9_65 ();
 FILLCELL_X8 FILLER_9_81 ();
 FILLCELL_X4 FILLER_9_108 ();
 FILLCELL_X2 FILLER_9_112 ();
 FILLCELL_X1 FILLER_9_114 ();
 FILLCELL_X1 FILLER_9_123 ();
 FILLCELL_X4 FILLER_9_158 ();
 FILLCELL_X2 FILLER_9_162 ();
 FILLCELL_X16 FILLER_9_172 ();
 FILLCELL_X1 FILLER_9_188 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X16 FILLER_10_65 ();
 FILLCELL_X8 FILLER_10_81 ();
 FILLCELL_X1 FILLER_10_89 ();
 FILLCELL_X8 FILLER_10_109 ();
 FILLCELL_X4 FILLER_10_117 ();
 FILLCELL_X2 FILLER_10_121 ();
 FILLCELL_X1 FILLER_10_123 ();
 FILLCELL_X8 FILLER_10_144 ();
 FILLCELL_X4 FILLER_10_152 ();
 FILLCELL_X2 FILLER_10_156 ();
 FILLCELL_X1 FILLER_10_158 ();
 FILLCELL_X2 FILLER_10_163 ();
 FILLCELL_X4 FILLER_10_182 ();
 FILLCELL_X2 FILLER_10_186 ();
 FILLCELL_X1 FILLER_10_188 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X16 FILLER_11_161 ();
 FILLCELL_X8 FILLER_11_177 ();
 FILLCELL_X4 FILLER_11_185 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X4 FILLER_12_129 ();
 FILLCELL_X2 FILLER_12_133 ();
 FILLCELL_X16 FILLER_12_140 ();
 FILLCELL_X1 FILLER_12_156 ();
 FILLCELL_X8 FILLER_12_174 ();
 FILLCELL_X4 FILLER_12_182 ();
 FILLCELL_X2 FILLER_12_186 ();
 FILLCELL_X1 FILLER_12_188 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X16 FILLER_13_129 ();
 FILLCELL_X8 FILLER_13_145 ();
 FILLCELL_X2 FILLER_13_153 ();
 FILLCELL_X1 FILLER_13_155 ();
 FILLCELL_X8 FILLER_13_178 ();
 FILLCELL_X2 FILLER_13_186 ();
 FILLCELL_X1 FILLER_13_188 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X2 FILLER_14_161 ();
 FILLCELL_X2 FILLER_14_183 ();
 FILLCELL_X1 FILLER_14_188 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X8 FILLER_15_161 ();
 FILLCELL_X4 FILLER_15_169 ();
 FILLCELL_X1 FILLER_15_173 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X16 FILLER_16_161 ();
 FILLCELL_X8 FILLER_16_177 ();
 FILLCELL_X4 FILLER_16_185 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X16 FILLER_17_161 ();
 FILLCELL_X8 FILLER_17_177 ();
 FILLCELL_X4 FILLER_17_185 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X16 FILLER_18_161 ();
 FILLCELL_X8 FILLER_18_177 ();
 FILLCELL_X4 FILLER_18_185 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X16 FILLER_19_161 ();
 FILLCELL_X8 FILLER_19_177 ();
 FILLCELL_X4 FILLER_19_185 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X16 FILLER_20_161 ();
 FILLCELL_X8 FILLER_20_177 ();
 FILLCELL_X4 FILLER_20_185 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X16 FILLER_21_161 ();
 FILLCELL_X8 FILLER_21_177 ();
 FILLCELL_X4 FILLER_21_185 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X16 FILLER_22_161 ();
 FILLCELL_X8 FILLER_22_177 ();
 FILLCELL_X4 FILLER_22_185 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X16 FILLER_23_161 ();
 FILLCELL_X8 FILLER_23_177 ();
 FILLCELL_X4 FILLER_23_185 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X16 FILLER_24_161 ();
 FILLCELL_X8 FILLER_24_177 ();
 FILLCELL_X4 FILLER_24_185 ();
endmodule
