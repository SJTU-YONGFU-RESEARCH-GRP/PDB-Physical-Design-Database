module dual_port_ram (clk,
    we_a,
    we_b,
    addr_a,
    addr_b,
    data_a,
    data_b,
    q_a,
    q_b);
 input clk;
 input we_a;
 input we_b;
 input [3:0] addr_a;
 input [3:0] addr_b;
 input [7:0] data_a;
 input [7:0] data_b;
 output [7:0] q_a;
 output [7:0] q_b;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire \ram[0][0] ;
 wire \ram[0][1] ;
 wire \ram[0][2] ;
 wire \ram[0][3] ;
 wire \ram[0][4] ;
 wire \ram[0][5] ;
 wire \ram[0][6] ;
 wire \ram[0][7] ;
 wire \ram[10][0] ;
 wire \ram[10][1] ;
 wire \ram[10][2] ;
 wire \ram[10][3] ;
 wire \ram[10][4] ;
 wire \ram[10][5] ;
 wire \ram[10][6] ;
 wire \ram[10][7] ;
 wire \ram[11][0] ;
 wire \ram[11][1] ;
 wire \ram[11][2] ;
 wire \ram[11][3] ;
 wire \ram[11][4] ;
 wire \ram[11][5] ;
 wire \ram[11][6] ;
 wire \ram[11][7] ;
 wire \ram[12][0] ;
 wire \ram[12][1] ;
 wire \ram[12][2] ;
 wire \ram[12][3] ;
 wire \ram[12][4] ;
 wire \ram[12][5] ;
 wire \ram[12][6] ;
 wire \ram[12][7] ;
 wire \ram[13][0] ;
 wire \ram[13][1] ;
 wire \ram[13][2] ;
 wire \ram[13][3] ;
 wire \ram[13][4] ;
 wire \ram[13][5] ;
 wire \ram[13][6] ;
 wire \ram[13][7] ;
 wire \ram[14][0] ;
 wire \ram[14][1] ;
 wire \ram[14][2] ;
 wire \ram[14][3] ;
 wire \ram[14][4] ;
 wire \ram[14][5] ;
 wire \ram[14][6] ;
 wire \ram[14][7] ;
 wire \ram[15][0] ;
 wire \ram[15][1] ;
 wire \ram[15][2] ;
 wire \ram[15][3] ;
 wire \ram[15][4] ;
 wire \ram[15][5] ;
 wire \ram[15][6] ;
 wire \ram[15][7] ;
 wire \ram[1][0] ;
 wire \ram[1][1] ;
 wire \ram[1][2] ;
 wire \ram[1][3] ;
 wire \ram[1][4] ;
 wire \ram[1][5] ;
 wire \ram[1][6] ;
 wire \ram[1][7] ;
 wire \ram[2][0] ;
 wire \ram[2][1] ;
 wire \ram[2][2] ;
 wire \ram[2][3] ;
 wire \ram[2][4] ;
 wire \ram[2][5] ;
 wire \ram[2][6] ;
 wire \ram[2][7] ;
 wire \ram[3][0] ;
 wire \ram[3][1] ;
 wire \ram[3][2] ;
 wire \ram[3][3] ;
 wire \ram[3][4] ;
 wire \ram[3][5] ;
 wire \ram[3][6] ;
 wire \ram[3][7] ;
 wire \ram[4][0] ;
 wire \ram[4][1] ;
 wire \ram[4][2] ;
 wire \ram[4][3] ;
 wire \ram[4][4] ;
 wire \ram[4][5] ;
 wire \ram[4][6] ;
 wire \ram[4][7] ;
 wire \ram[5][0] ;
 wire \ram[5][1] ;
 wire \ram[5][2] ;
 wire \ram[5][3] ;
 wire \ram[5][4] ;
 wire \ram[5][5] ;
 wire \ram[5][6] ;
 wire \ram[5][7] ;
 wire \ram[6][0] ;
 wire \ram[6][1] ;
 wire \ram[6][2] ;
 wire \ram[6][3] ;
 wire \ram[6][4] ;
 wire \ram[6][5] ;
 wire \ram[6][6] ;
 wire \ram[6][7] ;
 wire \ram[7][0] ;
 wire \ram[7][1] ;
 wire \ram[7][2] ;
 wire \ram[7][3] ;
 wire \ram[7][4] ;
 wire \ram[7][5] ;
 wire \ram[7][6] ;
 wire \ram[7][7] ;
 wire \ram[8][0] ;
 wire \ram[8][1] ;
 wire \ram[8][2] ;
 wire \ram[8][3] ;
 wire \ram[8][4] ;
 wire \ram[8][5] ;
 wire \ram[8][6] ;
 wire \ram[8][7] ;
 wire \ram[9][0] ;
 wire \ram[9][1] ;
 wire \ram[9][2] ;
 wire \ram[9][3] ;
 wire \ram[9][4] ;
 wire \ram[9][5] ;
 wire \ram[9][6] ;
 wire \ram[9][7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 sky130_fd_sc_hd__buf_4 _344_ (.A(addr_a[3]),
    .X(_160_));
 sky130_fd_sc_hd__nand2b_1 _345_ (.A_N(_160_),
    .B(net1),
    .Y(_161_));
 sky130_fd_sc_hd__buf_4 _346_ (.A(_161_),
    .X(_162_));
 sky130_fd_sc_hd__buf_4 _347_ (.A(addr_a[0]),
    .X(_163_));
 sky130_fd_sc_hd__buf_4 _348_ (.A(addr_a[2]),
    .X(_164_));
 sky130_fd_sc_hd__nand3_4 _349_ (.A(net20),
    .B(_163_),
    .C(_164_),
    .Y(_165_));
 sky130_fd_sc_hd__nand3b_4 _350_ (.A_N(net3),
    .B(net2),
    .C(net21),
    .Y(_166_));
 sky130_fd_sc_hd__buf_4 _351_ (.A(addr_b[0]),
    .X(_167_));
 sky130_fd_sc_hd__buf_6 _352_ (.A(_167_),
    .X(_168_));
 sky130_fd_sc_hd__buf_4 _353_ (.A(addr_b[1]),
    .X(_169_));
 sky130_fd_sc_hd__buf_4 _354_ (.A(_169_),
    .X(_170_));
 sky130_fd_sc_hd__nand2_4 _355_ (.A(_168_),
    .B(_170_),
    .Y(_171_));
 sky130_fd_sc_hd__o22ai_4 _356_ (.A1(_162_),
    .A2(_165_),
    .B1(_166_),
    .B2(_171_),
    .Y(_018_));
 sky130_fd_sc_hd__nand3b_4 _357_ (.A_N(net2),
    .B(net21),
    .C(net3),
    .Y(_172_));
 sky130_fd_sc_hd__or2_4 _358_ (.A(_168_),
    .B(_170_),
    .X(_173_));
 sky130_fd_sc_hd__buf_4 _359_ (.A(net1),
    .X(_174_));
 sky130_fd_sc_hd__nand2b_1 _360_ (.A_N(_174_),
    .B(_160_),
    .Y(_175_));
 sky130_fd_sc_hd__buf_4 _361_ (.A(_175_),
    .X(_176_));
 sky130_fd_sc_hd__nor3b_4 _362_ (.A(_163_),
    .B(_164_),
    .C_N(net20),
    .Y(_177_));
 sky130_fd_sc_hd__nand2b_1 _363_ (.A_N(_176_),
    .B(_177_),
    .Y(_178_));
 sky130_fd_sc_hd__buf_4 _364_ (.A(_178_),
    .X(_179_));
 sky130_fd_sc_hd__o21ai_4 _365_ (.A1(_172_),
    .A2(_173_),
    .B1(_179_),
    .Y(_017_));
 sky130_fd_sc_hd__nand3b_4 _366_ (.A_N(_164_),
    .B(_163_),
    .C(net20),
    .Y(_180_));
 sky130_fd_sc_hd__nand2b_4 _367_ (.A_N(_170_),
    .B(_168_),
    .Y(_181_));
 sky130_fd_sc_hd__o22ai_4 _368_ (.A1(_176_),
    .A2(_180_),
    .B1(_181_),
    .B2(_172_),
    .Y(_016_));
 sky130_fd_sc_hd__or3b_4 _369_ (.A(net3),
    .B(net2),
    .C_N(net21),
    .X(_182_));
 sky130_fd_sc_hd__nor2_2 _370_ (.A(_174_),
    .B(_160_),
    .Y(_183_));
 sky130_fd_sc_hd__nand2_8 _371_ (.A(_177_),
    .B(_183_),
    .Y(_184_));
 sky130_fd_sc_hd__o21ai_4 _372_ (.A1(_173_),
    .A2(_182_),
    .B1(_184_),
    .Y(_031_));
 sky130_fd_sc_hd__buf_4 _373_ (.A(_169_),
    .X(_185_));
 sky130_fd_sc_hd__nand2b_4 _374_ (.A_N(_168_),
    .B(_185_),
    .Y(_186_));
 sky130_fd_sc_hd__and3_1 _375_ (.A(_174_),
    .B(_160_),
    .C(_177_),
    .X(_187_));
 sky130_fd_sc_hd__clkbuf_4 _376_ (.A(_187_),
    .X(_188_));
 sky130_fd_sc_hd__o21bai_4 _377_ (.A1(_172_),
    .A2(_186_),
    .B1_N(_188_),
    .Y(_030_));
 sky130_fd_sc_hd__nand2_8 _378_ (.A(_174_),
    .B(_160_),
    .Y(_189_));
 sky130_fd_sc_hd__o22ai_4 _379_ (.A1(_171_),
    .A2(_172_),
    .B1(_180_),
    .B2(_189_),
    .Y(_029_));
 sky130_fd_sc_hd__nand3b_4 _380_ (.A_N(_163_),
    .B(_164_),
    .C(net20),
    .Y(_190_));
 sky130_fd_sc_hd__nand3_4 _381_ (.A(net3),
    .B(net2),
    .C(net21),
    .Y(_191_));
 sky130_fd_sc_hd__o22ai_4 _382_ (.A1(_176_),
    .A2(_190_),
    .B1(_191_),
    .B2(_173_),
    .Y(_028_));
 sky130_fd_sc_hd__o22ai_4 _383_ (.A1(_165_),
    .A2(_176_),
    .B1(_181_),
    .B2(_191_),
    .Y(_027_));
 sky130_fd_sc_hd__o22ai_4 _384_ (.A1(_189_),
    .A2(_190_),
    .B1(_191_),
    .B2(_186_),
    .Y(_026_));
 sky130_fd_sc_hd__o22ai_4 _385_ (.A1(_165_),
    .A2(_189_),
    .B1(_191_),
    .B2(_171_),
    .Y(_025_));
 sky130_fd_sc_hd__nand2b_1 _386_ (.A_N(_180_),
    .B(_183_),
    .Y(_192_));
 sky130_fd_sc_hd__buf_4 _387_ (.A(_192_),
    .X(_193_));
 sky130_fd_sc_hd__o21ai_4 _388_ (.A1(_181_),
    .A2(_182_),
    .B1(_193_),
    .Y(_024_));
 sky130_fd_sc_hd__nand2b_1 _389_ (.A_N(_162_),
    .B(_177_),
    .Y(_194_));
 sky130_fd_sc_hd__buf_4 _390_ (.A(_194_),
    .X(_195_));
 sky130_fd_sc_hd__o21ai_4 _391_ (.A1(_182_),
    .A2(_186_),
    .B1(_195_),
    .Y(_023_));
 sky130_fd_sc_hd__o22ai_4 _392_ (.A1(_162_),
    .A2(_180_),
    .B1(_182_),
    .B2(_171_),
    .Y(_022_));
 sky130_fd_sc_hd__or3_1 _393_ (.A(_174_),
    .B(_160_),
    .C(_190_),
    .X(_196_));
 sky130_fd_sc_hd__buf_6 _394_ (.A(_196_),
    .X(_197_));
 sky130_fd_sc_hd__o21ai_4 _395_ (.A1(_166_),
    .A2(_173_),
    .B1(_197_),
    .Y(_021_));
 sky130_fd_sc_hd__nand2b_1 _396_ (.A_N(_165_),
    .B(_183_),
    .Y(_198_));
 sky130_fd_sc_hd__buf_4 _397_ (.A(_198_),
    .X(_199_));
 sky130_fd_sc_hd__o21ai_4 _398_ (.A1(_166_),
    .A2(_181_),
    .B1(_199_),
    .Y(_020_));
 sky130_fd_sc_hd__o22ai_4 _399_ (.A1(_166_),
    .A2(_186_),
    .B1(_190_),
    .B2(_162_),
    .Y(_019_));
 sky130_fd_sc_hd__clkbuf_4 _400_ (.A(net10),
    .X(_200_));
 sky130_fd_sc_hd__mux2_1 _401_ (.A0(_200_),
    .A1(net18),
    .S(_184_),
    .X(_038_));
 sky130_fd_sc_hd__clkbuf_4 _402_ (.A(net11),
    .X(_201_));
 sky130_fd_sc_hd__mux2_1 _403_ (.A0(_201_),
    .A1(net19),
    .S(_184_),
    .X(_039_));
 sky130_fd_sc_hd__clkbuf_4 _404_ (.A(net4),
    .X(_202_));
 sky130_fd_sc_hd__mux2_1 _405_ (.A0(_202_),
    .A1(net12),
    .S(_193_),
    .X(_088_));
 sky130_fd_sc_hd__buf_4 _406_ (.A(net5),
    .X(_203_));
 sky130_fd_sc_hd__mux2_1 _407_ (.A0(_203_),
    .A1(net13),
    .S(_193_),
    .X(_089_));
 sky130_fd_sc_hd__buf_2 _408_ (.A(net6),
    .X(_204_));
 sky130_fd_sc_hd__mux2_1 _409_ (.A0(_204_),
    .A1(net14),
    .S(_193_),
    .X(_090_));
 sky130_fd_sc_hd__clkbuf_4 _410_ (.A(net7),
    .X(_205_));
 sky130_fd_sc_hd__mux2_1 _411_ (.A0(_205_),
    .A1(net15),
    .S(_193_),
    .X(_091_));
 sky130_fd_sc_hd__clkbuf_4 _412_ (.A(net8),
    .X(_206_));
 sky130_fd_sc_hd__mux2_1 _413_ (.A0(_206_),
    .A1(net16),
    .S(_193_),
    .X(_092_));
 sky130_fd_sc_hd__clkbuf_4 _414_ (.A(net9),
    .X(_207_));
 sky130_fd_sc_hd__mux2_1 _415_ (.A0(_207_),
    .A1(net17),
    .S(_193_),
    .X(_093_));
 sky130_fd_sc_hd__mux2_1 _416_ (.A0(_200_),
    .A1(net18),
    .S(_193_),
    .X(_094_));
 sky130_fd_sc_hd__mux2_1 _417_ (.A0(_201_),
    .A1(net19),
    .S(_193_),
    .X(_095_));
 sky130_fd_sc_hd__mux2_1 _418_ (.A0(_202_),
    .A1(net12),
    .S(_195_),
    .X(_096_));
 sky130_fd_sc_hd__mux2_1 _419_ (.A0(_203_),
    .A1(net13),
    .S(_195_),
    .X(_097_));
 sky130_fd_sc_hd__mux2_1 _420_ (.A0(_204_),
    .A1(net14),
    .S(_195_),
    .X(_098_));
 sky130_fd_sc_hd__mux2_1 _421_ (.A0(_205_),
    .A1(net15),
    .S(_195_),
    .X(_099_));
 sky130_fd_sc_hd__mux2_1 _422_ (.A0(_206_),
    .A1(net16),
    .S(_195_),
    .X(_100_));
 sky130_fd_sc_hd__mux2_1 _423_ (.A0(_207_),
    .A1(net17),
    .S(_195_),
    .X(_101_));
 sky130_fd_sc_hd__mux2_1 _424_ (.A0(_200_),
    .A1(net18),
    .S(_195_),
    .X(_102_));
 sky130_fd_sc_hd__mux2_1 _425_ (.A0(_201_),
    .A1(net19),
    .S(_195_),
    .X(_103_));
 sky130_fd_sc_hd__clkbuf_4 _426_ (.A(net12),
    .X(_208_));
 sky130_fd_sc_hd__nor2_4 _427_ (.A(_162_),
    .B(_180_),
    .Y(_209_));
 sky130_fd_sc_hd__mux2_1 _428_ (.A0(_208_),
    .A1(_202_),
    .S(_209_),
    .X(_104_));
 sky130_fd_sc_hd__clkbuf_4 _429_ (.A(net13),
    .X(_210_));
 sky130_fd_sc_hd__mux2_1 _430_ (.A0(_210_),
    .A1(_203_),
    .S(_209_),
    .X(_105_));
 sky130_fd_sc_hd__buf_2 _431_ (.A(net14),
    .X(_211_));
 sky130_fd_sc_hd__mux2_1 _432_ (.A0(_211_),
    .A1(_204_),
    .S(_209_),
    .X(_106_));
 sky130_fd_sc_hd__clkbuf_4 _433_ (.A(net15),
    .X(_212_));
 sky130_fd_sc_hd__mux2_1 _434_ (.A0(_212_),
    .A1(_205_),
    .S(_209_),
    .X(_107_));
 sky130_fd_sc_hd__clkbuf_4 _435_ (.A(net16),
    .X(_213_));
 sky130_fd_sc_hd__mux2_1 _436_ (.A0(_213_),
    .A1(_206_),
    .S(_209_),
    .X(_108_));
 sky130_fd_sc_hd__clkbuf_4 _437_ (.A(net17),
    .X(_214_));
 sky130_fd_sc_hd__mux2_1 _438_ (.A0(_214_),
    .A1(_207_),
    .S(_209_),
    .X(_109_));
 sky130_fd_sc_hd__clkbuf_4 _439_ (.A(net18),
    .X(_215_));
 sky130_fd_sc_hd__mux2_1 _440_ (.A0(_215_),
    .A1(_200_),
    .S(_209_),
    .X(_110_));
 sky130_fd_sc_hd__clkbuf_4 _441_ (.A(net19),
    .X(_216_));
 sky130_fd_sc_hd__mux2_1 _442_ (.A0(_216_),
    .A1(_201_),
    .S(_209_),
    .X(_111_));
 sky130_fd_sc_hd__mux2_1 _443_ (.A0(_202_),
    .A1(net12),
    .S(_197_),
    .X(_112_));
 sky130_fd_sc_hd__mux2_1 _444_ (.A0(_203_),
    .A1(net13),
    .S(_197_),
    .X(_113_));
 sky130_fd_sc_hd__mux2_1 _445_ (.A0(_204_),
    .A1(net14),
    .S(_197_),
    .X(_114_));
 sky130_fd_sc_hd__mux2_1 _446_ (.A0(_205_),
    .A1(net15),
    .S(_197_),
    .X(_115_));
 sky130_fd_sc_hd__mux2_1 _447_ (.A0(_206_),
    .A1(net16),
    .S(_197_),
    .X(_116_));
 sky130_fd_sc_hd__mux2_1 _448_ (.A0(_207_),
    .A1(net17),
    .S(_197_),
    .X(_117_));
 sky130_fd_sc_hd__mux2_1 _449_ (.A0(_200_),
    .A1(net18),
    .S(_197_),
    .X(_118_));
 sky130_fd_sc_hd__mux2_1 _450_ (.A0(_201_),
    .A1(net19),
    .S(_197_),
    .X(_119_));
 sky130_fd_sc_hd__mux2_1 _451_ (.A0(_202_),
    .A1(net12),
    .S(_199_),
    .X(_120_));
 sky130_fd_sc_hd__mux2_1 _452_ (.A0(_203_),
    .A1(net13),
    .S(_199_),
    .X(_121_));
 sky130_fd_sc_hd__mux2_1 _453_ (.A0(_204_),
    .A1(net14),
    .S(_199_),
    .X(_122_));
 sky130_fd_sc_hd__mux2_1 _454_ (.A0(_205_),
    .A1(net15),
    .S(_199_),
    .X(_123_));
 sky130_fd_sc_hd__mux2_1 _455_ (.A0(_206_),
    .A1(net16),
    .S(_199_),
    .X(_124_));
 sky130_fd_sc_hd__mux2_1 _456_ (.A0(_207_),
    .A1(net17),
    .S(_199_),
    .X(_125_));
 sky130_fd_sc_hd__mux2_1 _457_ (.A0(_200_),
    .A1(net18),
    .S(_199_),
    .X(_126_));
 sky130_fd_sc_hd__mux2_1 _458_ (.A0(_201_),
    .A1(net19),
    .S(_199_),
    .X(_127_));
 sky130_fd_sc_hd__nor2_4 _459_ (.A(_162_),
    .B(_190_),
    .Y(_217_));
 sky130_fd_sc_hd__mux2_1 _460_ (.A0(_208_),
    .A1(_202_),
    .S(_217_),
    .X(_128_));
 sky130_fd_sc_hd__mux2_1 _461_ (.A0(_210_),
    .A1(_203_),
    .S(_217_),
    .X(_129_));
 sky130_fd_sc_hd__mux2_1 _462_ (.A0(_211_),
    .A1(_204_),
    .S(_217_),
    .X(_130_));
 sky130_fd_sc_hd__mux2_1 _463_ (.A0(_212_),
    .A1(_205_),
    .S(_217_),
    .X(_131_));
 sky130_fd_sc_hd__mux2_1 _464_ (.A0(_213_),
    .A1(_206_),
    .S(_217_),
    .X(_132_));
 sky130_fd_sc_hd__mux2_1 _465_ (.A0(_214_),
    .A1(_207_),
    .S(_217_),
    .X(_133_));
 sky130_fd_sc_hd__mux2_1 _466_ (.A0(_215_),
    .A1(_200_),
    .S(_217_),
    .X(_134_));
 sky130_fd_sc_hd__mux2_1 _467_ (.A0(_216_),
    .A1(_201_),
    .S(_217_),
    .X(_135_));
 sky130_fd_sc_hd__nor2_4 _468_ (.A(_162_),
    .B(_165_),
    .Y(_218_));
 sky130_fd_sc_hd__mux2_1 _469_ (.A0(_208_),
    .A1(_202_),
    .S(_218_),
    .X(_136_));
 sky130_fd_sc_hd__mux2_1 _470_ (.A0(_210_),
    .A1(_203_),
    .S(_218_),
    .X(_137_));
 sky130_fd_sc_hd__mux2_1 _471_ (.A0(_211_),
    .A1(_204_),
    .S(_218_),
    .X(_138_));
 sky130_fd_sc_hd__mux2_1 _472_ (.A0(_212_),
    .A1(_205_),
    .S(_218_),
    .X(_139_));
 sky130_fd_sc_hd__mux2_1 _473_ (.A0(_213_),
    .A1(_206_),
    .S(_218_),
    .X(_140_));
 sky130_fd_sc_hd__mux2_1 _474_ (.A0(_214_),
    .A1(_207_),
    .S(_218_),
    .X(_141_));
 sky130_fd_sc_hd__mux2_1 _475_ (.A0(_215_),
    .A1(_200_),
    .S(_218_),
    .X(_142_));
 sky130_fd_sc_hd__mux2_1 _476_ (.A0(_216_),
    .A1(_201_),
    .S(_218_),
    .X(_143_));
 sky130_fd_sc_hd__mux2_1 _477_ (.A0(_202_),
    .A1(net12),
    .S(_179_),
    .X(_144_));
 sky130_fd_sc_hd__mux2_1 _478_ (.A0(_203_),
    .A1(net13),
    .S(_179_),
    .X(_145_));
 sky130_fd_sc_hd__mux2_1 _479_ (.A0(_204_),
    .A1(net14),
    .S(_179_),
    .X(_146_));
 sky130_fd_sc_hd__mux2_1 _480_ (.A0(_205_),
    .A1(net15),
    .S(_179_),
    .X(_147_));
 sky130_fd_sc_hd__mux2_1 _481_ (.A0(_206_),
    .A1(net16),
    .S(_179_),
    .X(_148_));
 sky130_fd_sc_hd__mux2_1 _482_ (.A0(_207_),
    .A1(net17),
    .S(_179_),
    .X(_149_));
 sky130_fd_sc_hd__mux2_1 _483_ (.A0(_200_),
    .A1(net18),
    .S(_179_),
    .X(_150_));
 sky130_fd_sc_hd__mux2_1 _484_ (.A0(_201_),
    .A1(net19),
    .S(_179_),
    .X(_151_));
 sky130_fd_sc_hd__nor2_4 _485_ (.A(_176_),
    .B(_180_),
    .Y(_219_));
 sky130_fd_sc_hd__mux2_1 _486_ (.A0(_208_),
    .A1(_202_),
    .S(_219_),
    .X(_152_));
 sky130_fd_sc_hd__mux2_1 _487_ (.A0(_210_),
    .A1(_203_),
    .S(_219_),
    .X(_153_));
 sky130_fd_sc_hd__mux2_1 _488_ (.A0(_211_),
    .A1(_204_),
    .S(_219_),
    .X(_154_));
 sky130_fd_sc_hd__mux2_1 _489_ (.A0(_212_),
    .A1(_205_),
    .S(_219_),
    .X(_155_));
 sky130_fd_sc_hd__mux2_1 _490_ (.A0(_213_),
    .A1(_206_),
    .S(_219_),
    .X(_156_));
 sky130_fd_sc_hd__mux2_1 _491_ (.A0(_214_),
    .A1(_207_),
    .S(_219_),
    .X(_157_));
 sky130_fd_sc_hd__mux2_1 _492_ (.A0(_215_),
    .A1(_200_),
    .S(_219_),
    .X(_158_));
 sky130_fd_sc_hd__mux2_1 _493_ (.A0(_216_),
    .A1(_201_),
    .S(_219_),
    .X(_159_));
 sky130_fd_sc_hd__mux2_1 _494_ (.A0(_208_),
    .A1(net4),
    .S(_188_),
    .X(_040_));
 sky130_fd_sc_hd__mux2_1 _495_ (.A0(_210_),
    .A1(net5),
    .S(_188_),
    .X(_041_));
 sky130_fd_sc_hd__mux2_1 _496_ (.A0(_211_),
    .A1(net6),
    .S(_188_),
    .X(_042_));
 sky130_fd_sc_hd__mux2_1 _497_ (.A0(_212_),
    .A1(net7),
    .S(_188_),
    .X(_043_));
 sky130_fd_sc_hd__mux2_1 _498_ (.A0(_213_),
    .A1(net8),
    .S(_188_),
    .X(_044_));
 sky130_fd_sc_hd__mux2_1 _499_ (.A0(_214_),
    .A1(net9),
    .S(_188_),
    .X(_045_));
 sky130_fd_sc_hd__mux2_1 _500_ (.A0(_215_),
    .A1(net10),
    .S(_188_),
    .X(_046_));
 sky130_fd_sc_hd__mux2_1 _501_ (.A0(_216_),
    .A1(net11),
    .S(_188_),
    .X(_047_));
 sky130_fd_sc_hd__nor2_4 _502_ (.A(_180_),
    .B(_189_),
    .Y(_220_));
 sky130_fd_sc_hd__mux2_1 _503_ (.A0(_208_),
    .A1(net4),
    .S(_220_),
    .X(_048_));
 sky130_fd_sc_hd__mux2_1 _504_ (.A0(_210_),
    .A1(net5),
    .S(_220_),
    .X(_049_));
 sky130_fd_sc_hd__mux2_1 _505_ (.A0(_211_),
    .A1(net6),
    .S(_220_),
    .X(_050_));
 sky130_fd_sc_hd__mux2_1 _506_ (.A0(_212_),
    .A1(net7),
    .S(_220_),
    .X(_051_));
 sky130_fd_sc_hd__mux2_1 _507_ (.A0(_213_),
    .A1(net8),
    .S(_220_),
    .X(_052_));
 sky130_fd_sc_hd__mux2_1 _508_ (.A0(_214_),
    .A1(net9),
    .S(_220_),
    .X(_053_));
 sky130_fd_sc_hd__mux2_1 _509_ (.A0(_215_),
    .A1(net10),
    .S(_220_),
    .X(_054_));
 sky130_fd_sc_hd__mux2_1 _510_ (.A0(_216_),
    .A1(net11),
    .S(_220_),
    .X(_055_));
 sky130_fd_sc_hd__nor2_4 _511_ (.A(_176_),
    .B(_190_),
    .Y(_221_));
 sky130_fd_sc_hd__mux2_1 _512_ (.A0(_208_),
    .A1(net4),
    .S(_221_),
    .X(_056_));
 sky130_fd_sc_hd__mux2_1 _513_ (.A0(_210_),
    .A1(net5),
    .S(_221_),
    .X(_057_));
 sky130_fd_sc_hd__mux2_1 _514_ (.A0(_211_),
    .A1(net6),
    .S(_221_),
    .X(_058_));
 sky130_fd_sc_hd__mux2_1 _515_ (.A0(_212_),
    .A1(net7),
    .S(_221_),
    .X(_059_));
 sky130_fd_sc_hd__mux2_1 _516_ (.A0(_213_),
    .A1(net8),
    .S(_221_),
    .X(_060_));
 sky130_fd_sc_hd__mux2_1 _517_ (.A0(_214_),
    .A1(net9),
    .S(_221_),
    .X(_061_));
 sky130_fd_sc_hd__mux2_1 _518_ (.A0(_215_),
    .A1(net10),
    .S(_221_),
    .X(_062_));
 sky130_fd_sc_hd__mux2_1 _519_ (.A0(_216_),
    .A1(net11),
    .S(_221_),
    .X(_063_));
 sky130_fd_sc_hd__nor2_4 _520_ (.A(_165_),
    .B(_176_),
    .Y(_222_));
 sky130_fd_sc_hd__mux2_1 _521_ (.A0(_208_),
    .A1(net4),
    .S(_222_),
    .X(_064_));
 sky130_fd_sc_hd__mux2_1 _522_ (.A0(_210_),
    .A1(net5),
    .S(_222_),
    .X(_065_));
 sky130_fd_sc_hd__mux2_1 _523_ (.A0(_211_),
    .A1(net6),
    .S(_222_),
    .X(_066_));
 sky130_fd_sc_hd__mux2_1 _524_ (.A0(_212_),
    .A1(net7),
    .S(_222_),
    .X(_067_));
 sky130_fd_sc_hd__mux2_1 _525_ (.A0(_213_),
    .A1(net8),
    .S(_222_),
    .X(_068_));
 sky130_fd_sc_hd__mux2_1 _526_ (.A0(_214_),
    .A1(net9),
    .S(_222_),
    .X(_069_));
 sky130_fd_sc_hd__mux2_1 _527_ (.A0(_215_),
    .A1(net10),
    .S(_222_),
    .X(_070_));
 sky130_fd_sc_hd__mux2_1 _528_ (.A0(_216_),
    .A1(net11),
    .S(_222_),
    .X(_071_));
 sky130_fd_sc_hd__nor2_4 _529_ (.A(_189_),
    .B(_190_),
    .Y(_223_));
 sky130_fd_sc_hd__mux2_1 _530_ (.A0(_208_),
    .A1(net4),
    .S(_223_),
    .X(_072_));
 sky130_fd_sc_hd__mux2_1 _531_ (.A0(_210_),
    .A1(net5),
    .S(_223_),
    .X(_073_));
 sky130_fd_sc_hd__mux2_1 _532_ (.A0(_211_),
    .A1(net6),
    .S(_223_),
    .X(_074_));
 sky130_fd_sc_hd__mux2_1 _533_ (.A0(_212_),
    .A1(net7),
    .S(_223_),
    .X(_075_));
 sky130_fd_sc_hd__mux2_1 _534_ (.A0(_213_),
    .A1(net8),
    .S(_223_),
    .X(_076_));
 sky130_fd_sc_hd__mux2_1 _535_ (.A0(_214_),
    .A1(net9),
    .S(_223_),
    .X(_077_));
 sky130_fd_sc_hd__mux2_1 _536_ (.A0(_215_),
    .A1(net10),
    .S(_223_),
    .X(_078_));
 sky130_fd_sc_hd__mux2_1 _537_ (.A0(_216_),
    .A1(net11),
    .S(_223_),
    .X(_079_));
 sky130_fd_sc_hd__nor2_4 _538_ (.A(_165_),
    .B(_189_),
    .Y(_224_));
 sky130_fd_sc_hd__mux2_1 _539_ (.A0(_208_),
    .A1(net4),
    .S(_224_),
    .X(_080_));
 sky130_fd_sc_hd__mux2_1 _540_ (.A0(_210_),
    .A1(net5),
    .S(_224_),
    .X(_081_));
 sky130_fd_sc_hd__mux2_1 _541_ (.A0(_211_),
    .A1(net6),
    .S(_224_),
    .X(_082_));
 sky130_fd_sc_hd__mux2_1 _542_ (.A0(_212_),
    .A1(net7),
    .S(_224_),
    .X(_083_));
 sky130_fd_sc_hd__mux2_1 _543_ (.A0(_213_),
    .A1(net8),
    .S(_224_),
    .X(_084_));
 sky130_fd_sc_hd__mux2_1 _544_ (.A0(_214_),
    .A1(net9),
    .S(_224_),
    .X(_085_));
 sky130_fd_sc_hd__mux2_1 _545_ (.A0(_215_),
    .A1(net10),
    .S(_224_),
    .X(_086_));
 sky130_fd_sc_hd__mux2_1 _546_ (.A0(_216_),
    .A1(net11),
    .S(_224_),
    .X(_087_));
 sky130_fd_sc_hd__buf_4 _547_ (.A(_167_),
    .X(_225_));
 sky130_fd_sc_hd__clkbuf_4 _548_ (.A(_169_),
    .X(_226_));
 sky130_fd_sc_hd__mux4_1 _549_ (.A0(\ram[4][0] ),
    .A1(\ram[5][0] ),
    .A2(\ram[6][0] ),
    .A3(\ram[7][0] ),
    .S0(_225_),
    .S1(_226_),
    .X(_227_));
 sky130_fd_sc_hd__nor2b_1 _550_ (.A(net3),
    .B_N(net2),
    .Y(_228_));
 sky130_fd_sc_hd__clkbuf_4 _551_ (.A(_228_),
    .X(_229_));
 sky130_fd_sc_hd__mux4_1 _552_ (.A0(\ram[12][0] ),
    .A1(\ram[13][0] ),
    .A2(\ram[14][0] ),
    .A3(\ram[15][0] ),
    .S0(_168_),
    .S1(_170_),
    .X(_230_));
 sky130_fd_sc_hd__and2_0 _553_ (.A(net3),
    .B(net2),
    .X(_231_));
 sky130_fd_sc_hd__clkbuf_4 _554_ (.A(_231_),
    .X(_232_));
 sky130_fd_sc_hd__a22oi_1 _555_ (.A1(_227_),
    .A2(_229_),
    .B1(_230_),
    .B2(_232_),
    .Y(_233_));
 sky130_fd_sc_hd__mux4_1 _556_ (.A0(\ram[0][0] ),
    .A1(\ram[1][0] ),
    .A2(\ram[2][0] ),
    .A3(\ram[3][0] ),
    .S0(_225_),
    .S1(_226_),
    .X(_234_));
 sky130_fd_sc_hd__nor2_4 _557_ (.A(net3),
    .B(net2),
    .Y(_235_));
 sky130_fd_sc_hd__clkbuf_8 _558_ (.A(_167_),
    .X(_236_));
 sky130_fd_sc_hd__mux4_2 _559_ (.A0(\ram[8][0] ),
    .A1(\ram[9][0] ),
    .A2(\ram[10][0] ),
    .A3(\ram[11][0] ),
    .S0(_236_),
    .S1(_185_),
    .X(_237_));
 sky130_fd_sc_hd__nor2b_1 _560_ (.A(net2),
    .B_N(net3),
    .Y(_238_));
 sky130_fd_sc_hd__clkbuf_4 _561_ (.A(_238_),
    .X(_239_));
 sky130_fd_sc_hd__a22oi_2 _562_ (.A1(_234_),
    .A2(_235_),
    .B1(_237_),
    .B2(_239_),
    .Y(_240_));
 sky130_fd_sc_hd__nand2_1 _563_ (.A(_233_),
    .B(_240_),
    .Y(_000_));
 sky130_fd_sc_hd__mux4_1 _564_ (.A0(\ram[4][1] ),
    .A1(\ram[5][1] ),
    .A2(\ram[6][1] ),
    .A3(\ram[7][1] ),
    .S0(_225_),
    .S1(_226_),
    .X(_241_));
 sky130_fd_sc_hd__mux4_1 _565_ (.A0(\ram[12][1] ),
    .A1(\ram[13][1] ),
    .A2(\ram[14][1] ),
    .A3(\ram[15][1] ),
    .S0(_168_),
    .S1(_170_),
    .X(_242_));
 sky130_fd_sc_hd__a22oi_1 _566_ (.A1(_229_),
    .A2(_241_),
    .B1(_242_),
    .B2(_232_),
    .Y(_243_));
 sky130_fd_sc_hd__mux4_1 _567_ (.A0(\ram[0][1] ),
    .A1(\ram[1][1] ),
    .A2(\ram[2][1] ),
    .A3(\ram[3][1] ),
    .S0(_225_),
    .S1(_226_),
    .X(_244_));
 sky130_fd_sc_hd__mux4_2 _568_ (.A0(\ram[8][1] ),
    .A1(\ram[9][1] ),
    .A2(\ram[10][1] ),
    .A3(\ram[11][1] ),
    .S0(_236_),
    .S1(_185_),
    .X(_245_));
 sky130_fd_sc_hd__a22oi_2 _569_ (.A1(_235_),
    .A2(_244_),
    .B1(_245_),
    .B2(_239_),
    .Y(_246_));
 sky130_fd_sc_hd__nand2_1 _570_ (.A(_243_),
    .B(_246_),
    .Y(_001_));
 sky130_fd_sc_hd__mux4_1 _571_ (.A0(\ram[4][2] ),
    .A1(\ram[5][2] ),
    .A2(\ram[6][2] ),
    .A3(\ram[7][2] ),
    .S0(_225_),
    .S1(_226_),
    .X(_247_));
 sky130_fd_sc_hd__mux4_1 _572_ (.A0(\ram[12][2] ),
    .A1(\ram[13][2] ),
    .A2(\ram[14][2] ),
    .A3(\ram[15][2] ),
    .S0(_168_),
    .S1(_170_),
    .X(_248_));
 sky130_fd_sc_hd__a22oi_1 _573_ (.A1(_229_),
    .A2(_247_),
    .B1(_248_),
    .B2(_232_),
    .Y(_249_));
 sky130_fd_sc_hd__mux4_1 _574_ (.A0(\ram[0][2] ),
    .A1(\ram[1][2] ),
    .A2(\ram[2][2] ),
    .A3(\ram[3][2] ),
    .S0(_167_),
    .S1(_169_),
    .X(_250_));
 sky130_fd_sc_hd__mux4_1 _575_ (.A0(\ram[8][2] ),
    .A1(\ram[9][2] ),
    .A2(\ram[10][2] ),
    .A3(\ram[11][2] ),
    .S0(_236_),
    .S1(_185_),
    .X(_251_));
 sky130_fd_sc_hd__a22oi_2 _576_ (.A1(_235_),
    .A2(_250_),
    .B1(_251_),
    .B2(_239_),
    .Y(_252_));
 sky130_fd_sc_hd__nand2_1 _577_ (.A(_249_),
    .B(_252_),
    .Y(_002_));
 sky130_fd_sc_hd__mux4_1 _578_ (.A0(\ram[4][3] ),
    .A1(\ram[5][3] ),
    .A2(\ram[6][3] ),
    .A3(\ram[7][3] ),
    .S0(_225_),
    .S1(_226_),
    .X(_253_));
 sky130_fd_sc_hd__mux4_4 _579_ (.A0(\ram[12][3] ),
    .A1(\ram[13][3] ),
    .A2(\ram[14][3] ),
    .A3(\ram[15][3] ),
    .S0(_168_),
    .S1(_170_),
    .X(_254_));
 sky130_fd_sc_hd__a22oi_2 _580_ (.A1(_229_),
    .A2(_253_),
    .B1(_254_),
    .B2(_232_),
    .Y(_255_));
 sky130_fd_sc_hd__mux4_1 _581_ (.A0(\ram[0][3] ),
    .A1(\ram[1][3] ),
    .A2(\ram[2][3] ),
    .A3(\ram[3][3] ),
    .S0(_167_),
    .S1(_169_),
    .X(_256_));
 sky130_fd_sc_hd__mux4_2 _582_ (.A0(\ram[8][3] ),
    .A1(\ram[9][3] ),
    .A2(\ram[10][3] ),
    .A3(\ram[11][3] ),
    .S0(_236_),
    .S1(_185_),
    .X(_257_));
 sky130_fd_sc_hd__a22oi_1 _583_ (.A1(_235_),
    .A2(_256_),
    .B1(_257_),
    .B2(_239_),
    .Y(_258_));
 sky130_fd_sc_hd__nand2_1 _584_ (.A(_255_),
    .B(_258_),
    .Y(_003_));
 sky130_fd_sc_hd__mux4_1 _585_ (.A0(\ram[4][4] ),
    .A1(\ram[5][4] ),
    .A2(\ram[6][4] ),
    .A3(\ram[7][4] ),
    .S0(_225_),
    .S1(_226_),
    .X(_259_));
 sky130_fd_sc_hd__mux4_2 _586_ (.A0(\ram[12][4] ),
    .A1(\ram[13][4] ),
    .A2(\ram[14][4] ),
    .A3(\ram[15][4] ),
    .S0(_168_),
    .S1(_170_),
    .X(_260_));
 sky130_fd_sc_hd__a22oi_1 _587_ (.A1(_229_),
    .A2(_259_),
    .B1(_260_),
    .B2(_232_),
    .Y(_261_));
 sky130_fd_sc_hd__mux4_1 _588_ (.A0(\ram[0][4] ),
    .A1(\ram[1][4] ),
    .A2(\ram[2][4] ),
    .A3(\ram[3][4] ),
    .S0(_167_),
    .S1(_169_),
    .X(_262_));
 sky130_fd_sc_hd__mux4_4 _589_ (.A0(\ram[8][4] ),
    .A1(\ram[9][4] ),
    .A2(\ram[10][4] ),
    .A3(\ram[11][4] ),
    .S0(_236_),
    .S1(_185_),
    .X(_263_));
 sky130_fd_sc_hd__a22oi_2 _590_ (.A1(_235_),
    .A2(_262_),
    .B1(_263_),
    .B2(_239_),
    .Y(_264_));
 sky130_fd_sc_hd__nand2_1 _591_ (.A(_261_),
    .B(_264_),
    .Y(_004_));
 sky130_fd_sc_hd__mux4_1 _592_ (.A0(\ram[4][5] ),
    .A1(\ram[5][5] ),
    .A2(\ram[6][5] ),
    .A3(\ram[7][5] ),
    .S0(_225_),
    .S1(_226_),
    .X(_265_));
 sky130_fd_sc_hd__mux4_2 _593_ (.A0(\ram[12][5] ),
    .A1(\ram[13][5] ),
    .A2(\ram[14][5] ),
    .A3(\ram[15][5] ),
    .S0(_168_),
    .S1(_170_),
    .X(_266_));
 sky130_fd_sc_hd__a22oi_2 _594_ (.A1(_229_),
    .A2(_265_),
    .B1(_266_),
    .B2(_232_),
    .Y(_267_));
 sky130_fd_sc_hd__mux4_1 _595_ (.A0(\ram[0][5] ),
    .A1(\ram[1][5] ),
    .A2(\ram[2][5] ),
    .A3(\ram[3][5] ),
    .S0(_167_),
    .S1(_169_),
    .X(_268_));
 sky130_fd_sc_hd__mux4_1 _596_ (.A0(\ram[8][5] ),
    .A1(\ram[9][5] ),
    .A2(\ram[10][5] ),
    .A3(\ram[11][5] ),
    .S0(_236_),
    .S1(_185_),
    .X(_269_));
 sky130_fd_sc_hd__a22oi_1 _597_ (.A1(_235_),
    .A2(_268_),
    .B1(_269_),
    .B2(_239_),
    .Y(_270_));
 sky130_fd_sc_hd__nand2_1 _598_ (.A(_267_),
    .B(_270_),
    .Y(_005_));
 sky130_fd_sc_hd__mux4_1 _599_ (.A0(\ram[4][6] ),
    .A1(\ram[5][6] ),
    .A2(\ram[6][6] ),
    .A3(\ram[7][6] ),
    .S0(_225_),
    .S1(_226_),
    .X(_271_));
 sky130_fd_sc_hd__mux4_2 _600_ (.A0(\ram[12][6] ),
    .A1(\ram[13][6] ),
    .A2(\ram[14][6] ),
    .A3(\ram[15][6] ),
    .S0(_236_),
    .S1(_170_),
    .X(_272_));
 sky130_fd_sc_hd__a22oi_2 _601_ (.A1(_229_),
    .A2(_271_),
    .B1(_272_),
    .B2(_232_),
    .Y(_273_));
 sky130_fd_sc_hd__mux4_1 _602_ (.A0(\ram[0][6] ),
    .A1(\ram[1][6] ),
    .A2(\ram[2][6] ),
    .A3(\ram[3][6] ),
    .S0(_167_),
    .S1(_169_),
    .X(_274_));
 sky130_fd_sc_hd__mux4_1 _603_ (.A0(\ram[8][6] ),
    .A1(\ram[9][6] ),
    .A2(\ram[10][6] ),
    .A3(\ram[11][6] ),
    .S0(_236_),
    .S1(_185_),
    .X(_275_));
 sky130_fd_sc_hd__a22oi_1 _604_ (.A1(_235_),
    .A2(_274_),
    .B1(_275_),
    .B2(_239_),
    .Y(_276_));
 sky130_fd_sc_hd__nand2_1 _605_ (.A(_273_),
    .B(_276_),
    .Y(_006_));
 sky130_fd_sc_hd__mux4_1 _606_ (.A0(\ram[4][7] ),
    .A1(\ram[5][7] ),
    .A2(\ram[6][7] ),
    .A3(\ram[7][7] ),
    .S0(_225_),
    .S1(_226_),
    .X(_277_));
 sky130_fd_sc_hd__mux4_2 _607_ (.A0(\ram[12][7] ),
    .A1(\ram[13][7] ),
    .A2(\ram[14][7] ),
    .A3(\ram[15][7] ),
    .S0(_236_),
    .S1(_185_),
    .X(_278_));
 sky130_fd_sc_hd__a22oi_2 _608_ (.A1(_229_),
    .A2(_277_),
    .B1(_278_),
    .B2(_232_),
    .Y(_279_));
 sky130_fd_sc_hd__mux4_1 _609_ (.A0(\ram[0][7] ),
    .A1(\ram[1][7] ),
    .A2(\ram[2][7] ),
    .A3(\ram[3][7] ),
    .S0(_167_),
    .S1(_169_),
    .X(_280_));
 sky130_fd_sc_hd__mux4_1 _610_ (.A0(\ram[8][7] ),
    .A1(\ram[9][7] ),
    .A2(\ram[10][7] ),
    .A3(\ram[11][7] ),
    .S0(_236_),
    .S1(_185_),
    .X(_281_));
 sky130_fd_sc_hd__a22oi_1 _611_ (.A1(_235_),
    .A2(_280_),
    .B1(_281_),
    .B2(_239_),
    .Y(_282_));
 sky130_fd_sc_hd__nand2_1 _612_ (.A(_279_),
    .B(_282_),
    .Y(_007_));
 sky130_fd_sc_hd__buf_6 _613_ (.A(_163_),
    .X(_283_));
 sky130_fd_sc_hd__buf_4 _614_ (.A(_174_),
    .X(_284_));
 sky130_fd_sc_hd__mux4_1 _615_ (.A0(\ram[4][0] ),
    .A1(\ram[5][0] ),
    .A2(\ram[6][0] ),
    .A3(\ram[7][0] ),
    .S0(_283_),
    .S1(_284_),
    .X(_285_));
 sky130_fd_sc_hd__nor2b_1 _616_ (.A(_160_),
    .B_N(_164_),
    .Y(_286_));
 sky130_fd_sc_hd__clkbuf_4 _617_ (.A(_286_),
    .X(_287_));
 sky130_fd_sc_hd__buf_6 _618_ (.A(_163_),
    .X(_288_));
 sky130_fd_sc_hd__buf_4 _619_ (.A(_174_),
    .X(_289_));
 sky130_fd_sc_hd__mux4_1 _620_ (.A0(\ram[12][0] ),
    .A1(\ram[13][0] ),
    .A2(\ram[14][0] ),
    .A3(\ram[15][0] ),
    .S0(_288_),
    .S1(_289_),
    .X(_290_));
 sky130_fd_sc_hd__and2_0 _621_ (.A(_160_),
    .B(_164_),
    .X(_291_));
 sky130_fd_sc_hd__clkbuf_4 _622_ (.A(_291_),
    .X(_292_));
 sky130_fd_sc_hd__a22oi_1 _623_ (.A1(_285_),
    .A2(_287_),
    .B1(_290_),
    .B2(_292_),
    .Y(_293_));
 sky130_fd_sc_hd__mux4_1 _624_ (.A0(\ram[0][0] ),
    .A1(\ram[1][0] ),
    .A2(\ram[2][0] ),
    .A3(\ram[3][0] ),
    .S0(_283_),
    .S1(_284_),
    .X(_294_));
 sky130_fd_sc_hd__nor2_4 _625_ (.A(_160_),
    .B(_164_),
    .Y(_295_));
 sky130_fd_sc_hd__mux4_2 _626_ (.A0(\ram[8][0] ),
    .A1(\ram[9][0] ),
    .A2(\ram[10][0] ),
    .A3(\ram[11][0] ),
    .S0(_288_),
    .S1(_289_),
    .X(_296_));
 sky130_fd_sc_hd__nor2b_1 _627_ (.A(_164_),
    .B_N(_160_),
    .Y(_297_));
 sky130_fd_sc_hd__clkbuf_4 _628_ (.A(_297_),
    .X(_298_));
 sky130_fd_sc_hd__a22oi_2 _629_ (.A1(_294_),
    .A2(_295_),
    .B1(_296_),
    .B2(_298_),
    .Y(_299_));
 sky130_fd_sc_hd__nand2_1 _630_ (.A(_293_),
    .B(_299_),
    .Y(_008_));
 sky130_fd_sc_hd__mux4_1 _631_ (.A0(\ram[4][1] ),
    .A1(\ram[5][1] ),
    .A2(\ram[6][1] ),
    .A3(\ram[7][1] ),
    .S0(_283_),
    .S1(_284_),
    .X(_300_));
 sky130_fd_sc_hd__mux4_1 _632_ (.A0(\ram[12][1] ),
    .A1(\ram[13][1] ),
    .A2(\ram[14][1] ),
    .A3(\ram[15][1] ),
    .S0(_288_),
    .S1(_289_),
    .X(_301_));
 sky130_fd_sc_hd__a22oi_1 _633_ (.A1(_287_),
    .A2(_300_),
    .B1(_301_),
    .B2(_292_),
    .Y(_302_));
 sky130_fd_sc_hd__buf_4 _634_ (.A(_163_),
    .X(_303_));
 sky130_fd_sc_hd__buf_4 _635_ (.A(_174_),
    .X(_304_));
 sky130_fd_sc_hd__mux4_1 _636_ (.A0(\ram[0][1] ),
    .A1(\ram[1][1] ),
    .A2(\ram[2][1] ),
    .A3(\ram[3][1] ),
    .S0(_303_),
    .S1(_304_),
    .X(_305_));
 sky130_fd_sc_hd__mux4_2 _637_ (.A0(\ram[8][1] ),
    .A1(\ram[9][1] ),
    .A2(\ram[10][1] ),
    .A3(\ram[11][1] ),
    .S0(_288_),
    .S1(_289_),
    .X(_306_));
 sky130_fd_sc_hd__a22oi_2 _638_ (.A1(_295_),
    .A2(_305_),
    .B1(_306_),
    .B2(_298_),
    .Y(_307_));
 sky130_fd_sc_hd__nand2_1 _639_ (.A(_302_),
    .B(_307_),
    .Y(_009_));
 sky130_fd_sc_hd__mux4_1 _640_ (.A0(\ram[4][2] ),
    .A1(\ram[5][2] ),
    .A2(\ram[6][2] ),
    .A3(\ram[7][2] ),
    .S0(_283_),
    .S1(_284_),
    .X(_308_));
 sky130_fd_sc_hd__mux4_1 _641_ (.A0(\ram[12][2] ),
    .A1(\ram[13][2] ),
    .A2(\ram[14][2] ),
    .A3(\ram[15][2] ),
    .S0(_288_),
    .S1(_289_),
    .X(_309_));
 sky130_fd_sc_hd__a22oi_1 _642_ (.A1(_287_),
    .A2(_308_),
    .B1(_309_),
    .B2(_292_),
    .Y(_310_));
 sky130_fd_sc_hd__mux4_1 _643_ (.A0(\ram[0][2] ),
    .A1(\ram[1][2] ),
    .A2(\ram[2][2] ),
    .A3(\ram[3][2] ),
    .S0(_303_),
    .S1(_304_),
    .X(_311_));
 sky130_fd_sc_hd__mux4_1 _644_ (.A0(\ram[8][2] ),
    .A1(\ram[9][2] ),
    .A2(\ram[10][2] ),
    .A3(\ram[11][2] ),
    .S0(_283_),
    .S1(_284_),
    .X(_312_));
 sky130_fd_sc_hd__a22oi_2 _645_ (.A1(_295_),
    .A2(_311_),
    .B1(_312_),
    .B2(_298_),
    .Y(_313_));
 sky130_fd_sc_hd__nand2_1 _646_ (.A(_310_),
    .B(_313_),
    .Y(_010_));
 sky130_fd_sc_hd__mux4_1 _647_ (.A0(\ram[4][3] ),
    .A1(\ram[5][3] ),
    .A2(\ram[6][3] ),
    .A3(\ram[7][3] ),
    .S0(_303_),
    .S1(_304_),
    .X(_314_));
 sky130_fd_sc_hd__mux4_2 _648_ (.A0(\ram[12][3] ),
    .A1(\ram[13][3] ),
    .A2(\ram[14][3] ),
    .A3(\ram[15][3] ),
    .S0(_288_),
    .S1(_289_),
    .X(_315_));
 sky130_fd_sc_hd__a22oi_1 _649_ (.A1(_287_),
    .A2(_314_),
    .B1(_315_),
    .B2(_292_),
    .Y(_316_));
 sky130_fd_sc_hd__mux4_1 _650_ (.A0(\ram[0][3] ),
    .A1(\ram[1][3] ),
    .A2(\ram[2][3] ),
    .A3(\ram[3][3] ),
    .S0(_303_),
    .S1(_304_),
    .X(_317_));
 sky130_fd_sc_hd__mux4_2 _651_ (.A0(\ram[8][3] ),
    .A1(\ram[9][3] ),
    .A2(\ram[10][3] ),
    .A3(\ram[11][3] ),
    .S0(_283_),
    .S1(_284_),
    .X(_318_));
 sky130_fd_sc_hd__a22oi_2 _652_ (.A1(_295_),
    .A2(_317_),
    .B1(_318_),
    .B2(_298_),
    .Y(_319_));
 sky130_fd_sc_hd__nand2_1 _653_ (.A(_316_),
    .B(_319_),
    .Y(_011_));
 sky130_fd_sc_hd__mux4_1 _654_ (.A0(\ram[4][4] ),
    .A1(\ram[5][4] ),
    .A2(\ram[6][4] ),
    .A3(\ram[7][4] ),
    .S0(_303_),
    .S1(_304_),
    .X(_320_));
 sky130_fd_sc_hd__mux4_2 _655_ (.A0(\ram[12][4] ),
    .A1(\ram[13][4] ),
    .A2(\ram[14][4] ),
    .A3(\ram[15][4] ),
    .S0(_288_),
    .S1(_289_),
    .X(_321_));
 sky130_fd_sc_hd__a22oi_1 _656_ (.A1(_287_),
    .A2(_320_),
    .B1(_321_),
    .B2(_292_),
    .Y(_322_));
 sky130_fd_sc_hd__mux4_1 _657_ (.A0(\ram[0][4] ),
    .A1(\ram[1][4] ),
    .A2(\ram[2][4] ),
    .A3(\ram[3][4] ),
    .S0(_303_),
    .S1(_304_),
    .X(_323_));
 sky130_fd_sc_hd__mux4_4 _658_ (.A0(\ram[8][4] ),
    .A1(\ram[9][4] ),
    .A2(\ram[10][4] ),
    .A3(\ram[11][4] ),
    .S0(_283_),
    .S1(_284_),
    .X(_324_));
 sky130_fd_sc_hd__a22oi_2 _659_ (.A1(_295_),
    .A2(_323_),
    .B1(_324_),
    .B2(_298_),
    .Y(_325_));
 sky130_fd_sc_hd__nand2_1 _660_ (.A(_322_),
    .B(_325_),
    .Y(_012_));
 sky130_fd_sc_hd__mux4_1 _661_ (.A0(\ram[4][5] ),
    .A1(\ram[5][5] ),
    .A2(\ram[6][5] ),
    .A3(\ram[7][5] ),
    .S0(_303_),
    .S1(_304_),
    .X(_326_));
 sky130_fd_sc_hd__mux4_2 _662_ (.A0(\ram[12][5] ),
    .A1(\ram[13][5] ),
    .A2(\ram[14][5] ),
    .A3(\ram[15][5] ),
    .S0(_288_),
    .S1(_289_),
    .X(_327_));
 sky130_fd_sc_hd__a22oi_2 _663_ (.A1(_287_),
    .A2(_326_),
    .B1(_327_),
    .B2(_292_),
    .Y(_328_));
 sky130_fd_sc_hd__mux4_1 _664_ (.A0(\ram[0][5] ),
    .A1(\ram[1][5] ),
    .A2(\ram[2][5] ),
    .A3(\ram[3][5] ),
    .S0(_303_),
    .S1(_304_),
    .X(_329_));
 sky130_fd_sc_hd__mux4_1 _665_ (.A0(\ram[8][5] ),
    .A1(\ram[9][5] ),
    .A2(\ram[10][5] ),
    .A3(\ram[11][5] ),
    .S0(_283_),
    .S1(_284_),
    .X(_330_));
 sky130_fd_sc_hd__a22oi_1 _666_ (.A1(_295_),
    .A2(_329_),
    .B1(_330_),
    .B2(_298_),
    .Y(_331_));
 sky130_fd_sc_hd__nand2_1 _667_ (.A(_328_),
    .B(_331_),
    .Y(_013_));
 sky130_fd_sc_hd__mux4_1 _668_ (.A0(\ram[4][6] ),
    .A1(\ram[5][6] ),
    .A2(\ram[6][6] ),
    .A3(\ram[7][6] ),
    .S0(_303_),
    .S1(_304_),
    .X(_332_));
 sky130_fd_sc_hd__mux4_2 _669_ (.A0(\ram[12][6] ),
    .A1(\ram[13][6] ),
    .A2(\ram[14][6] ),
    .A3(\ram[15][6] ),
    .S0(_288_),
    .S1(_289_),
    .X(_333_));
 sky130_fd_sc_hd__a22oi_2 _670_ (.A1(_287_),
    .A2(_332_),
    .B1(_333_),
    .B2(_292_),
    .Y(_334_));
 sky130_fd_sc_hd__mux4_1 _671_ (.A0(\ram[0][6] ),
    .A1(\ram[1][6] ),
    .A2(\ram[2][6] ),
    .A3(\ram[3][6] ),
    .S0(_163_),
    .S1(_174_),
    .X(_335_));
 sky130_fd_sc_hd__mux4_1 _672_ (.A0(\ram[8][6] ),
    .A1(\ram[9][6] ),
    .A2(\ram[10][6] ),
    .A3(\ram[11][6] ),
    .S0(_283_),
    .S1(_284_),
    .X(_336_));
 sky130_fd_sc_hd__a22oi_1 _673_ (.A1(_295_),
    .A2(_335_),
    .B1(_336_),
    .B2(_298_),
    .Y(_337_));
 sky130_fd_sc_hd__nand2_1 _674_ (.A(_334_),
    .B(_337_),
    .Y(_014_));
 sky130_fd_sc_hd__mux4_1 _675_ (.A0(\ram[4][7] ),
    .A1(\ram[5][7] ),
    .A2(\ram[6][7] ),
    .A3(\ram[7][7] ),
    .S0(_303_),
    .S1(_304_),
    .X(_338_));
 sky130_fd_sc_hd__mux4_2 _676_ (.A0(\ram[12][7] ),
    .A1(\ram[13][7] ),
    .A2(\ram[14][7] ),
    .A3(\ram[15][7] ),
    .S0(_288_),
    .S1(_289_),
    .X(_339_));
 sky130_fd_sc_hd__a22oi_2 _677_ (.A1(_287_),
    .A2(_338_),
    .B1(_339_),
    .B2(_292_),
    .Y(_340_));
 sky130_fd_sc_hd__mux4_1 _678_ (.A0(\ram[0][7] ),
    .A1(\ram[1][7] ),
    .A2(\ram[2][7] ),
    .A3(\ram[3][7] ),
    .S0(_163_),
    .S1(_174_),
    .X(_341_));
 sky130_fd_sc_hd__mux4_1 _679_ (.A0(\ram[8][7] ),
    .A1(\ram[9][7] ),
    .A2(\ram[10][7] ),
    .A3(\ram[11][7] ),
    .S0(_283_),
    .S1(_284_),
    .X(_342_));
 sky130_fd_sc_hd__a22oi_1 _680_ (.A1(_295_),
    .A2(_341_),
    .B1(_342_),
    .B2(_298_),
    .Y(_343_));
 sky130_fd_sc_hd__nand2_1 _681_ (.A(_340_),
    .B(_343_),
    .Y(_015_));
 sky130_fd_sc_hd__mux2_1 _682_ (.A0(_202_),
    .A1(net12),
    .S(_184_),
    .X(_032_));
 sky130_fd_sc_hd__mux2_1 _683_ (.A0(_203_),
    .A1(net13),
    .S(_184_),
    .X(_033_));
 sky130_fd_sc_hd__mux2_1 _684_ (.A0(_204_),
    .A1(net14),
    .S(_184_),
    .X(_034_));
 sky130_fd_sc_hd__mux2_1 _685_ (.A0(_205_),
    .A1(net15),
    .S(_184_),
    .X(_035_));
 sky130_fd_sc_hd__mux2_1 _686_ (.A0(_206_),
    .A1(net16),
    .S(_184_),
    .X(_036_));
 sky130_fd_sc_hd__mux2_1 _687_ (.A0(_207_),
    .A1(net17),
    .S(_184_),
    .X(_037_));
 sky130_fd_sc_hd__dfxtp_1 \q_a[0]$_DFF_P_  (.D(_008_),
    .Q(net22),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \q_a[1]$_DFF_P_  (.D(_009_),
    .Q(net23),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \q_a[2]$_DFF_P_  (.D(_010_),
    .Q(net24),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \q_a[3]$_DFF_P_  (.D(_011_),
    .Q(net25),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \q_a[4]$_DFF_P_  (.D(_012_),
    .Q(net26),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \q_a[5]$_DFF_P_  (.D(_013_),
    .Q(net27),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \q_a[6]$_DFF_P_  (.D(_014_),
    .Q(net28),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \q_a[7]$_DFF_P_  (.D(_015_),
    .Q(net29),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \q_b[0]$_DFF_P_  (.D(_000_),
    .Q(net30),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \q_b[1]$_DFF_P_  (.D(_001_),
    .Q(net31),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \q_b[2]$_DFF_P_  (.D(_002_),
    .Q(net32),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \q_b[3]$_DFF_P_  (.D(_003_),
    .Q(net33),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \q_b[4]$_DFF_P_  (.D(_004_),
    .Q(net34),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \q_b[5]$_DFF_P_  (.D(_005_),
    .Q(net35),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \q_b[6]$_DFF_P_  (.D(_006_),
    .Q(net36),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \q_b[7]$_DFF_P_  (.D(_007_),
    .Q(net37),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[0][0]$_DFFE_PP_  (.D(_032_),
    .DE(_031_),
    .Q(\ram[0][0] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[0][1]$_DFFE_PP_  (.D(_033_),
    .DE(_031_),
    .Q(\ram[0][1] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[0][2]$_DFFE_PP_  (.D(_034_),
    .DE(_031_),
    .Q(\ram[0][2] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[0][3]$_DFFE_PP_  (.D(_035_),
    .DE(_031_),
    .Q(\ram[0][3] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[0][4]$_DFFE_PP_  (.D(_036_),
    .DE(_031_),
    .Q(\ram[0][4] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[0][5]$_DFFE_PP_  (.D(_037_),
    .DE(_031_),
    .Q(\ram[0][5] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[0][6]$_DFFE_PP_  (.D(_038_),
    .DE(_031_),
    .Q(\ram[0][6] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[0][7]$_DFFE_PP_  (.D(_039_),
    .DE(_031_),
    .Q(\ram[0][7] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[10][0]$_DFFE_PP_  (.D(_040_),
    .DE(_030_),
    .Q(\ram[10][0] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[10][1]$_DFFE_PP_  (.D(_041_),
    .DE(_030_),
    .Q(\ram[10][1] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[10][2]$_DFFE_PP_  (.D(_042_),
    .DE(_030_),
    .Q(\ram[10][2] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[10][3]$_DFFE_PP_  (.D(_043_),
    .DE(_030_),
    .Q(\ram[10][3] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[10][4]$_DFFE_PP_  (.D(_044_),
    .DE(_030_),
    .Q(\ram[10][4] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[10][5]$_DFFE_PP_  (.D(_045_),
    .DE(_030_),
    .Q(\ram[10][5] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[10][6]$_DFFE_PP_  (.D(_046_),
    .DE(_030_),
    .Q(\ram[10][6] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[10][7]$_DFFE_PP_  (.D(_047_),
    .DE(_030_),
    .Q(\ram[10][7] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[11][0]$_DFFE_PP_  (.D(_048_),
    .DE(_029_),
    .Q(\ram[11][0] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[11][1]$_DFFE_PP_  (.D(_049_),
    .DE(_029_),
    .Q(\ram[11][1] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[11][2]$_DFFE_PP_  (.D(_050_),
    .DE(_029_),
    .Q(\ram[11][2] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[11][3]$_DFFE_PP_  (.D(_051_),
    .DE(_029_),
    .Q(\ram[11][3] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[11][4]$_DFFE_PP_  (.D(_052_),
    .DE(_029_),
    .Q(\ram[11][4] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[11][5]$_DFFE_PP_  (.D(_053_),
    .DE(_029_),
    .Q(\ram[11][5] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[11][6]$_DFFE_PP_  (.D(_054_),
    .DE(_029_),
    .Q(\ram[11][6] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[11][7]$_DFFE_PP_  (.D(_055_),
    .DE(_029_),
    .Q(\ram[11][7] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[12][0]$_DFFE_PP_  (.D(_056_),
    .DE(_028_),
    .Q(\ram[12][0] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[12][1]$_DFFE_PP_  (.D(_057_),
    .DE(_028_),
    .Q(\ram[12][1] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[12][2]$_DFFE_PP_  (.D(_058_),
    .DE(_028_),
    .Q(\ram[12][2] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[12][3]$_DFFE_PP_  (.D(_059_),
    .DE(_028_),
    .Q(\ram[12][3] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[12][4]$_DFFE_PP_  (.D(_060_),
    .DE(_028_),
    .Q(\ram[12][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[12][5]$_DFFE_PP_  (.D(_061_),
    .DE(_028_),
    .Q(\ram[12][5] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[12][6]$_DFFE_PP_  (.D(_062_),
    .DE(_028_),
    .Q(\ram[12][6] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[12][7]$_DFFE_PP_  (.D(_063_),
    .DE(_028_),
    .Q(\ram[12][7] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[13][0]$_DFFE_PP_  (.D(_064_),
    .DE(_027_),
    .Q(\ram[13][0] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[13][1]$_DFFE_PP_  (.D(_065_),
    .DE(_027_),
    .Q(\ram[13][1] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[13][2]$_DFFE_PP_  (.D(_066_),
    .DE(_027_),
    .Q(\ram[13][2] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[13][3]$_DFFE_PP_  (.D(_067_),
    .DE(_027_),
    .Q(\ram[13][3] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[13][4]$_DFFE_PP_  (.D(_068_),
    .DE(_027_),
    .Q(\ram[13][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[13][5]$_DFFE_PP_  (.D(_069_),
    .DE(_027_),
    .Q(\ram[13][5] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[13][6]$_DFFE_PP_  (.D(_070_),
    .DE(_027_),
    .Q(\ram[13][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[13][7]$_DFFE_PP_  (.D(_071_),
    .DE(_027_),
    .Q(\ram[13][7] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[14][0]$_DFFE_PP_  (.D(_072_),
    .DE(_026_),
    .Q(\ram[14][0] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[14][1]$_DFFE_PP_  (.D(_073_),
    .DE(_026_),
    .Q(\ram[14][1] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[14][2]$_DFFE_PP_  (.D(_074_),
    .DE(_026_),
    .Q(\ram[14][2] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[14][3]$_DFFE_PP_  (.D(_075_),
    .DE(_026_),
    .Q(\ram[14][3] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[14][4]$_DFFE_PP_  (.D(_076_),
    .DE(_026_),
    .Q(\ram[14][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[14][5]$_DFFE_PP_  (.D(_077_),
    .DE(_026_),
    .Q(\ram[14][5] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[14][6]$_DFFE_PP_  (.D(_078_),
    .DE(_026_),
    .Q(\ram[14][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[14][7]$_DFFE_PP_  (.D(_079_),
    .DE(_026_),
    .Q(\ram[14][7] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[15][0]$_DFFE_PP_  (.D(_080_),
    .DE(_025_),
    .Q(\ram[15][0] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[15][1]$_DFFE_PP_  (.D(_081_),
    .DE(_025_),
    .Q(\ram[15][1] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[15][2]$_DFFE_PP_  (.D(_082_),
    .DE(_025_),
    .Q(\ram[15][2] ),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[15][3]$_DFFE_PP_  (.D(_083_),
    .DE(_025_),
    .Q(\ram[15][3] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[15][4]$_DFFE_PP_  (.D(_084_),
    .DE(_025_),
    .Q(\ram[15][4] ),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[15][5]$_DFFE_PP_  (.D(_085_),
    .DE(_025_),
    .Q(\ram[15][5] ),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[15][6]$_DFFE_PP_  (.D(_086_),
    .DE(_025_),
    .Q(\ram[15][6] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[15][7]$_DFFE_PP_  (.D(_087_),
    .DE(_025_),
    .Q(\ram[15][7] ),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[1][0]$_DFFE_PP_  (.D(_088_),
    .DE(_024_),
    .Q(\ram[1][0] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[1][1]$_DFFE_PP_  (.D(_089_),
    .DE(_024_),
    .Q(\ram[1][1] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[1][2]$_DFFE_PP_  (.D(_090_),
    .DE(_024_),
    .Q(\ram[1][2] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[1][3]$_DFFE_PP_  (.D(_091_),
    .DE(_024_),
    .Q(\ram[1][3] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[1][4]$_DFFE_PP_  (.D(_092_),
    .DE(_024_),
    .Q(\ram[1][4] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[1][5]$_DFFE_PP_  (.D(_093_),
    .DE(_024_),
    .Q(\ram[1][5] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[1][6]$_DFFE_PP_  (.D(_094_),
    .DE(_024_),
    .Q(\ram[1][6] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[1][7]$_DFFE_PP_  (.D(_095_),
    .DE(_024_),
    .Q(\ram[1][7] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[2][0]$_DFFE_PP_  (.D(_096_),
    .DE(_023_),
    .Q(\ram[2][0] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[2][1]$_DFFE_PP_  (.D(_097_),
    .DE(_023_),
    .Q(\ram[2][1] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[2][2]$_DFFE_PP_  (.D(_098_),
    .DE(_023_),
    .Q(\ram[2][2] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[2][3]$_DFFE_PP_  (.D(_099_),
    .DE(_023_),
    .Q(\ram[2][3] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[2][4]$_DFFE_PP_  (.D(_100_),
    .DE(_023_),
    .Q(\ram[2][4] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[2][5]$_DFFE_PP_  (.D(_101_),
    .DE(_023_),
    .Q(\ram[2][5] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[2][6]$_DFFE_PP_  (.D(_102_),
    .DE(_023_),
    .Q(\ram[2][6] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[2][7]$_DFFE_PP_  (.D(_103_),
    .DE(_023_),
    .Q(\ram[2][7] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[3][0]$_DFFE_PP_  (.D(_104_),
    .DE(_022_),
    .Q(\ram[3][0] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[3][1]$_DFFE_PP_  (.D(_105_),
    .DE(_022_),
    .Q(\ram[3][1] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[3][2]$_DFFE_PP_  (.D(_106_),
    .DE(_022_),
    .Q(\ram[3][2] ),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[3][3]$_DFFE_PP_  (.D(_107_),
    .DE(_022_),
    .Q(\ram[3][3] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[3][4]$_DFFE_PP_  (.D(_108_),
    .DE(_022_),
    .Q(\ram[3][4] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[3][5]$_DFFE_PP_  (.D(_109_),
    .DE(_022_),
    .Q(\ram[3][5] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[3][6]$_DFFE_PP_  (.D(_110_),
    .DE(_022_),
    .Q(\ram[3][6] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[3][7]$_DFFE_PP_  (.D(_111_),
    .DE(_022_),
    .Q(\ram[3][7] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[4][0]$_DFFE_PP_  (.D(_112_),
    .DE(_021_),
    .Q(\ram[4][0] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[4][1]$_DFFE_PP_  (.D(_113_),
    .DE(_021_),
    .Q(\ram[4][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[4][2]$_DFFE_PP_  (.D(_114_),
    .DE(_021_),
    .Q(\ram[4][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[4][3]$_DFFE_PP_  (.D(_115_),
    .DE(_021_),
    .Q(\ram[4][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[4][4]$_DFFE_PP_  (.D(_116_),
    .DE(_021_),
    .Q(\ram[4][4] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[4][5]$_DFFE_PP_  (.D(_117_),
    .DE(_021_),
    .Q(\ram[4][5] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[4][6]$_DFFE_PP_  (.D(_118_),
    .DE(_021_),
    .Q(\ram[4][6] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[4][7]$_DFFE_PP_  (.D(_119_),
    .DE(_021_),
    .Q(\ram[4][7] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[5][0]$_DFFE_PP_  (.D(_120_),
    .DE(_020_),
    .Q(\ram[5][0] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[5][1]$_DFFE_PP_  (.D(_121_),
    .DE(_020_),
    .Q(\ram[5][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[5][2]$_DFFE_PP_  (.D(_122_),
    .DE(_020_),
    .Q(\ram[5][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[5][3]$_DFFE_PP_  (.D(_123_),
    .DE(_020_),
    .Q(\ram[5][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[5][4]$_DFFE_PP_  (.D(_124_),
    .DE(_020_),
    .Q(\ram[5][4] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[5][5]$_DFFE_PP_  (.D(_125_),
    .DE(_020_),
    .Q(\ram[5][5] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[5][6]$_DFFE_PP_  (.D(_126_),
    .DE(_020_),
    .Q(\ram[5][6] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[5][7]$_DFFE_PP_  (.D(_127_),
    .DE(_020_),
    .Q(\ram[5][7] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[6][0]$_DFFE_PP_  (.D(_128_),
    .DE(_019_),
    .Q(\ram[6][0] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[6][1]$_DFFE_PP_  (.D(_129_),
    .DE(_019_),
    .Q(\ram[6][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[6][2]$_DFFE_PP_  (.D(_130_),
    .DE(_019_),
    .Q(\ram[6][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[6][3]$_DFFE_PP_  (.D(_131_),
    .DE(_019_),
    .Q(\ram[6][3] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[6][4]$_DFFE_PP_  (.D(_132_),
    .DE(_019_),
    .Q(\ram[6][4] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[6][5]$_DFFE_PP_  (.D(_133_),
    .DE(_019_),
    .Q(\ram[6][5] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[6][6]$_DFFE_PP_  (.D(_134_),
    .DE(_019_),
    .Q(\ram[6][6] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[6][7]$_DFFE_PP_  (.D(_135_),
    .DE(_019_),
    .Q(\ram[6][7] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[7][0]$_DFFE_PP_  (.D(_136_),
    .DE(_018_),
    .Q(\ram[7][0] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[7][1]$_DFFE_PP_  (.D(_137_),
    .DE(_018_),
    .Q(\ram[7][1] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[7][2]$_DFFE_PP_  (.D(_138_),
    .DE(_018_),
    .Q(\ram[7][2] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[7][3]$_DFFE_PP_  (.D(_139_),
    .DE(_018_),
    .Q(\ram[7][3] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[7][4]$_DFFE_PP_  (.D(_140_),
    .DE(_018_),
    .Q(\ram[7][4] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[7][5]$_DFFE_PP_  (.D(_141_),
    .DE(_018_),
    .Q(\ram[7][5] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[7][6]$_DFFE_PP_  (.D(_142_),
    .DE(_018_),
    .Q(\ram[7][6] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[7][7]$_DFFE_PP_  (.D(_143_),
    .DE(_018_),
    .Q(\ram[7][7] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[8][0]$_DFFE_PP_  (.D(_144_),
    .DE(_017_),
    .Q(\ram[8][0] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[8][1]$_DFFE_PP_  (.D(_145_),
    .DE(_017_),
    .Q(\ram[8][1] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[8][2]$_DFFE_PP_  (.D(_146_),
    .DE(_017_),
    .Q(\ram[8][2] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[8][3]$_DFFE_PP_  (.D(_147_),
    .DE(_017_),
    .Q(\ram[8][3] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[8][4]$_DFFE_PP_  (.D(_148_),
    .DE(_017_),
    .Q(\ram[8][4] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[8][5]$_DFFE_PP_  (.D(_149_),
    .DE(_017_),
    .Q(\ram[8][5] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[8][6]$_DFFE_PP_  (.D(_150_),
    .DE(_017_),
    .Q(\ram[8][6] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[8][7]$_DFFE_PP_  (.D(_151_),
    .DE(_017_),
    .Q(\ram[8][7] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[9][0]$_DFFE_PP_  (.D(_152_),
    .DE(_016_),
    .Q(\ram[9][0] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[9][1]$_DFFE_PP_  (.D(_153_),
    .DE(_016_),
    .Q(\ram[9][1] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[9][2]$_DFFE_PP_  (.D(_154_),
    .DE(_016_),
    .Q(\ram[9][2] ),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[9][3]$_DFFE_PP_  (.D(_155_),
    .DE(_016_),
    .Q(\ram[9][3] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[9][4]$_DFFE_PP_  (.D(_156_),
    .DE(_016_),
    .Q(\ram[9][4] ),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[9][5]$_DFFE_PP_  (.D(_157_),
    .DE(_016_),
    .Q(\ram[9][5] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[9][6]$_DFFE_PP_  (.D(_158_),
    .DE(_016_),
    .Q(\ram[9][6] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \ram[9][7]$_DFFE_PP_  (.D(_159_),
    .DE(_016_),
    .Q(\ram[9][7] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_179 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(addr_a[1]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(addr_b[2]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(addr_b[3]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(data_a[0]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(data_a[1]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(data_a[2]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(data_a[3]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(data_a[4]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input9 (.A(data_a[5]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(data_a[6]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 input11 (.A(data_a[7]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(data_b[0]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(data_b[1]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(data_b[2]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(data_b[3]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(data_b[4]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(data_b[5]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(data_b[6]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(data_b[7]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(we_a),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(we_b),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net22),
    .X(q_a[0]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net23),
    .X(q_a[1]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net24),
    .X(q_a[2]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net25),
    .X(q_a[3]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net26),
    .X(q_a[4]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net27),
    .X(q_a[5]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net28),
    .X(q_a[6]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net29),
    .X(q_a[7]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net30),
    .X(q_b[0]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net31),
    .X(q_b[1]));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(net32),
    .X(q_b[2]));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net33),
    .X(q_b[3]));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net34),
    .X(q_b[4]));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(net35),
    .X(q_b[5]));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net36),
    .X(q_b[6]));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(net37),
    .X(q_b[7]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload1 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload2 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload3 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload4 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload5 (.A(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload6 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload7 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload8 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload9 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload10 (.A(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload11 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload12 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload13 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload14 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_30 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_210 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_54 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_25 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_126 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_258 ();
endmodule
