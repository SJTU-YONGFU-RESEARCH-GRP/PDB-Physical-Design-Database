module barrel_shifter (rotate,
    shift_direction,
    data_in,
    data_out,
    shift_amount);
 input rotate;
 input shift_direction;
 input [31:0] data_in;
 output [31:0] data_out;
 input [4:0] shift_amount;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;

 sky130_fd_sc_hd__buf_6 _0924_ (.A(net33),
    .X(_0672_));
 sky130_fd_sc_hd__buf_6 _0925_ (.A(_0672_),
    .X(_0683_));
 sky130_fd_sc_hd__clkinv_2 _0926_ (.A(_0683_),
    .Y(_0693_));
 sky130_fd_sc_hd__buf_6 _0927_ (.A(_0693_),
    .X(_0704_));
 sky130_fd_sc_hd__buf_4 _0928_ (.A(_0704_),
    .X(_0920_));
 sky130_fd_sc_hd__buf_4 _0929_ (.A(net34),
    .X(_0724_));
 sky130_fd_sc_hd__buf_6 _0930_ (.A(_0724_),
    .X(_0734_));
 sky130_fd_sc_hd__buf_4 _0931_ (.A(_0734_),
    .X(_0745_));
 sky130_fd_sc_hd__clkinv_2 _0932_ (.A(_0745_),
    .Y(_0921_));
 sky130_fd_sc_hd__buf_6 _0933_ (.A(_0672_),
    .X(_0765_));
 sky130_fd_sc_hd__buf_6 _0934_ (.A(_0765_),
    .X(_0775_));
 sky130_fd_sc_hd__buf_6 _0935_ (.A(_0775_),
    .X(_0785_));
 sky130_fd_sc_hd__nor2b_2 _0936_ (.A(_0785_),
    .B_N(net1),
    .Y(_0796_));
 sky130_fd_sc_hd__buf_6 _0937_ (.A(_0923_),
    .X(_0806_));
 sky130_fd_sc_hd__buf_6 _0938_ (.A(_0806_),
    .X(_0816_));
 sky130_fd_sc_hd__buf_4 _0939_ (.A(_0816_),
    .X(_0826_));
 sky130_fd_sc_hd__buf_4 _0940_ (.A(_0826_),
    .X(_0837_));
 sky130_fd_sc_hd__buf_4 _0941_ (.A(_0837_),
    .X(_0847_));
 sky130_fd_sc_hd__buf_4 _0942_ (.A(_0922_),
    .X(_0858_));
 sky130_fd_sc_hd__buf_4 _0943_ (.A(shift_amount[3]),
    .X(_0868_));
 sky130_fd_sc_hd__nor4_4 _0944_ (.A(_0868_),
    .B(net35),
    .C(net33),
    .D(net34),
    .Y(_0879_));
 sky130_fd_sc_hd__nor2_2 _0945_ (.A(_0672_),
    .B(_0724_),
    .Y(_0889_));
 sky130_fd_sc_hd__buf_6 _0946_ (.A(net35),
    .X(_0899_));
 sky130_fd_sc_hd__nand2b_1 _0947_ (.A_N(_0899_),
    .B(_0922_),
    .Y(_0910_));
 sky130_fd_sc_hd__nand2b_1 _0948_ (.A_N(_0858_),
    .B(_0899_),
    .Y(_0000_));
 sky130_fd_sc_hd__o21ai_1 _0949_ (.A1(_0889_),
    .A2(_0910_),
    .B1(_0000_),
    .Y(_0010_));
 sky130_fd_sc_hd__buf_6 _0950_ (.A(_0868_),
    .X(_0020_));
 sky130_fd_sc_hd__a22oi_4 _0951_ (.A1(_0858_),
    .A2(_0879_),
    .B1(_0010_),
    .B2(_0020_),
    .Y(_0030_));
 sky130_fd_sc_hd__buf_6 _0952_ (.A(shift_amount[4]),
    .X(_0031_));
 sky130_fd_sc_hd__or4_4 _0953_ (.A(_0031_),
    .B(_0868_),
    .C(_0899_),
    .D(_0724_),
    .X(_0032_));
 sky130_fd_sc_hd__o21a_2 _0954_ (.A1(_0775_),
    .A2(_0032_),
    .B1(net32),
    .X(_0033_));
 sky130_fd_sc_hd__inv_4 _0955_ (.A(_0031_),
    .Y(_0034_));
 sky130_fd_sc_hd__nor3b_4 _0956_ (.A(_0868_),
    .B(_0899_),
    .C_N(_0858_),
    .Y(_0035_));
 sky130_fd_sc_hd__xnor2_4 _0957_ (.A(_0034_),
    .B(_0035_),
    .Y(_0036_));
 sky130_fd_sc_hd__nand2_4 _0958_ (.A(_0033_),
    .B(_0036_),
    .Y(_0037_));
 sky130_fd_sc_hd__buf_4 _0959_ (.A(_0037_),
    .X(_0038_));
 sky130_fd_sc_hd__nor3_1 _0960_ (.A(_0847_),
    .B(_0030_),
    .C(_0038_),
    .Y(_0039_));
 sky130_fd_sc_hd__buf_4 _0961_ (.A(shift_direction),
    .X(_0040_));
 sky130_fd_sc_hd__buf_2 _0962_ (.A(_0040_),
    .X(_0041_));
 sky130_fd_sc_hd__buf_2 _0963_ (.A(_0041_),
    .X(_0042_));
 sky130_fd_sc_hd__buf_2 _0964_ (.A(_0031_),
    .X(_0043_));
 sky130_fd_sc_hd__clkbuf_4 _0965_ (.A(_0043_),
    .X(_0044_));
 sky130_fd_sc_hd__buf_2 _0966_ (.A(_0020_),
    .X(_0045_));
 sky130_fd_sc_hd__clkbuf_4 _0967_ (.A(_0045_),
    .X(_0046_));
 sky130_fd_sc_hd__buf_2 _0968_ (.A(net18),
    .X(_0047_));
 sky130_fd_sc_hd__buf_2 _0969_ (.A(net20),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _0970_ (.A0(_0047_),
    .A1(_0048_),
    .S(_0724_),
    .X(_0049_));
 sky130_fd_sc_hd__buf_2 _0971_ (.A(net17),
    .X(_0050_));
 sky130_fd_sc_hd__buf_2 _0972_ (.A(net19),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _0973_ (.A0(_0050_),
    .A1(_0051_),
    .S(_0724_),
    .X(_0052_));
 sky130_fd_sc_hd__buf_6 _0974_ (.A(_0693_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2i_4 _0975_ (.A0(_0049_),
    .A1(_0052_),
    .S(_0053_),
    .Y(_0054_));
 sky130_fd_sc_hd__buf_2 _0976_ (.A(net22),
    .X(_0055_));
 sky130_fd_sc_hd__buf_4 _0977_ (.A(data_in[31]),
    .X(_0056_));
 sky130_fd_sc_hd__mux2i_2 _0978_ (.A0(_0055_),
    .A1(_0056_),
    .S(_0734_),
    .Y(_0057_));
 sky130_fd_sc_hd__buf_2 _0979_ (.A(net21),
    .X(_0058_));
 sky130_fd_sc_hd__clkbuf_4 _0980_ (.A(net24),
    .X(_0059_));
 sky130_fd_sc_hd__clkbuf_4 _0981_ (.A(_0724_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2i_1 _0982_ (.A0(_0058_),
    .A1(_0059_),
    .S(_0060_),
    .Y(_0061_));
 sky130_fd_sc_hd__mux2_4 _0983_ (.A0(_0057_),
    .A1(_0061_),
    .S(_0053_),
    .X(_0062_));
 sky130_fd_sc_hd__buf_4 _0984_ (.A(_0899_),
    .X(_0063_));
 sky130_fd_sc_hd__buf_4 _0985_ (.A(_0063_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2i_4 _0986_ (.A0(_0054_),
    .A1(_0062_),
    .S(_0064_),
    .Y(_0065_));
 sky130_fd_sc_hd__clkbuf_4 _0987_ (.A(_0020_),
    .X(_0066_));
 sky130_fd_sc_hd__mux4_4 _0988_ (.A0(net13),
    .A1(net14),
    .A2(net15),
    .A3(net16),
    .S0(_0683_),
    .S1(_0734_),
    .X(_0067_));
 sky130_fd_sc_hd__clkbuf_4 _0989_ (.A(net8),
    .X(_0068_));
 sky130_fd_sc_hd__buf_2 _0990_ (.A(net9),
    .X(_0069_));
 sky130_fd_sc_hd__buf_2 _0991_ (.A(net10),
    .X(_0070_));
 sky130_fd_sc_hd__buf_2 _0992_ (.A(net11),
    .X(_0071_));
 sky130_fd_sc_hd__buf_4 _0993_ (.A(_0672_),
    .X(_0072_));
 sky130_fd_sc_hd__mux4_4 _0994_ (.A0(_0068_),
    .A1(_0069_),
    .A2(_0070_),
    .A3(_0071_),
    .S0(_0072_),
    .S1(_0745_),
    .X(_0073_));
 sky130_fd_sc_hd__inv_1 _0995_ (.A(_0063_),
    .Y(_0074_));
 sky130_fd_sc_hd__buf_6 _0996_ (.A(_0074_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2i_4 _0997_ (.A0(_0067_),
    .A1(_0073_),
    .S(_0075_),
    .Y(_0076_));
 sky130_fd_sc_hd__nor2_1 _0998_ (.A(_0066_),
    .B(_0076_),
    .Y(_0077_));
 sky130_fd_sc_hd__a21oi_1 _0999_ (.A1(_0046_),
    .A2(_0065_),
    .B1(_0077_),
    .Y(_0078_));
 sky130_fd_sc_hd__clkbuf_4 _1000_ (.A(net26),
    .X(_0079_));
 sky130_fd_sc_hd__clkbuf_4 _1001_ (.A(net27),
    .X(_0080_));
 sky130_fd_sc_hd__buf_2 _1002_ (.A(net28),
    .X(_0081_));
 sky130_fd_sc_hd__clkbuf_4 _1003_ (.A(net29),
    .X(_0082_));
 sky130_fd_sc_hd__buf_6 _1004_ (.A(_0683_),
    .X(_0083_));
 sky130_fd_sc_hd__clkbuf_4 _1005_ (.A(_0734_),
    .X(_0084_));
 sky130_fd_sc_hd__mux4_1 _1006_ (.A0(_0079_),
    .A1(_0080_),
    .A2(_0081_),
    .A3(_0082_),
    .S0(_0083_),
    .S1(_0084_),
    .X(_0085_));
 sky130_fd_sc_hd__nor2_1 _1007_ (.A(_0075_),
    .B(_0085_),
    .Y(_0086_));
 sky130_fd_sc_hd__buf_2 _1008_ (.A(_0063_),
    .X(_0087_));
 sky130_fd_sc_hd__clkbuf_4 _1009_ (.A(net23),
    .X(_0088_));
 sky130_fd_sc_hd__clkbuf_4 _1010_ (.A(net25),
    .X(_0089_));
 sky130_fd_sc_hd__clkbuf_4 _1011_ (.A(_0060_),
    .X(_0090_));
 sky130_fd_sc_hd__mux4_1 _1012_ (.A0(net1),
    .A1(net12),
    .A2(_0088_),
    .A3(_0089_),
    .S0(_0775_),
    .S1(_0090_),
    .X(_0091_));
 sky130_fd_sc_hd__nor2_1 _1013_ (.A(_0087_),
    .B(_0091_),
    .Y(_0092_));
 sky130_fd_sc_hd__buf_4 _1014_ (.A(net5),
    .X(_0093_));
 sky130_fd_sc_hd__buf_4 _1015_ (.A(net6),
    .X(_0094_));
 sky130_fd_sc_hd__clkbuf_4 _1016_ (.A(net7),
    .X(_0095_));
 sky130_fd_sc_hd__buf_4 _1017_ (.A(_0672_),
    .X(_0096_));
 sky130_fd_sc_hd__clkbuf_4 _1018_ (.A(_0724_),
    .X(_0097_));
 sky130_fd_sc_hd__mux4_2 _1019_ (.A0(net4),
    .A1(_0093_),
    .A2(_0094_),
    .A3(_0095_),
    .S0(_0096_),
    .S1(_0097_),
    .X(_0098_));
 sky130_fd_sc_hd__buf_2 _1020_ (.A(net3),
    .X(_0099_));
 sky130_fd_sc_hd__mux4_1 _1021_ (.A0(net30),
    .A1(net31),
    .A2(net2),
    .A3(_0099_),
    .S0(_0096_),
    .S1(_0097_),
    .X(_0100_));
 sky130_fd_sc_hd__buf_4 _1022_ (.A(_0074_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _1023_ (.A0(_0098_),
    .A1(_0100_),
    .S(_0101_),
    .X(_0102_));
 sky130_fd_sc_hd__nand2_1 _1024_ (.A(_0066_),
    .B(_0102_),
    .Y(_0103_));
 sky130_fd_sc_hd__o311a_1 _1025_ (.A1(_0045_),
    .A2(_0086_),
    .A3(_0092_),
    .B1(_0103_),
    .C1(_0034_),
    .X(_0104_));
 sky130_fd_sc_hd__a21oi_1 _1026_ (.A1(_0044_),
    .A2(_0078_),
    .B1(_0104_),
    .Y(_0105_));
 sky130_fd_sc_hd__a211oi_1 _1027_ (.A1(_0796_),
    .A2(_0039_),
    .B1(_0042_),
    .C1(_0105_),
    .Y(_0106_));
 sky130_fd_sc_hd__o21ai_4 _1028_ (.A1(_0775_),
    .A2(_0032_),
    .B1(net32),
    .Y(_0107_));
 sky130_fd_sc_hd__xnor2_4 _1029_ (.A(_0031_),
    .B(_0035_),
    .Y(_0108_));
 sky130_fd_sc_hd__nor2_1 _1030_ (.A(_0107_),
    .B(_0108_),
    .Y(_0109_));
 sky130_fd_sc_hd__buf_6 _1031_ (.A(_0109_),
    .X(_0110_));
 sky130_fd_sc_hd__buf_4 _1032_ (.A(_0110_),
    .X(_0111_));
 sky130_fd_sc_hd__xnor2_4 _1033_ (.A(_0899_),
    .B(_0858_),
    .Y(_0112_));
 sky130_fd_sc_hd__buf_4 _1034_ (.A(_0112_),
    .X(_0113_));
 sky130_fd_sc_hd__clkbuf_4 _1035_ (.A(_0113_),
    .X(_0114_));
 sky130_fd_sc_hd__clkbuf_4 _1036_ (.A(net31),
    .X(_0115_));
 sky130_fd_sc_hd__mux2i_2 _1037_ (.A0(_0115_),
    .A1(_0099_),
    .S(_0826_),
    .Y(_0116_));
 sky130_fd_sc_hd__clkbuf_4 _1038_ (.A(net30),
    .X(_0117_));
 sky130_fd_sc_hd__clkbuf_4 _1039_ (.A(net2),
    .X(_0118_));
 sky130_fd_sc_hd__nand2b_1 _1040_ (.A_N(_0118_),
    .B(_0837_),
    .Y(_0119_));
 sky130_fd_sc_hd__clkbuf_4 _1041_ (.A(_0053_),
    .X(_0120_));
 sky130_fd_sc_hd__o211ai_2 _1042_ (.A1(_0117_),
    .A2(_0847_),
    .B1(_0119_),
    .C1(_0120_),
    .Y(_0121_));
 sky130_fd_sc_hd__o21ai_4 _1043_ (.A1(_0920_),
    .A2(_0116_),
    .B1(_0121_),
    .Y(_0122_));
 sky130_fd_sc_hd__buf_6 _1044_ (.A(_0672_),
    .X(_0123_));
 sky130_fd_sc_hd__buf_6 _1045_ (.A(_0123_),
    .X(_0124_));
 sky130_fd_sc_hd__mux4_1 _1046_ (.A0(net1),
    .A1(net12),
    .A2(_0088_),
    .A3(_0089_),
    .S0(_0124_),
    .S1(_0847_),
    .X(_0125_));
 sky130_fd_sc_hd__o31a_1 _1047_ (.A1(_0899_),
    .A2(_0672_),
    .A3(net34),
    .B1(_0868_),
    .X(_0126_));
 sky130_fd_sc_hd__or2_0 _1048_ (.A(_0879_),
    .B(_0126_),
    .X(_0127_));
 sky130_fd_sc_hd__buf_6 _1049_ (.A(_0127_),
    .X(_0128_));
 sky130_fd_sc_hd__buf_4 _1050_ (.A(_0128_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2i_2 _1051_ (.A0(_0122_),
    .A1(_0125_),
    .S(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hd__buf_6 _1052_ (.A(_0128_),
    .X(_0131_));
 sky130_fd_sc_hd__buf_6 _1053_ (.A(_0131_),
    .X(_0132_));
 sky130_fd_sc_hd__buf_4 _1054_ (.A(_0816_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2i_2 _1055_ (.A0(_0093_),
    .A1(_0095_),
    .S(_0133_),
    .Y(_0134_));
 sky130_fd_sc_hd__clkbuf_4 _1056_ (.A(net4),
    .X(_0135_));
 sky130_fd_sc_hd__mux2i_2 _1057_ (.A0(_0135_),
    .A1(_0094_),
    .S(_0837_),
    .Y(_0136_));
 sky130_fd_sc_hd__mux2i_4 _1058_ (.A0(_0134_),
    .A1(_0136_),
    .S(_0704_),
    .Y(_0137_));
 sky130_fd_sc_hd__buf_4 _1059_ (.A(_0133_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2i_2 _1060_ (.A0(_0080_),
    .A1(_0082_),
    .S(_0138_),
    .Y(_0139_));
 sky130_fd_sc_hd__mux2i_1 _1061_ (.A0(_0079_),
    .A1(_0081_),
    .S(_0837_),
    .Y(_0140_));
 sky130_fd_sc_hd__nand2b_1 _1062_ (.A_N(_0140_),
    .B(_0704_),
    .Y(_0141_));
 sky130_fd_sc_hd__o211ai_2 _1063_ (.A1(_0920_),
    .A2(_0139_),
    .B1(_0141_),
    .C1(_0129_),
    .Y(_0142_));
 sky130_fd_sc_hd__buf_4 _1064_ (.A(_0112_),
    .X(_0143_));
 sky130_fd_sc_hd__buf_4 _1065_ (.A(_0143_),
    .X(_0144_));
 sky130_fd_sc_hd__o211ai_1 _1066_ (.A1(_0132_),
    .A2(_0137_),
    .B1(_0142_),
    .C1(_0144_),
    .Y(_0145_));
 sky130_fd_sc_hd__o21ai_1 _1067_ (.A1(_0114_),
    .A2(_0130_),
    .B1(_0145_),
    .Y(_0146_));
 sky130_fd_sc_hd__nor2_4 _1068_ (.A(_0107_),
    .B(_0036_),
    .Y(_0147_));
 sky130_fd_sc_hd__clkbuf_4 _1069_ (.A(_0147_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2i_4 _1070_ (.A0(net14),
    .A1(net16),
    .S(_0816_),
    .Y(_0149_));
 sky130_fd_sc_hd__buf_2 _1071_ (.A(net13),
    .X(_0150_));
 sky130_fd_sc_hd__buf_2 _1072_ (.A(net15),
    .X(_0151_));
 sky130_fd_sc_hd__mux2i_2 _1073_ (.A0(_0150_),
    .A1(_0151_),
    .S(_0826_),
    .Y(_0152_));
 sky130_fd_sc_hd__mux2i_4 _1074_ (.A0(_0149_),
    .A1(_0152_),
    .S(_0053_),
    .Y(_0153_));
 sky130_fd_sc_hd__mux2i_4 _1075_ (.A0(net9),
    .A1(net11),
    .S(_0816_),
    .Y(_0154_));
 sky130_fd_sc_hd__mux2i_2 _1076_ (.A0(_0068_),
    .A1(_0070_),
    .S(_0826_),
    .Y(_0155_));
 sky130_fd_sc_hd__mux2i_4 _1077_ (.A0(_0154_),
    .A1(_0155_),
    .S(_0053_),
    .Y(_0156_));
 sky130_fd_sc_hd__xor2_4 _1078_ (.A(net35),
    .B(_0922_),
    .X(_0157_));
 sky130_fd_sc_hd__buf_6 _1079_ (.A(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__buf_4 _1080_ (.A(_0158_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2i_2 _1081_ (.A0(_0153_),
    .A1(_0156_),
    .S(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__mux4_4 _1082_ (.A0(net21),
    .A1(net22),
    .A2(net24),
    .A3(_0056_),
    .S0(_0672_),
    .S1(_0816_),
    .X(_0161_));
 sky130_fd_sc_hd__mux4_4 _1083_ (.A0(net17),
    .A1(net18),
    .A2(net19),
    .A3(net20),
    .S0(_0672_),
    .S1(_0816_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_2 _1084_ (.A0(_0161_),
    .A1(_0162_),
    .S(_0158_),
    .X(_0163_));
 sky130_fd_sc_hd__nor2_1 _1085_ (.A(_0131_),
    .B(_0163_),
    .Y(_0164_));
 sky130_fd_sc_hd__a21oi_2 _1086_ (.A1(_0131_),
    .A2(_0160_),
    .B1(_0164_),
    .Y(_0165_));
 sky130_fd_sc_hd__nand2b_2 _1087_ (.A_N(_0123_),
    .B(net1),
    .Y(_0166_));
 sky130_fd_sc_hd__clkbuf_4 _1088_ (.A(_0040_),
    .X(_0167_));
 sky130_fd_sc_hd__o21ai_0 _1089_ (.A1(_0166_),
    .A2(_0032_),
    .B1(_0167_),
    .Y(_0168_));
 sky130_fd_sc_hd__a221oi_1 _1090_ (.A1(_0111_),
    .A2(_0146_),
    .B1(_0148_),
    .B2(_0165_),
    .C1(_0168_),
    .Y(_0169_));
 sky130_fd_sc_hd__nor2_1 _1091_ (.A(_0106_),
    .B(_0169_),
    .Y(net36));
 sky130_fd_sc_hd__clkbuf_4 _1092_ (.A(_0034_),
    .X(_0170_));
 sky130_fd_sc_hd__mux4_2 _1093_ (.A0(net15),
    .A1(net16),
    .A2(net17),
    .A3(_0047_),
    .S0(_0683_),
    .S1(_0734_),
    .X(_0171_));
 sky130_fd_sc_hd__buf_2 _1094_ (.A(net14),
    .X(_0172_));
 sky130_fd_sc_hd__mux4_1 _1095_ (.A0(_0070_),
    .A1(_0071_),
    .A2(_0150_),
    .A3(_0172_),
    .S0(_0083_),
    .S1(_0084_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2i_1 _1096_ (.A0(_0171_),
    .A1(_0173_),
    .S(_0075_),
    .Y(_0174_));
 sky130_fd_sc_hd__mux4_2 _1097_ (.A0(net6),
    .A1(net7),
    .A2(net8),
    .A3(net9),
    .S0(_0765_),
    .S1(_0060_),
    .X(_0175_));
 sky130_fd_sc_hd__mux4_2 _1098_ (.A0(net2),
    .A1(net3),
    .A2(net4),
    .A3(net5),
    .S0(_0683_),
    .S1(_0060_),
    .X(_0176_));
 sky130_fd_sc_hd__buf_6 _1099_ (.A(_0074_),
    .X(_0177_));
 sky130_fd_sc_hd__clkbuf_4 _1100_ (.A(_0177_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2i_1 _1101_ (.A0(_0175_),
    .A1(_0176_),
    .S(_0178_),
    .Y(_0179_));
 sky130_fd_sc_hd__inv_2 _1102_ (.A(_0020_),
    .Y(_0180_));
 sky130_fd_sc_hd__buf_4 _1103_ (.A(_0180_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2i_1 _1104_ (.A0(_0174_),
    .A1(_0179_),
    .S(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__mux2_2 _1105_ (.A0(net19),
    .A1(net21),
    .S(_0724_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _1106_ (.A0(net20),
    .A1(_0055_),
    .S(_0724_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2i_4 _1107_ (.A0(_0183_),
    .A1(_0184_),
    .S(_0124_),
    .Y(_0185_));
 sky130_fd_sc_hd__nand2_2 _1108_ (.A(_0063_),
    .B(_0921_),
    .Y(_0186_));
 sky130_fd_sc_hd__mux2i_4 _1109_ (.A0(_0059_),
    .A1(_0056_),
    .S(_0775_),
    .Y(_0187_));
 sky130_fd_sc_hd__o22ai_4 _1110_ (.A1(_0064_),
    .A2(_0185_),
    .B1(_0186_),
    .B2(_0187_),
    .Y(_0188_));
 sky130_fd_sc_hd__nor2_4 _1111_ (.A(_0034_),
    .B(_0020_),
    .Y(_0189_));
 sky130_fd_sc_hd__a22oi_1 _1112_ (.A1(_0170_),
    .A2(_0182_),
    .B1(_0188_),
    .B2(_0189_),
    .Y(_0190_));
 sky130_fd_sc_hd__clkbuf_4 _1113_ (.A(_0110_),
    .X(_0191_));
 sky130_fd_sc_hd__nor2_2 _1114_ (.A(_0879_),
    .B(_0126_),
    .Y(_0192_));
 sky130_fd_sc_hd__buf_4 _1115_ (.A(_0192_),
    .X(_0193_));
 sky130_fd_sc_hd__clkbuf_4 _1116_ (.A(_0193_),
    .X(_0194_));
 sky130_fd_sc_hd__buf_6 _1117_ (.A(_0785_),
    .X(_0195_));
 sky130_fd_sc_hd__buf_6 _1118_ (.A(_0806_),
    .X(_0196_));
 sky130_fd_sc_hd__mux2i_4 _1119_ (.A0(_0080_),
    .A1(_0089_),
    .S(_0196_),
    .Y(_0197_));
 sky130_fd_sc_hd__mux2i_4 _1120_ (.A0(_0115_),
    .A1(_0082_),
    .S(_0196_),
    .Y(_0198_));
 sky130_fd_sc_hd__mux2i_4 _1121_ (.A0(_0197_),
    .A1(_0198_),
    .S(_0158_),
    .Y(_0199_));
 sky130_fd_sc_hd__mux2i_4 _1122_ (.A0(net28),
    .A1(net26),
    .S(_0806_),
    .Y(_0200_));
 sky130_fd_sc_hd__mux2_1 _1123_ (.A0(_0118_),
    .A1(_0117_),
    .S(_0196_),
    .X(_0201_));
 sky130_fd_sc_hd__nor2_1 _1124_ (.A(_0112_),
    .B(_0201_),
    .Y(_0202_));
 sky130_fd_sc_hd__a211oi_1 _1125_ (.A1(_0143_),
    .A2(_0200_),
    .B1(_0202_),
    .C1(_0195_),
    .Y(_0203_));
 sky130_fd_sc_hd__a21oi_2 _1126_ (.A1(_0195_),
    .A2(_0199_),
    .B1(_0203_),
    .Y(_0204_));
 sky130_fd_sc_hd__nand2_2 _1127_ (.A(net12),
    .B(_0124_),
    .Y(_0205_));
 sky130_fd_sc_hd__mux2i_4 _1128_ (.A0(net23),
    .A1(net1),
    .S(_0806_),
    .Y(_0206_));
 sky130_fd_sc_hd__buf_6 _1129_ (.A(_0765_),
    .X(_0207_));
 sky130_fd_sc_hd__buf_6 _1130_ (.A(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__o22ai_4 _1131_ (.A1(_0837_),
    .A2(_0205_),
    .B1(_0206_),
    .B2(_0208_),
    .Y(_0209_));
 sky130_fd_sc_hd__nor3_2 _1132_ (.A(_0879_),
    .B(_0126_),
    .C(_0112_),
    .Y(_0210_));
 sky130_fd_sc_hd__nand2_1 _1133_ (.A(_0209_),
    .B(_0210_),
    .Y(_0211_));
 sky130_fd_sc_hd__o21ai_1 _1134_ (.A1(_0194_),
    .A2(_0204_),
    .B1(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__clkbuf_4 _1135_ (.A(_0041_),
    .X(_0213_));
 sky130_fd_sc_hd__a21oi_1 _1136_ (.A1(_0191_),
    .A2(_0212_),
    .B1(_0213_),
    .Y(_0214_));
 sky130_fd_sc_hd__clkbuf_4 _1137_ (.A(_0033_),
    .X(_0215_));
 sky130_fd_sc_hd__clkbuf_4 _1138_ (.A(_0108_),
    .X(_0216_));
 sky130_fd_sc_hd__buf_4 _1139_ (.A(_0196_),
    .X(_0217_));
 sky130_fd_sc_hd__mux4_2 _1140_ (.A0(net10),
    .A1(net11),
    .A2(net13),
    .A3(_0172_),
    .S0(_0096_),
    .S1(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__mux4_1 _1141_ (.A0(_0118_),
    .A1(_0099_),
    .A2(_0135_),
    .A3(_0093_),
    .S0(_0083_),
    .S1(_0837_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2i_1 _1142_ (.A0(_0218_),
    .A1(_0219_),
    .S(_0129_),
    .Y(_0220_));
 sky130_fd_sc_hd__clkbuf_4 _1143_ (.A(_0112_),
    .X(_0221_));
 sky130_fd_sc_hd__mux4_1 _1144_ (.A0(_0051_),
    .A1(_0048_),
    .A2(_0058_),
    .A3(_0055_),
    .S0(_0096_),
    .S1(_0133_),
    .X(_0222_));
 sky130_fd_sc_hd__o21ai_0 _1145_ (.A1(_0847_),
    .A2(_0187_),
    .B1(_0221_),
    .Y(_0223_));
 sky130_fd_sc_hd__o21ai_1 _1146_ (.A1(_0221_),
    .A2(_0222_),
    .B1(_0223_),
    .Y(_0224_));
 sky130_fd_sc_hd__nand2_1 _1147_ (.A(_0108_),
    .B(_0131_),
    .Y(_0225_));
 sky130_fd_sc_hd__o32ai_1 _1148_ (.A1(_0216_),
    .A2(_0144_),
    .A3(_0220_),
    .B1(_0224_),
    .B2(_0225_),
    .Y(_0226_));
 sky130_fd_sc_hd__mux2i_1 _1149_ (.A0(_0080_),
    .A1(_0089_),
    .S(_0734_),
    .Y(_0227_));
 sky130_fd_sc_hd__mux2i_1 _1150_ (.A0(_0081_),
    .A1(_0079_),
    .S(_0745_),
    .Y(_0228_));
 sky130_fd_sc_hd__mux2i_2 _1151_ (.A0(_0227_),
    .A1(_0228_),
    .S(_0704_),
    .Y(_0229_));
 sky130_fd_sc_hd__mux4_1 _1152_ (.A0(net2),
    .A1(net31),
    .A2(net30),
    .A3(net29),
    .S0(_0096_),
    .S1(_0097_),
    .X(_0230_));
 sky130_fd_sc_hd__clkbuf_4 _1153_ (.A(_0101_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2i_1 _1154_ (.A0(_0229_),
    .A1(_0230_),
    .S(_0231_),
    .Y(_0232_));
 sky130_fd_sc_hd__mux2i_2 _1155_ (.A0(_0088_),
    .A1(net1),
    .S(_0734_),
    .Y(_0233_));
 sky130_fd_sc_hd__o22a_1 _1156_ (.A1(_0195_),
    .A2(_0233_),
    .B1(_0205_),
    .B2(_0090_),
    .X(_0234_));
 sky130_fd_sc_hd__nand2b_2 _1157_ (.A_N(_0899_),
    .B(_0868_),
    .Y(_0235_));
 sky130_fd_sc_hd__o22ai_1 _1158_ (.A1(_0066_),
    .A2(_0232_),
    .B1(_0234_),
    .B2(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__buf_4 _1159_ (.A(_0158_),
    .X(_0237_));
 sky130_fd_sc_hd__clkbuf_4 _1160_ (.A(_0237_),
    .X(_0238_));
 sky130_fd_sc_hd__buf_2 _1161_ (.A(net16),
    .X(_0239_));
 sky130_fd_sc_hd__mux4_2 _1162_ (.A0(net15),
    .A1(_0239_),
    .A2(_0050_),
    .A3(_0047_),
    .S0(_0683_),
    .S1(_0133_),
    .X(_0240_));
 sky130_fd_sc_hd__nor2_1 _1163_ (.A(_0132_),
    .B(_0240_),
    .Y(_0241_));
 sky130_fd_sc_hd__mux4_2 _1164_ (.A0(_0094_),
    .A1(_0095_),
    .A2(_0068_),
    .A3(_0069_),
    .S0(_0072_),
    .S1(_0217_),
    .X(_0242_));
 sky130_fd_sc_hd__nor2_1 _1165_ (.A(_0194_),
    .B(_0242_),
    .Y(_0243_));
 sky130_fd_sc_hd__o41ai_1 _1166_ (.A1(_0037_),
    .A2(_0238_),
    .A3(_0241_),
    .A4(_0243_),
    .B1(_0167_),
    .Y(_0244_));
 sky130_fd_sc_hd__a221oi_1 _1167_ (.A1(_0215_),
    .A2(_0226_),
    .B1(_0236_),
    .B2(_0170_),
    .C1(_0244_),
    .Y(_0245_));
 sky130_fd_sc_hd__a21oi_1 _1168_ (.A1(_0190_),
    .A2(_0214_),
    .B1(_0245_),
    .Y(net37));
 sky130_fd_sc_hd__clkbuf_4 _1169_ (.A(_0131_),
    .X(_0246_));
 sky130_fd_sc_hd__mux4_2 _1170_ (.A0(net7),
    .A1(net8),
    .A2(net9),
    .A3(net10),
    .S0(_0683_),
    .S1(_0133_),
    .X(_0247_));
 sky130_fd_sc_hd__mux4_1 _1171_ (.A0(_0099_),
    .A1(_0135_),
    .A2(_0093_),
    .A3(_0094_),
    .S0(_0775_),
    .S1(_0138_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2i_4 _1172_ (.A0(_0247_),
    .A1(_0248_),
    .S(_0237_),
    .Y(_0249_));
 sky130_fd_sc_hd__nor2b_2 _1173_ (.A(_0672_),
    .B_N(_0056_),
    .Y(_0250_));
 sky130_fd_sc_hd__nand2b_1 _1174_ (.A_N(_0826_),
    .B(_0250_),
    .Y(_0251_));
 sky130_fd_sc_hd__mux4_1 _1175_ (.A0(net20),
    .A1(net21),
    .A2(net22),
    .A3(_0059_),
    .S0(_0683_),
    .S1(_0826_),
    .X(_0252_));
 sky130_fd_sc_hd__nor2_1 _1176_ (.A(_0221_),
    .B(_0252_),
    .Y(_0253_));
 sky130_fd_sc_hd__a21oi_2 _1177_ (.A1(_0113_),
    .A2(_0251_),
    .B1(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hd__nand2_1 _1178_ (.A(_0216_),
    .B(_0254_),
    .Y(_0255_));
 sky130_fd_sc_hd__o21ai_0 _1179_ (.A1(_0216_),
    .A2(_0249_),
    .B1(_0255_),
    .Y(_0256_));
 sky130_fd_sc_hd__buf_4 _1180_ (.A(_0031_),
    .X(_0257_));
 sky130_fd_sc_hd__clkbuf_4 _1181_ (.A(_0020_),
    .X(_0258_));
 sky130_fd_sc_hd__mux4_2 _1182_ (.A0(_0082_),
    .A1(_0081_),
    .A2(_0080_),
    .A3(_0079_),
    .S0(_0123_),
    .S1(_0084_),
    .X(_0259_));
 sky130_fd_sc_hd__mux4_2 _1183_ (.A0(_0099_),
    .A1(_0118_),
    .A2(_0115_),
    .A3(_0117_),
    .S0(_0123_),
    .S1(_0084_),
    .X(_0260_));
 sky130_fd_sc_hd__mux2i_4 _1184_ (.A0(_0259_),
    .A1(_0260_),
    .S(_0177_),
    .Y(_0261_));
 sky130_fd_sc_hd__mux2i_1 _1185_ (.A0(_0089_),
    .A1(net12),
    .S(_0734_),
    .Y(_0262_));
 sky130_fd_sc_hd__mux2_4 _1186_ (.A0(_0233_),
    .A1(_0262_),
    .S(_0053_),
    .X(_0263_));
 sky130_fd_sc_hd__o22a_1 _1187_ (.A1(_0258_),
    .A2(_0261_),
    .B1(_0263_),
    .B2(_0235_),
    .X(_0264_));
 sky130_fd_sc_hd__clkbuf_4 _1188_ (.A(_0193_),
    .X(_0265_));
 sky130_fd_sc_hd__nand2_1 _1189_ (.A(_0110_),
    .B(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__mux4_2 _1190_ (.A0(_0239_),
    .A1(net17),
    .A2(net18),
    .A3(net19),
    .S0(_0683_),
    .S1(_0826_),
    .X(_0267_));
 sky130_fd_sc_hd__mux4_2 _1191_ (.A0(net11),
    .A1(net13),
    .A2(net14),
    .A3(net15),
    .S0(_0683_),
    .S1(_0826_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2i_4 _1192_ (.A0(_0267_),
    .A1(_0268_),
    .S(_0237_),
    .Y(_0269_));
 sky130_fd_sc_hd__o221ai_1 _1193_ (.A1(_0257_),
    .A2(_0264_),
    .B1(_0266_),
    .B2(_0269_),
    .C1(_0167_),
    .Y(_0270_));
 sky130_fd_sc_hd__a31oi_1 _1194_ (.A1(_0215_),
    .A2(_0246_),
    .A3(_0256_),
    .B1(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__buf_4 _1195_ (.A(_0131_),
    .X(_0272_));
 sky130_fd_sc_hd__mux2i_2 _1196_ (.A0(net25),
    .A1(net12),
    .S(_0806_),
    .Y(_0273_));
 sky130_fd_sc_hd__nor2_1 _1197_ (.A(_0785_),
    .B(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__nor2_1 _1198_ (.A(_0120_),
    .B(_0206_),
    .Y(_0275_));
 sky130_fd_sc_hd__nor2_2 _1199_ (.A(_0274_),
    .B(_0275_),
    .Y(_0276_));
 sky130_fd_sc_hd__mux2i_4 _1200_ (.A0(net29),
    .A1(net27),
    .S(_0806_),
    .Y(_0277_));
 sky130_fd_sc_hd__mux2i_2 _1201_ (.A0(_0200_),
    .A1(_0277_),
    .S(_0920_),
    .Y(_0278_));
 sky130_fd_sc_hd__mux2_1 _1202_ (.A0(_0099_),
    .A1(_0115_),
    .S(_0196_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2i_4 _1203_ (.A0(_0201_),
    .A1(_0279_),
    .S(_0704_),
    .Y(_0280_));
 sky130_fd_sc_hd__nand2_1 _1204_ (.A(_0238_),
    .B(_0280_),
    .Y(_0281_));
 sky130_fd_sc_hd__o211ai_1 _1205_ (.A1(_0238_),
    .A2(_0278_),
    .B1(_0281_),
    .C1(_0272_),
    .Y(_0282_));
 sky130_fd_sc_hd__o31ai_2 _1206_ (.A1(_0272_),
    .A2(_0144_),
    .A3(_0276_),
    .B1(_0282_),
    .Y(_0283_));
 sky130_fd_sc_hd__mux4_1 _1207_ (.A0(_0239_),
    .A1(_0050_),
    .A2(_0047_),
    .A3(_0051_),
    .S0(_0765_),
    .S1(_0097_),
    .X(_0284_));
 sky130_fd_sc_hd__nor2_1 _1208_ (.A(_0075_),
    .B(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__clkbuf_4 _1209_ (.A(_0734_),
    .X(_0286_));
 sky130_fd_sc_hd__mux4_1 _1210_ (.A0(_0071_),
    .A1(_0150_),
    .A2(_0172_),
    .A3(_0151_),
    .S0(_0083_),
    .S1(_0286_),
    .X(_0287_));
 sky130_fd_sc_hd__nor2_1 _1211_ (.A(_0064_),
    .B(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__nor2_2 _1212_ (.A(_0285_),
    .B(_0288_),
    .Y(_0289_));
 sky130_fd_sc_hd__mux4_2 _1213_ (.A0(_0095_),
    .A1(_0068_),
    .A2(_0069_),
    .A3(_0070_),
    .S0(_0207_),
    .S1(_0090_),
    .X(_0290_));
 sky130_fd_sc_hd__mux4_2 _1214_ (.A0(_0099_),
    .A1(_0135_),
    .A2(_0093_),
    .A3(_0094_),
    .S0(_0207_),
    .S1(_0286_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2i_2 _1215_ (.A0(_0290_),
    .A1(_0291_),
    .S(_0075_),
    .Y(_0292_));
 sky130_fd_sc_hd__nor2_1 _1216_ (.A(_0066_),
    .B(_0292_),
    .Y(_0293_));
 sky130_fd_sc_hd__a21oi_1 _1217_ (.A1(_0046_),
    .A2(_0289_),
    .B1(_0293_),
    .Y(_0294_));
 sky130_fd_sc_hd__buf_4 _1218_ (.A(_0208_),
    .X(_0295_));
 sky130_fd_sc_hd__inv_1 _1219_ (.A(_0056_),
    .Y(_0296_));
 sky130_fd_sc_hd__o2bb2ai_1 _1220_ (.A1_N(_0101_),
    .A2_N(_0184_),
    .B1(_0186_),
    .B2(_0296_),
    .Y(_0297_));
 sky130_fd_sc_hd__clkbuf_4 _1221_ (.A(_0063_),
    .X(_0298_));
 sky130_fd_sc_hd__o21ai_1 _1222_ (.A1(_0298_),
    .A2(_0061_),
    .B1(_0295_),
    .Y(_0299_));
 sky130_fd_sc_hd__o21ai_4 _1223_ (.A1(_0295_),
    .A2(_0297_),
    .B1(_0299_),
    .Y(_0300_));
 sky130_fd_sc_hd__nand2_4 _1224_ (.A(_0031_),
    .B(_0180_),
    .Y(_0301_));
 sky130_fd_sc_hd__o22ai_2 _1225_ (.A1(_0257_),
    .A2(_0294_),
    .B1(_0300_),
    .B2(_0301_),
    .Y(_0302_));
 sky130_fd_sc_hd__a211oi_1 _1226_ (.A1(_0191_),
    .A2(_0283_),
    .B1(_0302_),
    .C1(_0213_),
    .Y(_0303_));
 sky130_fd_sc_hd__nor2_1 _1227_ (.A(_0271_),
    .B(_0303_),
    .Y(net38));
 sky130_fd_sc_hd__nor2_1 _1228_ (.A(_0053_),
    .B(_0273_),
    .Y(_0304_));
 sky130_fd_sc_hd__mux2i_4 _1229_ (.A0(_0079_),
    .A1(_0088_),
    .S(_0196_),
    .Y(_0305_));
 sky130_fd_sc_hd__nor2_1 _1230_ (.A(_0124_),
    .B(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__o21ai_4 _1231_ (.A1(_0304_),
    .A2(_0306_),
    .B1(_0158_),
    .Y(_0307_));
 sky130_fd_sc_hd__mux2i_1 _1232_ (.A0(_0099_),
    .A1(_0115_),
    .S(_0826_),
    .Y(_0308_));
 sky130_fd_sc_hd__mux2i_1 _1233_ (.A0(_0277_),
    .A1(_0308_),
    .S(_0158_),
    .Y(_0309_));
 sky130_fd_sc_hd__mux2i_4 _1234_ (.A0(_0117_),
    .A1(net28),
    .S(_0196_),
    .Y(_0310_));
 sky130_fd_sc_hd__mux2i_4 _1235_ (.A0(net4),
    .A1(_0118_),
    .S(_0816_),
    .Y(_0311_));
 sky130_fd_sc_hd__mux2i_1 _1236_ (.A0(_0310_),
    .A1(_0311_),
    .S(_0158_),
    .Y(_0312_));
 sky130_fd_sc_hd__mux2_2 _1237_ (.A0(_0309_),
    .A1(_0312_),
    .S(_0053_),
    .X(_0313_));
 sky130_fd_sc_hd__nand2_1 _1238_ (.A(_0132_),
    .B(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__nor2_4 _1239_ (.A(_0217_),
    .B(_0166_),
    .Y(_0315_));
 sky130_fd_sc_hd__nor2_4 _1240_ (.A(_0063_),
    .B(_0745_),
    .Y(_0316_));
 sky130_fd_sc_hd__xnor2_2 _1241_ (.A(_0020_),
    .B(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__nand3_1 _1242_ (.A(_0113_),
    .B(_0315_),
    .C(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__o211ai_2 _1243_ (.A1(_0132_),
    .A2(_0307_),
    .B1(_0314_),
    .C1(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__clkbuf_4 _1244_ (.A(_0298_),
    .X(_0320_));
 sky130_fd_sc_hd__nor3_1 _1245_ (.A(_0320_),
    .B(_0062_),
    .C(_0301_),
    .Y(_0321_));
 sky130_fd_sc_hd__nor2_1 _1246_ (.A(_0063_),
    .B(_0067_),
    .Y(_0322_));
 sky130_fd_sc_hd__a21o_1 _1247_ (.A1(_0298_),
    .A2(_0054_),
    .B1(_0322_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2i_4 _1248_ (.A0(_0073_),
    .A1(_0098_),
    .S(_0101_),
    .Y(_0324_));
 sky130_fd_sc_hd__mux2_1 _1249_ (.A0(_0323_),
    .A1(_0324_),
    .S(_0180_),
    .X(_0325_));
 sky130_fd_sc_hd__nor2_1 _1250_ (.A(_0043_),
    .B(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__clkbuf_4 _1251_ (.A(_0041_),
    .X(_0327_));
 sky130_fd_sc_hd__a2111oi_1 _1252_ (.A1(_0111_),
    .A2(_0319_),
    .B1(_0321_),
    .C1(_0326_),
    .D1(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hd__clkbuf_4 _1253_ (.A(_0237_),
    .X(_0329_));
 sky130_fd_sc_hd__nor2_1 _1254_ (.A(_0329_),
    .B(_0162_),
    .Y(_0330_));
 sky130_fd_sc_hd__nor2_1 _1255_ (.A(_0114_),
    .B(_0153_),
    .Y(_0331_));
 sky130_fd_sc_hd__nor2_4 _1256_ (.A(_0108_),
    .B(_0128_),
    .Y(_0332_));
 sky130_fd_sc_hd__o21ai_0 _1257_ (.A1(_0330_),
    .A2(_0331_),
    .B1(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__a21oi_1 _1258_ (.A1(_0114_),
    .A2(_0156_),
    .B1(_0265_),
    .Y(_0334_));
 sky130_fd_sc_hd__nand2_1 _1259_ (.A(_0036_),
    .B(_0137_),
    .Y(_0335_));
 sky130_fd_sc_hd__nand3_1 _1260_ (.A(_0216_),
    .B(_0132_),
    .C(_0161_),
    .Y(_0336_));
 sky130_fd_sc_hd__a21oi_1 _1261_ (.A1(_0335_),
    .A2(_0336_),
    .B1(_0144_),
    .Y(_0337_));
 sky130_fd_sc_hd__o21bai_1 _1262_ (.A1(_0216_),
    .A2(_0334_),
    .B1_N(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__mux4_4 _1263_ (.A0(net26),
    .A1(net25),
    .A2(_0088_),
    .A3(net12),
    .S0(_0096_),
    .S1(_0745_),
    .X(_0339_));
 sky130_fd_sc_hd__a2bb2oi_2 _1264_ (.A1_N(_0166_),
    .A2_N(_0186_),
    .B1(_0339_),
    .B2(_0177_),
    .Y(_0340_));
 sky130_fd_sc_hd__mux4_4 _1265_ (.A0(_0117_),
    .A1(_0082_),
    .A2(_0081_),
    .A3(_0080_),
    .S0(_0072_),
    .S1(_0084_),
    .X(_0341_));
 sky130_fd_sc_hd__mux4_2 _1266_ (.A0(_0135_),
    .A1(_0099_),
    .A2(_0118_),
    .A3(_0115_),
    .S0(_0072_),
    .S1(_0745_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2i_4 _1267_ (.A0(_0341_),
    .A1(_0342_),
    .S(_0177_),
    .Y(_0343_));
 sky130_fd_sc_hd__mux2_1 _1268_ (.A0(_0340_),
    .A1(_0343_),
    .S(_0180_),
    .X(_0344_));
 sky130_fd_sc_hd__o21ai_1 _1269_ (.A1(_0044_),
    .A2(_0344_),
    .B1(_0327_),
    .Y(_0345_));
 sky130_fd_sc_hd__a31oi_1 _1270_ (.A1(_0215_),
    .A2(_0333_),
    .A3(_0338_),
    .B1(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__nor2_1 _1271_ (.A(_0328_),
    .B(_0346_),
    .Y(net39));
 sky130_fd_sc_hd__mux2i_1 _1272_ (.A0(net15),
    .A1(net17),
    .S(_0816_),
    .Y(_0347_));
 sky130_fd_sc_hd__mux2_2 _1273_ (.A0(_0149_),
    .A1(_0347_),
    .S(_0072_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _1274_ (.A0(net18),
    .A1(net20),
    .S(_0806_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _1275_ (.A0(net19),
    .A1(net21),
    .S(_0806_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2i_1 _1276_ (.A0(_0349_),
    .A1(_0350_),
    .S(_0785_),
    .Y(_0351_));
 sky130_fd_sc_hd__mux2_1 _1277_ (.A0(_0348_),
    .A1(_0351_),
    .S(_0112_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2i_1 _1278_ (.A0(_0094_),
    .A1(_0068_),
    .S(_0133_),
    .Y(_0353_));
 sky130_fd_sc_hd__mux2_2 _1279_ (.A0(_0134_),
    .A1(_0353_),
    .S(_0208_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _1280_ (.A0(net22),
    .A1(_0056_),
    .S(_0806_),
    .X(_0355_));
 sky130_fd_sc_hd__nor2b_1 _1281_ (.A(_0806_),
    .B_N(net24),
    .Y(_0356_));
 sky130_fd_sc_hd__mux2i_4 _1282_ (.A0(_0355_),
    .A1(_0356_),
    .S(_0208_),
    .Y(_0357_));
 sky130_fd_sc_hd__o22ai_1 _1283_ (.A1(_0216_),
    .A2(_0354_),
    .B1(_0357_),
    .B2(_0225_),
    .Y(_0358_));
 sky130_fd_sc_hd__mux2i_1 _1284_ (.A0(net10),
    .A1(net13),
    .S(_0816_),
    .Y(_0359_));
 sky130_fd_sc_hd__mux2_2 _1285_ (.A0(_0154_),
    .A1(_0359_),
    .S(_0096_),
    .X(_0360_));
 sky130_fd_sc_hd__o21ai_0 _1286_ (.A1(_0237_),
    .A2(_0360_),
    .B1(_0129_),
    .Y(_0361_));
 sky130_fd_sc_hd__clkbuf_4 _1287_ (.A(_0036_),
    .X(_0362_));
 sky130_fd_sc_hd__a22oi_1 _1288_ (.A1(_0238_),
    .A2(_0358_),
    .B1(_0361_),
    .B2(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__a211o_1 _1289_ (.A1(_0332_),
    .A2(_0352_),
    .B1(_0363_),
    .C1(_0107_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2i_4 _1290_ (.A0(net12),
    .A1(net1),
    .S(_0123_),
    .Y(_0365_));
 sky130_fd_sc_hd__mux2i_1 _1291_ (.A0(_0079_),
    .A1(_0088_),
    .S(_0060_),
    .Y(_0366_));
 sky130_fd_sc_hd__mux2_1 _1292_ (.A0(_0227_),
    .A1(_0366_),
    .S(_0124_),
    .X(_0367_));
 sky130_fd_sc_hd__o22a_2 _1293_ (.A1(_0186_),
    .A2(_0365_),
    .B1(_0367_),
    .B2(_0064_),
    .X(_0368_));
 sky130_fd_sc_hd__mux4_2 _1294_ (.A0(_0115_),
    .A1(_0117_),
    .A2(_0082_),
    .A3(_0081_),
    .S0(_0083_),
    .S1(_0286_),
    .X(_0369_));
 sky130_fd_sc_hd__mux4_4 _1295_ (.A0(_0093_),
    .A1(_0135_),
    .A2(_0099_),
    .A3(_0118_),
    .S0(_0207_),
    .S1(_0286_),
    .X(_0370_));
 sky130_fd_sc_hd__mux2i_4 _1296_ (.A0(_0369_),
    .A1(_0370_),
    .S(_0075_),
    .Y(_0371_));
 sky130_fd_sc_hd__mux2i_2 _1297_ (.A0(_0368_),
    .A1(_0371_),
    .S(_0181_),
    .Y(_0372_));
 sky130_fd_sc_hd__nand2_1 _1298_ (.A(_0170_),
    .B(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__mux2i_1 _1299_ (.A0(_0198_),
    .A1(_0310_),
    .S(_0208_),
    .Y(_0374_));
 sky130_fd_sc_hd__mux2i_4 _1300_ (.A0(_0093_),
    .A1(net3),
    .S(_0816_),
    .Y(_0375_));
 sky130_fd_sc_hd__mux2i_1 _1301_ (.A0(_0311_),
    .A1(_0375_),
    .S(_0704_),
    .Y(_0376_));
 sky130_fd_sc_hd__mux2_2 _1302_ (.A0(_0374_),
    .A1(_0376_),
    .S(_0159_),
    .X(_0377_));
 sky130_fd_sc_hd__mux2i_2 _1303_ (.A0(_0197_),
    .A1(_0305_),
    .S(_0785_),
    .Y(_0378_));
 sky130_fd_sc_hd__o21ai_1 _1304_ (.A1(_0138_),
    .A2(_0365_),
    .B1(_0143_),
    .Y(_0379_));
 sky130_fd_sc_hd__o211ai_1 _1305_ (.A1(_0221_),
    .A2(_0378_),
    .B1(_0379_),
    .C1(_0193_),
    .Y(_0380_));
 sky130_fd_sc_hd__a21boi_2 _1306_ (.A1(_0132_),
    .A2(_0377_),
    .B1_N(_0380_),
    .Y(_0381_));
 sky130_fd_sc_hd__mux2i_4 _1307_ (.A0(_0049_),
    .A1(_0183_),
    .S(_0208_),
    .Y(_0382_));
 sky130_fd_sc_hd__mux4_2 _1308_ (.A0(_0172_),
    .A1(_0151_),
    .A2(_0239_),
    .A3(_0050_),
    .S0(_0123_),
    .S1(_0084_),
    .X(_0383_));
 sky130_fd_sc_hd__nor2_1 _1309_ (.A(_0064_),
    .B(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__a21oi_1 _1310_ (.A1(_0087_),
    .A2(_0382_),
    .B1(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__mux4_4 _1311_ (.A0(_0069_),
    .A1(_0070_),
    .A2(_0071_),
    .A3(_0150_),
    .S0(_0123_),
    .S1(_0084_),
    .X(_0386_));
 sky130_fd_sc_hd__mux4_2 _1312_ (.A0(_0093_),
    .A1(net6),
    .A2(net7),
    .A3(_0068_),
    .S0(_0765_),
    .S1(_0097_),
    .X(_0387_));
 sky130_fd_sc_hd__mux2i_4 _1313_ (.A0(_0386_),
    .A1(_0387_),
    .S(_0177_),
    .Y(_0388_));
 sky130_fd_sc_hd__nor2_1 _1314_ (.A(_0066_),
    .B(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__a21oi_1 _1315_ (.A1(_0046_),
    .A2(_0385_),
    .B1(_0389_),
    .Y(_0390_));
 sky130_fd_sc_hd__clkbuf_4 _1316_ (.A(_0181_),
    .X(_0391_));
 sky130_fd_sc_hd__nand3b_1 _1317_ (.A_N(_0097_),
    .B(_0059_),
    .C(_0124_),
    .Y(_0392_));
 sky130_fd_sc_hd__o21ai_4 _1318_ (.A1(_0124_),
    .A2(_0057_),
    .B1(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__nand4_1 _1319_ (.A(_0257_),
    .B(_0391_),
    .C(_0178_),
    .D(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__o221ai_1 _1320_ (.A1(_0038_),
    .A2(_0381_),
    .B1(_0390_),
    .B2(_0044_),
    .C1(_0394_),
    .Y(_0395_));
 sky130_fd_sc_hd__nor2_1 _1321_ (.A(_0213_),
    .B(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__a31oi_2 _1322_ (.A1(_0213_),
    .A2(_0364_),
    .A3(_0373_),
    .B1(_0396_),
    .Y(net40));
 sky130_fd_sc_hd__nor2_1 _1323_ (.A(_0704_),
    .B(_0198_),
    .Y(_0397_));
 sky130_fd_sc_hd__a21oi_1 _1324_ (.A1(_0120_),
    .A2(_0201_),
    .B1(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__inv_1 _1325_ (.A(_0858_),
    .Y(_0399_));
 sky130_fd_sc_hd__or2_0 _1326_ (.A(_0899_),
    .B(_0858_),
    .X(_0400_));
 sky130_fd_sc_hd__nand2_1 _1327_ (.A(_0899_),
    .B(_0858_),
    .Y(_0401_));
 sky130_fd_sc_hd__o21ai_0 _1328_ (.A1(_0889_),
    .A2(_0400_),
    .B1(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__a22o_2 _1329_ (.A1(_0399_),
    .A2(_0879_),
    .B1(_0402_),
    .B2(_0868_),
    .X(_0403_));
 sky130_fd_sc_hd__and2_1 _1330_ (.A(_0398_),
    .B(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__mux2i_2 _1331_ (.A0(_0200_),
    .A1(_0197_),
    .S(_0208_),
    .Y(_0405_));
 sky130_fd_sc_hd__mux2i_4 _1332_ (.A0(_0209_),
    .A1(_0405_),
    .S(_0159_),
    .Y(_0406_));
 sky130_fd_sc_hd__mux2i_4 _1333_ (.A0(_0094_),
    .A1(_0135_),
    .S(_0826_),
    .Y(_0407_));
 sky130_fd_sc_hd__mux2i_4 _1334_ (.A0(_0375_),
    .A1(_0407_),
    .S(_0704_),
    .Y(_0408_));
 sky130_fd_sc_hd__o2bb2ai_2 _1335_ (.A1_N(_0193_),
    .A2_N(_0406_),
    .B1(_0408_),
    .B2(_0030_),
    .Y(_0409_));
 sky130_fd_sc_hd__nor2_1 _1336_ (.A(_0404_),
    .B(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__nand2_1 _1337_ (.A(_0111_),
    .B(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__mux2_1 _1338_ (.A0(_0059_),
    .A1(_0056_),
    .S(_0785_),
    .X(_0412_));
 sky130_fd_sc_hd__nor3_2 _1339_ (.A(_0298_),
    .B(_0090_),
    .C(_0301_),
    .Y(_0413_));
 sky130_fd_sc_hd__a21oi_1 _1340_ (.A1(_0412_),
    .A2(_0413_),
    .B1(_0040_),
    .Y(_0414_));
 sky130_fd_sc_hd__buf_2 _1341_ (.A(_0258_),
    .X(_0415_));
 sky130_fd_sc_hd__nor2_1 _1342_ (.A(_0178_),
    .B(_0173_),
    .Y(_0416_));
 sky130_fd_sc_hd__nor2_1 _1343_ (.A(_0320_),
    .B(_0175_),
    .Y(_0417_));
 sky130_fd_sc_hd__nor2_1 _1344_ (.A(_0416_),
    .B(_0417_),
    .Y(_0418_));
 sky130_fd_sc_hd__nand2_1 _1345_ (.A(_0298_),
    .B(_0185_),
    .Y(_0419_));
 sky130_fd_sc_hd__o21ai_1 _1346_ (.A1(_0063_),
    .A2(_0171_),
    .B1(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__nand2_1 _1347_ (.A(_0415_),
    .B(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__o21ai_0 _1348_ (.A1(_0415_),
    .A2(_0418_),
    .B1(_0421_),
    .Y(_0422_));
 sky130_fd_sc_hd__nor2_2 _1349_ (.A(_0108_),
    .B(_0192_),
    .Y(_0423_));
 sky130_fd_sc_hd__mux2i_2 _1350_ (.A0(_0218_),
    .A1(_0242_),
    .S(_0159_),
    .Y(_0424_));
 sky130_fd_sc_hd__nand2_1 _1351_ (.A(_0423_),
    .B(_0424_),
    .Y(_0425_));
 sky130_fd_sc_hd__mux2i_1 _1352_ (.A0(_0222_),
    .A1(_0240_),
    .S(_0159_),
    .Y(_0426_));
 sky130_fd_sc_hd__nor2_1 _1353_ (.A(_0138_),
    .B(_0187_),
    .Y(_0427_));
 sky130_fd_sc_hd__o21ai_0 _1354_ (.A1(_0207_),
    .A2(_0734_),
    .B1(_0858_),
    .Y(_0428_));
 sky130_fd_sc_hd__nand3b_1 _1355_ (.A_N(_0858_),
    .B(_0063_),
    .C(_0868_),
    .Y(_0429_));
 sky130_fd_sc_hd__or3b_1 _1356_ (.A(_0765_),
    .B(_0724_),
    .C_N(_0031_),
    .X(_0430_));
 sky130_fd_sc_hd__o211ai_2 _1357_ (.A1(_0235_),
    .A2(_0428_),
    .B1(_0429_),
    .C1(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__a21oi_1 _1358_ (.A1(_0427_),
    .A2(_0431_),
    .B1(_0036_),
    .Y(_0432_));
 sky130_fd_sc_hd__a21oi_1 _1359_ (.A1(_0332_),
    .A2(_0426_),
    .B1(_0432_),
    .Y(_0433_));
 sky130_fd_sc_hd__clkinv_2 _1360_ (.A(_0040_),
    .Y(_0434_));
 sky130_fd_sc_hd__a31o_1 _1361_ (.A1(_0215_),
    .A2(_0425_),
    .A3(_0433_),
    .B1(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__o31ai_1 _1362_ (.A1(_0037_),
    .A2(_0404_),
    .A3(_0409_),
    .B1(_0414_),
    .Y(_0436_));
 sky130_fd_sc_hd__a21oi_1 _1363_ (.A1(_0435_),
    .A2(_0436_),
    .B1(_0170_),
    .Y(_0437_));
 sky130_fd_sc_hd__o22ai_2 _1364_ (.A1(_0785_),
    .A2(_0233_),
    .B1(_0205_),
    .B2(_0090_),
    .Y(_0438_));
 sky130_fd_sc_hd__mux2i_2 _1365_ (.A0(_0229_),
    .A1(_0438_),
    .S(_0298_),
    .Y(_0439_));
 sky130_fd_sc_hd__nor2_1 _1366_ (.A(_0391_),
    .B(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__mux4_2 _1367_ (.A0(net6),
    .A1(net5),
    .A2(net4),
    .A3(net3),
    .S0(_0765_),
    .S1(_0060_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2i_2 _1368_ (.A0(_0230_),
    .A1(_0441_),
    .S(_0101_),
    .Y(_0442_));
 sky130_fd_sc_hd__nor2_1 _1369_ (.A(_0415_),
    .B(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__nor3_1 _1370_ (.A(_0435_),
    .B(_0440_),
    .C(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__a311oi_2 _1371_ (.A1(_0411_),
    .A2(_0414_),
    .A3(_0422_),
    .B1(_0437_),
    .C1(_0444_),
    .Y(net41));
 sky130_fd_sc_hd__nor2_1 _1372_ (.A(_0159_),
    .B(_0252_),
    .Y(_0445_));
 sky130_fd_sc_hd__nor2_1 _1373_ (.A(_0112_),
    .B(_0267_),
    .Y(_0446_));
 sky130_fd_sc_hd__nor2_1 _1374_ (.A(_0445_),
    .B(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__nor3_1 _1375_ (.A(_0216_),
    .B(_0131_),
    .C(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__nor2b_1 _1376_ (.A(_0251_),
    .B_N(_0431_),
    .Y(_0449_));
 sky130_fd_sc_hd__nor2_1 _1377_ (.A(_0159_),
    .B(_0268_),
    .Y(_0450_));
 sky130_fd_sc_hd__nor2_1 _1378_ (.A(_0112_),
    .B(_0247_),
    .Y(_0451_));
 sky130_fd_sc_hd__nor2_1 _1379_ (.A(_0450_),
    .B(_0451_),
    .Y(_0452_));
 sky130_fd_sc_hd__nand2_1 _1380_ (.A(_0036_),
    .B(_0131_),
    .Y(_0453_));
 sky130_fd_sc_hd__o22ai_1 _1381_ (.A1(_0036_),
    .A2(_0449_),
    .B1(_0452_),
    .B2(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__o31a_1 _1382_ (.A1(_0107_),
    .A2(_0448_),
    .A3(_0454_),
    .B1(_0041_),
    .X(_0455_));
 sky130_fd_sc_hd__nor2_1 _1383_ (.A(_0298_),
    .B(_0259_),
    .Y(_0456_));
 sky130_fd_sc_hd__a21oi_2 _1384_ (.A1(_0064_),
    .A2(_0263_),
    .B1(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__mux4_2 _1385_ (.A0(_0095_),
    .A1(_0094_),
    .A2(_0093_),
    .A3(_0135_),
    .S0(_0123_),
    .S1(_0084_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2i_2 _1386_ (.A0(_0260_),
    .A1(_0458_),
    .S(_0177_),
    .Y(_0459_));
 sky130_fd_sc_hd__nor2_1 _1387_ (.A(_0258_),
    .B(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__a21oi_1 _1388_ (.A1(_0066_),
    .A2(_0457_),
    .B1(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__mux2i_4 _1389_ (.A0(_0095_),
    .A1(_0093_),
    .S(_0133_),
    .Y(_0462_));
 sky130_fd_sc_hd__mux2i_4 _1390_ (.A0(_0407_),
    .A1(_0462_),
    .S(_0053_),
    .Y(_0463_));
 sky130_fd_sc_hd__inv_1 _1391_ (.A(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__a22o_2 _1392_ (.A1(_0858_),
    .A2(_0879_),
    .B1(_0010_),
    .B2(_0868_),
    .X(_0465_));
 sky130_fd_sc_hd__mux4_4 _1393_ (.A0(_0206_),
    .A1(_0200_),
    .A2(_0273_),
    .A3(_0277_),
    .S0(_0157_),
    .S1(_0693_),
    .X(_0466_));
 sky130_fd_sc_hd__and2_0 _1394_ (.A(_0192_),
    .B(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__a221oi_4 _1395_ (.A1(_0280_),
    .A2(_0403_),
    .B1(_0464_),
    .B2(_0465_),
    .C1(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__a221oi_2 _1396_ (.A1(_0250_),
    .A2(_0413_),
    .B1(_0468_),
    .B2(_0110_),
    .C1(_0041_),
    .Y(_0469_));
 sky130_fd_sc_hd__buf_2 _1397_ (.A(_0045_),
    .X(_0470_));
 sky130_fd_sc_hd__nor2_1 _1398_ (.A(_0231_),
    .B(_0287_),
    .Y(_0471_));
 sky130_fd_sc_hd__nor2_1 _1399_ (.A(_0087_),
    .B(_0290_),
    .Y(_0472_));
 sky130_fd_sc_hd__nor2_1 _1400_ (.A(_0471_),
    .B(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__mux4_1 _1401_ (.A0(_0048_),
    .A1(_0058_),
    .A2(_0055_),
    .A3(_0059_),
    .S0(_0096_),
    .S1(_0097_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2i_2 _1402_ (.A0(_0284_),
    .A1(_0474_),
    .S(_0063_),
    .Y(_0475_));
 sky130_fd_sc_hd__nand2_1 _1403_ (.A(_0470_),
    .B(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__o21ai_0 _1404_ (.A1(_0470_),
    .A2(_0473_),
    .B1(_0476_),
    .Y(_0477_));
 sky130_fd_sc_hd__a22oi_1 _1405_ (.A1(_0455_),
    .A2(_0461_),
    .B1(_0469_),
    .B2(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__clkbuf_4 _1406_ (.A(_0043_),
    .X(_0479_));
 sky130_fd_sc_hd__o21ai_0 _1407_ (.A1(_0455_),
    .A2(_0469_),
    .B1(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__and2_0 _1408_ (.A(_0478_),
    .B(_0480_),
    .X(net42));
 sky130_fd_sc_hd__mux2i_4 _1409_ (.A0(_0305_),
    .A1(_0310_),
    .S(_0158_),
    .Y(_0481_));
 sky130_fd_sc_hd__nor2_2 _1410_ (.A(_0295_),
    .B(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__nand2_1 _1411_ (.A(_0159_),
    .B(_0277_),
    .Y(_0483_));
 sky130_fd_sc_hd__nand2_1 _1412_ (.A(_0112_),
    .B(_0273_),
    .Y(_0484_));
 sky130_fd_sc_hd__a21oi_4 _1413_ (.A1(_0483_),
    .A2(_0484_),
    .B1(_0120_),
    .Y(_0485_));
 sky130_fd_sc_hd__a22oi_2 _1414_ (.A1(_0317_),
    .A2(_0482_),
    .B1(_0485_),
    .B2(_0193_),
    .Y(_0486_));
 sky130_fd_sc_hd__mux2i_4 _1415_ (.A0(_0068_),
    .A1(_0094_),
    .S(_0196_),
    .Y(_0487_));
 sky130_fd_sc_hd__mux2i_4 _1416_ (.A0(_0462_),
    .A1(_0487_),
    .S(_0053_),
    .Y(_0488_));
 sky130_fd_sc_hd__nor2_1 _1417_ (.A(_0295_),
    .B(_0311_),
    .Y(_0489_));
 sky130_fd_sc_hd__a21oi_2 _1418_ (.A1(_0295_),
    .A2(_0279_),
    .B1(_0489_),
    .Y(_0490_));
 sky130_fd_sc_hd__a2bb2oi_1 _1419_ (.A1_N(_0030_),
    .A2_N(_0488_),
    .B1(_0403_),
    .B2(_0490_),
    .Y(_0491_));
 sky130_fd_sc_hd__a31o_1 _1420_ (.A1(_0465_),
    .A2(_0147_),
    .A3(_0315_),
    .B1(_0040_),
    .X(_0492_));
 sky130_fd_sc_hd__a31oi_4 _1421_ (.A1(_0110_),
    .A2(_0486_),
    .A3(_0491_),
    .B1(_0492_),
    .Y(_0493_));
 sky130_fd_sc_hd__a221oi_1 _1422_ (.A1(_0110_),
    .A2(_0165_),
    .B1(_0413_),
    .B2(_0796_),
    .C1(_0434_),
    .Y(_0494_));
 sky130_fd_sc_hd__nor2_1 _1423_ (.A(_0231_),
    .B(_0342_),
    .Y(_0495_));
 sky130_fd_sc_hd__mux4_2 _1424_ (.A0(net8),
    .A1(net7),
    .A2(net6),
    .A3(net5),
    .S0(_0765_),
    .S1(_0060_),
    .X(_0496_));
 sky130_fd_sc_hd__nor2_1 _1425_ (.A(_0087_),
    .B(_0496_),
    .Y(_0497_));
 sky130_fd_sc_hd__nor2_1 _1426_ (.A(_0495_),
    .B(_0497_),
    .Y(_0498_));
 sky130_fd_sc_hd__mux2i_4 _1427_ (.A0(_0339_),
    .A1(_0341_),
    .S(_0177_),
    .Y(_0499_));
 sky130_fd_sc_hd__nand2_1 _1428_ (.A(_0415_),
    .B(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__o21ai_0 _1429_ (.A1(_0415_),
    .A2(_0498_),
    .B1(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__o21a_1 _1430_ (.A1(_0493_),
    .A2(_0494_),
    .B1(_0479_),
    .X(_0502_));
 sky130_fd_sc_hd__a221oi_1 _1431_ (.A1(_0078_),
    .A2(_0493_),
    .B1(_0494_),
    .B2(_0501_),
    .C1(_0502_),
    .Y(net43));
 sky130_fd_sc_hd__mux2i_2 _1432_ (.A0(_0311_),
    .A1(_0487_),
    .S(_0158_),
    .Y(_0503_));
 sky130_fd_sc_hd__mux2i_2 _1433_ (.A0(_0069_),
    .A1(_0095_),
    .S(_0196_),
    .Y(_0504_));
 sky130_fd_sc_hd__mux2i_4 _1434_ (.A0(_0375_),
    .A1(_0504_),
    .S(_0158_),
    .Y(_0505_));
 sky130_fd_sc_hd__mux2i_4 _1435_ (.A0(_0503_),
    .A1(_0505_),
    .S(_0704_),
    .Y(_0506_));
 sky130_fd_sc_hd__mux2i_4 _1436_ (.A0(_0199_),
    .A1(_0481_),
    .S(_0785_),
    .Y(_0507_));
 sky130_fd_sc_hd__nor2_1 _1437_ (.A(_0138_),
    .B(_0365_),
    .Y(_0508_));
 sky130_fd_sc_hd__a21oi_1 _1438_ (.A1(_0508_),
    .A2(_0431_),
    .B1(_0036_),
    .Y(_0509_));
 sky130_fd_sc_hd__a221oi_4 _1439_ (.A1(_0423_),
    .A2(_0506_),
    .B1(_0507_),
    .B2(_0332_),
    .C1(_0509_),
    .Y(_0510_));
 sky130_fd_sc_hd__a21oi_1 _1440_ (.A1(_0215_),
    .A2(_0510_),
    .B1(_0040_),
    .Y(_0511_));
 sky130_fd_sc_hd__nand2_1 _1441_ (.A(_0298_),
    .B(_0393_),
    .Y(_0512_));
 sky130_fd_sc_hd__o21ai_2 _1442_ (.A1(_0298_),
    .A2(_0382_),
    .B1(_0512_),
    .Y(_0513_));
 sky130_fd_sc_hd__mux2i_4 _1443_ (.A0(_0383_),
    .A1(_0386_),
    .S(_0177_),
    .Y(_0514_));
 sky130_fd_sc_hd__nor2_1 _1444_ (.A(_0258_),
    .B(_0514_),
    .Y(_0515_));
 sky130_fd_sc_hd__a21oi_1 _1445_ (.A1(_0258_),
    .A2(_0513_),
    .B1(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__nand2_1 _1446_ (.A(_0316_),
    .B(_0189_),
    .Y(_0517_));
 sky130_fd_sc_hd__mux4_4 _1447_ (.A0(_0355_),
    .A1(_0349_),
    .A2(_0356_),
    .A3(_0350_),
    .S0(_0157_),
    .S1(_0072_),
    .X(_0518_));
 sky130_fd_sc_hd__nor2_1 _1448_ (.A(_0128_),
    .B(_0518_),
    .Y(_0519_));
 sky130_fd_sc_hd__a221o_2 _1449_ (.A1(_0465_),
    .A2(_0360_),
    .B1(_0348_),
    .B2(_0403_),
    .C1(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__o221ai_4 _1450_ (.A1(_0365_),
    .A2(_0517_),
    .B1(_0520_),
    .B2(_0037_),
    .C1(_0040_),
    .Y(_0521_));
 sky130_fd_sc_hd__nand2b_1 _1451_ (.A_N(_0511_),
    .B(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__nor2_1 _1452_ (.A(_0231_),
    .B(_0370_),
    .Y(_0523_));
 sky130_fd_sc_hd__mux4_2 _1453_ (.A0(_0069_),
    .A1(_0068_),
    .A2(_0095_),
    .A3(_0094_),
    .S0(_0207_),
    .S1(_0090_),
    .X(_0524_));
 sky130_fd_sc_hd__nor2_1 _1454_ (.A(_0087_),
    .B(_0524_),
    .Y(_0525_));
 sky130_fd_sc_hd__nor2_1 _1455_ (.A(_0523_),
    .B(_0525_),
    .Y(_0526_));
 sky130_fd_sc_hd__nand2_1 _1456_ (.A(_0064_),
    .B(_0367_),
    .Y(_0527_));
 sky130_fd_sc_hd__o21ai_2 _1457_ (.A1(_0064_),
    .A2(_0369_),
    .B1(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__nor2_1 _1458_ (.A(_0391_),
    .B(_0528_),
    .Y(_0529_));
 sky130_fd_sc_hd__a211oi_1 _1459_ (.A1(_0391_),
    .A2(_0526_),
    .B1(_0529_),
    .C1(_0521_),
    .Y(_0530_));
 sky130_fd_sc_hd__a221oi_1 _1460_ (.A1(_0511_),
    .A2(_0516_),
    .B1(_0522_),
    .B2(_0479_),
    .C1(_0530_),
    .Y(net44));
 sky130_fd_sc_hd__nor2_1 _1461_ (.A(_0391_),
    .B(_0232_),
    .Y(_0531_));
 sky130_fd_sc_hd__nor2_1 _1462_ (.A(_0178_),
    .B(_0441_),
    .Y(_0532_));
 sky130_fd_sc_hd__mux4_2 _1463_ (.A0(net10),
    .A1(_0069_),
    .A2(net8),
    .A3(_0095_),
    .S0(_0765_),
    .S1(_0097_),
    .X(_0533_));
 sky130_fd_sc_hd__nor2_1 _1464_ (.A(_0320_),
    .B(_0533_),
    .Y(_0534_));
 sky130_fd_sc_hd__nor3_1 _1465_ (.A(_0415_),
    .B(_0532_),
    .C(_0534_),
    .Y(_0535_));
 sky130_fd_sc_hd__o21ai_0 _1466_ (.A1(_0531_),
    .A2(_0535_),
    .B1(_0170_),
    .Y(_0536_));
 sky130_fd_sc_hd__nor2_1 _1467_ (.A(_0159_),
    .B(_0240_),
    .Y(_0537_));
 sky130_fd_sc_hd__nor2_1 _1468_ (.A(_0143_),
    .B(_0218_),
    .Y(_0538_));
 sky130_fd_sc_hd__or3_1 _1469_ (.A(_0193_),
    .B(_0537_),
    .C(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__o21ai_0 _1470_ (.A1(_0246_),
    .A2(_0224_),
    .B1(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__o31ai_1 _1471_ (.A1(_0320_),
    .A2(_0234_),
    .A3(_0301_),
    .B1(_0167_),
    .Y(_0541_));
 sky130_fd_sc_hd__a21oi_1 _1472_ (.A1(_0191_),
    .A2(_0540_),
    .B1(_0541_),
    .Y(_0542_));
 sky130_fd_sc_hd__nand2_1 _1473_ (.A(_0265_),
    .B(_0204_),
    .Y(_0543_));
 sky130_fd_sc_hd__mux2_1 _1474_ (.A0(_0070_),
    .A1(_0068_),
    .S(_0133_),
    .X(_0544_));
 sky130_fd_sc_hd__nor2_1 _1475_ (.A(_0221_),
    .B(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__a211oi_1 _1476_ (.A1(_0113_),
    .A2(_0407_),
    .B1(_0545_),
    .C1(_0195_),
    .Y(_0546_));
 sky130_fd_sc_hd__a21oi_2 _1477_ (.A1(_0195_),
    .A2(_0505_),
    .B1(_0546_),
    .Y(_0547_));
 sky130_fd_sc_hd__nand2_1 _1478_ (.A(_0246_),
    .B(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__nor2_1 _1479_ (.A(_0258_),
    .B(_0174_),
    .Y(_0549_));
 sky130_fd_sc_hd__a21oi_1 _1480_ (.A1(_0046_),
    .A2(_0188_),
    .B1(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__a31oi_1 _1481_ (.A1(_0465_),
    .A2(_0147_),
    .A3(_0209_),
    .B1(_0041_),
    .Y(_0551_));
 sky130_fd_sc_hd__o21ai_0 _1482_ (.A1(_0257_),
    .A2(_0550_),
    .B1(_0551_),
    .Y(_0552_));
 sky130_fd_sc_hd__a31oi_1 _1483_ (.A1(_0191_),
    .A2(_0543_),
    .A3(_0548_),
    .B1(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__a21oi_1 _1484_ (.A1(_0536_),
    .A2(_0542_),
    .B1(_0553_),
    .Y(net45));
 sky130_fd_sc_hd__nor2_1 _1485_ (.A(_0046_),
    .B(_0289_),
    .Y(_0554_));
 sky130_fd_sc_hd__a211oi_1 _1486_ (.A1(_0470_),
    .A2(_0300_),
    .B1(_0554_),
    .C1(_0043_),
    .Y(_0555_));
 sky130_fd_sc_hd__o21ai_1 _1487_ (.A1(_0238_),
    .A2(_0278_),
    .B1(_0281_),
    .Y(_0556_));
 sky130_fd_sc_hd__mux2_1 _1488_ (.A0(_0071_),
    .A1(_0069_),
    .S(_0196_),
    .X(_0557_));
 sky130_fd_sc_hd__mux2i_4 _1489_ (.A0(_0544_),
    .A1(_0557_),
    .S(_0120_),
    .Y(_0558_));
 sky130_fd_sc_hd__o22ai_1 _1490_ (.A1(_0225_),
    .A2(_0276_),
    .B1(_0558_),
    .B2(_0216_),
    .Y(_0559_));
 sky130_fd_sc_hd__nand2_1 _1491_ (.A(_0221_),
    .B(_0463_),
    .Y(_0560_));
 sky130_fd_sc_hd__a21oi_1 _1492_ (.A1(_0129_),
    .A2(_0560_),
    .B1(_0216_),
    .Y(_0561_));
 sky130_fd_sc_hd__a21oi_1 _1493_ (.A1(_0238_),
    .A2(_0559_),
    .B1(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__a211oi_4 _1494_ (.A1(_0556_),
    .A2(_0332_),
    .B1(_0562_),
    .C1(_0107_),
    .Y(_0563_));
 sky130_fd_sc_hd__nor2_1 _1495_ (.A(_0194_),
    .B(_0269_),
    .Y(_0564_));
 sky130_fd_sc_hd__a21oi_2 _1496_ (.A1(_0194_),
    .A2(_0254_),
    .B1(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__nor2_1 _1497_ (.A(_0181_),
    .B(_0261_),
    .Y(_0566_));
 sky130_fd_sc_hd__mux4_2 _1498_ (.A0(_0071_),
    .A1(_0070_),
    .A2(_0069_),
    .A3(_0068_),
    .S0(_0207_),
    .S1(_0286_),
    .X(_0567_));
 sky130_fd_sc_hd__mux2i_2 _1499_ (.A0(_0458_),
    .A1(_0567_),
    .S(_0231_),
    .Y(_0568_));
 sky130_fd_sc_hd__nor2_1 _1500_ (.A(_0046_),
    .B(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__nor2_1 _1501_ (.A(_0566_),
    .B(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__nor3_1 _1502_ (.A(_0320_),
    .B(_0301_),
    .C(_0263_),
    .Y(_0571_));
 sky130_fd_sc_hd__nor2_1 _1503_ (.A(_0434_),
    .B(_0571_),
    .Y(_0572_));
 sky130_fd_sc_hd__o221ai_1 _1504_ (.A1(_0038_),
    .A2(_0565_),
    .B1(_0570_),
    .B2(_0479_),
    .C1(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__o31a_1 _1505_ (.A1(_0327_),
    .A2(_0555_),
    .A3(_0563_),
    .B1(_0573_),
    .X(net46));
 sky130_fd_sc_hd__mux2i_1 _1506_ (.A0(_0080_),
    .A1(_0082_),
    .S(_0745_),
    .Y(_0574_));
 sky130_fd_sc_hd__mux2i_1 _1507_ (.A0(_0081_),
    .A1(_0117_),
    .S(_0060_),
    .Y(_0575_));
 sky130_fd_sc_hd__mux2i_2 _1508_ (.A0(_0574_),
    .A1(_0575_),
    .S(_0208_),
    .Y(_0576_));
 sky130_fd_sc_hd__nor2_1 _1509_ (.A(_0177_),
    .B(_0576_),
    .Y(_0577_));
 sky130_fd_sc_hd__mux4_1 _1510_ (.A0(net12),
    .A1(_0088_),
    .A2(_0089_),
    .A3(_0079_),
    .S0(_0083_),
    .S1(_0084_),
    .X(_0578_));
 sky130_fd_sc_hd__nor2_1 _1511_ (.A(_0064_),
    .B(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__nor2_1 _1512_ (.A(_0177_),
    .B(_0387_),
    .Y(_0580_));
 sky130_fd_sc_hd__mux4_2 _1513_ (.A0(net31),
    .A1(net2),
    .A2(net3),
    .A3(_0135_),
    .S0(_0096_),
    .S1(_0097_),
    .X(_0581_));
 sky130_fd_sc_hd__nor2_1 _1514_ (.A(_0298_),
    .B(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__nor2_1 _1515_ (.A(_0580_),
    .B(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__nand2_1 _1516_ (.A(_0045_),
    .B(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__o311a_1 _1517_ (.A1(_0020_),
    .A2(_0577_),
    .A3(_0579_),
    .B1(_0584_),
    .C1(_0034_),
    .X(_0585_));
 sky130_fd_sc_hd__a21oi_1 _1518_ (.A1(_0043_),
    .A2(_0516_),
    .B1(_0585_),
    .Y(_0586_));
 sky130_fd_sc_hd__nor4_1 _1519_ (.A(_0847_),
    .B(_0030_),
    .C(_0038_),
    .D(_0365_),
    .Y(_0587_));
 sky130_fd_sc_hd__o21ai_0 _1520_ (.A1(_0032_),
    .A2(_0365_),
    .B1(_0327_),
    .Y(_0588_));
 sky130_fd_sc_hd__nand2_1 _1521_ (.A(_0033_),
    .B(_0108_),
    .Y(_0589_));
 sky130_fd_sc_hd__mux2i_1 _1522_ (.A0(_0081_),
    .A1(_0117_),
    .S(_0138_),
    .Y(_0590_));
 sky130_fd_sc_hd__nand2_1 _1523_ (.A(_0195_),
    .B(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__nand2_1 _1524_ (.A(_0920_),
    .B(_0139_),
    .Y(_0592_));
 sky130_fd_sc_hd__nand3_1 _1525_ (.A(_0129_),
    .B(_0591_),
    .C(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__o21ai_1 _1526_ (.A1(_0129_),
    .A2(_0354_),
    .B1(_0593_),
    .Y(_0594_));
 sky130_fd_sc_hd__mux2i_1 _1527_ (.A0(_0118_),
    .A1(_0135_),
    .S(_0133_),
    .Y(_0595_));
 sky130_fd_sc_hd__mux2_1 _1528_ (.A0(_0116_),
    .A1(_0595_),
    .S(_0124_),
    .X(_0596_));
 sky130_fd_sc_hd__mux4_1 _1529_ (.A0(net12),
    .A1(_0088_),
    .A2(_0089_),
    .A3(_0079_),
    .S0(_0124_),
    .S1(_0847_),
    .X(_0597_));
 sky130_fd_sc_hd__nand2_1 _1530_ (.A(_0132_),
    .B(_0597_),
    .Y(_0598_));
 sky130_fd_sc_hd__o211ai_1 _1531_ (.A1(_0272_),
    .A2(_0596_),
    .B1(_0598_),
    .C1(_0329_),
    .Y(_0599_));
 sky130_fd_sc_hd__o21ai_0 _1532_ (.A1(_0329_),
    .A2(_0594_),
    .B1(_0599_),
    .Y(_0600_));
 sky130_fd_sc_hd__o22ai_1 _1533_ (.A1(_0589_),
    .A2(_0520_),
    .B1(_0600_),
    .B2(_0038_),
    .Y(_0601_));
 sky130_fd_sc_hd__o32a_1 _1534_ (.A1(_0167_),
    .A2(_0586_),
    .A3(_0587_),
    .B1(_0588_),
    .B2(_0601_),
    .X(net47));
 sky130_fd_sc_hd__nand3_4 _1535_ (.A(_0033_),
    .B(_0036_),
    .C(_0128_),
    .Y(_0602_));
 sky130_fd_sc_hd__nor2_1 _1536_ (.A(_0237_),
    .B(_0488_),
    .Y(_0603_));
 sky130_fd_sc_hd__mux2i_2 _1537_ (.A0(_0150_),
    .A1(_0070_),
    .S(_0217_),
    .Y(_0604_));
 sky130_fd_sc_hd__nand2_1 _1538_ (.A(_0785_),
    .B(_0557_),
    .Y(_0605_));
 sky130_fd_sc_hd__o21ai_4 _1539_ (.A1(_0785_),
    .A2(_0604_),
    .B1(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__nor2_1 _1540_ (.A(_0143_),
    .B(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__a31oi_1 _1541_ (.A1(_0109_),
    .A2(_0193_),
    .A3(_0313_),
    .B1(_0040_),
    .Y(_0608_));
 sky130_fd_sc_hd__nand2_1 _1542_ (.A(_0112_),
    .B(_0315_),
    .Y(_0609_));
 sky130_fd_sc_hd__a211o_1 _1543_ (.A1(_0307_),
    .A2(_0609_),
    .B1(_0192_),
    .C1(_0589_),
    .X(_0610_));
 sky130_fd_sc_hd__o311a_1 _1544_ (.A1(_0602_),
    .A2(_0603_),
    .A3(_0607_),
    .B1(_0608_),
    .C1(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__o221ai_1 _1545_ (.A1(_0062_),
    .A2(_0235_),
    .B1(_0323_),
    .B2(_0415_),
    .C1(_0611_),
    .Y(_0612_));
 sky130_fd_sc_hd__and2_0 _1546_ (.A(_0161_),
    .B(_0210_),
    .X(_0613_));
 sky130_fd_sc_hd__a221o_1 _1547_ (.A1(_0465_),
    .A2(_0153_),
    .B1(_0403_),
    .B2(_0162_),
    .C1(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__o21ai_0 _1548_ (.A1(_0301_),
    .A2(_0340_),
    .B1(_0040_),
    .Y(_0615_));
 sky130_fd_sc_hd__a21oi_1 _1549_ (.A1(_0110_),
    .A2(_0614_),
    .B1(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__mux4_2 _1550_ (.A0(net13),
    .A1(net11),
    .A2(net10),
    .A3(net9),
    .S0(_0765_),
    .S1(_0060_),
    .X(_0617_));
 sky130_fd_sc_hd__mux2_1 _1551_ (.A0(_0496_),
    .A1(_0617_),
    .S(_0101_),
    .X(_0618_));
 sky130_fd_sc_hd__nand2_1 _1552_ (.A(_0391_),
    .B(_0618_),
    .Y(_0619_));
 sky130_fd_sc_hd__o211ai_1 _1553_ (.A1(_0391_),
    .A2(_0343_),
    .B1(_0616_),
    .C1(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__o21ai_0 _1554_ (.A1(_0611_),
    .A2(_0616_),
    .B1(_0479_),
    .Y(_0621_));
 sky130_fd_sc_hd__and3_1 _1555_ (.A(_0612_),
    .B(_0620_),
    .C(_0621_),
    .X(net48));
 sky130_fd_sc_hd__mux4_2 _1556_ (.A0(_0172_),
    .A1(_0150_),
    .A2(_0071_),
    .A3(_0070_),
    .S0(_0207_),
    .S1(_0090_),
    .X(_0622_));
 sky130_fd_sc_hd__mux2i_2 _1557_ (.A0(_0524_),
    .A1(_0622_),
    .S(_0075_),
    .Y(_0623_));
 sky130_fd_sc_hd__mux2i_1 _1558_ (.A0(_0371_),
    .A1(_0623_),
    .S(_0391_),
    .Y(_0624_));
 sky130_fd_sc_hd__nor2_1 _1559_ (.A(_0301_),
    .B(_0368_),
    .Y(_0625_));
 sky130_fd_sc_hd__a21oi_1 _1560_ (.A1(_0170_),
    .A2(_0624_),
    .B1(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__or3_1 _1561_ (.A(_0131_),
    .B(_0143_),
    .C(_0357_),
    .X(_0627_));
 sky130_fd_sc_hd__o21ai_1 _1562_ (.A1(_0194_),
    .A2(_0352_),
    .B1(_0627_),
    .Y(_0628_));
 sky130_fd_sc_hd__clkbuf_4 _1563_ (.A(_0434_),
    .X(_0629_));
 sky130_fd_sc_hd__a21oi_1 _1564_ (.A1(_0191_),
    .A2(_0628_),
    .B1(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__o21ai_2 _1565_ (.A1(_0144_),
    .A2(_0378_),
    .B1(_0379_),
    .Y(_0631_));
 sky130_fd_sc_hd__or2_0 _1566_ (.A(_0120_),
    .B(_0487_),
    .X(_0632_));
 sky130_fd_sc_hd__mux2_1 _1567_ (.A0(_0069_),
    .A1(_0095_),
    .S(_0217_),
    .X(_0633_));
 sky130_fd_sc_hd__nand2_1 _1568_ (.A(_0920_),
    .B(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__mux4_1 _1569_ (.A0(_0172_),
    .A1(_0150_),
    .A2(_0071_),
    .A3(_0070_),
    .S0(_0775_),
    .S1(_0138_),
    .X(_0635_));
 sky130_fd_sc_hd__nor2_1 _1570_ (.A(_0221_),
    .B(_0635_),
    .Y(_0636_));
 sky130_fd_sc_hd__a31oi_2 _1571_ (.A1(_0113_),
    .A2(_0632_),
    .A3(_0634_),
    .B1(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__nand2_1 _1572_ (.A(_0362_),
    .B(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__o21ai_0 _1573_ (.A1(_0362_),
    .A2(_0631_),
    .B1(_0638_),
    .Y(_0639_));
 sky130_fd_sc_hd__nand3_1 _1574_ (.A(_0045_),
    .B(_0231_),
    .C(_0393_),
    .Y(_0640_));
 sky130_fd_sc_hd__a21boi_2 _1575_ (.A1(_0181_),
    .A2(_0385_),
    .B1_N(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__a31oi_1 _1576_ (.A1(_0111_),
    .A2(_0265_),
    .A3(_0377_),
    .B1(_0041_),
    .Y(_0642_));
 sky130_fd_sc_hd__o21ai_0 _1577_ (.A1(_0257_),
    .A2(_0641_),
    .B1(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__a31oi_1 _1578_ (.A1(_0215_),
    .A2(_0246_),
    .A3(_0639_),
    .B1(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__a21oi_1 _1579_ (.A1(_0626_),
    .A2(_0630_),
    .B1(_0644_),
    .Y(net49));
 sky130_fd_sc_hd__nand2_1 _1580_ (.A(_0020_),
    .B(_0316_),
    .Y(_0645_));
 sky130_fd_sc_hd__o22ai_1 _1581_ (.A1(_0020_),
    .A2(_0420_),
    .B1(_0645_),
    .B2(_0187_),
    .Y(_0646_));
 sky130_fd_sc_hd__mux4_1 _1582_ (.A0(_0151_),
    .A1(net14),
    .A2(net13),
    .A3(_0071_),
    .S0(_0072_),
    .S1(_0745_),
    .X(_0647_));
 sky130_fd_sc_hd__mux2i_1 _1583_ (.A0(_0533_),
    .A1(_0647_),
    .S(_0101_),
    .Y(_0648_));
 sky130_fd_sc_hd__mux2i_1 _1584_ (.A0(_0442_),
    .A1(_0648_),
    .S(_0180_),
    .Y(_0649_));
 sky130_fd_sc_hd__mux2_1 _1585_ (.A0(_0646_),
    .A1(_0649_),
    .S(_0040_),
    .X(_0650_));
 sky130_fd_sc_hd__clkbuf_4 _1586_ (.A(_0192_),
    .X(_0651_));
 sky130_fd_sc_hd__nor2_1 _1587_ (.A(_0651_),
    .B(_0426_),
    .Y(_0652_));
 sky130_fd_sc_hd__a31oi_2 _1588_ (.A1(_0651_),
    .A2(_0238_),
    .A3(_0427_),
    .B1(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__o22ai_1 _1589_ (.A1(_0301_),
    .A2(_0439_),
    .B1(_0653_),
    .B2(_0038_),
    .Y(_0654_));
 sky130_fd_sc_hd__nor2_1 _1590_ (.A(_0143_),
    .B(_0408_),
    .Y(_0655_));
 sky130_fd_sc_hd__a21oi_1 _1591_ (.A1(_0221_),
    .A2(_0398_),
    .B1(_0655_),
    .Y(_0656_));
 sky130_fd_sc_hd__nand2_1 _1592_ (.A(_0120_),
    .B(_0544_),
    .Y(_0657_));
 sky130_fd_sc_hd__nand2_1 _1593_ (.A(_0295_),
    .B(_0633_),
    .Y(_0658_));
 sky130_fd_sc_hd__mux4_1 _1594_ (.A0(_0151_),
    .A1(_0172_),
    .A2(_0150_),
    .A3(_0071_),
    .S0(_0123_),
    .S1(_0837_),
    .X(_0659_));
 sky130_fd_sc_hd__nor2_1 _1595_ (.A(_0143_),
    .B(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__a31oi_2 _1596_ (.A1(_0221_),
    .A2(_0657_),
    .A3(_0658_),
    .B1(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__nor2_1 _1597_ (.A(_0225_),
    .B(_0406_),
    .Y(_0662_));
 sky130_fd_sc_hd__a221oi_1 _1598_ (.A1(_0332_),
    .A2(_0656_),
    .B1(_0661_),
    .B2(_0423_),
    .C1(_0662_),
    .Y(_0663_));
 sky130_fd_sc_hd__nor3_1 _1599_ (.A(_0041_),
    .B(_0107_),
    .C(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__a221o_1 _1600_ (.A1(_0170_),
    .A2(_0650_),
    .B1(_0654_),
    .B2(_0167_),
    .C1(_0664_),
    .X(net50));
 sky130_fd_sc_hd__mux4_2 _1601_ (.A0(_0239_),
    .A1(_0151_),
    .A2(_0172_),
    .A3(_0150_),
    .S0(_0083_),
    .S1(_0286_),
    .X(_0665_));
 sky130_fd_sc_hd__mux2i_2 _1602_ (.A0(_0567_),
    .A1(_0665_),
    .S(_0075_),
    .Y(_0666_));
 sky130_fd_sc_hd__mux2i_1 _1603_ (.A0(_0459_),
    .A1(_0666_),
    .S(_0391_),
    .Y(_0667_));
 sky130_fd_sc_hd__nor2_1 _1604_ (.A(_0045_),
    .B(_0475_),
    .Y(_0668_));
 sky130_fd_sc_hd__a41oi_2 _1605_ (.A1(_0045_),
    .A2(_0231_),
    .A3(_0056_),
    .A4(_0889_),
    .B1(_0668_),
    .Y(_0669_));
 sky130_fd_sc_hd__nor2_1 _1606_ (.A(_0167_),
    .B(_0669_),
    .Y(_0670_));
 sky130_fd_sc_hd__a21oi_1 _1607_ (.A1(_0042_),
    .A2(_0667_),
    .B1(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__mux2i_2 _1608_ (.A0(_0239_),
    .A1(_0172_),
    .S(_0138_),
    .Y(_0673_));
 sky130_fd_sc_hd__nand2b_1 _1609_ (.A_N(_0150_),
    .B(_0217_),
    .Y(_0674_));
 sky130_fd_sc_hd__o211ai_1 _1610_ (.A1(_0151_),
    .A2(_0847_),
    .B1(_0674_),
    .C1(_0295_),
    .Y(_0675_));
 sky130_fd_sc_hd__o21ai_2 _1611_ (.A1(_0295_),
    .A2(_0673_),
    .B1(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__mux2i_2 _1612_ (.A0(_0463_),
    .A1(_0676_),
    .S(_0129_),
    .Y(_0677_));
 sky130_fd_sc_hd__nand2_1 _1613_ (.A(_0651_),
    .B(_0280_),
    .Y(_0678_));
 sky130_fd_sc_hd__nand2_1 _1614_ (.A(_0272_),
    .B(_0558_),
    .Y(_0679_));
 sky130_fd_sc_hd__nand3_1 _1615_ (.A(_0114_),
    .B(_0678_),
    .C(_0679_),
    .Y(_0680_));
 sky130_fd_sc_hd__o211ai_2 _1616_ (.A1(_0114_),
    .A2(_0677_),
    .B1(_0680_),
    .C1(_0362_),
    .Y(_0681_));
 sky130_fd_sc_hd__o21ai_0 _1617_ (.A1(_0265_),
    .A2(_0466_),
    .B1(_0216_),
    .Y(_0682_));
 sky130_fd_sc_hd__a31oi_1 _1618_ (.A1(_0215_),
    .A2(_0681_),
    .A3(_0682_),
    .B1(_0042_),
    .Y(_0684_));
 sky130_fd_sc_hd__nand2_1 _1619_ (.A(_0246_),
    .B(_0447_),
    .Y(_0685_));
 sky130_fd_sc_hd__o31ai_2 _1620_ (.A1(_0272_),
    .A2(_0144_),
    .A3(_0251_),
    .B1(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__a221oi_1 _1621_ (.A1(_0189_),
    .A2(_0457_),
    .B1(_0686_),
    .B2(_0111_),
    .C1(_0629_),
    .Y(_0687_));
 sky130_fd_sc_hd__o22ai_2 _1622_ (.A1(_0479_),
    .A2(_0671_),
    .B1(_0684_),
    .B2(_0687_),
    .Y(net51));
 sky130_fd_sc_hd__mux2_1 _1623_ (.A0(_0050_),
    .A1(_0151_),
    .S(_0217_),
    .X(_0688_));
 sky130_fd_sc_hd__nand2_1 _1624_ (.A(_0920_),
    .B(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__o21ai_1 _1625_ (.A1(_0920_),
    .A2(_0673_),
    .B1(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__mux2i_4 _1626_ (.A0(_0488_),
    .A1(_0690_),
    .S(_0132_),
    .Y(_0691_));
 sky130_fd_sc_hd__nor2_1 _1627_ (.A(_0114_),
    .B(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__nor2_1 _1628_ (.A(_0194_),
    .B(_0606_),
    .Y(_0694_));
 sky130_fd_sc_hd__a211oi_1 _1629_ (.A1(_0265_),
    .A2(_0490_),
    .B1(_0694_),
    .C1(_0329_),
    .Y(_0695_));
 sky130_fd_sc_hd__o21ai_0 _1630_ (.A1(_0692_),
    .A2(_0695_),
    .B1(_0191_),
    .Y(_0696_));
 sky130_fd_sc_hd__nor2_4 _1631_ (.A(_0031_),
    .B(_0045_),
    .Y(_0697_));
 sky130_fd_sc_hd__nand3_1 _1632_ (.A(_0237_),
    .B(_0315_),
    .C(_0317_),
    .Y(_0698_));
 sky130_fd_sc_hd__o31ai_1 _1633_ (.A1(_0194_),
    .A2(_0482_),
    .A3(_0485_),
    .B1(_0698_),
    .Y(_0699_));
 sky130_fd_sc_hd__a221oi_1 _1634_ (.A1(_0065_),
    .A2(_0697_),
    .B1(_0148_),
    .B2(_0699_),
    .C1(_0327_),
    .Y(_0700_));
 sky130_fd_sc_hd__nor2_1 _1635_ (.A(_0038_),
    .B(_0265_),
    .Y(_0701_));
 sky130_fd_sc_hd__nor2_1 _1636_ (.A(_0258_),
    .B(_0499_),
    .Y(_0702_));
 sky130_fd_sc_hd__a31oi_2 _1637_ (.A1(_0066_),
    .A2(_0796_),
    .A3(_0316_),
    .B1(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__nor2_1 _1638_ (.A(_0231_),
    .B(_0617_),
    .Y(_0705_));
 sky130_fd_sc_hd__mux4_1 _1639_ (.A0(_0050_),
    .A1(_0239_),
    .A2(_0151_),
    .A3(_0172_),
    .S0(_0123_),
    .S1(_0084_),
    .X(_0706_));
 sky130_fd_sc_hd__nor2_1 _1640_ (.A(_0087_),
    .B(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hd__nor3_1 _1641_ (.A(_0045_),
    .B(_0705_),
    .C(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__a211oi_1 _1642_ (.A1(_0046_),
    .A2(_0498_),
    .B1(_0708_),
    .C1(_0043_),
    .Y(_0709_));
 sky130_fd_sc_hd__a21oi_1 _1643_ (.A1(_0257_),
    .A2(_0703_),
    .B1(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__a211oi_1 _1644_ (.A1(_0163_),
    .A2(_0701_),
    .B1(_0710_),
    .C1(_0629_),
    .Y(_0711_));
 sky130_fd_sc_hd__a21oi_1 _1645_ (.A1(_0696_),
    .A2(_0700_),
    .B1(_0711_),
    .Y(net52));
 sky130_fd_sc_hd__o22ai_2 _1646_ (.A1(_0066_),
    .A2(_0528_),
    .B1(_0645_),
    .B2(_0365_),
    .Y(_0712_));
 sky130_fd_sc_hd__nor2_1 _1647_ (.A(_0178_),
    .B(_0622_),
    .Y(_0713_));
 sky130_fd_sc_hd__mux4_1 _1648_ (.A0(_0047_),
    .A1(_0050_),
    .A2(_0239_),
    .A3(_0151_),
    .S0(_0083_),
    .S1(_0286_),
    .X(_0714_));
 sky130_fd_sc_hd__nor2_1 _1649_ (.A(_0087_),
    .B(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__nor3_1 _1650_ (.A(_0066_),
    .B(_0713_),
    .C(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__a21oi_1 _1651_ (.A1(_0470_),
    .A2(_0526_),
    .B1(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__nor2_1 _1652_ (.A(_0044_),
    .B(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__a21oi_1 _1653_ (.A1(_0479_),
    .A2(_0712_),
    .B1(_0718_),
    .Y(_0719_));
 sky130_fd_sc_hd__nand2_1 _1654_ (.A(_0518_),
    .B(_0701_),
    .Y(_0720_));
 sky130_fd_sc_hd__mux2i_1 _1655_ (.A0(_0047_),
    .A1(_0239_),
    .S(_0217_),
    .Y(_0721_));
 sky130_fd_sc_hd__nor2_1 _1656_ (.A(_0295_),
    .B(_0721_),
    .Y(_0722_));
 sky130_fd_sc_hd__a21oi_1 _1657_ (.A1(_0195_),
    .A2(_0688_),
    .B1(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__nor2_1 _1658_ (.A(_0237_),
    .B(_0635_),
    .Y(_0725_));
 sky130_fd_sc_hd__a211o_1 _1659_ (.A1(_0238_),
    .A2(_0723_),
    .B1(_0725_),
    .C1(_0651_),
    .X(_0726_));
 sky130_fd_sc_hd__o21ai_1 _1660_ (.A1(_0246_),
    .A2(_0506_),
    .B1(_0726_),
    .Y(_0727_));
 sky130_fd_sc_hd__nand2_1 _1661_ (.A(_0210_),
    .B(_0508_),
    .Y(_0728_));
 sky130_fd_sc_hd__o21ai_2 _1662_ (.A1(_0193_),
    .A2(_0507_),
    .B1(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__a221o_1 _1663_ (.A1(_0697_),
    .A2(_0513_),
    .B1(_0729_),
    .B2(_0147_),
    .C1(_0041_),
    .X(_0730_));
 sky130_fd_sc_hd__a21oi_1 _1664_ (.A1(_0191_),
    .A2(_0727_),
    .B1(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__a31oi_1 _1665_ (.A1(_0213_),
    .A2(_0719_),
    .A3(_0720_),
    .B1(_0731_),
    .Y(net53));
 sky130_fd_sc_hd__nor2_1 _1666_ (.A(_0246_),
    .B(_0547_),
    .Y(_0732_));
 sky130_fd_sc_hd__mux2i_1 _1667_ (.A0(_0051_),
    .A1(_0050_),
    .S(_0217_),
    .Y(_0733_));
 sky130_fd_sc_hd__mux2_1 _1668_ (.A0(_0721_),
    .A1(_0733_),
    .S(_0704_),
    .X(_0735_));
 sky130_fd_sc_hd__nor2_1 _1669_ (.A(_0238_),
    .B(_0659_),
    .Y(_0736_));
 sky130_fd_sc_hd__a211oi_1 _1670_ (.A1(_0329_),
    .A2(_0735_),
    .B1(_0736_),
    .C1(_0265_),
    .Y(_0737_));
 sky130_fd_sc_hd__o21ai_0 _1671_ (.A1(_0732_),
    .A2(_0737_),
    .B1(_0191_),
    .Y(_0738_));
 sky130_fd_sc_hd__a221oi_1 _1672_ (.A1(_0697_),
    .A2(_0188_),
    .B1(_0212_),
    .B2(_0148_),
    .C1(_0327_),
    .Y(_0739_));
 sky130_fd_sc_hd__mux4_1 _1673_ (.A0(_0051_),
    .A1(_0047_),
    .A2(_0050_),
    .A3(_0239_),
    .S0(_0072_),
    .S1(_0745_),
    .X(_0740_));
 sky130_fd_sc_hd__mux4_1 _1674_ (.A0(_0441_),
    .A1(_0533_),
    .A2(_0647_),
    .A3(_0740_),
    .S0(_0101_),
    .S1(_0181_),
    .X(_0741_));
 sky130_fd_sc_hd__nand2_1 _1675_ (.A(_0170_),
    .B(_0741_),
    .Y(_0742_));
 sky130_fd_sc_hd__nand2_1 _1676_ (.A(_0044_),
    .B(_0236_),
    .Y(_0743_));
 sky130_fd_sc_hd__o2111a_1 _1677_ (.A1(_0224_),
    .A2(_0602_),
    .B1(_0742_),
    .C1(_0743_),
    .D1(_0327_),
    .X(_0744_));
 sky130_fd_sc_hd__a21oi_1 _1678_ (.A1(_0738_),
    .A2(_0739_),
    .B1(_0744_),
    .Y(net54));
 sky130_fd_sc_hd__nand2_1 _1679_ (.A(_0470_),
    .B(_0568_),
    .Y(_0746_));
 sky130_fd_sc_hd__nor2_1 _1680_ (.A(_0178_),
    .B(_0665_),
    .Y(_0747_));
 sky130_fd_sc_hd__mux4_1 _1681_ (.A0(_0048_),
    .A1(_0051_),
    .A2(_0047_),
    .A3(_0050_),
    .S0(_0083_),
    .S1(_0286_),
    .X(_0748_));
 sky130_fd_sc_hd__nor2_1 _1682_ (.A(_0320_),
    .B(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__o21ai_1 _1683_ (.A1(_0747_),
    .A2(_0749_),
    .B1(_0391_),
    .Y(_0750_));
 sky130_fd_sc_hd__nor2_1 _1684_ (.A(_0170_),
    .B(_0264_),
    .Y(_0751_));
 sky130_fd_sc_hd__a31oi_2 _1685_ (.A1(_0170_),
    .A2(_0746_),
    .A3(_0750_),
    .B1(_0751_),
    .Y(_0752_));
 sky130_fd_sc_hd__nand2_1 _1686_ (.A(_0254_),
    .B(_0701_),
    .Y(_0753_));
 sky130_fd_sc_hd__nand2_2 _1687_ (.A(_0034_),
    .B(_0181_),
    .Y(_0754_));
 sky130_fd_sc_hd__nor2_1 _1688_ (.A(_0754_),
    .B(_0300_),
    .Y(_0755_));
 sky130_fd_sc_hd__a211oi_1 _1689_ (.A1(_0148_),
    .A2(_0283_),
    .B1(_0755_),
    .C1(_0042_),
    .Y(_0756_));
 sky130_fd_sc_hd__nor2_1 _1690_ (.A(_0329_),
    .B(_0677_),
    .Y(_0757_));
 sky130_fd_sc_hd__nor2_1 _1691_ (.A(_0920_),
    .B(_0733_),
    .Y(_0758_));
 sky130_fd_sc_hd__mux2i_2 _1692_ (.A0(_0048_),
    .A1(_0047_),
    .S(_0847_),
    .Y(_0759_));
 sky130_fd_sc_hd__nor2_1 _1693_ (.A(_0195_),
    .B(_0759_),
    .Y(_0760_));
 sky130_fd_sc_hd__nand2_1 _1694_ (.A(_0651_),
    .B(_0558_),
    .Y(_0761_));
 sky130_fd_sc_hd__o31ai_1 _1695_ (.A1(_0651_),
    .A2(_0758_),
    .A3(_0760_),
    .B1(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__nor2_1 _1696_ (.A(_0114_),
    .B(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__o21ai_1 _1697_ (.A1(_0757_),
    .A2(_0763_),
    .B1(_0191_),
    .Y(_0764_));
 sky130_fd_sc_hd__a32oi_1 _1698_ (.A1(_0213_),
    .A2(_0752_),
    .A3(_0753_),
    .B1(_0756_),
    .B2(_0764_),
    .Y(net55));
 sky130_fd_sc_hd__o31ai_1 _1699_ (.A1(_0320_),
    .A2(_0062_),
    .A3(_0754_),
    .B1(_0629_),
    .Y(_0766_));
 sky130_fd_sc_hd__a21oi_1 _1700_ (.A1(_0148_),
    .A2(_0319_),
    .B1(_0766_),
    .Y(_0767_));
 sky130_fd_sc_hd__nor2_1 _1701_ (.A(_0329_),
    .B(_0691_),
    .Y(_0768_));
 sky130_fd_sc_hd__nor2_1 _1702_ (.A(_0246_),
    .B(_0606_),
    .Y(_0769_));
 sky130_fd_sc_hd__mux2i_2 _1703_ (.A0(_0058_),
    .A1(_0051_),
    .S(_0847_),
    .Y(_0770_));
 sky130_fd_sc_hd__mux2i_4 _1704_ (.A0(_0759_),
    .A1(_0770_),
    .S(_0920_),
    .Y(_0771_));
 sky130_fd_sc_hd__nor2_1 _1705_ (.A(_0265_),
    .B(_0771_),
    .Y(_0772_));
 sky130_fd_sc_hd__nor3_1 _1706_ (.A(_0114_),
    .B(_0769_),
    .C(_0772_),
    .Y(_0773_));
 sky130_fd_sc_hd__o21ai_1 _1707_ (.A1(_0768_),
    .A2(_0773_),
    .B1(_0191_),
    .Y(_0774_));
 sky130_fd_sc_hd__nor2_1 _1708_ (.A(_0030_),
    .B(_0038_),
    .Y(_0776_));
 sky130_fd_sc_hd__nor2_1 _1709_ (.A(_0075_),
    .B(_0706_),
    .Y(_0777_));
 sky130_fd_sc_hd__mux4_1 _1710_ (.A0(_0058_),
    .A1(_0048_),
    .A2(_0051_),
    .A3(_0047_),
    .S0(_0083_),
    .S1(_0286_),
    .X(_0778_));
 sky130_fd_sc_hd__nor2_1 _1711_ (.A(_0064_),
    .B(_0778_),
    .Y(_0779_));
 sky130_fd_sc_hd__nand2_1 _1712_ (.A(_0258_),
    .B(_0618_),
    .Y(_0780_));
 sky130_fd_sc_hd__o311a_1 _1713_ (.A1(_0045_),
    .A2(_0777_),
    .A3(_0779_),
    .B1(_0780_),
    .C1(_0034_),
    .X(_0781_));
 sky130_fd_sc_hd__a21oi_1 _1714_ (.A1(_0257_),
    .A2(_0344_),
    .B1(_0781_),
    .Y(_0782_));
 sky130_fd_sc_hd__a211oi_1 _1715_ (.A1(_0776_),
    .A2(_0161_),
    .B1(_0782_),
    .C1(_0629_),
    .Y(_0783_));
 sky130_fd_sc_hd__a21oi_1 _1716_ (.A1(_0767_),
    .A2(_0774_),
    .B1(_0783_),
    .Y(net56));
 sky130_fd_sc_hd__mux4_1 _1717_ (.A0(_0055_),
    .A1(_0058_),
    .A2(_0048_),
    .A3(_0051_),
    .S0(_0775_),
    .S1(_0138_),
    .X(_0784_));
 sky130_fd_sc_hd__nor2_1 _1718_ (.A(_0113_),
    .B(_0784_),
    .Y(_0786_));
 sky130_fd_sc_hd__a211oi_1 _1719_ (.A1(_0144_),
    .A2(_0723_),
    .B1(_0786_),
    .C1(_0651_),
    .Y(_0787_));
 sky130_fd_sc_hd__a21oi_1 _1720_ (.A1(_0265_),
    .A2(_0637_),
    .B1(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__o22a_1 _1721_ (.A1(_0589_),
    .A2(_0381_),
    .B1(_0788_),
    .B2(_0038_),
    .X(_0789_));
 sky130_fd_sc_hd__nor2_1 _1722_ (.A(_0320_),
    .B(_0754_),
    .Y(_0790_));
 sky130_fd_sc_hd__a21oi_1 _1723_ (.A1(_0790_),
    .A2(_0393_),
    .B1(_0213_),
    .Y(_0791_));
 sky130_fd_sc_hd__mux4_1 _1724_ (.A0(_0055_),
    .A1(net21),
    .A2(_0048_),
    .A3(_0051_),
    .S0(_0096_),
    .S1(_0097_),
    .X(_0792_));
 sky130_fd_sc_hd__and2_0 _1725_ (.A(_0101_),
    .B(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__a211oi_1 _1726_ (.A1(_0087_),
    .A2(_0714_),
    .B1(_0793_),
    .C1(_0258_),
    .Y(_0794_));
 sky130_fd_sc_hd__a211oi_1 _1727_ (.A1(_0046_),
    .A2(_0623_),
    .B1(_0794_),
    .C1(_0043_),
    .Y(_0795_));
 sky130_fd_sc_hd__nor3_1 _1728_ (.A(_0144_),
    .B(_0357_),
    .C(_0602_),
    .Y(_0797_));
 sky130_fd_sc_hd__a2111oi_0 _1729_ (.A1(_0257_),
    .A2(_0372_),
    .B1(_0795_),
    .C1(_0797_),
    .D1(_0629_),
    .Y(_0798_));
 sky130_fd_sc_hd__a21oi_1 _1730_ (.A1(_0789_),
    .A2(_0791_),
    .B1(_0798_),
    .Y(net57));
 sky130_fd_sc_hd__a21oi_1 _1731_ (.A1(_0438_),
    .A2(_0790_),
    .B1(_0629_),
    .Y(_0799_));
 sky130_fd_sc_hd__mux2i_1 _1732_ (.A0(_0089_),
    .A1(_0080_),
    .S(_0837_),
    .Y(_0800_));
 sky130_fd_sc_hd__nand2b_1 _1733_ (.A_N(_0079_),
    .B(_0133_),
    .Y(_0801_));
 sky130_fd_sc_hd__o211ai_1 _1734_ (.A1(_0088_),
    .A2(_0138_),
    .B1(_0801_),
    .C1(_0120_),
    .Y(_0802_));
 sky130_fd_sc_hd__o21ai_0 _1735_ (.A1(_0120_),
    .A2(_0800_),
    .B1(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__mux4_1 _1736_ (.A0(_0081_),
    .A1(_0082_),
    .A2(_0117_),
    .A3(_0115_),
    .S0(_0207_),
    .S1(_0837_),
    .X(_0804_));
 sky130_fd_sc_hd__mux4_1 _1737_ (.A0(_0219_),
    .A1(_0242_),
    .A2(_0803_),
    .A3(_0804_),
    .S0(_0143_),
    .S1(_0272_),
    .X(_0805_));
 sky130_fd_sc_hd__a22oi_1 _1738_ (.A1(_0148_),
    .A2(_0540_),
    .B1(_0805_),
    .B2(_0111_),
    .Y(_0807_));
 sky130_fd_sc_hd__mux2i_1 _1739_ (.A0(_0082_),
    .A1(_0115_),
    .S(_0060_),
    .Y(_0808_));
 sky130_fd_sc_hd__mux2i_1 _1740_ (.A0(_0575_),
    .A1(_0808_),
    .S(_0208_),
    .Y(_0809_));
 sky130_fd_sc_hd__mux4_1 _1741_ (.A0(_0088_),
    .A1(_0089_),
    .A2(net26),
    .A3(_0080_),
    .S0(_0072_),
    .S1(_0745_),
    .X(_0810_));
 sky130_fd_sc_hd__mux4_1 _1742_ (.A0(_0175_),
    .A1(_0176_),
    .A2(_0809_),
    .A3(_0810_),
    .S0(_0101_),
    .S1(_0180_),
    .X(_0811_));
 sky130_fd_sc_hd__nand2_1 _1743_ (.A(_0034_),
    .B(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__o21ai_0 _1744_ (.A1(_0034_),
    .A2(_0550_),
    .B1(_0812_),
    .Y(_0813_));
 sky130_fd_sc_hd__a211oi_1 _1745_ (.A1(_0776_),
    .A2(_0209_),
    .B1(_0813_),
    .C1(_0213_),
    .Y(_0814_));
 sky130_fd_sc_hd__a21oi_1 _1746_ (.A1(_0799_),
    .A2(_0807_),
    .B1(_0814_),
    .Y(net58));
 sky130_fd_sc_hd__mux4_1 _1747_ (.A0(_0059_),
    .A1(_0055_),
    .A2(_0058_),
    .A3(_0048_),
    .S0(_0775_),
    .S1(_0090_),
    .X(_0815_));
 sky130_fd_sc_hd__mux2i_1 _1748_ (.A0(_0740_),
    .A1(_0815_),
    .S(_0075_),
    .Y(_0817_));
 sky130_fd_sc_hd__mux4_1 _1749_ (.A0(_0439_),
    .A1(_0442_),
    .A2(_0648_),
    .A3(_0817_),
    .S0(_0180_),
    .S1(_0034_),
    .X(_0818_));
 sky130_fd_sc_hd__nand2_1 _1750_ (.A(_0039_),
    .B(_0412_),
    .Y(_0819_));
 sky130_fd_sc_hd__mux4_1 _1751_ (.A0(_0059_),
    .A1(_0055_),
    .A2(_0058_),
    .A3(_0048_),
    .S0(_0207_),
    .S1(_0837_),
    .X(_0820_));
 sky130_fd_sc_hd__nor2_1 _1752_ (.A(_0221_),
    .B(_0820_),
    .Y(_0821_));
 sky130_fd_sc_hd__a211oi_1 _1753_ (.A1(_0113_),
    .A2(_0735_),
    .B1(_0821_),
    .C1(_0651_),
    .Y(_0822_));
 sky130_fd_sc_hd__a21oi_1 _1754_ (.A1(_0194_),
    .A2(_0661_),
    .B1(_0822_),
    .Y(_0823_));
 sky130_fd_sc_hd__o221ai_1 _1755_ (.A1(_0032_),
    .A2(_0187_),
    .B1(_0823_),
    .B2(_0038_),
    .C1(_0629_),
    .Y(_0824_));
 sky130_fd_sc_hd__a21oi_1 _1756_ (.A1(_0148_),
    .A2(_0410_),
    .B1(_0824_),
    .Y(_0825_));
 sky130_fd_sc_hd__a31oi_2 _1757_ (.A1(_0213_),
    .A2(_0818_),
    .A3(_0819_),
    .B1(_0825_),
    .Y(net59));
 sky130_fd_sc_hd__a31oi_1 _1758_ (.A1(_0316_),
    .A2(_0697_),
    .A3(_0250_),
    .B1(_0042_),
    .Y(_0827_));
 sky130_fd_sc_hd__nor2_1 _1759_ (.A(_0329_),
    .B(_0762_),
    .Y(_0828_));
 sky130_fd_sc_hd__nor2_1 _1760_ (.A(_0246_),
    .B(_0676_),
    .Y(_0829_));
 sky130_fd_sc_hd__mux4_1 _1761_ (.A0(_0056_),
    .A1(_0059_),
    .A2(_0055_),
    .A3(_0058_),
    .S0(_0208_),
    .S1(_0847_),
    .X(_0830_));
 sky130_fd_sc_hd__nor2_1 _1762_ (.A(_0194_),
    .B(_0830_),
    .Y(_0831_));
 sky130_fd_sc_hd__nor3_1 _1763_ (.A(_0114_),
    .B(_0829_),
    .C(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__o21ai_2 _1764_ (.A1(_0828_),
    .A2(_0832_),
    .B1(_0111_),
    .Y(_0833_));
 sky130_fd_sc_hd__nand2_1 _1765_ (.A(_0148_),
    .B(_0468_),
    .Y(_0834_));
 sky130_fd_sc_hd__nand2_1 _1766_ (.A(_0066_),
    .B(_0666_),
    .Y(_0835_));
 sky130_fd_sc_hd__nor2_1 _1767_ (.A(_0231_),
    .B(_0748_),
    .Y(_0836_));
 sky130_fd_sc_hd__mux4_1 _1768_ (.A0(_0056_),
    .A1(_0059_),
    .A2(_0055_),
    .A3(_0058_),
    .S0(_0775_),
    .S1(_0090_),
    .X(_0838_));
 sky130_fd_sc_hd__nor2_1 _1769_ (.A(_0087_),
    .B(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hd__o21ai_0 _1770_ (.A1(_0836_),
    .A2(_0839_),
    .B1(_0181_),
    .Y(_0840_));
 sky130_fd_sc_hd__a21oi_1 _1771_ (.A1(_0835_),
    .A2(_0840_),
    .B1(_0043_),
    .Y(_0841_));
 sky130_fd_sc_hd__a21oi_1 _1772_ (.A1(_0257_),
    .A2(_0461_),
    .B1(_0841_),
    .Y(_0842_));
 sky130_fd_sc_hd__a211oi_1 _1773_ (.A1(_0039_),
    .A2(_0250_),
    .B1(_0842_),
    .C1(_0629_),
    .Y(_0843_));
 sky130_fd_sc_hd__a31oi_2 _1774_ (.A1(_0827_),
    .A2(_0833_),
    .A3(_0834_),
    .B1(_0843_),
    .Y(net60));
 sky130_fd_sc_hd__mux2i_1 _1775_ (.A0(_0292_),
    .A1(_0300_),
    .S(_0031_),
    .Y(_0844_));
 sky130_fd_sc_hd__nor3_1 _1776_ (.A(_0030_),
    .B(_0037_),
    .C(_0276_),
    .Y(_0845_));
 sky130_fd_sc_hd__or2_0 _1777_ (.A(_0286_),
    .B(_0117_),
    .X(_0846_));
 sky130_fd_sc_hd__o211ai_1 _1778_ (.A1(_0921_),
    .A2(_0118_),
    .B1(_0846_),
    .C1(_0195_),
    .Y(_0848_));
 sky130_fd_sc_hd__o21ai_2 _1779_ (.A1(_0195_),
    .A2(_0808_),
    .B1(_0848_),
    .Y(_0849_));
 sky130_fd_sc_hd__mux4_1 _1780_ (.A0(_0089_),
    .A1(_0079_),
    .A2(_0080_),
    .A3(_0081_),
    .S0(_0124_),
    .S1(_0090_),
    .X(_0850_));
 sky130_fd_sc_hd__mux2i_2 _1781_ (.A0(_0849_),
    .A1(_0850_),
    .S(_0178_),
    .Y(_0851_));
 sky130_fd_sc_hd__nand2_1 _1782_ (.A(_0189_),
    .B(_0289_),
    .Y(_0852_));
 sky130_fd_sc_hd__o21ai_0 _1783_ (.A1(_0754_),
    .A2(_0851_),
    .B1(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__a2111oi_0 _1784_ (.A1(_0415_),
    .A2(_0844_),
    .B1(_0845_),
    .C1(_0167_),
    .D1(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__nor2_1 _1785_ (.A(_0272_),
    .B(_0249_),
    .Y(_0855_));
 sky130_fd_sc_hd__nor2_1 _1786_ (.A(_0120_),
    .B(_0140_),
    .Y(_0856_));
 sky130_fd_sc_hd__nor2_1 _1787_ (.A(_0295_),
    .B(_0800_),
    .Y(_0857_));
 sky130_fd_sc_hd__mux4_1 _1788_ (.A0(_0082_),
    .A1(net30),
    .A2(_0115_),
    .A3(_0118_),
    .S0(_0072_),
    .S1(_0217_),
    .X(_0859_));
 sky130_fd_sc_hd__or2_0 _1789_ (.A(_0159_),
    .B(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__o311a_1 _1790_ (.A1(_0143_),
    .A2(_0856_),
    .A3(_0857_),
    .B1(_0860_),
    .C1(_0132_),
    .X(_0861_));
 sky130_fd_sc_hd__o21ai_1 _1791_ (.A1(_0855_),
    .A2(_0861_),
    .B1(_0362_),
    .Y(_0862_));
 sky130_fd_sc_hd__o21ai_1 _1792_ (.A1(_0362_),
    .A2(_0565_),
    .B1(_0862_),
    .Y(_0863_));
 sky130_fd_sc_hd__o31ai_1 _1793_ (.A1(_0320_),
    .A2(_0754_),
    .A3(_0263_),
    .B1(_0042_),
    .Y(_0864_));
 sky130_fd_sc_hd__a21oi_1 _1794_ (.A1(_0215_),
    .A2(_0863_),
    .B1(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__nor2_1 _1795_ (.A(_0854_),
    .B(_0865_),
    .Y(net61));
 sky130_fd_sc_hd__nor2_1 _1796_ (.A(_0178_),
    .B(_0100_),
    .Y(_0866_));
 sky130_fd_sc_hd__nor2_1 _1797_ (.A(_0320_),
    .B(_0085_),
    .Y(_0867_));
 sky130_fd_sc_hd__nor2_1 _1798_ (.A(_0866_),
    .B(_0867_),
    .Y(_0869_));
 sky130_fd_sc_hd__nor2_1 _1799_ (.A(_0470_),
    .B(_0869_),
    .Y(_0870_));
 sky130_fd_sc_hd__a21oi_1 _1800_ (.A1(_0415_),
    .A2(_0324_),
    .B1(_0870_),
    .Y(_0871_));
 sky130_fd_sc_hd__o221ai_1 _1801_ (.A1(_0062_),
    .A2(_0235_),
    .B1(_0323_),
    .B2(_0415_),
    .C1(_0044_),
    .Y(_0872_));
 sky130_fd_sc_hd__o21ai_0 _1802_ (.A1(_0479_),
    .A2(_0871_),
    .B1(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__a21oi_1 _1803_ (.A1(_0307_),
    .A2(_0609_),
    .B1(_0602_),
    .Y(_0874_));
 sky130_fd_sc_hd__nor2_1 _1804_ (.A(_0042_),
    .B(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__nand2_1 _1805_ (.A(_0148_),
    .B(_0614_),
    .Y(_0876_));
 sky130_fd_sc_hd__mux2i_1 _1806_ (.A0(_0156_),
    .A1(_0122_),
    .S(_0132_),
    .Y(_0877_));
 sky130_fd_sc_hd__o211ai_1 _1807_ (.A1(_0272_),
    .A2(_0137_),
    .B1(_0142_),
    .C1(_0329_),
    .Y(_0878_));
 sky130_fd_sc_hd__o21ai_1 _1808_ (.A1(_0329_),
    .A2(_0877_),
    .B1(_0878_),
    .Y(_0880_));
 sky130_fd_sc_hd__o21ai_0 _1809_ (.A1(_0754_),
    .A2(_0340_),
    .B1(_0167_),
    .Y(_0881_));
 sky130_fd_sc_hd__a21oi_1 _1810_ (.A1(_0111_),
    .A2(_0880_),
    .B1(_0881_),
    .Y(_0882_));
 sky130_fd_sc_hd__a22oi_1 _1811_ (.A1(_0873_),
    .A2(_0875_),
    .B1(_0876_),
    .B2(_0882_),
    .Y(net62));
 sky130_fd_sc_hd__nor2_1 _1812_ (.A(_0181_),
    .B(_0388_),
    .Y(_0883_));
 sky130_fd_sc_hd__nor2_1 _1813_ (.A(_0231_),
    .B(_0581_),
    .Y(_0884_));
 sky130_fd_sc_hd__nor2_1 _1814_ (.A(_0087_),
    .B(_0576_),
    .Y(_0885_));
 sky130_fd_sc_hd__nor3_1 _1815_ (.A(_0258_),
    .B(_0884_),
    .C(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__nor3_1 _1816_ (.A(_0043_),
    .B(_0883_),
    .C(_0886_),
    .Y(_0887_));
 sky130_fd_sc_hd__a21oi_2 _1817_ (.A1(_0257_),
    .A2(_0641_),
    .B1(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__nor2_1 _1818_ (.A(_0631_),
    .B(_0602_),
    .Y(_0890_));
 sky130_fd_sc_hd__mux2i_1 _1819_ (.A0(_0360_),
    .A1(_0596_),
    .S(_0131_),
    .Y(_0891_));
 sky130_fd_sc_hd__nand2b_1 _1820_ (.A_N(_0891_),
    .B(_0113_),
    .Y(_0892_));
 sky130_fd_sc_hd__o211ai_2 _1821_ (.A1(_0114_),
    .A2(_0594_),
    .B1(_0892_),
    .C1(_0111_),
    .Y(_0893_));
 sky130_fd_sc_hd__nand2_1 _1822_ (.A(_0148_),
    .B(_0628_),
    .Y(_0894_));
 sky130_fd_sc_hd__o2111ai_1 _1823_ (.A1(_0754_),
    .A2(_0368_),
    .B1(_0893_),
    .C1(_0894_),
    .D1(_0042_),
    .Y(_0895_));
 sky130_fd_sc_hd__o31a_1 _1824_ (.A1(_0327_),
    .A2(_0888_),
    .A3(_0890_),
    .B1(_0895_),
    .X(net63));
 sky130_fd_sc_hd__mux2i_1 _1825_ (.A0(_0176_),
    .A1(_0809_),
    .S(_0178_),
    .Y(_0896_));
 sky130_fd_sc_hd__nand2_1 _1826_ (.A(_0470_),
    .B(_0418_),
    .Y(_0897_));
 sky130_fd_sc_hd__o21ai_0 _1827_ (.A1(_0470_),
    .A2(_0896_),
    .B1(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__o211ai_1 _1828_ (.A1(_0406_),
    .A2(_0602_),
    .B1(_0044_),
    .C1(_0629_),
    .Y(_0900_));
 sky130_fd_sc_hd__o32ai_1 _1829_ (.A1(_0479_),
    .A2(_0167_),
    .A3(_0898_),
    .B1(_0900_),
    .B2(_0646_),
    .Y(_0901_));
 sky130_fd_sc_hd__nor2_1 _1830_ (.A(_0272_),
    .B(_0424_),
    .Y(_0902_));
 sky130_fd_sc_hd__nor2_1 _1831_ (.A(_0237_),
    .B(_0219_),
    .Y(_0903_));
 sky130_fd_sc_hd__nor2_1 _1832_ (.A(_0113_),
    .B(_0804_),
    .Y(_0904_));
 sky130_fd_sc_hd__nor3_1 _1833_ (.A(_0651_),
    .B(_0903_),
    .C(_0904_),
    .Y(_0905_));
 sky130_fd_sc_hd__o21ai_0 _1834_ (.A1(_0902_),
    .A2(_0905_),
    .B1(_0362_),
    .Y(_0906_));
 sky130_fd_sc_hd__o21ai_1 _1835_ (.A1(_0362_),
    .A2(_0653_),
    .B1(_0906_),
    .Y(_0907_));
 sky130_fd_sc_hd__o21ai_0 _1836_ (.A1(_0754_),
    .A2(_0439_),
    .B1(_0327_),
    .Y(_0908_));
 sky130_fd_sc_hd__a21oi_1 _1837_ (.A1(_0215_),
    .A2(_0907_),
    .B1(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__nor2_1 _1838_ (.A(_0901_),
    .B(_0909_),
    .Y(net64));
 sky130_fd_sc_hd__nand2_1 _1839_ (.A(_0697_),
    .B(_0457_),
    .Y(_0911_));
 sky130_fd_sc_hd__nor2_1 _1840_ (.A(_0237_),
    .B(_0248_),
    .Y(_0912_));
 sky130_fd_sc_hd__nor2_1 _1841_ (.A(_0113_),
    .B(_0859_),
    .Y(_0913_));
 sky130_fd_sc_hd__nand2_1 _1842_ (.A(_0194_),
    .B(_0452_),
    .Y(_0914_));
 sky130_fd_sc_hd__o311ai_2 _1843_ (.A1(_0651_),
    .A2(_0912_),
    .A3(_0913_),
    .B1(_0914_),
    .C1(_0362_),
    .Y(_0915_));
 sky130_fd_sc_hd__o211ai_1 _1844_ (.A1(_0362_),
    .A2(_0686_),
    .B1(_0915_),
    .C1(_0215_),
    .Y(_0916_));
 sky130_fd_sc_hd__mux2i_2 _1845_ (.A0(_0291_),
    .A1(_0849_),
    .S(_0178_),
    .Y(_0917_));
 sky130_fd_sc_hd__nor3_1 _1846_ (.A(_0031_),
    .B(_0181_),
    .C(_0473_),
    .Y(_0918_));
 sky130_fd_sc_hd__a221oi_2 _1847_ (.A1(_0043_),
    .A2(_0669_),
    .B1(_0917_),
    .B2(_0697_),
    .C1(_0918_),
    .Y(_0919_));
 sky130_fd_sc_hd__nor2_1 _1848_ (.A(_0466_),
    .B(_0602_),
    .Y(_0001_));
 sky130_fd_sc_hd__nor3_1 _1849_ (.A(_0042_),
    .B(_0919_),
    .C(_0001_),
    .Y(_0002_));
 sky130_fd_sc_hd__a31oi_2 _1850_ (.A1(_0213_),
    .A2(_0911_),
    .A3(_0916_),
    .B1(_0002_),
    .Y(net65));
 sky130_fd_sc_hd__nor2_1 _1851_ (.A(_0129_),
    .B(_0153_),
    .Y(_0003_));
 sky130_fd_sc_hd__nor2_1 _1852_ (.A(_0193_),
    .B(_0137_),
    .Y(_0004_));
 sky130_fd_sc_hd__o21ai_1 _1853_ (.A1(_0003_),
    .A2(_0004_),
    .B1(_0144_),
    .Y(_0005_));
 sky130_fd_sc_hd__nand2b_1 _1854_ (.A_N(_0156_),
    .B(_0210_),
    .Y(_0006_));
 sky130_fd_sc_hd__o2111ai_4 _1855_ (.A1(_0030_),
    .A2(_0122_),
    .B1(_0005_),
    .C1(_0006_),
    .D1(_0111_),
    .Y(_0007_));
 sky130_fd_sc_hd__nand3_1 _1856_ (.A(_0246_),
    .B(_0163_),
    .C(_0147_),
    .Y(_0008_));
 sky130_fd_sc_hd__o2111ai_1 _1857_ (.A1(_0044_),
    .A2(_0703_),
    .B1(_0007_),
    .C1(_0008_),
    .D1(_0327_),
    .Y(_0009_));
 sky130_fd_sc_hd__nand2_1 _1858_ (.A(_0470_),
    .B(_0076_),
    .Y(_0011_));
 sky130_fd_sc_hd__o21ai_1 _1859_ (.A1(_0470_),
    .A2(_0102_),
    .B1(_0011_),
    .Y(_0012_));
 sky130_fd_sc_hd__nor3_1 _1860_ (.A(_0482_),
    .B(_0485_),
    .C(_0602_),
    .Y(_0013_));
 sky130_fd_sc_hd__o21ai_0 _1861_ (.A1(_0037_),
    .A2(_0698_),
    .B1(_0434_),
    .Y(_0014_));
 sky130_fd_sc_hd__a211oi_1 _1862_ (.A1(_0065_),
    .A2(_0189_),
    .B1(_0013_),
    .C1(_0014_),
    .Y(_0015_));
 sky130_fd_sc_hd__o21ai_0 _1863_ (.A1(_0044_),
    .A2(_0012_),
    .B1(_0015_),
    .Y(_0016_));
 sky130_fd_sc_hd__and2_0 _1864_ (.A(_0009_),
    .B(_0016_),
    .X(net66));
 sky130_fd_sc_hd__nand3_1 _1865_ (.A(_0272_),
    .B(_0147_),
    .C(_0518_),
    .Y(_0017_));
 sky130_fd_sc_hd__nand2_1 _1866_ (.A(_0193_),
    .B(_0348_),
    .Y(_0018_));
 sky130_fd_sc_hd__nand2_1 _1867_ (.A(_0129_),
    .B(_0354_),
    .Y(_0019_));
 sky130_fd_sc_hd__nand4_1 _1868_ (.A(_0110_),
    .B(_0144_),
    .C(_0018_),
    .D(_0019_),
    .Y(_0021_));
 sky130_fd_sc_hd__nand2_1 _1869_ (.A(_0017_),
    .B(_0021_),
    .Y(_0022_));
 sky130_fd_sc_hd__and3_1 _1870_ (.A(_0110_),
    .B(_0238_),
    .C(_0891_),
    .X(_0023_));
 sky130_fd_sc_hd__nor2_1 _1871_ (.A(_0022_),
    .B(_0023_),
    .Y(_0024_));
 sky130_fd_sc_hd__nor4_1 _1872_ (.A(_0434_),
    .B(_0712_),
    .C(_0022_),
    .D(_0023_),
    .Y(_0025_));
 sky130_fd_sc_hd__nand2_1 _1873_ (.A(_0046_),
    .B(_0514_),
    .Y(_0026_));
 sky130_fd_sc_hd__o21ai_1 _1874_ (.A1(_0046_),
    .A2(_0583_),
    .B1(_0026_),
    .Y(_0027_));
 sky130_fd_sc_hd__a221oi_1 _1875_ (.A1(_0189_),
    .A2(_0513_),
    .B1(_0729_),
    .B2(_0110_),
    .C1(_0041_),
    .Y(_0028_));
 sky130_fd_sc_hd__o21a_1 _1876_ (.A1(_0044_),
    .A2(_0027_),
    .B1(_0028_),
    .X(_0029_));
 sky130_fd_sc_hd__a311oi_1 _1877_ (.A1(_0479_),
    .A2(_0042_),
    .A3(_0024_),
    .B1(_0025_),
    .C1(_0029_),
    .Y(net67));
 sky130_fd_sc_hd__ha_2 _1878_ (.A(_0920_),
    .B(_0921_),
    .COUT(_0922_),
    .SUM(_0923_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_171 ();
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(data_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(data_in[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(data_in[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input4 (.A(data_in[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(data_in[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(data_in[14]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(data_in[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(data_in[16]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(data_in[17]),
    .X(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(data_in[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(data_in[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(data_in[1]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(data_in[20]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(data_in[21]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(data_in[22]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(data_in[23]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(data_in[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(data_in[25]),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(data_in[26]),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 input20 (.A(data_in[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(data_in[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(data_in[29]),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(data_in[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(data_in[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(data_in[3]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(data_in[4]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(data_in[5]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(data_in[6]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(data_in[7]),
    .X(net29));
 sky130_fd_sc_hd__dlymetal6s2s_1 input30 (.A(data_in[8]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(data_in[9]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input32 (.A(rotate),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(shift_amount[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input34 (.A(shift_amount[1]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 input35 (.A(shift_amount[2]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net36),
    .X(data_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(net37),
    .X(data_out[10]));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net38),
    .X(data_out[11]));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(net39),
    .X(data_out[12]));
 sky130_fd_sc_hd__clkbuf_1 output40 (.A(net40),
    .X(data_out[13]));
 sky130_fd_sc_hd__clkbuf_1 output41 (.A(net41),
    .X(data_out[14]));
 sky130_fd_sc_hd__clkbuf_1 output42 (.A(net42),
    .X(data_out[15]));
 sky130_fd_sc_hd__clkbuf_1 output43 (.A(net43),
    .X(data_out[16]));
 sky130_fd_sc_hd__clkbuf_1 output44 (.A(net44),
    .X(data_out[17]));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(net45),
    .X(data_out[18]));
 sky130_fd_sc_hd__clkbuf_1 output46 (.A(net46),
    .X(data_out[19]));
 sky130_fd_sc_hd__clkbuf_1 output47 (.A(net47),
    .X(data_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output48 (.A(net48),
    .X(data_out[20]));
 sky130_fd_sc_hd__clkbuf_1 output49 (.A(net49),
    .X(data_out[21]));
 sky130_fd_sc_hd__clkbuf_1 output50 (.A(net50),
    .X(data_out[22]));
 sky130_fd_sc_hd__clkbuf_1 output51 (.A(net51),
    .X(data_out[23]));
 sky130_fd_sc_hd__clkbuf_1 output52 (.A(net52),
    .X(data_out[24]));
 sky130_fd_sc_hd__clkbuf_1 output53 (.A(net53),
    .X(data_out[25]));
 sky130_fd_sc_hd__clkbuf_1 output54 (.A(net54),
    .X(data_out[26]));
 sky130_fd_sc_hd__clkbuf_1 output55 (.A(net55),
    .X(data_out[27]));
 sky130_fd_sc_hd__clkbuf_1 output56 (.A(net56),
    .X(data_out[28]));
 sky130_fd_sc_hd__clkbuf_1 output57 (.A(net57),
    .X(data_out[29]));
 sky130_fd_sc_hd__clkbuf_1 output58 (.A(net58),
    .X(data_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output59 (.A(net59),
    .X(data_out[30]));
 sky130_fd_sc_hd__clkbuf_1 output60 (.A(net60),
    .X(data_out[31]));
 sky130_fd_sc_hd__clkbuf_1 output61 (.A(net61),
    .X(data_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output62 (.A(net62),
    .X(data_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output63 (.A(net63),
    .X(data_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output64 (.A(net64),
    .X(data_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output65 (.A(net65),
    .X(data_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net66),
    .X(data_out[8]));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net67),
    .X(data_out[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0161_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0161_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(data_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(data_in[13]));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_126 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_234 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_224 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_234 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_241 ();
endmodule
