module smart_fifo (almost_empty,
    almost_full,
    clear_errors,
    clk,
    empty,
    error_detected,
    full,
    overflow_detected,
    rd_en,
    rd_valid,
    rst_n,
    underflow_detected,
    wr_en,
    wr_ready,
    data_count,
    error_count,
    rd_data,
    wr_data);
 output almost_empty;
 output almost_full;
 input clear_errors;
 input clk;
 output empty;
 output error_detected;
 output full;
 output overflow_detected;
 input rd_en;
 output rd_valid;
 input rst_n;
 output underflow_detected;
 input wr_en;
 output wr_ready;
 output [4:0] data_count;
 output [15:0] error_count;
 output [31:0] rd_data;
 input [31:0] wr_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire _0629_;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire _0633_;
 wire clknet_3_0__leaf_clk;
 wire _0635_;
 wire _0636_;
 wire clknet_0_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_11_clk;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_7_clk;
 wire _0711_;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_4_clk;
 wire _0715_;
 wire _0716_;
 wire clknet_leaf_3_clk;
 wire _0718_;
 wire net207;
 wire net206;
 wire net201;
 wire net198;
 wire _0723_;
 wire net197;
 wire net173;
 wire net172;
 wire _0727_;
 wire clknet_leaf_0_clk;
 wire net210;
 wire net178;
 wire _0731_;
 wire net174;
 wire net209;
 wire net204;
 wire _0735_;
 wire net203;
 wire net192;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_1_clk;
 wire _0740_;
 wire net208;
 wire net205;
 wire net200;
 wire net199;
 wire _0745_;
 wire net196;
 wire net195;
 wire net194;
 wire net202;
 wire _0750_;
 wire _0751_;
 wire net191;
 wire net190;
 wire net189;
 wire net188;
 wire _0756_;
 wire net187;
 wire net186;
 wire net185;
 wire net184;
 wire _0761_;
 wire net183;
 wire net182;
 wire net181;
 wire net180;
 wire _0766_;
 wire net179;
 wire net177;
 wire net193;
 wire net176;
 wire _0771_;
 wire net175;
 wire _0775_;
 wire _0780_;
 wire _0782_;
 wire _0783_;
 wire _0785_;
 wire _0787_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0801_;
 wire _0802_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0809_;
 wire _0810_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0872_;
 wire _0873_;
 wire _0877_;
 wire _0880_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0902_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0910_;
 wire _0913_;
 wire _0916_;
 wire _0917_;
 wire _0920_;
 wire _0922_;
 wire _0924_;
 wire _0926_;
 wire _0928_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1028_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1067_;
 wire _1068_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire net36;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire net35;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire net34;
 wire _1105_;
 wire net33;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire net32;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire net31;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire net30;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire net29;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire net28;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire net27;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire net26;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire net25;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire net24;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire net23;
 wire _1219_;
 wire net22;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire net21;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire net20;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire net19;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire net18;
 wire _1258_;
 wire _1259_;
 wire net17;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire net16;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire net15;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire net14;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire net13;
 wire _1296_;
 wire net12;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire net11;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire net10;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire net9;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire net8;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire net7;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire net6;
 wire _1530_;
 wire net5;
 wire _1532_;
 wire _1533_;
 wire net4;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire net3;
 wire _1553_;
 wire net2;
 wire _1555_;
 wire _1556_;
 wire net1;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire \last_valid_data[0] ;
 wire \last_valid_data[10] ;
 wire \last_valid_data[11] ;
 wire \last_valid_data[12] ;
 wire \last_valid_data[13] ;
 wire \last_valid_data[14] ;
 wire \last_valid_data[15] ;
 wire \last_valid_data[16] ;
 wire \last_valid_data[17] ;
 wire \last_valid_data[18] ;
 wire \last_valid_data[19] ;
 wire \last_valid_data[1] ;
 wire \last_valid_data[20] ;
 wire \last_valid_data[21] ;
 wire \last_valid_data[22] ;
 wire \last_valid_data[23] ;
 wire \last_valid_data[24] ;
 wire \last_valid_data[25] ;
 wire \last_valid_data[26] ;
 wire \last_valid_data[27] ;
 wire \last_valid_data[28] ;
 wire \last_valid_data[29] ;
 wire \last_valid_data[2] ;
 wire \last_valid_data[30] ;
 wire \last_valid_data[31] ;
 wire \last_valid_data[3] ;
 wire \last_valid_data[4] ;
 wire \last_valid_data[5] ;
 wire \last_valid_data[6] ;
 wire \last_valid_data[7] ;
 wire \last_valid_data[8] ;
 wire \last_valid_data[9] ;
 wire last_valid_data_available;
 wire \mem[0][0] ;
 wire \mem[0][10] ;
 wire \mem[0][11] ;
 wire \mem[0][12] ;
 wire \mem[0][13] ;
 wire \mem[0][14] ;
 wire \mem[0][15] ;
 wire \mem[0][16] ;
 wire \mem[0][17] ;
 wire \mem[0][18] ;
 wire \mem[0][19] ;
 wire \mem[0][1] ;
 wire \mem[0][20] ;
 wire \mem[0][21] ;
 wire \mem[0][22] ;
 wire \mem[0][23] ;
 wire \mem[0][24] ;
 wire \mem[0][25] ;
 wire \mem[0][26] ;
 wire \mem[0][27] ;
 wire \mem[0][28] ;
 wire \mem[0][29] ;
 wire \mem[0][2] ;
 wire \mem[0][30] ;
 wire \mem[0][31] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[0][8] ;
 wire \mem[0][9] ;
 wire \mem[10][0] ;
 wire \mem[10][10] ;
 wire \mem[10][11] ;
 wire \mem[10][12] ;
 wire \mem[10][13] ;
 wire \mem[10][14] ;
 wire \mem[10][15] ;
 wire \mem[10][16] ;
 wire \mem[10][17] ;
 wire \mem[10][18] ;
 wire \mem[10][19] ;
 wire \mem[10][1] ;
 wire \mem[10][20] ;
 wire \mem[10][21] ;
 wire \mem[10][22] ;
 wire \mem[10][23] ;
 wire \mem[10][24] ;
 wire \mem[10][25] ;
 wire \mem[10][26] ;
 wire \mem[10][27] ;
 wire \mem[10][28] ;
 wire \mem[10][29] ;
 wire \mem[10][2] ;
 wire \mem[10][30] ;
 wire \mem[10][31] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[10][8] ;
 wire \mem[10][9] ;
 wire \mem[11][0] ;
 wire \mem[11][10] ;
 wire \mem[11][11] ;
 wire \mem[11][12] ;
 wire \mem[11][13] ;
 wire \mem[11][14] ;
 wire \mem[11][15] ;
 wire \mem[11][16] ;
 wire \mem[11][17] ;
 wire \mem[11][18] ;
 wire \mem[11][19] ;
 wire \mem[11][1] ;
 wire \mem[11][20] ;
 wire \mem[11][21] ;
 wire \mem[11][22] ;
 wire \mem[11][23] ;
 wire \mem[11][24] ;
 wire \mem[11][25] ;
 wire \mem[11][26] ;
 wire \mem[11][27] ;
 wire \mem[11][28] ;
 wire \mem[11][29] ;
 wire \mem[11][2] ;
 wire \mem[11][30] ;
 wire \mem[11][31] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[11][8] ;
 wire \mem[11][9] ;
 wire \mem[12][0] ;
 wire \mem[12][10] ;
 wire \mem[12][11] ;
 wire \mem[12][12] ;
 wire \mem[12][13] ;
 wire \mem[12][14] ;
 wire \mem[12][15] ;
 wire \mem[12][16] ;
 wire \mem[12][17] ;
 wire \mem[12][18] ;
 wire \mem[12][19] ;
 wire \mem[12][1] ;
 wire \mem[12][20] ;
 wire \mem[12][21] ;
 wire \mem[12][22] ;
 wire \mem[12][23] ;
 wire \mem[12][24] ;
 wire \mem[12][25] ;
 wire \mem[12][26] ;
 wire \mem[12][27] ;
 wire \mem[12][28] ;
 wire \mem[12][29] ;
 wire \mem[12][2] ;
 wire \mem[12][30] ;
 wire \mem[12][31] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[12][8] ;
 wire \mem[12][9] ;
 wire \mem[13][0] ;
 wire \mem[13][10] ;
 wire \mem[13][11] ;
 wire \mem[13][12] ;
 wire \mem[13][13] ;
 wire \mem[13][14] ;
 wire \mem[13][15] ;
 wire \mem[13][16] ;
 wire \mem[13][17] ;
 wire \mem[13][18] ;
 wire \mem[13][19] ;
 wire \mem[13][1] ;
 wire \mem[13][20] ;
 wire \mem[13][21] ;
 wire \mem[13][22] ;
 wire \mem[13][23] ;
 wire \mem[13][24] ;
 wire \mem[13][25] ;
 wire \mem[13][26] ;
 wire \mem[13][27] ;
 wire \mem[13][28] ;
 wire \mem[13][29] ;
 wire \mem[13][2] ;
 wire \mem[13][30] ;
 wire \mem[13][31] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[13][8] ;
 wire \mem[13][9] ;
 wire \mem[14][0] ;
 wire \mem[14][10] ;
 wire \mem[14][11] ;
 wire \mem[14][12] ;
 wire \mem[14][13] ;
 wire \mem[14][14] ;
 wire \mem[14][15] ;
 wire \mem[14][16] ;
 wire \mem[14][17] ;
 wire \mem[14][18] ;
 wire \mem[14][19] ;
 wire \mem[14][1] ;
 wire \mem[14][20] ;
 wire \mem[14][21] ;
 wire \mem[14][22] ;
 wire \mem[14][23] ;
 wire \mem[14][24] ;
 wire \mem[14][25] ;
 wire \mem[14][26] ;
 wire \mem[14][27] ;
 wire \mem[14][28] ;
 wire \mem[14][29] ;
 wire \mem[14][2] ;
 wire \mem[14][30] ;
 wire \mem[14][31] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[14][8] ;
 wire \mem[14][9] ;
 wire \mem[15][0] ;
 wire \mem[15][10] ;
 wire \mem[15][11] ;
 wire \mem[15][12] ;
 wire \mem[15][13] ;
 wire \mem[15][14] ;
 wire \mem[15][15] ;
 wire \mem[15][16] ;
 wire \mem[15][17] ;
 wire \mem[15][18] ;
 wire \mem[15][19] ;
 wire \mem[15][1] ;
 wire \mem[15][20] ;
 wire \mem[15][21] ;
 wire \mem[15][22] ;
 wire \mem[15][23] ;
 wire \mem[15][24] ;
 wire \mem[15][25] ;
 wire \mem[15][26] ;
 wire \mem[15][27] ;
 wire \mem[15][28] ;
 wire \mem[15][29] ;
 wire \mem[15][2] ;
 wire \mem[15][30] ;
 wire \mem[15][31] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[15][8] ;
 wire \mem[15][9] ;
 wire \mem[1][0] ;
 wire \mem[1][10] ;
 wire \mem[1][11] ;
 wire \mem[1][12] ;
 wire \mem[1][13] ;
 wire \mem[1][14] ;
 wire \mem[1][15] ;
 wire \mem[1][16] ;
 wire \mem[1][17] ;
 wire \mem[1][18] ;
 wire \mem[1][19] ;
 wire \mem[1][1] ;
 wire \mem[1][20] ;
 wire \mem[1][21] ;
 wire \mem[1][22] ;
 wire \mem[1][23] ;
 wire \mem[1][24] ;
 wire \mem[1][25] ;
 wire \mem[1][26] ;
 wire \mem[1][27] ;
 wire \mem[1][28] ;
 wire \mem[1][29] ;
 wire \mem[1][2] ;
 wire \mem[1][30] ;
 wire \mem[1][31] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[1][8] ;
 wire \mem[1][9] ;
 wire \mem[2][0] ;
 wire \mem[2][10] ;
 wire \mem[2][11] ;
 wire \mem[2][12] ;
 wire \mem[2][13] ;
 wire \mem[2][14] ;
 wire \mem[2][15] ;
 wire \mem[2][16] ;
 wire \mem[2][17] ;
 wire \mem[2][18] ;
 wire \mem[2][19] ;
 wire \mem[2][1] ;
 wire \mem[2][20] ;
 wire \mem[2][21] ;
 wire \mem[2][22] ;
 wire \mem[2][23] ;
 wire \mem[2][24] ;
 wire \mem[2][25] ;
 wire \mem[2][26] ;
 wire \mem[2][27] ;
 wire \mem[2][28] ;
 wire \mem[2][29] ;
 wire \mem[2][2] ;
 wire \mem[2][30] ;
 wire \mem[2][31] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[2][8] ;
 wire \mem[2][9] ;
 wire \mem[3][0] ;
 wire \mem[3][10] ;
 wire \mem[3][11] ;
 wire \mem[3][12] ;
 wire \mem[3][13] ;
 wire \mem[3][14] ;
 wire \mem[3][15] ;
 wire \mem[3][16] ;
 wire \mem[3][17] ;
 wire \mem[3][18] ;
 wire \mem[3][19] ;
 wire \mem[3][1] ;
 wire \mem[3][20] ;
 wire \mem[3][21] ;
 wire \mem[3][22] ;
 wire \mem[3][23] ;
 wire \mem[3][24] ;
 wire \mem[3][25] ;
 wire \mem[3][26] ;
 wire \mem[3][27] ;
 wire \mem[3][28] ;
 wire \mem[3][29] ;
 wire \mem[3][2] ;
 wire \mem[3][30] ;
 wire \mem[3][31] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[3][8] ;
 wire \mem[3][9] ;
 wire \mem[4][0] ;
 wire \mem[4][10] ;
 wire \mem[4][11] ;
 wire \mem[4][12] ;
 wire \mem[4][13] ;
 wire \mem[4][14] ;
 wire \mem[4][15] ;
 wire \mem[4][16] ;
 wire \mem[4][17] ;
 wire \mem[4][18] ;
 wire \mem[4][19] ;
 wire \mem[4][1] ;
 wire \mem[4][20] ;
 wire \mem[4][21] ;
 wire \mem[4][22] ;
 wire \mem[4][23] ;
 wire \mem[4][24] ;
 wire \mem[4][25] ;
 wire \mem[4][26] ;
 wire \mem[4][27] ;
 wire \mem[4][28] ;
 wire \mem[4][29] ;
 wire \mem[4][2] ;
 wire \mem[4][30] ;
 wire \mem[4][31] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[4][8] ;
 wire \mem[4][9] ;
 wire \mem[5][0] ;
 wire \mem[5][10] ;
 wire \mem[5][11] ;
 wire \mem[5][12] ;
 wire \mem[5][13] ;
 wire \mem[5][14] ;
 wire \mem[5][15] ;
 wire \mem[5][16] ;
 wire \mem[5][17] ;
 wire \mem[5][18] ;
 wire \mem[5][19] ;
 wire \mem[5][1] ;
 wire \mem[5][20] ;
 wire \mem[5][21] ;
 wire \mem[5][22] ;
 wire \mem[5][23] ;
 wire \mem[5][24] ;
 wire \mem[5][25] ;
 wire \mem[5][26] ;
 wire \mem[5][27] ;
 wire \mem[5][28] ;
 wire \mem[5][29] ;
 wire \mem[5][2] ;
 wire \mem[5][30] ;
 wire \mem[5][31] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[5][8] ;
 wire \mem[5][9] ;
 wire \mem[6][0] ;
 wire \mem[6][10] ;
 wire \mem[6][11] ;
 wire \mem[6][12] ;
 wire \mem[6][13] ;
 wire \mem[6][14] ;
 wire \mem[6][15] ;
 wire \mem[6][16] ;
 wire \mem[6][17] ;
 wire \mem[6][18] ;
 wire \mem[6][19] ;
 wire \mem[6][1] ;
 wire \mem[6][20] ;
 wire \mem[6][21] ;
 wire \mem[6][22] ;
 wire \mem[6][23] ;
 wire \mem[6][24] ;
 wire \mem[6][25] ;
 wire \mem[6][26] ;
 wire \mem[6][27] ;
 wire \mem[6][28] ;
 wire \mem[6][29] ;
 wire \mem[6][2] ;
 wire \mem[6][30] ;
 wire \mem[6][31] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[6][8] ;
 wire \mem[6][9] ;
 wire \mem[7][0] ;
 wire \mem[7][10] ;
 wire \mem[7][11] ;
 wire \mem[7][12] ;
 wire \mem[7][13] ;
 wire \mem[7][14] ;
 wire \mem[7][15] ;
 wire \mem[7][16] ;
 wire \mem[7][17] ;
 wire \mem[7][18] ;
 wire \mem[7][19] ;
 wire \mem[7][1] ;
 wire \mem[7][20] ;
 wire \mem[7][21] ;
 wire \mem[7][22] ;
 wire \mem[7][23] ;
 wire \mem[7][24] ;
 wire \mem[7][25] ;
 wire \mem[7][26] ;
 wire \mem[7][27] ;
 wire \mem[7][28] ;
 wire \mem[7][29] ;
 wire \mem[7][2] ;
 wire \mem[7][30] ;
 wire \mem[7][31] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[7][8] ;
 wire \mem[7][9] ;
 wire \mem[8][0] ;
 wire \mem[8][10] ;
 wire \mem[8][11] ;
 wire \mem[8][12] ;
 wire \mem[8][13] ;
 wire \mem[8][14] ;
 wire \mem[8][15] ;
 wire \mem[8][16] ;
 wire \mem[8][17] ;
 wire \mem[8][18] ;
 wire \mem[8][19] ;
 wire \mem[8][1] ;
 wire \mem[8][20] ;
 wire \mem[8][21] ;
 wire \mem[8][22] ;
 wire \mem[8][23] ;
 wire \mem[8][24] ;
 wire \mem[8][25] ;
 wire \mem[8][26] ;
 wire \mem[8][27] ;
 wire \mem[8][28] ;
 wire \mem[8][29] ;
 wire \mem[8][2] ;
 wire \mem[8][30] ;
 wire \mem[8][31] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[8][8] ;
 wire \mem[8][9] ;
 wire \mem[9][0] ;
 wire \mem[9][10] ;
 wire \mem[9][11] ;
 wire \mem[9][12] ;
 wire \mem[9][13] ;
 wire \mem[9][14] ;
 wire \mem[9][15] ;
 wire \mem[9][16] ;
 wire \mem[9][17] ;
 wire \mem[9][18] ;
 wire \mem[9][19] ;
 wire \mem[9][1] ;
 wire \mem[9][20] ;
 wire \mem[9][21] ;
 wire \mem[9][22] ;
 wire \mem[9][23] ;
 wire \mem[9][24] ;
 wire \mem[9][25] ;
 wire \mem[9][26] ;
 wire \mem[9][27] ;
 wire \mem[9][28] ;
 wire \mem[9][29] ;
 wire \mem[9][2] ;
 wire \mem[9][30] ;
 wire \mem[9][31] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \mem[9][8] ;
 wire \mem[9][9] ;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire \rd_ptr[0] ;
 wire \rd_ptr[1] ;
 wire \rd_ptr[2] ;
 wire \rd_ptr[3] ;
 wire \rd_ptr[4] ;
 wire net96;
 wire net97;
 wire \wr_ptr[0] ;
 wire \wr_ptr[1] ;
 wire \wr_ptr[2] ;
 wire \wr_ptr[3] ;
 wire \wr_ptr[4] ;
 wire net98;

 CLKBUF_X3 clkload3 (.A(clknet_3_3__leaf_clk));
 INV_X1 _2158_ (.A(_0025_),
    .ZN(net39));
 INV_X2 clkload2 (.A(clknet_3_2__leaf_clk));
 XNOR2_X2 _2160_ (.A(_0009_),
    .B(_0007_),
    .ZN(_0604_));
 INV_X1 _2161_ (.A(_0604_),
    .ZN(net41));
 INV_X1 _2162_ (.A(_0024_),
    .ZN(_0006_));
 AND3_X1 _2163_ (.A1(_0009_),
    .A2(_0006_),
    .A3(_0011_),
    .ZN(_0605_));
 AOI21_X2 _2164_ (.A(_0008_),
    .B1(_0010_),
    .B2(_0009_),
    .ZN(_0606_));
 INV_X1 _2165_ (.A(_0606_),
    .ZN(_0607_));
 OAI21_X1 _2166_ (.A(_0013_),
    .B1(_0605_),
    .B2(_0607_),
    .ZN(_0608_));
 INV_X1 _2167_ (.A(_0013_),
    .ZN(_0609_));
 NAND3_X1 _2168_ (.A1(_0009_),
    .A2(_0006_),
    .A3(_0011_),
    .ZN(_0610_));
 NAND3_X1 _2169_ (.A1(_0609_),
    .A2(_0610_),
    .A3(_0606_),
    .ZN(_0611_));
 NAND2_X1 _2170_ (.A1(_0608_),
    .A2(_0611_),
    .ZN(_0612_));
 INV_X1 _2171_ (.A(_0612_),
    .ZN(net42));
 INV_X1 _2172_ (.A(_0012_),
    .ZN(_0613_));
 AOI21_X1 _2173_ (.A(_0008_),
    .B1(_0007_),
    .B2(_0009_),
    .ZN(_0614_));
 OAI21_X1 _2174_ (.A(_0613_),
    .B1(_0614_),
    .B2(_0609_),
    .ZN(_0615_));
 XOR2_X1 _2175_ (.A(\wr_ptr[4] ),
    .B(\rd_ptr[4] ),
    .Z(_0616_));
 XOR2_X2 _2176_ (.A(_0615_),
    .B(_0616_),
    .Z(_0617_));
 INV_X1 _2177_ (.A(_0617_),
    .ZN(net43));
 INV_X1 _2178_ (.A(net40),
    .ZN(_0618_));
 NAND4_X1 _2179_ (.A1(_0013_),
    .A2(_0618_),
    .A3(_0025_),
    .A4(_0604_),
    .ZN(_0619_));
 AOI21_X4 _2180_ (.A(_0619_),
    .B1(_0606_),
    .B2(_0610_),
    .ZN(_0620_));
 NAND4_X2 _2181_ (.A1(_0609_),
    .A2(_0618_),
    .A3(_0025_),
    .A4(_0604_),
    .ZN(_0621_));
 NOR3_X4 _2182_ (.A1(_0605_),
    .A2(_0607_),
    .A3(_0621_),
    .ZN(_0622_));
 OAI21_X2 _2183_ (.A(net43),
    .B1(_0620_),
    .B2(_0622_),
    .ZN(net98));
 INV_X1 _2184_ (.A(net98),
    .ZN(net62));
 OAI21_X4 _2185_ (.A(_0617_),
    .B1(_0620_),
    .B2(_0622_),
    .ZN(net96));
 INV_X8 _2186_ (.A(net96),
    .ZN(net44));
 CLKBUF_X3 clkload1 (.A(clknet_3_1__leaf_clk));
 INV_X2 clkload0 (.A(clknet_3_0__leaf_clk));
 CLKBUF_X3 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_7__leaf_clk));
 CLKBUF_X3 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_6__leaf_clk));
 CLKBUF_X3 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_5__leaf_clk));
 CLKBUF_X3 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_4__leaf_clk));
 INV_X1 _2193_ (.A(net2),
    .ZN(_0629_));
 NOR2_X1 _2194_ (.A1(_0629_),
    .A2(net96),
    .ZN(net97));
 CLKBUF_X3 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_3__leaf_clk));
 CLKBUF_X3 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_2__leaf_clk));
 CLKBUF_X3 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_1__leaf_clk));
 INV_X1 _2198_ (.A(net36),
    .ZN(_0633_));
 CLKBUF_X3 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_0__leaf_clk));
 NOR3_X1 _2200_ (.A1(_0633_),
    .A2(\wr_ptr[3] ),
    .A3(\wr_ptr[2] ),
    .ZN(_0635_));
 AND2_X1 _2201_ (.A1(_0019_),
    .A2(_0635_),
    .ZN(_0636_));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_leaf_76_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_76_clk));
 MUX2_X1 _2204_ (.A(\mem[0][0] ),
    .B(net4),
    .S(_0636_),
    .Z(_0080_));
 CLKBUF_X3 clkbuf_leaf_75_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_75_clk));
 CLKBUF_X3 clkbuf_leaf_74_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_74_clk));
 MUX2_X1 _2207_ (.A(\mem[0][10] ),
    .B(net5),
    .S(net196),
    .Z(_0081_));
 CLKBUF_X3 clkbuf_leaf_73_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_73_clk));
 CLKBUF_X3 clkbuf_leaf_72_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_72_clk));
 MUX2_X1 _2210_ (.A(\mem[0][11] ),
    .B(net6),
    .S(net196),
    .Z(_0082_));
 CLKBUF_X3 clkbuf_leaf_71_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_71_clk));
 CLKBUF_X3 clkbuf_leaf_70_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_70_clk));
 MUX2_X1 _2213_ (.A(\mem[0][12] ),
    .B(net7),
    .S(net196),
    .Z(_0083_));
 CLKBUF_X3 clkbuf_leaf_69_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_69_clk));
 CLKBUF_X3 clkbuf_leaf_68_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_68_clk));
 MUX2_X1 _2216_ (.A(\mem[0][13] ),
    .B(net8),
    .S(net196),
    .Z(_0084_));
 CLKBUF_X3 clkbuf_leaf_67_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_67_clk));
 CLKBUF_X3 clkbuf_leaf_66_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_66_clk));
 MUX2_X1 _2219_ (.A(\mem[0][14] ),
    .B(net9),
    .S(net196),
    .Z(_0085_));
 CLKBUF_X3 clkbuf_leaf_65_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_65_clk));
 CLKBUF_X3 clkbuf_leaf_64_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_64_clk));
 MUX2_X1 _2222_ (.A(\mem[0][15] ),
    .B(net10),
    .S(net196),
    .Z(_0086_));
 CLKBUF_X3 clkbuf_leaf_63_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_63_clk));
 CLKBUF_X3 clkbuf_leaf_62_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_62_clk));
 MUX2_X1 _2225_ (.A(\mem[0][16] ),
    .B(net11),
    .S(net196),
    .Z(_0087_));
 CLKBUF_X3 clkbuf_leaf_61_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_61_clk));
 CLKBUF_X3 clkbuf_leaf_60_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_60_clk));
 MUX2_X1 _2228_ (.A(\mem[0][17] ),
    .B(net12),
    .S(_0636_),
    .Z(_0088_));
 CLKBUF_X3 clkbuf_leaf_59_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_59_clk));
 CLKBUF_X3 clkbuf_leaf_58_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_58_clk));
 MUX2_X1 _2231_ (.A(\mem[0][18] ),
    .B(net13),
    .S(_0636_),
    .Z(_0089_));
 CLKBUF_X3 clkbuf_leaf_57_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_57_clk));
 CLKBUF_X3 clkbuf_leaf_56_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_56_clk));
 CLKBUF_X3 clkbuf_leaf_55_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_55_clk));
 MUX2_X1 _2235_ (.A(\mem[0][19] ),
    .B(net14),
    .S(net197),
    .Z(_0090_));
 CLKBUF_X3 clkbuf_leaf_54_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_54_clk));
 CLKBUF_X3 clkbuf_leaf_53_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_53_clk));
 MUX2_X1 _2238_ (.A(\mem[0][1] ),
    .B(net15),
    .S(_0636_),
    .Z(_0091_));
 CLKBUF_X3 clkbuf_leaf_52_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_52_clk));
 CLKBUF_X3 clkbuf_leaf_51_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_51_clk));
 MUX2_X1 _2241_ (.A(\mem[0][20] ),
    .B(net16),
    .S(_0636_),
    .Z(_0092_));
 CLKBUF_X3 clkbuf_leaf_50_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_50_clk));
 CLKBUF_X3 clkbuf_leaf_49_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_49_clk));
 MUX2_X1 _2244_ (.A(\mem[0][21] ),
    .B(net17),
    .S(_0636_),
    .Z(_0093_));
 CLKBUF_X3 clkbuf_leaf_48_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_48_clk));
 CLKBUF_X3 clkbuf_leaf_47_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_47_clk));
 MUX2_X1 _2247_ (.A(\mem[0][22] ),
    .B(net18),
    .S(_0636_),
    .Z(_0094_));
 CLKBUF_X3 clkbuf_leaf_46_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_46_clk));
 CLKBUF_X3 clkbuf_leaf_45_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_45_clk));
 MUX2_X1 _2250_ (.A(\mem[0][23] ),
    .B(net19),
    .S(_0636_),
    .Z(_0095_));
 CLKBUF_X3 clkbuf_leaf_44_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_44_clk));
 CLKBUF_X3 clkbuf_leaf_43_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_43_clk));
 MUX2_X1 _2253_ (.A(\mem[0][24] ),
    .B(net20),
    .S(_0636_),
    .Z(_0096_));
 CLKBUF_X3 clkbuf_leaf_42_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_42_clk));
 CLKBUF_X3 clkbuf_leaf_41_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_41_clk));
 MUX2_X1 _2256_ (.A(\mem[0][25] ),
    .B(net21),
    .S(net197),
    .Z(_0097_));
 CLKBUF_X3 clkbuf_leaf_40_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_40_clk));
 CLKBUF_X3 clkbuf_leaf_39_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_39_clk));
 MUX2_X1 _2259_ (.A(\mem[0][26] ),
    .B(net22),
    .S(net197),
    .Z(_0098_));
 CLKBUF_X3 clkbuf_leaf_38_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_38_clk));
 CLKBUF_X3 clkbuf_leaf_37_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_37_clk));
 MUX2_X1 _2262_ (.A(\mem[0][27] ),
    .B(net23),
    .S(net197),
    .Z(_0099_));
 CLKBUF_X3 clkbuf_leaf_36_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_36_clk));
 CLKBUF_X3 clkbuf_leaf_35_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_35_clk));
 CLKBUF_X3 clkbuf_leaf_34_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_34_clk));
 MUX2_X1 _2266_ (.A(\mem[0][28] ),
    .B(net24),
    .S(net197),
    .Z(_0100_));
 CLKBUF_X3 clkbuf_leaf_33_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_33_clk));
 CLKBUF_X3 clkbuf_leaf_32_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_32_clk));
 MUX2_X1 _2269_ (.A(\mem[0][29] ),
    .B(net25),
    .S(net197),
    .Z(_0101_));
 CLKBUF_X3 clkbuf_leaf_31_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_31_clk));
 CLKBUF_X3 clkbuf_leaf_30_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_30_clk));
 MUX2_X1 _2272_ (.A(\mem[0][2] ),
    .B(net26),
    .S(net197),
    .Z(_0102_));
 CLKBUF_X3 clkbuf_leaf_29_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_29_clk));
 CLKBUF_X3 clkbuf_leaf_28_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_28_clk));
 MUX2_X1 _2275_ (.A(\mem[0][30] ),
    .B(net27),
    .S(net197),
    .Z(_0103_));
 CLKBUF_X3 clkbuf_leaf_27_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_27_clk));
 CLKBUF_X3 clkbuf_leaf_26_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_26_clk));
 MUX2_X1 _2278_ (.A(\mem[0][31] ),
    .B(net28),
    .S(net197),
    .Z(_0104_));
 CLKBUF_X3 clkbuf_leaf_25_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_25_clk));
 CLKBUF_X3 clkbuf_leaf_24_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_24_clk));
 MUX2_X1 _2281_ (.A(\mem[0][3] ),
    .B(net29),
    .S(net197),
    .Z(_0105_));
 CLKBUF_X3 clkbuf_leaf_23_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_23_clk));
 CLKBUF_X3 clkbuf_leaf_22_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_22_clk));
 MUX2_X1 _2284_ (.A(\mem[0][4] ),
    .B(net30),
    .S(net197),
    .Z(_0106_));
 CLKBUF_X3 clkbuf_leaf_21_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_21_clk));
 CLKBUF_X3 clkbuf_leaf_20_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_20_clk));
 MUX2_X1 _2287_ (.A(\mem[0][5] ),
    .B(net31),
    .S(_0636_),
    .Z(_0107_));
 CLKBUF_X3 clkbuf_leaf_19_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_19_clk));
 CLKBUF_X3 clkbuf_leaf_18_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_18_clk));
 MUX2_X1 _2290_ (.A(\mem[0][6] ),
    .B(net32),
    .S(_0636_),
    .Z(_0108_));
 CLKBUF_X3 clkbuf_leaf_17_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_17_clk));
 CLKBUF_X3 clkbuf_leaf_16_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_16_clk));
 MUX2_X1 _2293_ (.A(\mem[0][7] ),
    .B(net33),
    .S(net196),
    .Z(_0109_));
 CLKBUF_X3 clkbuf_leaf_15_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_15_clk));
 CLKBUF_X3 clkbuf_leaf_14_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_14_clk));
 MUX2_X1 _2296_ (.A(\mem[0][8] ),
    .B(net34),
    .S(_0636_),
    .Z(_0110_));
 CLKBUF_X3 clkbuf_leaf_13_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_13_clk));
 CLKBUF_X3 clkbuf_leaf_12_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_12_clk));
 MUX2_X1 _2299_ (.A(\mem[0][9] ),
    .B(net35),
    .S(net196),
    .Z(_0111_));
 CLKBUF_X3 clkbuf_leaf_11_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_11_clk));
 INV_X1 _2301_ (.A(\wr_ptr[3] ),
    .ZN(_0704_));
 NOR3_X1 _2302_ (.A1(_0633_),
    .A2(_0704_),
    .A3(\wr_ptr[2] ),
    .ZN(_0705_));
 NAND2_X2 _2303_ (.A1(_0021_),
    .A2(net195),
    .ZN(_0706_));
 CLKBUF_X3 clkbuf_leaf_10_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_10_clk));
 MUX2_X1 _2305_ (.A(net4),
    .B(\mem[10][0] ),
    .S(_0706_),
    .Z(_0112_));
 MUX2_X1 _2306_ (.A(net5),
    .B(\mem[10][10] ),
    .S(_0706_),
    .Z(_0113_));
 MUX2_X1 _2307_ (.A(net6),
    .B(\mem[10][11] ),
    .S(_0706_),
    .Z(_0114_));
 MUX2_X1 _2308_ (.A(net7),
    .B(\mem[10][12] ),
    .S(_0706_),
    .Z(_0115_));
 MUX2_X1 _2309_ (.A(net8),
    .B(\mem[10][13] ),
    .S(_0706_),
    .Z(_0116_));
 MUX2_X1 _2310_ (.A(net9),
    .B(\mem[10][14] ),
    .S(_0706_),
    .Z(_0117_));
 MUX2_X1 _2311_ (.A(net10),
    .B(\mem[10][15] ),
    .S(_0706_),
    .Z(_0118_));
 MUX2_X1 _2312_ (.A(net11),
    .B(\mem[10][16] ),
    .S(_0706_),
    .Z(_0119_));
 MUX2_X1 _2313_ (.A(net12),
    .B(\mem[10][17] ),
    .S(_0706_),
    .Z(_0120_));
 MUX2_X1 _2314_ (.A(net13),
    .B(\mem[10][18] ),
    .S(_0706_),
    .Z(_0121_));
 CLKBUF_X3 clkbuf_leaf_9_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_9_clk));
 MUX2_X1 _2316_ (.A(net14),
    .B(\mem[10][19] ),
    .S(_0706_),
    .Z(_0122_));
 MUX2_X1 _2317_ (.A(net15),
    .B(\mem[10][1] ),
    .S(net187),
    .Z(_0123_));
 MUX2_X1 _2318_ (.A(net16),
    .B(\mem[10][20] ),
    .S(net187),
    .Z(_0124_));
 MUX2_X1 _2319_ (.A(net17),
    .B(\mem[10][21] ),
    .S(net187),
    .Z(_0125_));
 MUX2_X1 _2320_ (.A(net18),
    .B(\mem[10][22] ),
    .S(net187),
    .Z(_0126_));
 MUX2_X1 _2321_ (.A(net19),
    .B(\mem[10][23] ),
    .S(net187),
    .Z(_0127_));
 MUX2_X1 _2322_ (.A(net20),
    .B(\mem[10][24] ),
    .S(net187),
    .Z(_0128_));
 MUX2_X1 _2323_ (.A(net21),
    .B(\mem[10][25] ),
    .S(_0706_),
    .Z(_0129_));
 MUX2_X1 _2324_ (.A(net22),
    .B(\mem[10][26] ),
    .S(net187),
    .Z(_0130_));
 MUX2_X1 _2325_ (.A(net23),
    .B(\mem[10][27] ),
    .S(_0706_),
    .Z(_0131_));
 CLKBUF_X3 clkbuf_leaf_8_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_8_clk));
 MUX2_X1 _2327_ (.A(net24),
    .B(\mem[10][28] ),
    .S(net187),
    .Z(_0132_));
 MUX2_X1 _2328_ (.A(net25),
    .B(\mem[10][29] ),
    .S(net187),
    .Z(_0133_));
 MUX2_X1 _2329_ (.A(net26),
    .B(\mem[10][2] ),
    .S(net187),
    .Z(_0134_));
 MUX2_X1 _2330_ (.A(net27),
    .B(\mem[10][30] ),
    .S(net187),
    .Z(_0135_));
 MUX2_X1 _2331_ (.A(net28),
    .B(\mem[10][31] ),
    .S(_0706_),
    .Z(_0136_));
 MUX2_X1 _2332_ (.A(net29),
    .B(\mem[10][3] ),
    .S(net187),
    .Z(_0137_));
 MUX2_X1 _2333_ (.A(net30),
    .B(\mem[10][4] ),
    .S(_0706_),
    .Z(_0138_));
 MUX2_X1 _2334_ (.A(net31),
    .B(\mem[10][5] ),
    .S(_0706_),
    .Z(_0139_));
 MUX2_X1 _2335_ (.A(net32),
    .B(\mem[10][6] ),
    .S(_0706_),
    .Z(_0140_));
 MUX2_X1 _2336_ (.A(net33),
    .B(\mem[10][7] ),
    .S(_0706_),
    .Z(_0141_));
 MUX2_X1 _2337_ (.A(net34),
    .B(\mem[10][8] ),
    .S(_0706_),
    .Z(_0142_));
 MUX2_X1 _2338_ (.A(net35),
    .B(\mem[10][9] ),
    .S(_0706_),
    .Z(_0143_));
 CLKBUF_X3 clkbuf_leaf_7_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_7_clk));
 NAND2_X2 _2340_ (.A1(_0023_),
    .A2(net195),
    .ZN(_0711_));
 CLKBUF_X3 clkbuf_leaf_6_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_6_clk));
 MUX2_X1 _2342_ (.A(net4),
    .B(\mem[11][0] ),
    .S(net186),
    .Z(_0144_));
 MUX2_X1 _2343_ (.A(net5),
    .B(\mem[11][10] ),
    .S(net186),
    .Z(_0145_));
 MUX2_X1 _2344_ (.A(net6),
    .B(\mem[11][11] ),
    .S(net186),
    .Z(_0146_));
 MUX2_X1 _2345_ (.A(net7),
    .B(\mem[11][12] ),
    .S(net186),
    .Z(_0147_));
 MUX2_X1 _2346_ (.A(net8),
    .B(\mem[11][13] ),
    .S(net186),
    .Z(_0148_));
 MUX2_X1 _2347_ (.A(net9),
    .B(\mem[11][14] ),
    .S(net186),
    .Z(_0149_));
 MUX2_X1 _2348_ (.A(net10),
    .B(\mem[11][15] ),
    .S(net186),
    .Z(_0150_));
 MUX2_X1 _2349_ (.A(net11),
    .B(\mem[11][16] ),
    .S(net186),
    .Z(_0151_));
 MUX2_X1 _2350_ (.A(net12),
    .B(\mem[11][17] ),
    .S(net186),
    .Z(_0152_));
 MUX2_X1 _2351_ (.A(net13),
    .B(\mem[11][18] ),
    .S(net186),
    .Z(_0153_));
 CLKBUF_X3 clkbuf_leaf_5_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_5_clk));
 MUX2_X1 _2353_ (.A(net14),
    .B(\mem[11][19] ),
    .S(_0711_),
    .Z(_0154_));
 MUX2_X1 _2354_ (.A(net15),
    .B(\mem[11][1] ),
    .S(_0711_),
    .Z(_0155_));
 MUX2_X1 _2355_ (.A(net16),
    .B(\mem[11][20] ),
    .S(_0711_),
    .Z(_0156_));
 MUX2_X1 _2356_ (.A(net17),
    .B(\mem[11][21] ),
    .S(_0711_),
    .Z(_0157_));
 MUX2_X1 _2357_ (.A(net18),
    .B(\mem[11][22] ),
    .S(_0711_),
    .Z(_0158_));
 MUX2_X1 _2358_ (.A(net19),
    .B(\mem[11][23] ),
    .S(_0711_),
    .Z(_0159_));
 MUX2_X1 _2359_ (.A(net20),
    .B(\mem[11][24] ),
    .S(_0711_),
    .Z(_0160_));
 MUX2_X1 _2360_ (.A(net21),
    .B(\mem[11][25] ),
    .S(_0711_),
    .Z(_0161_));
 MUX2_X1 _2361_ (.A(net22),
    .B(\mem[11][26] ),
    .S(_0711_),
    .Z(_0162_));
 MUX2_X1 _2362_ (.A(net23),
    .B(\mem[11][27] ),
    .S(_0711_),
    .Z(_0163_));
 CLKBUF_X3 clkbuf_leaf_4_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_4_clk));
 MUX2_X1 _2364_ (.A(net24),
    .B(\mem[11][28] ),
    .S(_0711_),
    .Z(_0164_));
 MUX2_X1 _2365_ (.A(net25),
    .B(\mem[11][29] ),
    .S(_0711_),
    .Z(_0165_));
 MUX2_X1 _2366_ (.A(net26),
    .B(\mem[11][2] ),
    .S(_0711_),
    .Z(_0166_));
 MUX2_X1 _2367_ (.A(net27),
    .B(\mem[11][30] ),
    .S(_0711_),
    .Z(_0167_));
 MUX2_X1 _2368_ (.A(net28),
    .B(\mem[11][31] ),
    .S(_0711_),
    .Z(_0168_));
 MUX2_X1 _2369_ (.A(net29),
    .B(\mem[11][3] ),
    .S(_0711_),
    .Z(_0169_));
 MUX2_X1 _2370_ (.A(net30),
    .B(\mem[11][4] ),
    .S(_0711_),
    .Z(_0170_));
 MUX2_X1 _2371_ (.A(net31),
    .B(\mem[11][5] ),
    .S(_0711_),
    .Z(_0171_));
 MUX2_X1 _2372_ (.A(net32),
    .B(\mem[11][6] ),
    .S(_0711_),
    .Z(_0172_));
 MUX2_X1 _2373_ (.A(net33),
    .B(\mem[11][7] ),
    .S(net186),
    .Z(_0173_));
 MUX2_X1 _2374_ (.A(net34),
    .B(\mem[11][8] ),
    .S(_0711_),
    .Z(_0174_));
 MUX2_X1 _2375_ (.A(net35),
    .B(\mem[11][9] ),
    .S(net186),
    .Z(_0175_));
 AND2_X1 _2376_ (.A1(net36),
    .A2(\wr_ptr[2] ),
    .ZN(_0715_));
 AND2_X1 _2377_ (.A1(\wr_ptr[3] ),
    .A2(_0715_),
    .ZN(_0716_));
 CLKBUF_X3 clkbuf_leaf_3_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_3_clk));
 NAND2_X2 _2379_ (.A1(_0019_),
    .A2(_0716_),
    .ZN(_0718_));
 BUF_X4 place207 (.A(_0000_),
    .Z(net207));
 MUX2_X1 _2381_ (.A(net4),
    .B(\mem[12][0] ),
    .S(_0718_),
    .Z(_0176_));
 MUX2_X1 _2382_ (.A(net5),
    .B(\mem[12][10] ),
    .S(_0718_),
    .Z(_0177_));
 MUX2_X1 _2383_ (.A(net6),
    .B(\mem[12][11] ),
    .S(_0718_),
    .Z(_0178_));
 MUX2_X1 _2384_ (.A(net7),
    .B(\mem[12][12] ),
    .S(_0718_),
    .Z(_0179_));
 MUX2_X1 _2385_ (.A(net8),
    .B(\mem[12][13] ),
    .S(_0718_),
    .Z(_0180_));
 MUX2_X1 _2386_ (.A(net9),
    .B(\mem[12][14] ),
    .S(_0718_),
    .Z(_0181_));
 MUX2_X1 _2387_ (.A(net10),
    .B(\mem[12][15] ),
    .S(_0718_),
    .Z(_0182_));
 MUX2_X1 _2388_ (.A(net11),
    .B(\mem[12][16] ),
    .S(_0718_),
    .Z(_0183_));
 MUX2_X1 _2389_ (.A(net12),
    .B(\mem[12][17] ),
    .S(_0718_),
    .Z(_0184_));
 MUX2_X1 _2390_ (.A(net13),
    .B(\mem[12][18] ),
    .S(_0718_),
    .Z(_0185_));
 BUF_X4 place206 (.A(_0000_),
    .Z(net206));
 MUX2_X1 _2392_ (.A(net14),
    .B(\mem[12][19] ),
    .S(_0718_),
    .Z(_0186_));
 MUX2_X1 _2393_ (.A(net15),
    .B(\mem[12][1] ),
    .S(net185),
    .Z(_0187_));
 MUX2_X1 _2394_ (.A(net16),
    .B(\mem[12][20] ),
    .S(net185),
    .Z(_0188_));
 MUX2_X1 _2395_ (.A(net17),
    .B(\mem[12][21] ),
    .S(net185),
    .Z(_0189_));
 MUX2_X1 _2396_ (.A(net18),
    .B(\mem[12][22] ),
    .S(net185),
    .Z(_0190_));
 MUX2_X1 _2397_ (.A(net19),
    .B(\mem[12][23] ),
    .S(net185),
    .Z(_0191_));
 MUX2_X1 _2398_ (.A(net20),
    .B(\mem[12][24] ),
    .S(net185),
    .Z(_0192_));
 MUX2_X1 _2399_ (.A(net21),
    .B(\mem[12][25] ),
    .S(net185),
    .Z(_0193_));
 MUX2_X1 _2400_ (.A(net22),
    .B(\mem[12][26] ),
    .S(net185),
    .Z(_0194_));
 MUX2_X1 _2401_ (.A(net23),
    .B(\mem[12][27] ),
    .S(net185),
    .Z(_0195_));
 BUF_X4 place201 (.A(_0002_),
    .Z(net201));
 MUX2_X1 _2403_ (.A(net24),
    .B(\mem[12][28] ),
    .S(net185),
    .Z(_0196_));
 MUX2_X1 _2404_ (.A(net25),
    .B(\mem[12][29] ),
    .S(net185),
    .Z(_0197_));
 MUX2_X1 _2405_ (.A(net26),
    .B(\mem[12][2] ),
    .S(net185),
    .Z(_0198_));
 MUX2_X1 _2406_ (.A(net27),
    .B(\mem[12][30] ),
    .S(net185),
    .Z(_0199_));
 MUX2_X1 _2407_ (.A(net28),
    .B(\mem[12][31] ),
    .S(_0718_),
    .Z(_0200_));
 MUX2_X1 _2408_ (.A(net29),
    .B(\mem[12][3] ),
    .S(_0718_),
    .Z(_0201_));
 MUX2_X1 _2409_ (.A(net30),
    .B(\mem[12][4] ),
    .S(_0718_),
    .Z(_0202_));
 MUX2_X1 _2410_ (.A(net31),
    .B(\mem[12][5] ),
    .S(_0718_),
    .Z(_0203_));
 MUX2_X1 _2411_ (.A(net32),
    .B(\mem[12][6] ),
    .S(_0718_),
    .Z(_0204_));
 MUX2_X1 _2412_ (.A(net33),
    .B(\mem[12][7] ),
    .S(_0718_),
    .Z(_0205_));
 MUX2_X1 _2413_ (.A(net34),
    .B(\mem[12][8] ),
    .S(_0718_),
    .Z(_0206_));
 MUX2_X1 _2414_ (.A(net35),
    .B(\mem[12][9] ),
    .S(_0718_),
    .Z(_0207_));
 BUF_X2 place198 (.A(_0880_),
    .Z(net198));
 NAND2_X2 _2416_ (.A1(_0022_),
    .A2(_0716_),
    .ZN(_0723_));
 BUF_X1 place197 (.A(_0636_),
    .Z(net197));
 MUX2_X1 _2418_ (.A(net4),
    .B(\mem[13][0] ),
    .S(_0723_),
    .Z(_0208_));
 MUX2_X1 _2419_ (.A(net5),
    .B(\mem[13][10] ),
    .S(net184),
    .Z(_0209_));
 MUX2_X1 _2420_ (.A(net6),
    .B(\mem[13][11] ),
    .S(net184),
    .Z(_0210_));
 MUX2_X1 _2421_ (.A(net7),
    .B(\mem[13][12] ),
    .S(net184),
    .Z(_0211_));
 MUX2_X1 _2422_ (.A(net8),
    .B(\mem[13][13] ),
    .S(net184),
    .Z(_0212_));
 MUX2_X1 _2423_ (.A(net9),
    .B(\mem[13][14] ),
    .S(net184),
    .Z(_0213_));
 MUX2_X1 _2424_ (.A(net10),
    .B(\mem[13][15] ),
    .S(net184),
    .Z(_0214_));
 MUX2_X1 _2425_ (.A(net11),
    .B(\mem[13][16] ),
    .S(net184),
    .Z(_0215_));
 MUX2_X1 _2426_ (.A(net12),
    .B(\mem[13][17] ),
    .S(_0723_),
    .Z(_0216_));
 MUX2_X1 _2427_ (.A(net13),
    .B(\mem[13][18] ),
    .S(_0723_),
    .Z(_0217_));
 BUF_X2 place173 (.A(net96),
    .Z(net173));
 MUX2_X1 _2429_ (.A(net14),
    .B(\mem[13][19] ),
    .S(_0723_),
    .Z(_0218_));
 MUX2_X1 _2430_ (.A(net15),
    .B(\mem[13][1] ),
    .S(_0723_),
    .Z(_0219_));
 MUX2_X1 _2431_ (.A(net16),
    .B(\mem[13][20] ),
    .S(_0723_),
    .Z(_0220_));
 MUX2_X1 _2432_ (.A(net17),
    .B(\mem[13][21] ),
    .S(_0723_),
    .Z(_0221_));
 MUX2_X1 _2433_ (.A(net18),
    .B(\mem[13][22] ),
    .S(_0723_),
    .Z(_0222_));
 MUX2_X1 _2434_ (.A(net19),
    .B(\mem[13][23] ),
    .S(_0723_),
    .Z(_0223_));
 MUX2_X1 _2435_ (.A(net20),
    .B(\mem[13][24] ),
    .S(_0723_),
    .Z(_0224_));
 MUX2_X1 _2436_ (.A(net21),
    .B(\mem[13][25] ),
    .S(_0723_),
    .Z(_0225_));
 MUX2_X1 _2437_ (.A(net22),
    .B(\mem[13][26] ),
    .S(_0723_),
    .Z(_0226_));
 MUX2_X1 _2438_ (.A(net23),
    .B(\mem[13][27] ),
    .S(_0723_),
    .Z(_0227_));
 BUF_X8 place172 (.A(net44),
    .Z(net172));
 MUX2_X1 _2440_ (.A(net24),
    .B(\mem[13][28] ),
    .S(_0723_),
    .Z(_0228_));
 MUX2_X1 _2441_ (.A(net25),
    .B(\mem[13][29] ),
    .S(_0723_),
    .Z(_0229_));
 MUX2_X1 _2442_ (.A(net26),
    .B(\mem[13][2] ),
    .S(_0723_),
    .Z(_0230_));
 MUX2_X1 _2443_ (.A(net27),
    .B(\mem[13][30] ),
    .S(_0723_),
    .Z(_0231_));
 MUX2_X1 _2444_ (.A(net28),
    .B(\mem[13][31] ),
    .S(_0723_),
    .Z(_0232_));
 MUX2_X1 _2445_ (.A(net29),
    .B(\mem[13][3] ),
    .S(_0723_),
    .Z(_0233_));
 MUX2_X1 _2446_ (.A(net30),
    .B(\mem[13][4] ),
    .S(_0723_),
    .Z(_0234_));
 MUX2_X1 _2447_ (.A(net31),
    .B(\mem[13][5] ),
    .S(_0723_),
    .Z(_0235_));
 MUX2_X1 _2448_ (.A(net32),
    .B(\mem[13][6] ),
    .S(_0723_),
    .Z(_0236_));
 MUX2_X1 _2449_ (.A(net33),
    .B(\mem[13][7] ),
    .S(net184),
    .Z(_0237_));
 MUX2_X1 _2450_ (.A(net34),
    .B(\mem[13][8] ),
    .S(_0723_),
    .Z(_0238_));
 MUX2_X1 _2451_ (.A(net35),
    .B(\mem[13][9] ),
    .S(net184),
    .Z(_0239_));
 NAND2_X2 _2452_ (.A1(_0021_),
    .A2(_0716_),
    .ZN(_0727_));
 CLKBUF_X3 clkbuf_leaf_0_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_0_clk));
 MUX2_X1 _2454_ (.A(net4),
    .B(\mem[14][0] ),
    .S(net183),
    .Z(_0240_));
 MUX2_X1 _2455_ (.A(net5),
    .B(\mem[14][10] ),
    .S(net183),
    .Z(_0241_));
 MUX2_X1 _2456_ (.A(net6),
    .B(\mem[14][11] ),
    .S(net183),
    .Z(_0242_));
 MUX2_X1 _2457_ (.A(net7),
    .B(\mem[14][12] ),
    .S(net183),
    .Z(_0243_));
 MUX2_X1 _2458_ (.A(net8),
    .B(\mem[14][13] ),
    .S(net183),
    .Z(_0244_));
 MUX2_X1 _2459_ (.A(net9),
    .B(\mem[14][14] ),
    .S(net183),
    .Z(_0245_));
 MUX2_X1 _2460_ (.A(net10),
    .B(\mem[14][15] ),
    .S(net183),
    .Z(_0246_));
 MUX2_X1 _2461_ (.A(net11),
    .B(\mem[14][16] ),
    .S(net183),
    .Z(_0247_));
 MUX2_X1 _2462_ (.A(net12),
    .B(\mem[14][17] ),
    .S(net183),
    .Z(_0248_));
 MUX2_X1 _2463_ (.A(net13),
    .B(\mem[14][18] ),
    .S(net183),
    .Z(_0249_));
 BUF_X2 place210 (.A(net2),
    .Z(net210));
 MUX2_X1 _2465_ (.A(net14),
    .B(\mem[14][19] ),
    .S(_0727_),
    .Z(_0250_));
 MUX2_X1 _2466_ (.A(net15),
    .B(\mem[14][1] ),
    .S(_0727_),
    .Z(_0251_));
 MUX2_X1 _2467_ (.A(net16),
    .B(\mem[14][20] ),
    .S(_0727_),
    .Z(_0252_));
 MUX2_X1 _2468_ (.A(net17),
    .B(\mem[14][21] ),
    .S(_0727_),
    .Z(_0253_));
 MUX2_X1 _2469_ (.A(net18),
    .B(\mem[14][22] ),
    .S(_0727_),
    .Z(_0254_));
 MUX2_X1 _2470_ (.A(net19),
    .B(\mem[14][23] ),
    .S(_0727_),
    .Z(_0255_));
 MUX2_X1 _2471_ (.A(net20),
    .B(\mem[14][24] ),
    .S(_0727_),
    .Z(_0256_));
 MUX2_X1 _2472_ (.A(net21),
    .B(\mem[14][25] ),
    .S(_0727_),
    .Z(_0257_));
 MUX2_X1 _2473_ (.A(net22),
    .B(\mem[14][26] ),
    .S(_0727_),
    .Z(_0258_));
 MUX2_X1 _2474_ (.A(net23),
    .B(\mem[14][27] ),
    .S(_0727_),
    .Z(_0259_));
 BUF_X1 place178 (.A(_0766_),
    .Z(net178));
 MUX2_X1 _2476_ (.A(net24),
    .B(\mem[14][28] ),
    .S(_0727_),
    .Z(_0260_));
 MUX2_X1 _2477_ (.A(net25),
    .B(\mem[14][29] ),
    .S(_0727_),
    .Z(_0261_));
 MUX2_X1 _2478_ (.A(net26),
    .B(\mem[14][2] ),
    .S(_0727_),
    .Z(_0262_));
 MUX2_X1 _2479_ (.A(net27),
    .B(\mem[14][30] ),
    .S(_0727_),
    .Z(_0263_));
 MUX2_X1 _2480_ (.A(net28),
    .B(\mem[14][31] ),
    .S(net183),
    .Z(_0264_));
 MUX2_X1 _2481_ (.A(net29),
    .B(\mem[14][3] ),
    .S(_0727_),
    .Z(_0265_));
 MUX2_X1 _2482_ (.A(net30),
    .B(\mem[14][4] ),
    .S(net183),
    .Z(_0266_));
 MUX2_X1 _2483_ (.A(net31),
    .B(\mem[14][5] ),
    .S(net183),
    .Z(_0267_));
 MUX2_X1 _2484_ (.A(net32),
    .B(\mem[14][6] ),
    .S(net183),
    .Z(_0268_));
 MUX2_X1 _2485_ (.A(net33),
    .B(\mem[14][7] ),
    .S(net183),
    .Z(_0269_));
 MUX2_X1 _2486_ (.A(net34),
    .B(\mem[14][8] ),
    .S(net183),
    .Z(_0270_));
 MUX2_X1 _2487_ (.A(net35),
    .B(\mem[14][9] ),
    .S(net183),
    .Z(_0271_));
 NAND2_X2 _2488_ (.A1(_0023_),
    .A2(_0716_),
    .ZN(_0731_));
 BUF_X2 place174 (.A(net96),
    .Z(net174));
 MUX2_X1 _2490_ (.A(net4),
    .B(\mem[15][0] ),
    .S(net182),
    .Z(_0272_));
 MUX2_X1 _2491_ (.A(net5),
    .B(\mem[15][10] ),
    .S(net182),
    .Z(_0273_));
 MUX2_X1 _2492_ (.A(net6),
    .B(\mem[15][11] ),
    .S(net182),
    .Z(_0274_));
 MUX2_X1 _2493_ (.A(net7),
    .B(\mem[15][12] ),
    .S(net182),
    .Z(_0275_));
 MUX2_X1 _2494_ (.A(net8),
    .B(\mem[15][13] ),
    .S(net182),
    .Z(_0276_));
 MUX2_X1 _2495_ (.A(net9),
    .B(\mem[15][14] ),
    .S(net182),
    .Z(_0277_));
 MUX2_X1 _2496_ (.A(net10),
    .B(\mem[15][15] ),
    .S(net182),
    .Z(_0278_));
 MUX2_X1 _2497_ (.A(net11),
    .B(\mem[15][16] ),
    .S(net182),
    .Z(_0279_));
 MUX2_X1 _2498_ (.A(net12),
    .B(\mem[15][17] ),
    .S(net182),
    .Z(_0280_));
 MUX2_X1 _2499_ (.A(net13),
    .B(\mem[15][18] ),
    .S(net182),
    .Z(_0281_));
 BUF_X1 place209 (.A(_0629_),
    .Z(net209));
 MUX2_X1 _2501_ (.A(net14),
    .B(\mem[15][19] ),
    .S(_0731_),
    .Z(_0282_));
 MUX2_X1 _2502_ (.A(net15),
    .B(\mem[15][1] ),
    .S(_0731_),
    .Z(_0283_));
 MUX2_X1 _2503_ (.A(net16),
    .B(\mem[15][20] ),
    .S(_0731_),
    .Z(_0284_));
 MUX2_X1 _2504_ (.A(net17),
    .B(\mem[15][21] ),
    .S(_0731_),
    .Z(_0285_));
 MUX2_X1 _2505_ (.A(net18),
    .B(\mem[15][22] ),
    .S(_0731_),
    .Z(_0286_));
 MUX2_X1 _2506_ (.A(net19),
    .B(\mem[15][23] ),
    .S(_0731_),
    .Z(_0287_));
 MUX2_X1 _2507_ (.A(net20),
    .B(\mem[15][24] ),
    .S(_0731_),
    .Z(_0288_));
 MUX2_X1 _2508_ (.A(net21),
    .B(\mem[15][25] ),
    .S(_0731_),
    .Z(_0289_));
 MUX2_X1 _2509_ (.A(net22),
    .B(\mem[15][26] ),
    .S(_0731_),
    .Z(_0290_));
 MUX2_X1 _2510_ (.A(net23),
    .B(\mem[15][27] ),
    .S(_0731_),
    .Z(_0291_));
 BUF_X8 place204 (.A(_0002_),
    .Z(net204));
 MUX2_X1 _2512_ (.A(net24),
    .B(\mem[15][28] ),
    .S(_0731_),
    .Z(_0292_));
 MUX2_X1 _2513_ (.A(net25),
    .B(\mem[15][29] ),
    .S(_0731_),
    .Z(_0293_));
 MUX2_X1 _2514_ (.A(net26),
    .B(\mem[15][2] ),
    .S(_0731_),
    .Z(_0294_));
 MUX2_X1 _2515_ (.A(net27),
    .B(\mem[15][30] ),
    .S(_0731_),
    .Z(_0295_));
 MUX2_X1 _2516_ (.A(net28),
    .B(\mem[15][31] ),
    .S(_0731_),
    .Z(_0296_));
 MUX2_X1 _2517_ (.A(net29),
    .B(\mem[15][3] ),
    .S(_0731_),
    .Z(_0297_));
 MUX2_X1 _2518_ (.A(net30),
    .B(\mem[15][4] ),
    .S(_0731_),
    .Z(_0298_));
 MUX2_X1 _2519_ (.A(net31),
    .B(\mem[15][5] ),
    .S(_0731_),
    .Z(_0299_));
 MUX2_X1 _2520_ (.A(net32),
    .B(\mem[15][6] ),
    .S(net182),
    .Z(_0300_));
 MUX2_X1 _2521_ (.A(net33),
    .B(\mem[15][7] ),
    .S(net182),
    .Z(_0301_));
 MUX2_X1 _2522_ (.A(net34),
    .B(\mem[15][8] ),
    .S(_0731_),
    .Z(_0302_));
 MUX2_X1 _2523_ (.A(net35),
    .B(\mem[15][9] ),
    .S(net182),
    .Z(_0303_));
 AND2_X1 _2524_ (.A1(_0022_),
    .A2(_0635_),
    .ZN(_0735_));
 BUF_X8 place203 (.A(_0002_),
    .Z(net203));
 BUF_X1 place192 (.A(_0745_),
    .Z(net192));
 MUX2_X1 _2527_ (.A(\mem[1][0] ),
    .B(net4),
    .S(net194),
    .Z(_0304_));
 MUX2_X1 _2528_ (.A(\mem[1][10] ),
    .B(net5),
    .S(net194),
    .Z(_0305_));
 MUX2_X1 _2529_ (.A(\mem[1][11] ),
    .B(net6),
    .S(net194),
    .Z(_0306_));
 MUX2_X1 _2530_ (.A(\mem[1][12] ),
    .B(net7),
    .S(net194),
    .Z(_0307_));
 MUX2_X1 _2531_ (.A(\mem[1][13] ),
    .B(net8),
    .S(net194),
    .Z(_0308_));
 MUX2_X1 _2532_ (.A(\mem[1][14] ),
    .B(net9),
    .S(net194),
    .Z(_0309_));
 MUX2_X1 _2533_ (.A(\mem[1][15] ),
    .B(net10),
    .S(net194),
    .Z(_0310_));
 MUX2_X1 _2534_ (.A(\mem[1][16] ),
    .B(net11),
    .S(net194),
    .Z(_0311_));
 MUX2_X1 _2535_ (.A(\mem[1][17] ),
    .B(net12),
    .S(net194),
    .Z(_0312_));
 MUX2_X1 _2536_ (.A(\mem[1][18] ),
    .B(net13),
    .S(net194),
    .Z(_0313_));
 CLKBUF_X3 clkbuf_leaf_2_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_2_clk));
 MUX2_X1 _2538_ (.A(\mem[1][19] ),
    .B(net14),
    .S(net194),
    .Z(_0314_));
 MUX2_X1 _2539_ (.A(\mem[1][1] ),
    .B(net15),
    .S(net194),
    .Z(_0315_));
 MUX2_X1 _2540_ (.A(\mem[1][20] ),
    .B(net16),
    .S(net194),
    .Z(_0316_));
 MUX2_X1 _2541_ (.A(\mem[1][21] ),
    .B(net17),
    .S(net194),
    .Z(_0317_));
 MUX2_X1 _2542_ (.A(\mem[1][22] ),
    .B(net18),
    .S(net194),
    .Z(_0318_));
 MUX2_X1 _2543_ (.A(\mem[1][23] ),
    .B(net19),
    .S(net194),
    .Z(_0319_));
 MUX2_X1 _2544_ (.A(\mem[1][24] ),
    .B(net20),
    .S(net194),
    .Z(_0320_));
 MUX2_X1 _2545_ (.A(\mem[1][25] ),
    .B(net21),
    .S(net194),
    .Z(_0321_));
 MUX2_X1 _2546_ (.A(\mem[1][26] ),
    .B(net22),
    .S(net194),
    .Z(_0322_));
 MUX2_X1 _2547_ (.A(\mem[1][27] ),
    .B(net23),
    .S(net194),
    .Z(_0323_));
 CLKBUF_X3 clkbuf_leaf_1_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_1_clk));
 MUX2_X1 _2549_ (.A(\mem[1][28] ),
    .B(net24),
    .S(net194),
    .Z(_0324_));
 MUX2_X1 _2550_ (.A(\mem[1][29] ),
    .B(net25),
    .S(net194),
    .Z(_0325_));
 MUX2_X1 _2551_ (.A(\mem[1][2] ),
    .B(net26),
    .S(net194),
    .Z(_0326_));
 MUX2_X1 _2552_ (.A(\mem[1][30] ),
    .B(net27),
    .S(net194),
    .Z(_0327_));
 MUX2_X1 _2553_ (.A(\mem[1][31] ),
    .B(net28),
    .S(net194),
    .Z(_0328_));
 MUX2_X1 _2554_ (.A(\mem[1][3] ),
    .B(net29),
    .S(net194),
    .Z(_0329_));
 MUX2_X1 _2555_ (.A(\mem[1][4] ),
    .B(net30),
    .S(net194),
    .Z(_0330_));
 MUX2_X1 _2556_ (.A(\mem[1][5] ),
    .B(net31),
    .S(net194),
    .Z(_0331_));
 MUX2_X1 _2557_ (.A(\mem[1][6] ),
    .B(net32),
    .S(net194),
    .Z(_0332_));
 MUX2_X1 _2558_ (.A(\mem[1][7] ),
    .B(net33),
    .S(net194),
    .Z(_0333_));
 MUX2_X1 _2559_ (.A(\mem[1][8] ),
    .B(net34),
    .S(net194),
    .Z(_0334_));
 MUX2_X1 _2560_ (.A(\mem[1][9] ),
    .B(net35),
    .S(net194),
    .Z(_0335_));
 AND2_X1 _2561_ (.A1(_0021_),
    .A2(_0635_),
    .ZN(_0740_));
 BUF_X2 place208 (.A(_0783_),
    .Z(net208));
 BUF_X2 place205 (.A(_0000_),
    .Z(net205));
 MUX2_X1 _2564_ (.A(\mem[2][0] ),
    .B(net4),
    .S(net193),
    .Z(_0336_));
 MUX2_X1 _2565_ (.A(\mem[2][10] ),
    .B(net5),
    .S(_0740_),
    .Z(_0337_));
 MUX2_X1 _2566_ (.A(\mem[2][11] ),
    .B(net6),
    .S(_0740_),
    .Z(_0338_));
 MUX2_X1 _2567_ (.A(\mem[2][12] ),
    .B(net7),
    .S(_0740_),
    .Z(_0339_));
 MUX2_X1 _2568_ (.A(\mem[2][13] ),
    .B(net8),
    .S(net193),
    .Z(_0340_));
 MUX2_X1 _2569_ (.A(\mem[2][14] ),
    .B(net9),
    .S(_0740_),
    .Z(_0341_));
 MUX2_X1 _2570_ (.A(\mem[2][15] ),
    .B(net10),
    .S(_0740_),
    .Z(_0342_));
 MUX2_X1 _2571_ (.A(\mem[2][16] ),
    .B(net11),
    .S(_0740_),
    .Z(_0343_));
 MUX2_X1 _2572_ (.A(\mem[2][17] ),
    .B(net12),
    .S(net193),
    .Z(_0344_));
 MUX2_X1 _2573_ (.A(\mem[2][18] ),
    .B(net13),
    .S(net193),
    .Z(_0345_));
 BUF_X2 place200 (.A(_0002_),
    .Z(net200));
 MUX2_X1 _2575_ (.A(\mem[2][19] ),
    .B(net14),
    .S(net193),
    .Z(_0346_));
 MUX2_X1 _2576_ (.A(\mem[2][1] ),
    .B(net15),
    .S(_0740_),
    .Z(_0347_));
 MUX2_X1 _2577_ (.A(\mem[2][20] ),
    .B(net16),
    .S(_0740_),
    .Z(_0348_));
 MUX2_X1 _2578_ (.A(\mem[2][21] ),
    .B(net17),
    .S(_0740_),
    .Z(_0349_));
 MUX2_X1 _2579_ (.A(\mem[2][22] ),
    .B(net18),
    .S(_0740_),
    .Z(_0350_));
 MUX2_X1 _2580_ (.A(\mem[2][23] ),
    .B(net19),
    .S(_0740_),
    .Z(_0351_));
 MUX2_X1 _2581_ (.A(\mem[2][24] ),
    .B(net20),
    .S(_0740_),
    .Z(_0352_));
 MUX2_X1 _2582_ (.A(\mem[2][25] ),
    .B(net21),
    .S(net193),
    .Z(_0353_));
 MUX2_X1 _2583_ (.A(\mem[2][26] ),
    .B(net22),
    .S(_0740_),
    .Z(_0354_));
 MUX2_X1 _2584_ (.A(\mem[2][27] ),
    .B(net23),
    .S(net193),
    .Z(_0355_));
 BUF_X1 place199 (.A(last_valid_data_available),
    .Z(net199));
 MUX2_X1 _2586_ (.A(\mem[2][28] ),
    .B(net24),
    .S(_0740_),
    .Z(_0356_));
 MUX2_X1 _2587_ (.A(\mem[2][29] ),
    .B(net25),
    .S(net193),
    .Z(_0357_));
 MUX2_X1 _2588_ (.A(\mem[2][2] ),
    .B(net26),
    .S(net193),
    .Z(_0358_));
 MUX2_X1 _2589_ (.A(\mem[2][30] ),
    .B(net27),
    .S(net193),
    .Z(_0359_));
 MUX2_X1 _2590_ (.A(\mem[2][31] ),
    .B(net28),
    .S(net193),
    .Z(_0360_));
 MUX2_X1 _2591_ (.A(\mem[2][3] ),
    .B(net29),
    .S(net193),
    .Z(_0361_));
 MUX2_X1 _2592_ (.A(\mem[2][4] ),
    .B(net30),
    .S(net193),
    .Z(_0362_));
 MUX2_X1 _2593_ (.A(\mem[2][5] ),
    .B(net31),
    .S(net193),
    .Z(_0363_));
 MUX2_X1 _2594_ (.A(\mem[2][6] ),
    .B(net32),
    .S(net193),
    .Z(_0364_));
 MUX2_X1 _2595_ (.A(\mem[2][7] ),
    .B(net33),
    .S(net193),
    .Z(_0365_));
 MUX2_X1 _2596_ (.A(\mem[2][8] ),
    .B(net34),
    .S(net193),
    .Z(_0366_));
 MUX2_X1 _2597_ (.A(\mem[2][9] ),
    .B(net35),
    .S(net193),
    .Z(_0367_));
 AND2_X1 _2598_ (.A1(_0023_),
    .A2(_0635_),
    .ZN(_0745_));
 BUF_X1 place196 (.A(_0636_),
    .Z(net196));
 BUF_X1 place195 (.A(_0705_),
    .Z(net195));
 MUX2_X1 _2601_ (.A(\mem[3][0] ),
    .B(net4),
    .S(net191),
    .Z(_0368_));
 MUX2_X1 _2602_ (.A(\mem[3][10] ),
    .B(net5),
    .S(_0745_),
    .Z(_0369_));
 MUX2_X1 _2603_ (.A(\mem[3][11] ),
    .B(net6),
    .S(net191),
    .Z(_0370_));
 MUX2_X1 _2604_ (.A(\mem[3][12] ),
    .B(net7),
    .S(_0745_),
    .Z(_0371_));
 MUX2_X1 _2605_ (.A(\mem[3][13] ),
    .B(net8),
    .S(net191),
    .Z(_0372_));
 MUX2_X1 _2606_ (.A(\mem[3][14] ),
    .B(net9),
    .S(_0745_),
    .Z(_0373_));
 MUX2_X1 _2607_ (.A(\mem[3][15] ),
    .B(net10),
    .S(_0745_),
    .Z(_0374_));
 MUX2_X1 _2608_ (.A(\mem[3][16] ),
    .B(net11),
    .S(_0745_),
    .Z(_0375_));
 MUX2_X1 _2609_ (.A(\mem[3][17] ),
    .B(net12),
    .S(net192),
    .Z(_0376_));
 MUX2_X1 _2610_ (.A(\mem[3][18] ),
    .B(net13),
    .S(net191),
    .Z(_0377_));
 BUF_X4 place194 (.A(_0735_),
    .Z(net194));
 MUX2_X1 _2612_ (.A(\mem[3][19] ),
    .B(net14),
    .S(net192),
    .Z(_0378_));
 MUX2_X1 _2613_ (.A(\mem[3][1] ),
    .B(net15),
    .S(_0745_),
    .Z(_0379_));
 MUX2_X1 _2614_ (.A(\mem[3][20] ),
    .B(net16),
    .S(_0745_),
    .Z(_0380_));
 MUX2_X1 _2615_ (.A(\mem[3][21] ),
    .B(net17),
    .S(_0745_),
    .Z(_0381_));
 MUX2_X1 _2616_ (.A(\mem[3][22] ),
    .B(net18),
    .S(_0745_),
    .Z(_0382_));
 MUX2_X1 _2617_ (.A(\mem[3][23] ),
    .B(net19),
    .S(_0745_),
    .Z(_0383_));
 MUX2_X1 _2618_ (.A(\mem[3][24] ),
    .B(net20),
    .S(_0745_),
    .Z(_0384_));
 MUX2_X1 _2619_ (.A(\mem[3][25] ),
    .B(net21),
    .S(net192),
    .Z(_0385_));
 MUX2_X1 _2620_ (.A(\mem[3][26] ),
    .B(net22),
    .S(_0745_),
    .Z(_0386_));
 MUX2_X1 _2621_ (.A(\mem[3][27] ),
    .B(net23),
    .S(net192),
    .Z(_0387_));
 BUF_X1 place202 (.A(_0002_),
    .Z(net202));
 MUX2_X1 _2623_ (.A(\mem[3][28] ),
    .B(net24),
    .S(_0745_),
    .Z(_0388_));
 MUX2_X1 _2624_ (.A(\mem[3][29] ),
    .B(net25),
    .S(net192),
    .Z(_0389_));
 MUX2_X1 _2625_ (.A(\mem[3][2] ),
    .B(net26),
    .S(net192),
    .Z(_0390_));
 MUX2_X1 _2626_ (.A(\mem[3][30] ),
    .B(net27),
    .S(net192),
    .Z(_0391_));
 MUX2_X1 _2627_ (.A(\mem[3][31] ),
    .B(net28),
    .S(net192),
    .Z(_0392_));
 MUX2_X1 _2628_ (.A(\mem[3][3] ),
    .B(net29),
    .S(net192),
    .Z(_0393_));
 MUX2_X1 _2629_ (.A(\mem[3][4] ),
    .B(net30),
    .S(net192),
    .Z(_0394_));
 MUX2_X1 _2630_ (.A(\mem[3][5] ),
    .B(net31),
    .S(net191),
    .Z(_0395_));
 MUX2_X1 _2631_ (.A(\mem[3][6] ),
    .B(net32),
    .S(net191),
    .Z(_0396_));
 MUX2_X1 _2632_ (.A(\mem[3][7] ),
    .B(net33),
    .S(net191),
    .Z(_0397_));
 MUX2_X1 _2633_ (.A(\mem[3][8] ),
    .B(net34),
    .S(net191),
    .Z(_0398_));
 MUX2_X1 _2634_ (.A(\mem[3][9] ),
    .B(net35),
    .S(net191),
    .Z(_0399_));
 AND2_X1 _2635_ (.A1(_0704_),
    .A2(_0715_),
    .ZN(_0750_));
 AND2_X1 _2636_ (.A1(_0019_),
    .A2(_0750_),
    .ZN(_0751_));
 BUF_X1 place191 (.A(_0745_),
    .Z(net191));
 BUF_X2 place190 (.A(_0883_),
    .Z(net190));
 MUX2_X1 _2639_ (.A(\mem[4][0] ),
    .B(net4),
    .S(net181),
    .Z(_0400_));
 MUX2_X1 _2640_ (.A(\mem[4][10] ),
    .B(net5),
    .S(net181),
    .Z(_0401_));
 MUX2_X1 _2641_ (.A(\mem[4][11] ),
    .B(net6),
    .S(net181),
    .Z(_0402_));
 MUX2_X1 _2642_ (.A(\mem[4][12] ),
    .B(net7),
    .S(net181),
    .Z(_0403_));
 MUX2_X1 _2643_ (.A(\mem[4][13] ),
    .B(net8),
    .S(net181),
    .Z(_0404_));
 MUX2_X1 _2644_ (.A(\mem[4][14] ),
    .B(net9),
    .S(net181),
    .Z(_0405_));
 MUX2_X1 _2645_ (.A(\mem[4][15] ),
    .B(net10),
    .S(net181),
    .Z(_0406_));
 MUX2_X1 _2646_ (.A(\mem[4][16] ),
    .B(net11),
    .S(net181),
    .Z(_0407_));
 MUX2_X1 _2647_ (.A(\mem[4][17] ),
    .B(net12),
    .S(net181),
    .Z(_0408_));
 MUX2_X1 _2648_ (.A(\mem[4][18] ),
    .B(net13),
    .S(net181),
    .Z(_0409_));
 BUF_X2 place189 (.A(_0892_),
    .Z(net189));
 MUX2_X1 _2650_ (.A(\mem[4][19] ),
    .B(net14),
    .S(net181),
    .Z(_0410_));
 MUX2_X1 _2651_ (.A(\mem[4][1] ),
    .B(net15),
    .S(net181),
    .Z(_0411_));
 MUX2_X1 _2652_ (.A(\mem[4][20] ),
    .B(net16),
    .S(net181),
    .Z(_0412_));
 MUX2_X1 _2653_ (.A(\mem[4][21] ),
    .B(net17),
    .S(net181),
    .Z(_0413_));
 MUX2_X1 _2654_ (.A(\mem[4][22] ),
    .B(net18),
    .S(net181),
    .Z(_0414_));
 MUX2_X1 _2655_ (.A(\mem[4][23] ),
    .B(net19),
    .S(net181),
    .Z(_0415_));
 MUX2_X1 _2656_ (.A(\mem[4][24] ),
    .B(net20),
    .S(net181),
    .Z(_0416_));
 MUX2_X1 _2657_ (.A(\mem[4][25] ),
    .B(net21),
    .S(net181),
    .Z(_0417_));
 MUX2_X1 _2658_ (.A(\mem[4][26] ),
    .B(net22),
    .S(net181),
    .Z(_0418_));
 MUX2_X1 _2659_ (.A(\mem[4][27] ),
    .B(net23),
    .S(net181),
    .Z(_0419_));
 BUF_X2 place188 (.A(_0894_),
    .Z(net188));
 MUX2_X1 _2661_ (.A(\mem[4][28] ),
    .B(net24),
    .S(net181),
    .Z(_0420_));
 MUX2_X1 _2662_ (.A(\mem[4][29] ),
    .B(net25),
    .S(net181),
    .Z(_0421_));
 MUX2_X1 _2663_ (.A(\mem[4][2] ),
    .B(net26),
    .S(net181),
    .Z(_0422_));
 MUX2_X1 _2664_ (.A(\mem[4][30] ),
    .B(net27),
    .S(net181),
    .Z(_0423_));
 MUX2_X1 _2665_ (.A(\mem[4][31] ),
    .B(net28),
    .S(net181),
    .Z(_0424_));
 MUX2_X1 _2666_ (.A(\mem[4][3] ),
    .B(net29),
    .S(net181),
    .Z(_0425_));
 MUX2_X1 _2667_ (.A(\mem[4][4] ),
    .B(net30),
    .S(net181),
    .Z(_0426_));
 MUX2_X1 _2668_ (.A(\mem[4][5] ),
    .B(net31),
    .S(net181),
    .Z(_0427_));
 MUX2_X1 _2669_ (.A(\mem[4][6] ),
    .B(net32),
    .S(net181),
    .Z(_0428_));
 MUX2_X1 _2670_ (.A(\mem[4][7] ),
    .B(net33),
    .S(net181),
    .Z(_0429_));
 MUX2_X1 _2671_ (.A(\mem[4][8] ),
    .B(net34),
    .S(net181),
    .Z(_0430_));
 MUX2_X1 _2672_ (.A(\mem[4][9] ),
    .B(net35),
    .S(net181),
    .Z(_0431_));
 AND2_X1 _2673_ (.A1(_0022_),
    .A2(_0750_),
    .ZN(_0756_));
 BUF_X1 place187 (.A(_0706_),
    .Z(net187));
 BUF_X1 place186 (.A(_0711_),
    .Z(net186));
 MUX2_X1 _2676_ (.A(\mem[5][0] ),
    .B(net4),
    .S(net180),
    .Z(_0432_));
 MUX2_X1 _2677_ (.A(\mem[5][10] ),
    .B(net5),
    .S(net180),
    .Z(_0433_));
 MUX2_X1 _2678_ (.A(\mem[5][11] ),
    .B(net6),
    .S(net180),
    .Z(_0434_));
 MUX2_X1 _2679_ (.A(\mem[5][12] ),
    .B(net7),
    .S(net180),
    .Z(_0435_));
 MUX2_X1 _2680_ (.A(\mem[5][13] ),
    .B(net8),
    .S(net180),
    .Z(_0436_));
 MUX2_X1 _2681_ (.A(\mem[5][14] ),
    .B(net9),
    .S(net180),
    .Z(_0437_));
 MUX2_X1 _2682_ (.A(\mem[5][15] ),
    .B(net10),
    .S(net180),
    .Z(_0438_));
 MUX2_X1 _2683_ (.A(\mem[5][16] ),
    .B(net11),
    .S(net180),
    .Z(_0439_));
 MUX2_X1 _2684_ (.A(\mem[5][17] ),
    .B(net12),
    .S(net180),
    .Z(_0440_));
 MUX2_X1 _2685_ (.A(\mem[5][18] ),
    .B(net13),
    .S(net180),
    .Z(_0441_));
 BUF_X1 place185 (.A(_0718_),
    .Z(net185));
 MUX2_X1 _2687_ (.A(\mem[5][19] ),
    .B(net14),
    .S(net180),
    .Z(_0442_));
 MUX2_X1 _2688_ (.A(\mem[5][1] ),
    .B(net15),
    .S(net180),
    .Z(_0443_));
 MUX2_X1 _2689_ (.A(\mem[5][20] ),
    .B(net16),
    .S(net180),
    .Z(_0444_));
 MUX2_X1 _2690_ (.A(\mem[5][21] ),
    .B(net17),
    .S(net180),
    .Z(_0445_));
 MUX2_X1 _2691_ (.A(\mem[5][22] ),
    .B(net18),
    .S(net180),
    .Z(_0446_));
 MUX2_X1 _2692_ (.A(\mem[5][23] ),
    .B(net19),
    .S(net180),
    .Z(_0447_));
 MUX2_X1 _2693_ (.A(\mem[5][24] ),
    .B(net20),
    .S(net180),
    .Z(_0448_));
 MUX2_X1 _2694_ (.A(\mem[5][25] ),
    .B(net21),
    .S(net180),
    .Z(_0449_));
 MUX2_X1 _2695_ (.A(\mem[5][26] ),
    .B(net22),
    .S(net180),
    .Z(_0450_));
 MUX2_X1 _2696_ (.A(\mem[5][27] ),
    .B(net23),
    .S(net180),
    .Z(_0451_));
 BUF_X1 place184 (.A(_0723_),
    .Z(net184));
 MUX2_X1 _2698_ (.A(\mem[5][28] ),
    .B(net24),
    .S(net180),
    .Z(_0452_));
 MUX2_X1 _2699_ (.A(\mem[5][29] ),
    .B(net25),
    .S(net180),
    .Z(_0453_));
 MUX2_X1 _2700_ (.A(\mem[5][2] ),
    .B(net26),
    .S(net180),
    .Z(_0454_));
 MUX2_X1 _2701_ (.A(\mem[5][30] ),
    .B(net27),
    .S(net180),
    .Z(_0455_));
 MUX2_X1 _2702_ (.A(\mem[5][31] ),
    .B(net28),
    .S(net180),
    .Z(_0456_));
 MUX2_X1 _2703_ (.A(\mem[5][3] ),
    .B(net29),
    .S(net180),
    .Z(_0457_));
 MUX2_X1 _2704_ (.A(\mem[5][4] ),
    .B(net30),
    .S(net180),
    .Z(_0458_));
 MUX2_X1 _2705_ (.A(\mem[5][5] ),
    .B(net31),
    .S(net180),
    .Z(_0459_));
 MUX2_X1 _2706_ (.A(\mem[5][6] ),
    .B(net32),
    .S(net180),
    .Z(_0460_));
 MUX2_X1 _2707_ (.A(\mem[5][7] ),
    .B(net33),
    .S(net180),
    .Z(_0461_));
 MUX2_X1 _2708_ (.A(\mem[5][8] ),
    .B(net34),
    .S(net180),
    .Z(_0462_));
 MUX2_X1 _2709_ (.A(\mem[5][9] ),
    .B(net35),
    .S(net180),
    .Z(_0463_));
 AND2_X1 _2710_ (.A1(_0021_),
    .A2(_0750_),
    .ZN(_0761_));
 BUF_X2 place183 (.A(_0727_),
    .Z(net183));
 BUF_X1 place182 (.A(_0731_),
    .Z(net182));
 MUX2_X1 _2713_ (.A(\mem[6][0] ),
    .B(net4),
    .S(net179),
    .Z(_0464_));
 MUX2_X1 _2714_ (.A(\mem[6][10] ),
    .B(net5),
    .S(net179),
    .Z(_0465_));
 MUX2_X1 _2715_ (.A(\mem[6][11] ),
    .B(net6),
    .S(net179),
    .Z(_0466_));
 MUX2_X1 _2716_ (.A(\mem[6][12] ),
    .B(net7),
    .S(net179),
    .Z(_0467_));
 MUX2_X1 _2717_ (.A(\mem[6][13] ),
    .B(net8),
    .S(net179),
    .Z(_0468_));
 MUX2_X1 _2718_ (.A(\mem[6][14] ),
    .B(net9),
    .S(net179),
    .Z(_0469_));
 MUX2_X1 _2719_ (.A(\mem[6][15] ),
    .B(net10),
    .S(net179),
    .Z(_0470_));
 MUX2_X1 _2720_ (.A(\mem[6][16] ),
    .B(net11),
    .S(net179),
    .Z(_0471_));
 MUX2_X1 _2721_ (.A(\mem[6][17] ),
    .B(net12),
    .S(net179),
    .Z(_0472_));
 MUX2_X1 _2722_ (.A(\mem[6][18] ),
    .B(net13),
    .S(net179),
    .Z(_0473_));
 BUF_X4 place181 (.A(_0751_),
    .Z(net181));
 MUX2_X1 _2724_ (.A(\mem[6][19] ),
    .B(net14),
    .S(net179),
    .Z(_0474_));
 MUX2_X1 _2725_ (.A(\mem[6][1] ),
    .B(net15),
    .S(_0761_),
    .Z(_0475_));
 MUX2_X1 _2726_ (.A(\mem[6][20] ),
    .B(net16),
    .S(_0761_),
    .Z(_0476_));
 MUX2_X1 _2727_ (.A(\mem[6][21] ),
    .B(net17),
    .S(_0761_),
    .Z(_0477_));
 MUX2_X1 _2728_ (.A(\mem[6][22] ),
    .B(net18),
    .S(_0761_),
    .Z(_0478_));
 MUX2_X1 _2729_ (.A(\mem[6][23] ),
    .B(net19),
    .S(_0761_),
    .Z(_0479_));
 MUX2_X1 _2730_ (.A(\mem[6][24] ),
    .B(net20),
    .S(_0761_),
    .Z(_0480_));
 MUX2_X1 _2731_ (.A(\mem[6][25] ),
    .B(net21),
    .S(_0761_),
    .Z(_0481_));
 MUX2_X1 _2732_ (.A(\mem[6][26] ),
    .B(net22),
    .S(_0761_),
    .Z(_0482_));
 MUX2_X1 _2733_ (.A(\mem[6][27] ),
    .B(net23),
    .S(net179),
    .Z(_0483_));
 BUF_X4 place180 (.A(_0756_),
    .Z(net180));
 MUX2_X1 _2735_ (.A(\mem[6][28] ),
    .B(net24),
    .S(_0761_),
    .Z(_0484_));
 MUX2_X1 _2736_ (.A(\mem[6][29] ),
    .B(net25),
    .S(_0761_),
    .Z(_0485_));
 MUX2_X1 _2737_ (.A(\mem[6][2] ),
    .B(net26),
    .S(_0761_),
    .Z(_0486_));
 MUX2_X1 _2738_ (.A(\mem[6][30] ),
    .B(net27),
    .S(_0761_),
    .Z(_0487_));
 MUX2_X1 _2739_ (.A(\mem[6][31] ),
    .B(net28),
    .S(net179),
    .Z(_0488_));
 MUX2_X1 _2740_ (.A(\mem[6][3] ),
    .B(net29),
    .S(net179),
    .Z(_0489_));
 MUX2_X1 _2741_ (.A(\mem[6][4] ),
    .B(net30),
    .S(net179),
    .Z(_0490_));
 MUX2_X1 _2742_ (.A(\mem[6][5] ),
    .B(net31),
    .S(net179),
    .Z(_0491_));
 MUX2_X1 _2743_ (.A(\mem[6][6] ),
    .B(net32),
    .S(net179),
    .Z(_0492_));
 MUX2_X1 _2744_ (.A(\mem[6][7] ),
    .B(net33),
    .S(net179),
    .Z(_0493_));
 MUX2_X1 _2745_ (.A(\mem[6][8] ),
    .B(net34),
    .S(net179),
    .Z(_0494_));
 MUX2_X1 _2746_ (.A(\mem[6][9] ),
    .B(net35),
    .S(net179),
    .Z(_0495_));
 AND2_X1 _2747_ (.A1(_0023_),
    .A2(_0750_),
    .ZN(_0766_));
 BUF_X2 place179 (.A(_0761_),
    .Z(net179));
 BUF_X1 place177 (.A(_0766_),
    .Z(net177));
 MUX2_X1 _2750_ (.A(\mem[7][0] ),
    .B(net4),
    .S(net177),
    .Z(_0496_));
 MUX2_X1 _2751_ (.A(\mem[7][10] ),
    .B(net5),
    .S(_0766_),
    .Z(_0497_));
 MUX2_X1 _2752_ (.A(\mem[7][11] ),
    .B(net6),
    .S(net177),
    .Z(_0498_));
 MUX2_X1 _2753_ (.A(\mem[7][12] ),
    .B(net7),
    .S(_0766_),
    .Z(_0499_));
 MUX2_X1 _2754_ (.A(\mem[7][13] ),
    .B(net8),
    .S(net177),
    .Z(_0500_));
 MUX2_X1 _2755_ (.A(\mem[7][14] ),
    .B(net9),
    .S(_0766_),
    .Z(_0501_));
 MUX2_X1 _2756_ (.A(\mem[7][15] ),
    .B(net10),
    .S(_0766_),
    .Z(_0502_));
 MUX2_X1 _2757_ (.A(\mem[7][16] ),
    .B(net11),
    .S(_0766_),
    .Z(_0503_));
 MUX2_X1 _2758_ (.A(\mem[7][17] ),
    .B(net12),
    .S(net178),
    .Z(_0504_));
 MUX2_X1 _2759_ (.A(\mem[7][18] ),
    .B(net13),
    .S(net177),
    .Z(_0505_));
 BUF_X2 place193 (.A(_0740_),
    .Z(net193));
 MUX2_X1 _2761_ (.A(\mem[7][19] ),
    .B(net14),
    .S(net178),
    .Z(_0506_));
 MUX2_X1 _2762_ (.A(\mem[7][1] ),
    .B(net15),
    .S(_0766_),
    .Z(_0507_));
 MUX2_X1 _2763_ (.A(\mem[7][20] ),
    .B(net16),
    .S(_0766_),
    .Z(_0508_));
 MUX2_X1 _2764_ (.A(\mem[7][21] ),
    .B(net17),
    .S(_0766_),
    .Z(_0509_));
 MUX2_X1 _2765_ (.A(\mem[7][22] ),
    .B(net18),
    .S(_0766_),
    .Z(_0510_));
 MUX2_X1 _2766_ (.A(\mem[7][23] ),
    .B(net19),
    .S(_0766_),
    .Z(_0511_));
 MUX2_X1 _2767_ (.A(\mem[7][24] ),
    .B(net20),
    .S(_0766_),
    .Z(_0512_));
 MUX2_X1 _2768_ (.A(\mem[7][25] ),
    .B(net21),
    .S(net178),
    .Z(_0513_));
 MUX2_X1 _2769_ (.A(\mem[7][26] ),
    .B(net22),
    .S(_0766_),
    .Z(_0514_));
 MUX2_X1 _2770_ (.A(\mem[7][27] ),
    .B(net23),
    .S(net178),
    .Z(_0515_));
 BUF_X1 place176 (.A(_0771_),
    .Z(net176));
 MUX2_X1 _2772_ (.A(\mem[7][28] ),
    .B(net24),
    .S(_0766_),
    .Z(_0516_));
 MUX2_X1 _2773_ (.A(\mem[7][29] ),
    .B(net25),
    .S(net178),
    .Z(_0517_));
 MUX2_X1 _2774_ (.A(\mem[7][2] ),
    .B(net26),
    .S(net178),
    .Z(_0518_));
 MUX2_X1 _2775_ (.A(\mem[7][30] ),
    .B(net27),
    .S(net178),
    .Z(_0519_));
 MUX2_X1 _2776_ (.A(\mem[7][31] ),
    .B(net28),
    .S(net178),
    .Z(_0520_));
 MUX2_X1 _2777_ (.A(\mem[7][3] ),
    .B(net29),
    .S(net178),
    .Z(_0521_));
 MUX2_X1 _2778_ (.A(\mem[7][4] ),
    .B(net30),
    .S(net178),
    .Z(_0522_));
 MUX2_X1 _2779_ (.A(\mem[7][5] ),
    .B(net31),
    .S(net177),
    .Z(_0523_));
 MUX2_X1 _2780_ (.A(\mem[7][6] ),
    .B(net32),
    .S(net177),
    .Z(_0524_));
 MUX2_X1 _2781_ (.A(\mem[7][7] ),
    .B(net33),
    .S(net177),
    .Z(_0525_));
 MUX2_X1 _2782_ (.A(\mem[7][8] ),
    .B(net34),
    .S(net177),
    .Z(_0526_));
 MUX2_X1 _2783_ (.A(\mem[7][9] ),
    .B(net35),
    .S(net177),
    .Z(_0527_));
 NAND2_X2 _2784_ (.A1(_0019_),
    .A2(net195),
    .ZN(_0771_));
 BUF_X1 place175 (.A(_0775_),
    .Z(net175));
 MUX2_X1 _2786_ (.A(net4),
    .B(\mem[8][0] ),
    .S(_0771_),
    .Z(_0528_));
 MUX2_X1 _2787_ (.A(net5),
    .B(\mem[8][10] ),
    .S(net176),
    .Z(_0529_));
 MUX2_X1 _2788_ (.A(net6),
    .B(\mem[8][11] ),
    .S(net176),
    .Z(_0530_));
 MUX2_X1 _2789_ (.A(net7),
    .B(\mem[8][12] ),
    .S(net176),
    .Z(_0531_));
 MUX2_X1 _2790_ (.A(net8),
    .B(\mem[8][13] ),
    .S(net176),
    .Z(_0532_));
 MUX2_X1 _2791_ (.A(net9),
    .B(\mem[8][14] ),
    .S(net176),
    .Z(_0533_));
 MUX2_X1 _2792_ (.A(net10),
    .B(\mem[8][15] ),
    .S(net176),
    .Z(_0534_));
 MUX2_X1 _2793_ (.A(net11),
    .B(\mem[8][16] ),
    .S(net176),
    .Z(_0535_));
 MUX2_X1 _2794_ (.A(net12),
    .B(\mem[8][17] ),
    .S(_0771_),
    .Z(_0536_));
 MUX2_X1 _2795_ (.A(net13),
    .B(\mem[8][18] ),
    .S(net176),
    .Z(_0537_));
 BUF_X1 output98 (.A(net98),
    .Z(wr_ready));
 MUX2_X1 _2797_ (.A(net14),
    .B(\mem[8][19] ),
    .S(_0771_),
    .Z(_0538_));
 MUX2_X1 _2798_ (.A(net15),
    .B(\mem[8][1] ),
    .S(_0771_),
    .Z(_0539_));
 MUX2_X1 _2799_ (.A(net16),
    .B(\mem[8][20] ),
    .S(_0771_),
    .Z(_0540_));
 MUX2_X1 _2800_ (.A(net17),
    .B(\mem[8][21] ),
    .S(_0771_),
    .Z(_0541_));
 MUX2_X1 _2801_ (.A(net18),
    .B(\mem[8][22] ),
    .S(_0771_),
    .Z(_0542_));
 MUX2_X1 _2802_ (.A(net19),
    .B(\mem[8][23] ),
    .S(_0771_),
    .Z(_0543_));
 MUX2_X1 _2803_ (.A(net20),
    .B(\mem[8][24] ),
    .S(_0771_),
    .Z(_0544_));
 MUX2_X1 _2804_ (.A(net21),
    .B(\mem[8][25] ),
    .S(_0771_),
    .Z(_0545_));
 MUX2_X1 _2805_ (.A(net22),
    .B(\mem[8][26] ),
    .S(_0771_),
    .Z(_0546_));
 MUX2_X1 _2806_ (.A(net23),
    .B(\mem[8][27] ),
    .S(_0771_),
    .Z(_0547_));
 BUF_X1 output97 (.A(net97),
    .Z(underflow_detected));
 MUX2_X1 _2808_ (.A(net24),
    .B(\mem[8][28] ),
    .S(_0771_),
    .Z(_0548_));
 MUX2_X1 _2809_ (.A(net25),
    .B(\mem[8][29] ),
    .S(_0771_),
    .Z(_0549_));
 MUX2_X1 _2810_ (.A(net26),
    .B(\mem[8][2] ),
    .S(_0771_),
    .Z(_0550_));
 MUX2_X1 _2811_ (.A(net27),
    .B(\mem[8][30] ),
    .S(_0771_),
    .Z(_0551_));
 MUX2_X1 _2812_ (.A(net28),
    .B(\mem[8][31] ),
    .S(_0771_),
    .Z(_0552_));
 MUX2_X1 _2813_ (.A(net29),
    .B(\mem[8][3] ),
    .S(_0771_),
    .Z(_0553_));
 MUX2_X1 _2814_ (.A(net30),
    .B(\mem[8][4] ),
    .S(_0771_),
    .Z(_0554_));
 MUX2_X1 _2815_ (.A(net31),
    .B(\mem[8][5] ),
    .S(_0771_),
    .Z(_0555_));
 MUX2_X1 _2816_ (.A(net32),
    .B(\mem[8][6] ),
    .S(_0771_),
    .Z(_0556_));
 MUX2_X1 _2817_ (.A(net33),
    .B(\mem[8][7] ),
    .S(net176),
    .Z(_0557_));
 MUX2_X1 _2818_ (.A(net34),
    .B(\mem[8][8] ),
    .S(_0771_),
    .Z(_0558_));
 MUX2_X1 _2819_ (.A(net35),
    .B(\mem[8][9] ),
    .S(net176),
    .Z(_0559_));
 NAND2_X2 _2820_ (.A1(_0022_),
    .A2(net195),
    .ZN(_0775_));
 BUF_X1 output96 (.A(net96),
    .Z(rd_valid));
 MUX2_X1 _2822_ (.A(net4),
    .B(\mem[9][0] ),
    .S(_0775_),
    .Z(_0560_));
 MUX2_X1 _2823_ (.A(net5),
    .B(\mem[9][10] ),
    .S(net175),
    .Z(_0561_));
 MUX2_X1 _2824_ (.A(net6),
    .B(\mem[9][11] ),
    .S(net175),
    .Z(_0562_));
 MUX2_X1 _2825_ (.A(net7),
    .B(\mem[9][12] ),
    .S(net175),
    .Z(_0563_));
 MUX2_X1 _2826_ (.A(net8),
    .B(\mem[9][13] ),
    .S(net175),
    .Z(_0564_));
 MUX2_X1 _2827_ (.A(net9),
    .B(\mem[9][14] ),
    .S(net175),
    .Z(_0565_));
 MUX2_X1 _2828_ (.A(net10),
    .B(\mem[9][15] ),
    .S(net175),
    .Z(_0566_));
 MUX2_X1 _2829_ (.A(net11),
    .B(\mem[9][16] ),
    .S(net175),
    .Z(_0567_));
 MUX2_X1 _2830_ (.A(net12),
    .B(\mem[9][17] ),
    .S(_0775_),
    .Z(_0568_));
 MUX2_X1 _2831_ (.A(net13),
    .B(\mem[9][18] ),
    .S(_0775_),
    .Z(_0569_));
 BUF_X1 output95 (.A(net95),
    .Z(rd_data[9]));
 MUX2_X1 _2833_ (.A(net14),
    .B(\mem[9][19] ),
    .S(_0775_),
    .Z(_0570_));
 MUX2_X1 _2834_ (.A(net15),
    .B(\mem[9][1] ),
    .S(_0775_),
    .Z(_0571_));
 MUX2_X1 _2835_ (.A(net16),
    .B(\mem[9][20] ),
    .S(_0775_),
    .Z(_0572_));
 MUX2_X1 _2836_ (.A(net17),
    .B(\mem[9][21] ),
    .S(_0775_),
    .Z(_0573_));
 MUX2_X1 _2837_ (.A(net18),
    .B(\mem[9][22] ),
    .S(_0775_),
    .Z(_0574_));
 MUX2_X1 _2838_ (.A(net19),
    .B(\mem[9][23] ),
    .S(_0775_),
    .Z(_0575_));
 MUX2_X1 _2839_ (.A(net20),
    .B(\mem[9][24] ),
    .S(_0775_),
    .Z(_0576_));
 MUX2_X1 _2840_ (.A(net21),
    .B(\mem[9][25] ),
    .S(_0775_),
    .Z(_0577_));
 MUX2_X1 _2841_ (.A(net22),
    .B(\mem[9][26] ),
    .S(_0775_),
    .Z(_0578_));
 MUX2_X1 _2842_ (.A(net23),
    .B(\mem[9][27] ),
    .S(_0775_),
    .Z(_0579_));
 BUF_X1 output94 (.A(net94),
    .Z(rd_data[8]));
 MUX2_X1 _2844_ (.A(net24),
    .B(\mem[9][28] ),
    .S(_0775_),
    .Z(_0580_));
 MUX2_X1 _2845_ (.A(net25),
    .B(\mem[9][29] ),
    .S(_0775_),
    .Z(_0581_));
 MUX2_X1 _2846_ (.A(net26),
    .B(\mem[9][2] ),
    .S(_0775_),
    .Z(_0582_));
 MUX2_X1 _2847_ (.A(net27),
    .B(\mem[9][30] ),
    .S(_0775_),
    .Z(_0583_));
 MUX2_X1 _2848_ (.A(net28),
    .B(\mem[9][31] ),
    .S(_0775_),
    .Z(_0584_));
 MUX2_X1 _2849_ (.A(net29),
    .B(\mem[9][3] ),
    .S(_0775_),
    .Z(_0585_));
 MUX2_X1 _2850_ (.A(net30),
    .B(\mem[9][4] ),
    .S(_0775_),
    .Z(_0586_));
 MUX2_X1 _2851_ (.A(net31),
    .B(\mem[9][5] ),
    .S(_0775_),
    .Z(_0587_));
 MUX2_X1 _2852_ (.A(net32),
    .B(\mem[9][6] ),
    .S(_0775_),
    .Z(_0588_));
 MUX2_X1 _2853_ (.A(net33),
    .B(\mem[9][7] ),
    .S(net175),
    .Z(_0589_));
 MUX2_X1 _2854_ (.A(net34),
    .B(\mem[9][8] ),
    .S(_0775_),
    .Z(_0590_));
 MUX2_X1 _2855_ (.A(net35),
    .B(\mem[9][9] ),
    .S(net175),
    .Z(_0591_));
 BUF_X1 output93 (.A(net93),
    .Z(rd_data[7]));
 AND2_X1 _2857_ (.A1(\rd_ptr[0] ),
    .A2(net3),
    .ZN(_0780_));
 BUF_X1 output92 (.A(net92),
    .Z(rd_data[6]));
 OAI21_X1 _2859_ (.A(_0780_),
    .B1(net172),
    .B2(_0629_),
    .ZN(_0782_));
 INV_X2 _2860_ (.A(net3),
    .ZN(_0783_));
 BUF_X1 output91 (.A(net91),
    .Z(rd_data[5]));
 OR2_X1 _2862_ (.A1(\rd_ptr[0] ),
    .A2(_0783_),
    .ZN(_0785_));
 BUF_X1 output90 (.A(net90),
    .Z(rd_data[4]));
 NAND2_X1 _2864_ (.A1(net210),
    .A2(net96),
    .ZN(_0787_));
 OAI21_X1 _2865_ (.A(_0782_),
    .B1(_0785_),
    .B2(_0787_),
    .ZN(_0026_));
 BUF_X1 output89 (.A(net89),
    .Z(rd_data[3]));
 BUF_X1 output88 (.A(net88),
    .Z(rd_data[31]));
 NAND3_X1 _2868_ (.A1(net210),
    .A2(_0015_),
    .A3(net96),
    .ZN(_0790_));
 OAI21_X1 _2869_ (.A(\rd_ptr[1] ),
    .B1(net172),
    .B2(_0629_),
    .ZN(_0791_));
 AOI21_X1 _2870_ (.A(_0783_),
    .B1(_0790_),
    .B2(_0791_),
    .ZN(_0027_));
 NOR2_X1 _2871_ (.A1(\rd_ptr[2] ),
    .A2(_0783_),
    .ZN(_0792_));
 AND2_X1 _2872_ (.A1(\rd_ptr[2] ),
    .A2(net3),
    .ZN(_0793_));
 NAND3_X1 _2873_ (.A1(net210),
    .A2(_0014_),
    .A3(net96),
    .ZN(_0794_));
 MUX2_X1 _2874_ (.A(_0792_),
    .B(_0793_),
    .S(_0794_),
    .Z(_0028_));
 NAND4_X1 _2875_ (.A1(net210),
    .A2(\rd_ptr[0] ),
    .A3(\rd_ptr[1] ),
    .A4(\rd_ptr[2] ),
    .ZN(_0795_));
 OAI21_X1 _2876_ (.A(\rd_ptr[3] ),
    .B1(net172),
    .B2(_0795_),
    .ZN(_0796_));
 OR3_X1 _2877_ (.A1(\rd_ptr[3] ),
    .A2(net172),
    .A3(_0795_),
    .ZN(_0797_));
 AOI21_X1 _2878_ (.A(net208),
    .B1(_0796_),
    .B2(_0797_),
    .ZN(_0029_));
 BUF_X1 output87 (.A(net87),
    .Z(rd_data[30]));
 BUF_X1 output86 (.A(net86),
    .Z(rd_data[2]));
 BUF_X1 output85 (.A(net85),
    .Z(rd_data[29]));
 NAND4_X1 _2882_ (.A1(net2),
    .A2(_0005_),
    .A3(net3),
    .A4(net44),
    .ZN(_0801_));
 NAND2_X1 _2883_ (.A1(net45),
    .A2(net3),
    .ZN(_0802_));
 OAI21_X1 _2884_ (.A(_0801_),
    .B1(_0802_),
    .B2(net97),
    .ZN(_0030_));
 BUF_X1 output84 (.A(net84),
    .Z(rd_data[28]));
 AND2_X1 _2886_ (.A1(net46),
    .A2(net3),
    .ZN(_0804_));
 NOR2_X1 _2887_ (.A1(net46),
    .A2(_0783_),
    .ZN(_0805_));
 INV_X1 _2888_ (.A(net60),
    .ZN(_0806_));
 BUF_X1 output83 (.A(net83),
    .Z(rd_data[27]));
 BUF_X1 output82 (.A(net82),
    .Z(rd_data[26]));
 NAND4_X2 _2891_ (.A1(net56),
    .A2(net57),
    .A3(net58),
    .A4(net59),
    .ZN(_0809_));
 NAND2_X1 _2892_ (.A1(net2),
    .A2(net53),
    .ZN(_0810_));
 BUF_X1 output81 (.A(net81),
    .Z(rd_data[25]));
 BUF_X1 output80 (.A(net80),
    .Z(rd_data[24]));
 NAND3_X1 _2895_ (.A1(_0016_),
    .A2(net54),
    .A3(net55),
    .ZN(_0813_));
 OR2_X1 _2896_ (.A1(_0810_),
    .A2(_0813_),
    .ZN(_0814_));
 NOR4_X4 _2897_ (.A1(_0806_),
    .A2(net96),
    .A3(_0809_),
    .A4(_0814_),
    .ZN(_0815_));
 MUX2_X1 _2898_ (.A(_0804_),
    .B(_0805_),
    .S(_0815_),
    .Z(_0031_));
 AND2_X1 _2899_ (.A1(net2),
    .A2(net53),
    .ZN(_0816_));
 AND4_X1 _2900_ (.A1(net52),
    .A2(net45),
    .A3(net54),
    .A4(net55),
    .ZN(_0817_));
 NAND2_X1 _2901_ (.A1(_0816_),
    .A2(_0817_),
    .ZN(_0818_));
 INV_X1 _2902_ (.A(_0818_),
    .ZN(_0819_));
 OAI211_X2 _2903_ (.A(_0617_),
    .B(_0819_),
    .C1(_0622_),
    .C2(_0620_),
    .ZN(_0820_));
 NOR2_X1 _2904_ (.A1(_0806_),
    .A2(_0809_),
    .ZN(_0821_));
 NAND2_X1 _2905_ (.A1(net46),
    .A2(_0821_),
    .ZN(_0822_));
 OAI21_X1 _2906_ (.A(net47),
    .B1(_0820_),
    .B2(_0822_),
    .ZN(_0823_));
 OR3_X1 _2907_ (.A1(net47),
    .A2(_0820_),
    .A3(_0822_),
    .ZN(_0824_));
 AOI21_X1 _2908_ (.A(_0783_),
    .B1(_0823_),
    .B2(_0824_),
    .ZN(_0032_));
 AND2_X1 _2909_ (.A1(net48),
    .A2(net3),
    .ZN(_0825_));
 NOR2_X1 _2910_ (.A1(net48),
    .A2(_0783_),
    .ZN(_0826_));
 NAND3_X1 _2911_ (.A1(net46),
    .A2(net47),
    .A3(_0821_),
    .ZN(_0827_));
 NOR3_X1 _2912_ (.A1(net96),
    .A2(_0814_),
    .A3(_0827_),
    .ZN(_0828_));
 MUX2_X1 _2913_ (.A(_0825_),
    .B(_0826_),
    .S(_0828_),
    .Z(_0033_));
 NAND4_X1 _2914_ (.A1(net46),
    .A2(net47),
    .A3(net48),
    .A4(_0821_),
    .ZN(_0829_));
 OAI21_X1 _2915_ (.A(net49),
    .B1(_0820_),
    .B2(_0829_),
    .ZN(_0830_));
 OR3_X1 _2916_ (.A1(net49),
    .A2(_0820_),
    .A3(_0829_),
    .ZN(_0831_));
 AOI21_X1 _2917_ (.A(_0783_),
    .B1(_0830_),
    .B2(_0831_),
    .ZN(_0034_));
 AND2_X1 _2918_ (.A1(net50),
    .A2(net3),
    .ZN(_0832_));
 NOR2_X1 _2919_ (.A1(net50),
    .A2(_0783_),
    .ZN(_0833_));
 INV_X1 _2920_ (.A(net49),
    .ZN(_0834_));
 NOR4_X4 _2921_ (.A1(_0834_),
    .A2(net96),
    .A3(_0814_),
    .A4(_0829_),
    .ZN(_0835_));
 MUX2_X1 _2922_ (.A(_0832_),
    .B(_0833_),
    .S(_0835_),
    .Z(_0035_));
 AND2_X1 _2923_ (.A1(net51),
    .A2(net3),
    .ZN(_0836_));
 NOR2_X1 _2924_ (.A1(net51),
    .A2(_0783_),
    .ZN(_0837_));
 NAND2_X1 _2925_ (.A1(net49),
    .A2(net50),
    .ZN(_0838_));
 NOR3_X1 _2926_ (.A1(_0820_),
    .A2(_0829_),
    .A3(_0838_),
    .ZN(_0839_));
 MUX2_X1 _2927_ (.A(_0836_),
    .B(_0837_),
    .S(_0839_),
    .Z(_0036_));
 NAND4_X1 _2928_ (.A1(net2),
    .A2(_0017_),
    .A3(net3),
    .A4(net44),
    .ZN(_0840_));
 NAND2_X1 _2929_ (.A1(net52),
    .A2(net3),
    .ZN(_0841_));
 OAI21_X1 _2930_ (.A(_0840_),
    .B1(_0841_),
    .B2(net97),
    .ZN(_0037_));
 NOR2_X1 _2931_ (.A1(net53),
    .A2(_0783_),
    .ZN(_0842_));
 AND2_X1 _2932_ (.A1(net53),
    .A2(net3),
    .ZN(_0843_));
 NAND3_X1 _2933_ (.A1(net2),
    .A2(_0016_),
    .A3(net44),
    .ZN(_0844_));
 MUX2_X1 _2934_ (.A(_0842_),
    .B(_0843_),
    .S(_0844_),
    .Z(_0038_));
 NAND2_X1 _2935_ (.A1(net52),
    .A2(net45),
    .ZN(_0845_));
 OAI211_X2 _2936_ (.A(_0617_),
    .B(_0816_),
    .C1(_0622_),
    .C2(_0620_),
    .ZN(_0846_));
 OAI21_X1 _2937_ (.A(net54),
    .B1(_0845_),
    .B2(_0846_),
    .ZN(_0847_));
 OR3_X1 _2938_ (.A1(net54),
    .A2(_0845_),
    .A3(_0846_),
    .ZN(_0848_));
 AOI21_X1 _2939_ (.A(_0783_),
    .B1(_0847_),
    .B2(_0848_),
    .ZN(_0039_));
 NAND2_X1 _2940_ (.A1(_0016_),
    .A2(net54),
    .ZN(_0849_));
 OAI21_X1 _2941_ (.A(net55),
    .B1(_0849_),
    .B2(_0846_),
    .ZN(_0850_));
 OR3_X1 _2942_ (.A1(net55),
    .A2(_0849_),
    .A3(_0846_),
    .ZN(_0851_));
 AOI21_X1 _2943_ (.A(_0783_),
    .B1(_0850_),
    .B2(_0851_),
    .ZN(_0040_));
 XOR2_X1 _2944_ (.A(net56),
    .B(_0820_),
    .Z(_0852_));
 NOR2_X1 _2945_ (.A1(_0783_),
    .A2(_0852_),
    .ZN(_0041_));
 NAND4_X1 _2946_ (.A1(_0016_),
    .A2(net54),
    .A3(net55),
    .A4(net56),
    .ZN(_0853_));
 OAI21_X1 _2947_ (.A(net57),
    .B1(_0846_),
    .B2(_0853_),
    .ZN(_0854_));
 OR3_X1 _2948_ (.A1(net57),
    .A2(_0846_),
    .A3(_0853_),
    .ZN(_0855_));
 AOI21_X1 _2949_ (.A(_0783_),
    .B1(_0854_),
    .B2(_0855_),
    .ZN(_0042_));
 NAND3_X1 _2950_ (.A1(net56),
    .A2(net57),
    .A3(_0817_),
    .ZN(_0856_));
 OAI21_X1 _2951_ (.A(net58),
    .B1(_0846_),
    .B2(_0856_),
    .ZN(_0857_));
 OR3_X1 _2952_ (.A1(net58),
    .A2(_0846_),
    .A3(_0856_),
    .ZN(_0858_));
 AOI21_X1 _2953_ (.A(_0783_),
    .B1(_0857_),
    .B2(_0858_),
    .ZN(_0043_));
 AND2_X1 _2954_ (.A1(net59),
    .A2(net3),
    .ZN(_0859_));
 NOR2_X1 _2955_ (.A1(net59),
    .A2(_0783_),
    .ZN(_0860_));
 NAND3_X1 _2956_ (.A1(net56),
    .A2(net57),
    .A3(net58),
    .ZN(_0861_));
 NOR4_X2 _2957_ (.A1(net96),
    .A2(_0861_),
    .A3(_0810_),
    .A4(_0813_),
    .ZN(_0862_));
 MUX2_X1 _2958_ (.A(_0859_),
    .B(_0860_),
    .S(_0862_),
    .Z(_0044_));
 BUF_X1 output79 (.A(net79),
    .Z(rd_data[23]));
 OAI21_X1 _2960_ (.A(net60),
    .B1(_0809_),
    .B2(_0820_),
    .ZN(_0864_));
 OR3_X1 _2961_ (.A1(net60),
    .A2(_0809_),
    .A3(_0820_),
    .ZN(_0865_));
 AOI21_X1 _2962_ (.A(_0783_),
    .B1(_0864_),
    .B2(_0865_),
    .ZN(_0045_));
 INV_X1 _2963_ (.A(net1),
    .ZN(_0866_));
 AOI22_X1 _2964_ (.A1(net61),
    .A2(_0866_),
    .B1(net44),
    .B2(net2),
    .ZN(_0867_));
 NOR2_X1 _2965_ (.A1(_0783_),
    .A2(_0867_),
    .ZN(_0046_));
 BUF_X1 output78 (.A(net78),
    .Z(rd_data[22]));
 BUF_X1 output77 (.A(net77),
    .Z(rd_data[21]));
 BUF_X1 output76 (.A(net76),
    .Z(rd_data[20]));
 BUF_X1 output75 (.A(net75),
    .Z(rd_data[1]));
 MUX2_X1 _2970_ (.A(\mem[0][0] ),
    .B(\mem[4][0] ),
    .S(net203),
    .Z(_0872_));
 MUX2_X1 _2971_ (.A(\mem[1][0] ),
    .B(\mem[5][0] ),
    .S(net203),
    .Z(_0873_));
 BUF_X1 output74 (.A(net74),
    .Z(rd_data[19]));
 BUF_X1 output73 (.A(net73),
    .Z(rd_data[18]));
 BUF_X1 output72 (.A(net72),
    .Z(rd_data[17]));
 MUX2_X1 _2975_ (.A(_0872_),
    .B(_0873_),
    .S(net206),
    .Z(_0877_));
 BUF_X1 output71 (.A(net71),
    .Z(rd_data[16]));
 BUF_X1 output70 (.A(net70),
    .Z(rd_data[15]));
 NOR2_X2 _2978_ (.A1(_0001_),
    .A2(_0003_),
    .ZN(_0880_));
 BUF_X1 output69 (.A(net69),
    .Z(rd_data[14]));
 INV_X1 _2980_ (.A(_0003_),
    .ZN(_0882_));
 NOR2_X2 _2981_ (.A1(_0001_),
    .A2(_0882_),
    .ZN(_0883_));
 MUX2_X1 _2982_ (.A(\mem[8][0] ),
    .B(\mem[12][0] ),
    .S(net203),
    .Z(_0884_));
 MUX2_X1 _2983_ (.A(\mem[9][0] ),
    .B(\mem[13][0] ),
    .S(net203),
    .Z(_0885_));
 MUX2_X1 _2984_ (.A(_0884_),
    .B(_0885_),
    .S(net206),
    .Z(_0886_));
 AOI22_X1 _2985_ (.A1(_0877_),
    .A2(net198),
    .B1(net190),
    .B2(_0886_),
    .ZN(_0887_));
 MUX2_X1 _2986_ (.A(\mem[2][0] ),
    .B(\mem[6][0] ),
    .S(net203),
    .Z(_0888_));
 MUX2_X1 _2987_ (.A(\mem[3][0] ),
    .B(\mem[7][0] ),
    .S(net203),
    .Z(_0889_));
 MUX2_X1 _2988_ (.A(_0888_),
    .B(_0889_),
    .S(net206),
    .Z(_0890_));
 INV_X1 _2989_ (.A(_0001_),
    .ZN(_0891_));
 NOR2_X2 _2990_ (.A1(_0891_),
    .A2(_0003_),
    .ZN(_0892_));
 BUF_X1 output68 (.A(net68),
    .Z(rd_data[13]));
 NOR2_X2 _2992_ (.A1(_0891_),
    .A2(_0882_),
    .ZN(_0894_));
 MUX2_X1 _2993_ (.A(\mem[10][0] ),
    .B(\mem[14][0] ),
    .S(net203),
    .Z(_0895_));
 MUX2_X1 _2994_ (.A(\mem[11][0] ),
    .B(\mem[15][0] ),
    .S(net203),
    .Z(_0896_));
 MUX2_X1 _2995_ (.A(_0895_),
    .B(_0896_),
    .S(net206),
    .Z(_0897_));
 AOI22_X1 _2996_ (.A1(_0890_),
    .A2(net189),
    .B1(net188),
    .B2(_0897_),
    .ZN(_0898_));
 NAND2_X1 _2997_ (.A1(_0887_),
    .A2(_0898_),
    .ZN(_0899_));
 NAND3_X1 _2998_ (.A1(net210),
    .A2(net173),
    .A3(_0899_),
    .ZN(_0900_));
 BUF_X1 output67 (.A(net67),
    .Z(rd_data[12]));
 OAI21_X1 _3000_ (.A(\last_valid_data[0] ),
    .B1(net44),
    .B2(net209),
    .ZN(_0902_));
 AOI21_X1 _3001_ (.A(net208),
    .B1(_0900_),
    .B2(_0902_),
    .ZN(_0047_));
 BUF_X1 output66 (.A(net66),
    .Z(rd_data[11]));
 BUF_X1 output65 (.A(net65),
    .Z(rd_data[10]));
 MUX2_X1 _3004_ (.A(\mem[8][10] ),
    .B(\mem[12][10] ),
    .S(net204),
    .Z(_0905_));
 MUX2_X1 _3005_ (.A(\mem[9][10] ),
    .B(\mem[13][10] ),
    .S(net204),
    .Z(_0906_));
 MUX2_X1 _3006_ (.A(_0905_),
    .B(_0906_),
    .S(_0000_),
    .Z(_0907_));
 BUF_X1 output64 (.A(net64),
    .Z(rd_data[0]));
 BUF_X1 output63 (.A(net63),
    .Z(overflow_detected));
 MUX2_X1 _3009_ (.A(\mem[0][10] ),
    .B(\mem[4][10] ),
    .S(net204),
    .Z(_0910_));
 BUF_X1 output62 (.A(net62),
    .Z(full));
 BUF_X1 output61 (.A(net61),
    .Z(error_detected));
 MUX2_X1 _3012_ (.A(\mem[1][10] ),
    .B(\mem[5][10] ),
    .S(net204),
    .Z(_0913_));
 BUF_X1 output60 (.A(net60),
    .Z(error_count[9]));
 BUF_X1 output59 (.A(net59),
    .Z(error_count[8]));
 MUX2_X1 _3015_ (.A(_0910_),
    .B(_0913_),
    .S(_0000_),
    .Z(_0916_));
 AOI22_X1 _3016_ (.A1(net190),
    .A2(_0907_),
    .B1(_0916_),
    .B2(net198),
    .ZN(_0917_));
 BUF_X1 output58 (.A(net58),
    .Z(error_count[7]));
 BUF_X1 output57 (.A(net57),
    .Z(error_count[6]));
 MUX2_X1 _3019_ (.A(\mem[10][10] ),
    .B(\mem[14][10] ),
    .S(net204),
    .Z(_0920_));
 BUF_X1 output56 (.A(net56),
    .Z(error_count[5]));
 MUX2_X1 _3021_ (.A(\mem[11][10] ),
    .B(\mem[15][10] ),
    .S(net204),
    .Z(_0922_));
 BUF_X1 output55 (.A(net55),
    .Z(error_count[4]));
 MUX2_X1 _3023_ (.A(_0920_),
    .B(_0922_),
    .S(_0000_),
    .Z(_0924_));
 BUF_X1 output54 (.A(net54),
    .Z(error_count[3]));
 MUX2_X1 _3025_ (.A(\mem[2][10] ),
    .B(\mem[6][10] ),
    .S(net204),
    .Z(_0926_));
 BUF_X1 output53 (.A(net53),
    .Z(error_count[2]));
 MUX2_X1 _3027_ (.A(\mem[3][10] ),
    .B(\mem[7][10] ),
    .S(net204),
    .Z(_0928_));
 BUF_X1 output52 (.A(net52),
    .Z(error_count[1]));
 MUX2_X1 _3029_ (.A(_0926_),
    .B(_0928_),
    .S(_0000_),
    .Z(_0930_));
 AOI22_X1 _3030_ (.A1(_0894_),
    .A2(_0924_),
    .B1(_0930_),
    .B2(net189),
    .ZN(_0931_));
 NAND2_X1 _3031_ (.A1(_0917_),
    .A2(_0931_),
    .ZN(_0932_));
 NAND3_X1 _3032_ (.A1(net2),
    .A2(net96),
    .A3(_0932_),
    .ZN(_0933_));
 OAI21_X1 _3033_ (.A(\last_valid_data[10] ),
    .B1(net44),
    .B2(_0629_),
    .ZN(_0934_));
 AOI21_X1 _3034_ (.A(net208),
    .B1(_0933_),
    .B2(_0934_),
    .ZN(_0048_));
 MUX2_X1 _3035_ (.A(\mem[8][11] ),
    .B(\mem[12][11] ),
    .S(net204),
    .Z(_0935_));
 MUX2_X1 _3036_ (.A(\mem[9][11] ),
    .B(\mem[13][11] ),
    .S(net204),
    .Z(_0936_));
 MUX2_X1 _3037_ (.A(_0935_),
    .B(_0936_),
    .S(net206),
    .Z(_0937_));
 BUF_X1 output51 (.A(net51),
    .Z(error_count[15]));
 MUX2_X1 _3039_ (.A(\mem[0][11] ),
    .B(\mem[4][11] ),
    .S(net204),
    .Z(_0939_));
 MUX2_X1 _3040_ (.A(\mem[1][11] ),
    .B(\mem[5][11] ),
    .S(net204),
    .Z(_0940_));
 MUX2_X1 _3041_ (.A(_0939_),
    .B(_0940_),
    .S(net206),
    .Z(_0941_));
 AOI22_X1 _3042_ (.A1(net190),
    .A2(_0937_),
    .B1(_0941_),
    .B2(net198),
    .ZN(_0942_));
 MUX2_X1 _3043_ (.A(\mem[10][11] ),
    .B(\mem[14][11] ),
    .S(net204),
    .Z(_0943_));
 MUX2_X1 _3044_ (.A(\mem[11][11] ),
    .B(\mem[15][11] ),
    .S(net204),
    .Z(_0944_));
 MUX2_X1 _3045_ (.A(_0943_),
    .B(_0944_),
    .S(net206),
    .Z(_0945_));
 MUX2_X1 _3046_ (.A(\mem[2][11] ),
    .B(\mem[6][11] ),
    .S(net204),
    .Z(_0946_));
 MUX2_X1 _3047_ (.A(\mem[3][11] ),
    .B(\mem[7][11] ),
    .S(net204),
    .Z(_0947_));
 MUX2_X1 _3048_ (.A(_0946_),
    .B(_0947_),
    .S(net206),
    .Z(_0948_));
 AOI22_X1 _3049_ (.A1(net188),
    .A2(_0945_),
    .B1(_0948_),
    .B2(net189),
    .ZN(_0949_));
 NAND2_X1 _3050_ (.A1(_0942_),
    .A2(_0949_),
    .ZN(_0950_));
 NAND3_X1 _3051_ (.A1(net210),
    .A2(net173),
    .A3(_0950_),
    .ZN(_0951_));
 OAI21_X1 _3052_ (.A(\last_valid_data[11] ),
    .B1(net44),
    .B2(net209),
    .ZN(_0952_));
 AOI21_X1 _3053_ (.A(net208),
    .B1(_0951_),
    .B2(_0952_),
    .ZN(_0049_));
 MUX2_X1 _3054_ (.A(\mem[8][12] ),
    .B(\mem[12][12] ),
    .S(net204),
    .Z(_0953_));
 MUX2_X1 _3055_ (.A(\mem[9][12] ),
    .B(\mem[13][12] ),
    .S(net204),
    .Z(_0954_));
 MUX2_X1 _3056_ (.A(_0953_),
    .B(_0954_),
    .S(_0000_),
    .Z(_0955_));
 MUX2_X1 _3057_ (.A(\mem[0][12] ),
    .B(\mem[4][12] ),
    .S(net204),
    .Z(_0956_));
 BUF_X1 output50 (.A(net50),
    .Z(error_count[14]));
 MUX2_X1 _3059_ (.A(\mem[1][12] ),
    .B(\mem[5][12] ),
    .S(net204),
    .Z(_0958_));
 MUX2_X1 _3060_ (.A(_0956_),
    .B(_0958_),
    .S(_0000_),
    .Z(_0959_));
 AOI22_X1 _3061_ (.A1(net190),
    .A2(_0955_),
    .B1(_0959_),
    .B2(net198),
    .ZN(_0960_));
 MUX2_X1 _3062_ (.A(\mem[10][12] ),
    .B(\mem[14][12] ),
    .S(net204),
    .Z(_0961_));
 MUX2_X1 _3063_ (.A(\mem[11][12] ),
    .B(\mem[15][12] ),
    .S(net204),
    .Z(_0962_));
 MUX2_X1 _3064_ (.A(_0961_),
    .B(_0962_),
    .S(_0000_),
    .Z(_0963_));
 MUX2_X1 _3065_ (.A(\mem[2][12] ),
    .B(\mem[6][12] ),
    .S(net204),
    .Z(_0964_));
 MUX2_X1 _3066_ (.A(\mem[3][12] ),
    .B(\mem[7][12] ),
    .S(net204),
    .Z(_0965_));
 MUX2_X1 _3067_ (.A(_0964_),
    .B(_0965_),
    .S(_0000_),
    .Z(_0966_));
 AOI22_X1 _3068_ (.A1(_0894_),
    .A2(_0963_),
    .B1(_0966_),
    .B2(net189),
    .ZN(_0967_));
 NAND2_X1 _3069_ (.A1(_0960_),
    .A2(_0967_),
    .ZN(_0968_));
 NAND3_X1 _3070_ (.A1(net2),
    .A2(net96),
    .A3(_0968_),
    .ZN(_0969_));
 OAI21_X1 _3071_ (.A(\last_valid_data[12] ),
    .B1(net44),
    .B2(_0629_),
    .ZN(_0970_));
 AOI21_X1 _3072_ (.A(net208),
    .B1(_0969_),
    .B2(_0970_),
    .ZN(_0050_));
 MUX2_X1 _3073_ (.A(\mem[8][13] ),
    .B(\mem[12][13] ),
    .S(net204),
    .Z(_0971_));
 MUX2_X1 _3074_ (.A(\mem[9][13] ),
    .B(\mem[13][13] ),
    .S(net204),
    .Z(_0972_));
 MUX2_X1 _3075_ (.A(_0971_),
    .B(_0972_),
    .S(net206),
    .Z(_0973_));
 MUX2_X1 _3076_ (.A(\mem[0][13] ),
    .B(\mem[4][13] ),
    .S(net204),
    .Z(_0974_));
 MUX2_X1 _3077_ (.A(\mem[1][13] ),
    .B(\mem[5][13] ),
    .S(net204),
    .Z(_0975_));
 MUX2_X1 _3078_ (.A(_0974_),
    .B(_0975_),
    .S(net206),
    .Z(_0976_));
 AOI22_X1 _3079_ (.A1(net190),
    .A2(_0973_),
    .B1(_0976_),
    .B2(net198),
    .ZN(_0977_));
 BUF_X1 output49 (.A(net49),
    .Z(error_count[13]));
 MUX2_X1 _3081_ (.A(\mem[10][13] ),
    .B(\mem[14][13] ),
    .S(net204),
    .Z(_0979_));
 MUX2_X1 _3082_ (.A(\mem[11][13] ),
    .B(\mem[15][13] ),
    .S(net204),
    .Z(_0980_));
 MUX2_X1 _3083_ (.A(_0979_),
    .B(_0980_),
    .S(net206),
    .Z(_0981_));
 MUX2_X1 _3084_ (.A(\mem[2][13] ),
    .B(\mem[6][13] ),
    .S(net203),
    .Z(_0982_));
 MUX2_X1 _3085_ (.A(\mem[3][13] ),
    .B(\mem[7][13] ),
    .S(net203),
    .Z(_0983_));
 MUX2_X1 _3086_ (.A(_0982_),
    .B(_0983_),
    .S(net206),
    .Z(_0984_));
 AOI22_X1 _3087_ (.A1(net188),
    .A2(_0981_),
    .B1(_0984_),
    .B2(net189),
    .ZN(_0985_));
 NAND2_X1 _3088_ (.A1(_0977_),
    .A2(_0985_),
    .ZN(_0986_));
 NAND3_X1 _3089_ (.A1(net210),
    .A2(net173),
    .A3(_0986_),
    .ZN(_0987_));
 BUF_X1 output48 (.A(net48),
    .Z(error_count[12]));
 OAI21_X1 _3091_ (.A(\last_valid_data[13] ),
    .B1(net44),
    .B2(net209),
    .ZN(_0989_));
 AOI21_X1 _3092_ (.A(net208),
    .B1(_0987_),
    .B2(_0989_),
    .ZN(_0051_));
 MUX2_X1 _3093_ (.A(\mem[8][14] ),
    .B(\mem[12][14] ),
    .S(net204),
    .Z(_0990_));
 MUX2_X1 _3094_ (.A(\mem[9][14] ),
    .B(\mem[13][14] ),
    .S(net204),
    .Z(_0991_));
 MUX2_X1 _3095_ (.A(_0990_),
    .B(_0991_),
    .S(net206),
    .Z(_0992_));
 MUX2_X1 _3096_ (.A(\mem[0][14] ),
    .B(\mem[4][14] ),
    .S(net204),
    .Z(_0993_));
 MUX2_X1 _3097_ (.A(\mem[1][14] ),
    .B(\mem[5][14] ),
    .S(net204),
    .Z(_0994_));
 MUX2_X1 _3098_ (.A(_0993_),
    .B(_0994_),
    .S(net206),
    .Z(_0995_));
 AOI22_X1 _3099_ (.A1(net190),
    .A2(_0992_),
    .B1(_0995_),
    .B2(net198),
    .ZN(_0996_));
 MUX2_X1 _3100_ (.A(\mem[10][14] ),
    .B(\mem[14][14] ),
    .S(net204),
    .Z(_0997_));
 BUF_X1 output47 (.A(net47),
    .Z(error_count[11]));
 MUX2_X1 _3102_ (.A(\mem[11][14] ),
    .B(\mem[15][14] ),
    .S(net204),
    .Z(_0999_));
 MUX2_X1 _3103_ (.A(_0997_),
    .B(_0999_),
    .S(net206),
    .Z(_1000_));
 MUX2_X1 _3104_ (.A(\mem[2][14] ),
    .B(\mem[6][14] ),
    .S(net204),
    .Z(_1001_));
 MUX2_X1 _3105_ (.A(\mem[3][14] ),
    .B(\mem[7][14] ),
    .S(net204),
    .Z(_1002_));
 MUX2_X1 _3106_ (.A(_1001_),
    .B(_1002_),
    .S(net206),
    .Z(_1003_));
 AOI22_X1 _3107_ (.A1(net188),
    .A2(_1000_),
    .B1(_1003_),
    .B2(net189),
    .ZN(_1004_));
 NAND2_X1 _3108_ (.A1(_0996_),
    .A2(_1004_),
    .ZN(_1005_));
 NAND3_X1 _3109_ (.A1(net210),
    .A2(net173),
    .A3(_1005_),
    .ZN(_1006_));
 OAI21_X1 _3110_ (.A(\last_valid_data[14] ),
    .B1(net44),
    .B2(net209),
    .ZN(_1007_));
 AOI21_X1 _3111_ (.A(net208),
    .B1(_1006_),
    .B2(_1007_),
    .ZN(_0052_));
 BUF_X1 output46 (.A(net46),
    .Z(error_count[10]));
 MUX2_X1 _3113_ (.A(\mem[8][15] ),
    .B(\mem[12][15] ),
    .S(net204),
    .Z(_1009_));
 MUX2_X1 _3114_ (.A(\mem[9][15] ),
    .B(\mem[13][15] ),
    .S(net204),
    .Z(_1010_));
 MUX2_X1 _3115_ (.A(_1009_),
    .B(_1010_),
    .S(net206),
    .Z(_1011_));
 MUX2_X1 _3116_ (.A(\mem[0][15] ),
    .B(\mem[4][15] ),
    .S(net204),
    .Z(_1012_));
 MUX2_X1 _3117_ (.A(\mem[1][15] ),
    .B(\mem[5][15] ),
    .S(net204),
    .Z(_1013_));
 MUX2_X1 _3118_ (.A(_1012_),
    .B(_1013_),
    .S(net206),
    .Z(_1014_));
 AOI22_X1 _3119_ (.A1(net190),
    .A2(_1011_),
    .B1(_1014_),
    .B2(net198),
    .ZN(_1015_));
 MUX2_X1 _3120_ (.A(\mem[10][15] ),
    .B(\mem[14][15] ),
    .S(net204),
    .Z(_1016_));
 MUX2_X1 _3121_ (.A(\mem[11][15] ),
    .B(\mem[15][15] ),
    .S(net204),
    .Z(_1017_));
 MUX2_X1 _3122_ (.A(_1016_),
    .B(_1017_),
    .S(net206),
    .Z(_1018_));
 MUX2_X1 _3123_ (.A(\mem[2][15] ),
    .B(\mem[6][15] ),
    .S(net204),
    .Z(_1019_));
 MUX2_X1 _3124_ (.A(\mem[3][15] ),
    .B(\mem[7][15] ),
    .S(net204),
    .Z(_1020_));
 BUF_X1 output45 (.A(net45),
    .Z(error_count[0]));
 MUX2_X1 _3126_ (.A(_1019_),
    .B(_1020_),
    .S(net206),
    .Z(_1022_));
 AOI22_X1 _3127_ (.A1(net188),
    .A2(_1018_),
    .B1(_1022_),
    .B2(net189),
    .ZN(_1023_));
 NAND2_X1 _3128_ (.A1(_1015_),
    .A2(_1023_),
    .ZN(_1024_));
 NAND3_X1 _3129_ (.A1(net210),
    .A2(net173),
    .A3(_1024_),
    .ZN(_1025_));
 OAI21_X1 _3130_ (.A(\last_valid_data[15] ),
    .B1(net44),
    .B2(net209),
    .ZN(_1026_));
 AOI21_X1 _3131_ (.A(net208),
    .B1(_1025_),
    .B2(_1026_),
    .ZN(_0053_));
 BUF_X1 output44 (.A(net44),
    .Z(empty));
 MUX2_X1 _3133_ (.A(\mem[8][16] ),
    .B(\mem[12][16] ),
    .S(net204),
    .Z(_1028_));
 BUF_X1 output43 (.A(net43),
    .Z(data_count[4]));
 MUX2_X1 _3135_ (.A(\mem[9][16] ),
    .B(\mem[13][16] ),
    .S(net204),
    .Z(_1030_));
 MUX2_X1 _3136_ (.A(_1028_),
    .B(_1030_),
    .S(_0000_),
    .Z(_1031_));
 MUX2_X1 _3137_ (.A(\mem[0][16] ),
    .B(\mem[4][16] ),
    .S(net204),
    .Z(_1032_));
 MUX2_X1 _3138_ (.A(\mem[1][16] ),
    .B(\mem[5][16] ),
    .S(net204),
    .Z(_1033_));
 BUF_X1 output42 (.A(net42),
    .Z(data_count[3]));
 MUX2_X1 _3140_ (.A(_1032_),
    .B(_1033_),
    .S(_0000_),
    .Z(_1035_));
 AOI22_X1 _3141_ (.A1(net190),
    .A2(_1031_),
    .B1(_1035_),
    .B2(net198),
    .ZN(_1036_));
 MUX2_X1 _3142_ (.A(\mem[10][16] ),
    .B(\mem[14][16] ),
    .S(net204),
    .Z(_1037_));
 MUX2_X1 _3143_ (.A(\mem[11][16] ),
    .B(\mem[15][16] ),
    .S(net204),
    .Z(_1038_));
 MUX2_X1 _3144_ (.A(_1037_),
    .B(_1038_),
    .S(_0000_),
    .Z(_1039_));
 MUX2_X1 _3145_ (.A(\mem[2][16] ),
    .B(\mem[6][16] ),
    .S(net204),
    .Z(_1040_));
 MUX2_X1 _3146_ (.A(\mem[3][16] ),
    .B(\mem[7][16] ),
    .S(net204),
    .Z(_1041_));
 MUX2_X1 _3147_ (.A(_1040_),
    .B(_1041_),
    .S(_0000_),
    .Z(_1042_));
 AOI22_X1 _3148_ (.A1(_0894_),
    .A2(_1039_),
    .B1(_1042_),
    .B2(net189),
    .ZN(_1043_));
 NAND2_X1 _3149_ (.A1(_1036_),
    .A2(_1043_),
    .ZN(_1044_));
 NAND3_X1 _3150_ (.A1(net2),
    .A2(net96),
    .A3(_1044_),
    .ZN(_1045_));
 OAI21_X1 _3151_ (.A(\last_valid_data[16] ),
    .B1(net44),
    .B2(_0629_),
    .ZN(_1046_));
 AOI21_X1 _3152_ (.A(net208),
    .B1(_1045_),
    .B2(_1046_),
    .ZN(_0054_));
 BUF_X1 output41 (.A(net41),
    .Z(data_count[2]));
 MUX2_X1 _3154_ (.A(\mem[8][17] ),
    .B(\mem[12][17] ),
    .S(net203),
    .Z(_1048_));
 MUX2_X1 _3155_ (.A(\mem[9][17] ),
    .B(\mem[13][17] ),
    .S(net203),
    .Z(_1049_));
 MUX2_X1 _3156_ (.A(_1048_),
    .B(_1049_),
    .S(_0000_),
    .Z(_1050_));
 MUX2_X1 _3157_ (.A(\mem[0][17] ),
    .B(\mem[4][17] ),
    .S(net203),
    .Z(_1051_));
 MUX2_X1 _3158_ (.A(\mem[1][17] ),
    .B(\mem[5][17] ),
    .S(net204),
    .Z(_1052_));
 MUX2_X1 _3159_ (.A(_1051_),
    .B(_1052_),
    .S(_0000_),
    .Z(_1053_));
 AOI22_X1 _3160_ (.A1(net190),
    .A2(_1050_),
    .B1(_1053_),
    .B2(net198),
    .ZN(_1054_));
 MUX2_X1 _3161_ (.A(\mem[10][17] ),
    .B(\mem[14][17] ),
    .S(net204),
    .Z(_1055_));
 MUX2_X1 _3162_ (.A(\mem[11][17] ),
    .B(\mem[15][17] ),
    .S(net204),
    .Z(_1056_));
 BUF_X1 output40 (.A(net40),
    .Z(data_count[1]));
 MUX2_X1 _3164_ (.A(_1055_),
    .B(_1056_),
    .S(_0000_),
    .Z(_1058_));
 MUX2_X1 _3165_ (.A(\mem[2][17] ),
    .B(\mem[6][17] ),
    .S(net203),
    .Z(_1059_));
 MUX2_X1 _3166_ (.A(\mem[3][17] ),
    .B(\mem[7][17] ),
    .S(net203),
    .Z(_1060_));
 MUX2_X1 _3167_ (.A(_1059_),
    .B(_1060_),
    .S(_0000_),
    .Z(_1061_));
 AOI22_X1 _3168_ (.A1(net188),
    .A2(_1058_),
    .B1(_1061_),
    .B2(net189),
    .ZN(_1062_));
 NAND2_X1 _3169_ (.A1(_1054_),
    .A2(_1062_),
    .ZN(_1063_));
 NAND3_X1 _3170_ (.A1(net210),
    .A2(net173),
    .A3(_1063_),
    .ZN(_1064_));
 OAI21_X1 _3171_ (.A(\last_valid_data[17] ),
    .B1(net44),
    .B2(net209),
    .ZN(_1065_));
 AOI21_X1 _3172_ (.A(net208),
    .B1(_1064_),
    .B2(_1065_),
    .ZN(_0055_));
 BUF_X1 output39 (.A(net39),
    .Z(data_count[0]));
 MUX2_X1 _3174_ (.A(\mem[8][18] ),
    .B(\mem[12][18] ),
    .S(net204),
    .Z(_1067_));
 MUX2_X1 _3175_ (.A(\mem[9][18] ),
    .B(\mem[13][18] ),
    .S(net204),
    .Z(_1068_));
 BUF_X1 output38 (.A(net38),
    .Z(almost_full));
 MUX2_X1 _3177_ (.A(_1067_),
    .B(_1068_),
    .S(net206),
    .Z(_1070_));
 MUX2_X1 _3178_ (.A(\mem[0][18] ),
    .B(\mem[4][18] ),
    .S(net204),
    .Z(_1071_));
 MUX2_X1 _3179_ (.A(\mem[1][18] ),
    .B(\mem[5][18] ),
    .S(net204),
    .Z(_1072_));
 MUX2_X1 _3180_ (.A(_1071_),
    .B(_1072_),
    .S(net206),
    .Z(_1073_));
 AOI22_X1 _3181_ (.A1(net190),
    .A2(_1070_),
    .B1(_1073_),
    .B2(net198),
    .ZN(_1074_));
 MUX2_X1 _3182_ (.A(\mem[10][18] ),
    .B(\mem[14][18] ),
    .S(net204),
    .Z(_1075_));
 MUX2_X1 _3183_ (.A(\mem[11][18] ),
    .B(\mem[15][18] ),
    .S(net204),
    .Z(_1076_));
 MUX2_X1 _3184_ (.A(_1075_),
    .B(_1076_),
    .S(net206),
    .Z(_1077_));
 MUX2_X1 _3185_ (.A(\mem[2][18] ),
    .B(\mem[6][18] ),
    .S(net204),
    .Z(_1078_));
 MUX2_X1 _3186_ (.A(\mem[3][18] ),
    .B(\mem[7][18] ),
    .S(net204),
    .Z(_1079_));
 MUX2_X1 _3187_ (.A(_1078_),
    .B(_1079_),
    .S(net206),
    .Z(_1080_));
 AOI22_X1 _3188_ (.A1(net188),
    .A2(_1077_),
    .B1(_1080_),
    .B2(net189),
    .ZN(_1081_));
 NAND2_X1 _3189_ (.A1(_1074_),
    .A2(_1081_),
    .ZN(_1082_));
 NAND3_X1 _3190_ (.A1(net210),
    .A2(net173),
    .A3(_1082_),
    .ZN(_1083_));
 OAI21_X1 _3191_ (.A(\last_valid_data[18] ),
    .B1(net44),
    .B2(net209),
    .ZN(_1084_));
 AOI21_X1 _3192_ (.A(net208),
    .B1(_1083_),
    .B2(_1084_),
    .ZN(_0056_));
 MUX2_X1 _3193_ (.A(\mem[8][19] ),
    .B(\mem[12][19] ),
    .S(net203),
    .Z(_1085_));
 MUX2_X1 _3194_ (.A(\mem[9][19] ),
    .B(\mem[13][19] ),
    .S(net203),
    .Z(_1086_));
 MUX2_X1 _3195_ (.A(_1085_),
    .B(_1086_),
    .S(net205),
    .Z(_1087_));
 MUX2_X1 _3196_ (.A(\mem[0][19] ),
    .B(\mem[4][19] ),
    .S(net201),
    .Z(_1088_));
 MUX2_X1 _3197_ (.A(\mem[1][19] ),
    .B(\mem[5][19] ),
    .S(net201),
    .Z(_1089_));
 MUX2_X1 _3198_ (.A(_1088_),
    .B(_1089_),
    .S(net205),
    .Z(_1090_));
 BUF_X1 output37 (.A(net37),
    .Z(almost_empty));
 AOI22_X1 _3200_ (.A1(net190),
    .A2(_1087_),
    .B1(_1090_),
    .B2(net198),
    .ZN(_1092_));
 MUX2_X1 _3201_ (.A(\mem[10][19] ),
    .B(\mem[14][19] ),
    .S(net203),
    .Z(_1093_));
 MUX2_X1 _3202_ (.A(\mem[11][19] ),
    .B(\mem[15][19] ),
    .S(net203),
    .Z(_1094_));
 MUX2_X1 _3203_ (.A(_1093_),
    .B(_1094_),
    .S(net205),
    .Z(_1095_));
 BUF_X1 input36 (.A(wr_en),
    .Z(net36));
 MUX2_X1 _3205_ (.A(\mem[2][19] ),
    .B(\mem[6][19] ),
    .S(net203),
    .Z(_1097_));
 MUX2_X1 _3206_ (.A(\mem[3][19] ),
    .B(\mem[7][19] ),
    .S(net203),
    .Z(_1098_));
 MUX2_X1 _3207_ (.A(_1097_),
    .B(_1098_),
    .S(net205),
    .Z(_1099_));
 BUF_X1 input35 (.A(wr_data[9]),
    .Z(net35));
 AOI22_X1 _3209_ (.A1(net188),
    .A2(_1095_),
    .B1(_1099_),
    .B2(net189),
    .ZN(_1101_));
 NAND2_X1 _3210_ (.A1(_1092_),
    .A2(_1101_),
    .ZN(_1102_));
 NAND3_X1 _3211_ (.A1(net210),
    .A2(net96),
    .A3(_1102_),
    .ZN(_1103_));
 BUF_X1 input34 (.A(wr_data[8]),
    .Z(net34));
 OAI21_X1 _3213_ (.A(\last_valid_data[19] ),
    .B1(net172),
    .B2(_0629_),
    .ZN(_1105_));
 AOI21_X1 _3214_ (.A(_0783_),
    .B1(_1103_),
    .B2(_1105_),
    .ZN(_0057_));
 BUF_X1 input33 (.A(wr_data[7]),
    .Z(net33));
 MUX2_X1 _3216_ (.A(\mem[8][1] ),
    .B(\mem[12][1] ),
    .S(net202),
    .Z(_1107_));
 MUX2_X1 _3217_ (.A(\mem[9][1] ),
    .B(\mem[13][1] ),
    .S(net202),
    .Z(_1108_));
 MUX2_X1 _3218_ (.A(_1107_),
    .B(_1108_),
    .S(net207),
    .Z(_1109_));
 MUX2_X1 _3219_ (.A(\mem[0][1] ),
    .B(\mem[4][1] ),
    .S(net202),
    .Z(_1110_));
 MUX2_X1 _3220_ (.A(\mem[1][1] ),
    .B(\mem[5][1] ),
    .S(net202),
    .Z(_1111_));
 MUX2_X1 _3221_ (.A(_1110_),
    .B(_1111_),
    .S(net207),
    .Z(_1112_));
 AOI22_X1 _3222_ (.A1(_0883_),
    .A2(_1109_),
    .B1(_1112_),
    .B2(_0880_),
    .ZN(_1113_));
 BUF_X1 input32 (.A(wr_data[6]),
    .Z(net32));
 MUX2_X1 _3224_ (.A(\mem[10][1] ),
    .B(\mem[14][1] ),
    .S(net202),
    .Z(_1115_));
 MUX2_X1 _3225_ (.A(\mem[11][1] ),
    .B(\mem[15][1] ),
    .S(net202),
    .Z(_1116_));
 MUX2_X1 _3226_ (.A(_1115_),
    .B(_1116_),
    .S(net207),
    .Z(_1117_));
 MUX2_X1 _3227_ (.A(\mem[2][1] ),
    .B(\mem[6][1] ),
    .S(net202),
    .Z(_1118_));
 BUF_X1 input31 (.A(wr_data[5]),
    .Z(net31));
 MUX2_X1 _3229_ (.A(\mem[3][1] ),
    .B(\mem[7][1] ),
    .S(net202),
    .Z(_1120_));
 MUX2_X1 _3230_ (.A(_1118_),
    .B(_1120_),
    .S(net207),
    .Z(_1121_));
 AOI22_X1 _3231_ (.A1(_0894_),
    .A2(_1117_),
    .B1(_1121_),
    .B2(_0892_),
    .ZN(_1122_));
 NAND2_X1 _3232_ (.A1(_1113_),
    .A2(_1122_),
    .ZN(_1123_));
 NAND3_X1 _3233_ (.A1(net210),
    .A2(net174),
    .A3(_1123_),
    .ZN(_1124_));
 OAI21_X1 _3234_ (.A(\last_valid_data[1] ),
    .B1(net172),
    .B2(_0629_),
    .ZN(_1125_));
 AOI21_X1 _3235_ (.A(_0783_),
    .B1(_1124_),
    .B2(_1125_),
    .ZN(_0058_));
 MUX2_X1 _3236_ (.A(\mem[8][20] ),
    .B(\mem[12][20] ),
    .S(net202),
    .Z(_1126_));
 MUX2_X1 _3237_ (.A(\mem[9][20] ),
    .B(\mem[13][20] ),
    .S(net202),
    .Z(_1127_));
 MUX2_X1 _3238_ (.A(_1126_),
    .B(_1127_),
    .S(net207),
    .Z(_1128_));
 BUF_X1 input30 (.A(wr_data[4]),
    .Z(net30));
 MUX2_X1 _3240_ (.A(\mem[0][20] ),
    .B(\mem[4][20] ),
    .S(_0002_),
    .Z(_1130_));
 MUX2_X1 _3241_ (.A(\mem[1][20] ),
    .B(\mem[5][20] ),
    .S(_0002_),
    .Z(_1131_));
 MUX2_X1 _3242_ (.A(_1130_),
    .B(_1131_),
    .S(net207),
    .Z(_1132_));
 AOI22_X1 _3243_ (.A1(_0883_),
    .A2(_1128_),
    .B1(_1132_),
    .B2(_0880_),
    .ZN(_1133_));
 MUX2_X1 _3244_ (.A(\mem[10][20] ),
    .B(\mem[14][20] ),
    .S(net202),
    .Z(_1134_));
 MUX2_X1 _3245_ (.A(\mem[11][20] ),
    .B(\mem[15][20] ),
    .S(net202),
    .Z(_1135_));
 MUX2_X1 _3246_ (.A(_1134_),
    .B(_1135_),
    .S(net207),
    .Z(_1136_));
 MUX2_X1 _3247_ (.A(\mem[2][20] ),
    .B(\mem[6][20] ),
    .S(_0002_),
    .Z(_1137_));
 MUX2_X1 _3248_ (.A(\mem[3][20] ),
    .B(\mem[7][20] ),
    .S(_0002_),
    .Z(_1138_));
 MUX2_X1 _3249_ (.A(_1137_),
    .B(_1138_),
    .S(net207),
    .Z(_1139_));
 AOI22_X1 _3250_ (.A1(_0894_),
    .A2(_1136_),
    .B1(_1139_),
    .B2(_0892_),
    .ZN(_1140_));
 NAND2_X1 _3251_ (.A1(_1133_),
    .A2(_1140_),
    .ZN(_1141_));
 NAND3_X1 _3252_ (.A1(net210),
    .A2(net96),
    .A3(_1141_),
    .ZN(_1142_));
 OAI21_X1 _3253_ (.A(\last_valid_data[20] ),
    .B1(net172),
    .B2(_0629_),
    .ZN(_1143_));
 AOI21_X1 _3254_ (.A(_0783_),
    .B1(_1142_),
    .B2(_1143_),
    .ZN(_0059_));
 MUX2_X1 _3255_ (.A(\mem[8][21] ),
    .B(\mem[12][21] ),
    .S(_0002_),
    .Z(_1144_));
 MUX2_X1 _3256_ (.A(\mem[9][21] ),
    .B(\mem[13][21] ),
    .S(_0002_),
    .Z(_1145_));
 MUX2_X1 _3257_ (.A(_1144_),
    .B(_1145_),
    .S(net207),
    .Z(_1146_));
 MUX2_X1 _3258_ (.A(\mem[0][21] ),
    .B(\mem[4][21] ),
    .S(_0002_),
    .Z(_1147_));
 BUF_X1 input29 (.A(wr_data[3]),
    .Z(net29));
 MUX2_X1 _3260_ (.A(\mem[1][21] ),
    .B(\mem[5][21] ),
    .S(_0002_),
    .Z(_1149_));
 MUX2_X1 _3261_ (.A(_1147_),
    .B(_1149_),
    .S(net207),
    .Z(_1150_));
 AOI22_X1 _3262_ (.A1(_0883_),
    .A2(_1146_),
    .B1(_1150_),
    .B2(_0880_),
    .ZN(_1151_));
 MUX2_X1 _3263_ (.A(\mem[10][21] ),
    .B(\mem[14][21] ),
    .S(_0002_),
    .Z(_1152_));
 MUX2_X1 _3264_ (.A(\mem[11][21] ),
    .B(\mem[15][21] ),
    .S(_0002_),
    .Z(_1153_));
 MUX2_X1 _3265_ (.A(_1152_),
    .B(_1153_),
    .S(net207),
    .Z(_1154_));
 MUX2_X1 _3266_ (.A(\mem[2][21] ),
    .B(\mem[6][21] ),
    .S(_0002_),
    .Z(_1155_));
 MUX2_X1 _3267_ (.A(\mem[3][21] ),
    .B(\mem[7][21] ),
    .S(_0002_),
    .Z(_1156_));
 MUX2_X1 _3268_ (.A(_1155_),
    .B(_1156_),
    .S(net207),
    .Z(_1157_));
 AOI22_X1 _3269_ (.A1(_0894_),
    .A2(_1154_),
    .B1(_1157_),
    .B2(_0892_),
    .ZN(_1158_));
 NAND2_X1 _3270_ (.A1(_1151_),
    .A2(_1158_),
    .ZN(_1159_));
 NAND3_X1 _3271_ (.A1(net210),
    .A2(net96),
    .A3(_1159_),
    .ZN(_1160_));
 OAI21_X1 _3272_ (.A(\last_valid_data[21] ),
    .B1(net172),
    .B2(_0629_),
    .ZN(_1161_));
 AOI21_X1 _3273_ (.A(_0783_),
    .B1(_1160_),
    .B2(_1161_),
    .ZN(_0060_));
 MUX2_X1 _3274_ (.A(\mem[8][22] ),
    .B(\mem[12][22] ),
    .S(_0002_),
    .Z(_1162_));
 MUX2_X1 _3275_ (.A(\mem[9][22] ),
    .B(\mem[13][22] ),
    .S(_0002_),
    .Z(_1163_));
 MUX2_X1 _3276_ (.A(_1162_),
    .B(_1163_),
    .S(net207),
    .Z(_1164_));
 MUX2_X1 _3277_ (.A(\mem[0][22] ),
    .B(\mem[4][22] ),
    .S(_0002_),
    .Z(_1165_));
 MUX2_X1 _3278_ (.A(\mem[1][22] ),
    .B(\mem[5][22] ),
    .S(_0002_),
    .Z(_1166_));
 MUX2_X1 _3279_ (.A(_1165_),
    .B(_1166_),
    .S(net207),
    .Z(_1167_));
 AOI22_X1 _3280_ (.A1(_0883_),
    .A2(_1164_),
    .B1(_1167_),
    .B2(_0880_),
    .ZN(_1168_));
 BUF_X1 input28 (.A(wr_data[31]),
    .Z(net28));
 MUX2_X1 _3282_ (.A(\mem[10][22] ),
    .B(\mem[14][22] ),
    .S(_0002_),
    .Z(_1170_));
 MUX2_X1 _3283_ (.A(\mem[11][22] ),
    .B(\mem[15][22] ),
    .S(_0002_),
    .Z(_1171_));
 MUX2_X1 _3284_ (.A(_1170_),
    .B(_1171_),
    .S(net207),
    .Z(_1172_));
 MUX2_X1 _3285_ (.A(\mem[2][22] ),
    .B(\mem[6][22] ),
    .S(_0002_),
    .Z(_1173_));
 MUX2_X1 _3286_ (.A(\mem[3][22] ),
    .B(\mem[7][22] ),
    .S(_0002_),
    .Z(_1174_));
 MUX2_X1 _3287_ (.A(_1173_),
    .B(_1174_),
    .S(net207),
    .Z(_1175_));
 AOI22_X1 _3288_ (.A1(_0894_),
    .A2(_1172_),
    .B1(_1175_),
    .B2(_0892_),
    .ZN(_1176_));
 NAND2_X1 _3289_ (.A1(_1168_),
    .A2(_1176_),
    .ZN(_1177_));
 NAND3_X1 _3290_ (.A1(net210),
    .A2(net174),
    .A3(_1177_),
    .ZN(_1178_));
 BUF_X1 input27 (.A(wr_data[30]),
    .Z(net27));
 OAI21_X1 _3292_ (.A(\last_valid_data[22] ),
    .B1(net172),
    .B2(_0629_),
    .ZN(_1180_));
 AOI21_X1 _3293_ (.A(_0783_),
    .B1(_1178_),
    .B2(_1180_),
    .ZN(_0061_));
 MUX2_X1 _3294_ (.A(\mem[8][23] ),
    .B(\mem[12][23] ),
    .S(net200),
    .Z(_1181_));
 MUX2_X1 _3295_ (.A(\mem[9][23] ),
    .B(\mem[13][23] ),
    .S(net200),
    .Z(_1182_));
 MUX2_X1 _3296_ (.A(_1181_),
    .B(_1182_),
    .S(net207),
    .Z(_1183_));
 MUX2_X1 _3297_ (.A(\mem[0][23] ),
    .B(\mem[4][23] ),
    .S(net200),
    .Z(_1184_));
 MUX2_X1 _3298_ (.A(\mem[1][23] ),
    .B(\mem[5][23] ),
    .S(net200),
    .Z(_1185_));
 MUX2_X1 _3299_ (.A(_1184_),
    .B(_1185_),
    .S(net207),
    .Z(_1186_));
 AOI22_X1 _3300_ (.A1(_0883_),
    .A2(_1183_),
    .B1(_1186_),
    .B2(_0880_),
    .ZN(_1187_));
 MUX2_X1 _3301_ (.A(\mem[10][23] ),
    .B(\mem[14][23] ),
    .S(net200),
    .Z(_1188_));
 BUF_X1 input26 (.A(wr_data[2]),
    .Z(net26));
 MUX2_X1 _3303_ (.A(\mem[11][23] ),
    .B(\mem[15][23] ),
    .S(net200),
    .Z(_1190_));
 MUX2_X1 _3304_ (.A(_1188_),
    .B(_1190_),
    .S(net207),
    .Z(_1191_));
 MUX2_X1 _3305_ (.A(\mem[2][23] ),
    .B(\mem[6][23] ),
    .S(net200),
    .Z(_1192_));
 MUX2_X1 _3306_ (.A(\mem[3][23] ),
    .B(\mem[7][23] ),
    .S(net200),
    .Z(_1193_));
 MUX2_X1 _3307_ (.A(_1192_),
    .B(_1193_),
    .S(net207),
    .Z(_1194_));
 AOI22_X1 _3308_ (.A1(_0894_),
    .A2(_1191_),
    .B1(_1194_),
    .B2(_0892_),
    .ZN(_1195_));
 NAND2_X1 _3309_ (.A1(_1187_),
    .A2(_1195_),
    .ZN(_1196_));
 NAND3_X1 _3310_ (.A1(net210),
    .A2(net174),
    .A3(_1196_),
    .ZN(_1197_));
 OAI21_X1 _3311_ (.A(\last_valid_data[23] ),
    .B1(net172),
    .B2(_0629_),
    .ZN(_1198_));
 AOI21_X1 _3312_ (.A(_0783_),
    .B1(_1197_),
    .B2(_1198_),
    .ZN(_0062_));
 BUF_X1 input25 (.A(wr_data[29]),
    .Z(net25));
 MUX2_X1 _3314_ (.A(\mem[8][24] ),
    .B(\mem[12][24] ),
    .S(net200),
    .Z(_1200_));
 MUX2_X1 _3315_ (.A(\mem[9][24] ),
    .B(\mem[13][24] ),
    .S(net200),
    .Z(_1201_));
 MUX2_X1 _3316_ (.A(_1200_),
    .B(_1201_),
    .S(net207),
    .Z(_1202_));
 MUX2_X1 _3317_ (.A(\mem[0][24] ),
    .B(\mem[4][24] ),
    .S(net200),
    .Z(_1203_));
 MUX2_X1 _3318_ (.A(\mem[1][24] ),
    .B(\mem[5][24] ),
    .S(net200),
    .Z(_1204_));
 MUX2_X1 _3319_ (.A(_1203_),
    .B(_1204_),
    .S(net207),
    .Z(_1205_));
 AOI22_X1 _3320_ (.A1(_0883_),
    .A2(_1202_),
    .B1(_1205_),
    .B2(_0880_),
    .ZN(_1206_));
 MUX2_X1 _3321_ (.A(\mem[10][24] ),
    .B(\mem[14][24] ),
    .S(net200),
    .Z(_1207_));
 MUX2_X1 _3322_ (.A(\mem[11][24] ),
    .B(\mem[15][24] ),
    .S(net200),
    .Z(_1208_));
 MUX2_X1 _3323_ (.A(_1207_),
    .B(_1208_),
    .S(net207),
    .Z(_1209_));
 MUX2_X1 _3324_ (.A(\mem[2][24] ),
    .B(\mem[6][24] ),
    .S(net200),
    .Z(_1210_));
 MUX2_X1 _3325_ (.A(\mem[3][24] ),
    .B(\mem[7][24] ),
    .S(net200),
    .Z(_1211_));
 BUF_X1 input24 (.A(wr_data[28]),
    .Z(net24));
 MUX2_X1 _3327_ (.A(_1210_),
    .B(_1211_),
    .S(net207),
    .Z(_1213_));
 AOI22_X1 _3328_ (.A1(_0894_),
    .A2(_1209_),
    .B1(_1213_),
    .B2(_0892_),
    .ZN(_1214_));
 NAND2_X1 _3329_ (.A1(_1206_),
    .A2(_1214_),
    .ZN(_1215_));
 NAND3_X1 _3330_ (.A1(net210),
    .A2(net174),
    .A3(_1215_),
    .ZN(_1216_));
 OAI21_X1 _3331_ (.A(\last_valid_data[24] ),
    .B1(net172),
    .B2(_0629_),
    .ZN(_1217_));
 AOI21_X1 _3332_ (.A(_0783_),
    .B1(_1216_),
    .B2(_1217_),
    .ZN(_0063_));
 BUF_X1 input23 (.A(wr_data[27]),
    .Z(net23));
 MUX2_X1 _3334_ (.A(\mem[8][25] ),
    .B(\mem[12][25] ),
    .S(_0002_),
    .Z(_1219_));
 BUF_X1 input22 (.A(wr_data[26]),
    .Z(net22));
 MUX2_X1 _3336_ (.A(\mem[9][25] ),
    .B(\mem[13][25] ),
    .S(net202),
    .Z(_1221_));
 MUX2_X1 _3337_ (.A(_1219_),
    .B(_1221_),
    .S(_0000_),
    .Z(_1222_));
 MUX2_X1 _3338_ (.A(\mem[0][25] ),
    .B(\mem[4][25] ),
    .S(_0002_),
    .Z(_1223_));
 MUX2_X1 _3339_ (.A(\mem[1][25] ),
    .B(\mem[5][25] ),
    .S(_0002_),
    .Z(_1224_));
 BUF_X1 input21 (.A(wr_data[25]),
    .Z(net21));
 MUX2_X1 _3341_ (.A(_1223_),
    .B(_1224_),
    .S(_0000_),
    .Z(_1226_));
 AOI22_X1 _3342_ (.A1(net190),
    .A2(_1222_),
    .B1(_1226_),
    .B2(net198),
    .ZN(_1227_));
 MUX2_X1 _3343_ (.A(\mem[10][25] ),
    .B(\mem[14][25] ),
    .S(_0002_),
    .Z(_1228_));
 MUX2_X1 _3344_ (.A(\mem[11][25] ),
    .B(\mem[15][25] ),
    .S(_0002_),
    .Z(_1229_));
 MUX2_X1 _3345_ (.A(_1228_),
    .B(_1229_),
    .S(_0000_),
    .Z(_1230_));
 MUX2_X1 _3346_ (.A(\mem[2][25] ),
    .B(\mem[6][25] ),
    .S(net200),
    .Z(_1231_));
 MUX2_X1 _3347_ (.A(\mem[3][25] ),
    .B(\mem[7][25] ),
    .S(net200),
    .Z(_1232_));
 MUX2_X1 _3348_ (.A(_1231_),
    .B(_1232_),
    .S(_0000_),
    .Z(_1233_));
 AOI22_X1 _3349_ (.A1(net188),
    .A2(_1230_),
    .B1(_1233_),
    .B2(net189),
    .ZN(_1234_));
 NAND2_X1 _3350_ (.A1(_1227_),
    .A2(_1234_),
    .ZN(_1235_));
 NAND3_X1 _3351_ (.A1(net210),
    .A2(net96),
    .A3(_1235_),
    .ZN(_1236_));
 OAI21_X1 _3352_ (.A(\last_valid_data[25] ),
    .B1(net172),
    .B2(_0629_),
    .ZN(_1237_));
 AOI21_X1 _3353_ (.A(_0783_),
    .B1(_1236_),
    .B2(_1237_),
    .ZN(_0064_));
 BUF_X1 input20 (.A(wr_data[24]),
    .Z(net20));
 MUX2_X1 _3355_ (.A(\mem[8][26] ),
    .B(\mem[12][26] ),
    .S(net200),
    .Z(_1239_));
 MUX2_X1 _3356_ (.A(\mem[9][26] ),
    .B(\mem[13][26] ),
    .S(net200),
    .Z(_1240_));
 MUX2_X1 _3357_ (.A(_1239_),
    .B(_1240_),
    .S(net207),
    .Z(_1241_));
 MUX2_X1 _3358_ (.A(\mem[0][26] ),
    .B(\mem[4][26] ),
    .S(net200),
    .Z(_1242_));
 MUX2_X1 _3359_ (.A(\mem[1][26] ),
    .B(\mem[5][26] ),
    .S(net200),
    .Z(_1243_));
 MUX2_X1 _3360_ (.A(_1242_),
    .B(_1243_),
    .S(net207),
    .Z(_1244_));
 AOI22_X1 _3361_ (.A1(net190),
    .A2(_1241_),
    .B1(_1244_),
    .B2(net198),
    .ZN(_1245_));
 MUX2_X1 _3362_ (.A(\mem[10][26] ),
    .B(\mem[14][26] ),
    .S(net200),
    .Z(_1246_));
 MUX2_X1 _3363_ (.A(\mem[11][26] ),
    .B(\mem[15][26] ),
    .S(net200),
    .Z(_1247_));
 BUF_X1 input19 (.A(wr_data[23]),
    .Z(net19));
 MUX2_X1 _3365_ (.A(_1246_),
    .B(_1247_),
    .S(net207),
    .Z(_1249_));
 MUX2_X1 _3366_ (.A(\mem[2][26] ),
    .B(\mem[6][26] ),
    .S(net200),
    .Z(_1250_));
 MUX2_X1 _3367_ (.A(\mem[3][26] ),
    .B(\mem[7][26] ),
    .S(net200),
    .Z(_1251_));
 MUX2_X1 _3368_ (.A(_1250_),
    .B(_1251_),
    .S(net207),
    .Z(_1252_));
 AOI22_X1 _3369_ (.A1(net188),
    .A2(_1249_),
    .B1(_1252_),
    .B2(net189),
    .ZN(_1253_));
 NAND2_X1 _3370_ (.A1(_1245_),
    .A2(_1253_),
    .ZN(_1254_));
 NAND3_X1 _3371_ (.A1(net210),
    .A2(net96),
    .A3(_1254_),
    .ZN(_1255_));
 OAI21_X1 _3372_ (.A(\last_valid_data[26] ),
    .B1(net172),
    .B2(_0629_),
    .ZN(_1256_));
 AOI21_X1 _3373_ (.A(_0783_),
    .B1(_1255_),
    .B2(_1256_),
    .ZN(_0065_));
 BUF_X1 input18 (.A(wr_data[22]),
    .Z(net18));
 MUX2_X1 _3375_ (.A(\mem[8][27] ),
    .B(\mem[12][27] ),
    .S(net201),
    .Z(_1258_));
 MUX2_X1 _3376_ (.A(\mem[9][27] ),
    .B(\mem[13][27] ),
    .S(net201),
    .Z(_1259_));
 BUF_X1 input17 (.A(wr_data[21]),
    .Z(net17));
 MUX2_X1 _3378_ (.A(_1258_),
    .B(_1259_),
    .S(net205),
    .Z(_1261_));
 MUX2_X1 _3379_ (.A(\mem[0][27] ),
    .B(\mem[4][27] ),
    .S(net201),
    .Z(_1262_));
 MUX2_X1 _3380_ (.A(\mem[1][27] ),
    .B(\mem[5][27] ),
    .S(net201),
    .Z(_1263_));
 MUX2_X1 _3381_ (.A(_1262_),
    .B(_1263_),
    .S(net205),
    .Z(_1264_));
 AOI22_X1 _3382_ (.A1(net190),
    .A2(_1261_),
    .B1(_1264_),
    .B2(net198),
    .ZN(_1265_));
 MUX2_X1 _3383_ (.A(\mem[10][27] ),
    .B(\mem[14][27] ),
    .S(net201),
    .Z(_1266_));
 MUX2_X1 _3384_ (.A(\mem[11][27] ),
    .B(\mem[15][27] ),
    .S(net201),
    .Z(_1267_));
 MUX2_X1 _3385_ (.A(_1266_),
    .B(_1267_),
    .S(net205),
    .Z(_1268_));
 MUX2_X1 _3386_ (.A(\mem[2][27] ),
    .B(\mem[6][27] ),
    .S(net201),
    .Z(_1269_));
 MUX2_X1 _3387_ (.A(\mem[3][27] ),
    .B(\mem[7][27] ),
    .S(net201),
    .Z(_1270_));
 MUX2_X1 _3388_ (.A(_1269_),
    .B(_1270_),
    .S(net205),
    .Z(_1271_));
 AOI22_X1 _3389_ (.A1(net188),
    .A2(_1268_),
    .B1(_1271_),
    .B2(net189),
    .ZN(_1272_));
 NAND2_X1 _3390_ (.A1(_1265_),
    .A2(_1272_),
    .ZN(_1273_));
 NAND3_X1 _3391_ (.A1(net210),
    .A2(net174),
    .A3(_1273_),
    .ZN(_1274_));
 OAI21_X1 _3392_ (.A(\last_valid_data[27] ),
    .B1(net172),
    .B2(_0629_),
    .ZN(_1275_));
 AOI21_X1 _3393_ (.A(_0783_),
    .B1(_1274_),
    .B2(_1275_),
    .ZN(_0066_));
 MUX2_X1 _3394_ (.A(\mem[8][28] ),
    .B(\mem[12][28] ),
    .S(net201),
    .Z(_1276_));
 MUX2_X1 _3395_ (.A(\mem[9][28] ),
    .B(\mem[13][28] ),
    .S(net201),
    .Z(_1277_));
 MUX2_X1 _3396_ (.A(_1276_),
    .B(_1277_),
    .S(net207),
    .Z(_1278_));
 MUX2_X1 _3397_ (.A(\mem[0][28] ),
    .B(\mem[4][28] ),
    .S(net201),
    .Z(_1279_));
 MUX2_X1 _3398_ (.A(\mem[1][28] ),
    .B(\mem[5][28] ),
    .S(net201),
    .Z(_1280_));
 MUX2_X1 _3399_ (.A(_1279_),
    .B(_1280_),
    .S(net207),
    .Z(_1281_));
 BUF_X1 input16 (.A(wr_data[20]),
    .Z(net16));
 AOI22_X1 _3401_ (.A1(_0883_),
    .A2(_1278_),
    .B1(_1281_),
    .B2(_0880_),
    .ZN(_1283_));
 MUX2_X1 _3402_ (.A(\mem[10][28] ),
    .B(\mem[14][28] ),
    .S(net201),
    .Z(_1284_));
 MUX2_X1 _3403_ (.A(\mem[11][28] ),
    .B(\mem[15][28] ),
    .S(net201),
    .Z(_1285_));
 MUX2_X1 _3404_ (.A(_1284_),
    .B(_1285_),
    .S(net207),
    .Z(_1286_));
 BUF_X1 input15 (.A(wr_data[1]),
    .Z(net15));
 MUX2_X1 _3406_ (.A(\mem[2][28] ),
    .B(\mem[6][28] ),
    .S(net201),
    .Z(_1288_));
 MUX2_X1 _3407_ (.A(\mem[3][28] ),
    .B(\mem[7][28] ),
    .S(net201),
    .Z(_1289_));
 MUX2_X1 _3408_ (.A(_1288_),
    .B(_1289_),
    .S(net207),
    .Z(_1290_));
 BUF_X1 input14 (.A(wr_data[19]),
    .Z(net14));
 AOI22_X1 _3410_ (.A1(_0894_),
    .A2(_1286_),
    .B1(_1290_),
    .B2(_0892_),
    .ZN(_1292_));
 NAND2_X1 _3411_ (.A1(_1283_),
    .A2(_1292_),
    .ZN(_1293_));
 NAND3_X1 _3412_ (.A1(net210),
    .A2(net174),
    .A3(_1293_),
    .ZN(_1294_));
 BUF_X1 input13 (.A(wr_data[18]),
    .Z(net13));
 OAI21_X1 _3414_ (.A(\last_valid_data[28] ),
    .B1(net172),
    .B2(net209),
    .ZN(_1296_));
 AOI21_X1 _3415_ (.A(net208),
    .B1(_1294_),
    .B2(_1296_),
    .ZN(_0067_));
 BUF_X1 input12 (.A(wr_data[17]),
    .Z(net12));
 MUX2_X1 _3417_ (.A(\mem[8][29] ),
    .B(\mem[12][29] ),
    .S(net201),
    .Z(_1298_));
 MUX2_X1 _3418_ (.A(\mem[9][29] ),
    .B(\mem[13][29] ),
    .S(net201),
    .Z(_1299_));
 MUX2_X1 _3419_ (.A(_1298_),
    .B(_1299_),
    .S(net207),
    .Z(_1300_));
 MUX2_X1 _3420_ (.A(\mem[0][29] ),
    .B(\mem[4][29] ),
    .S(net201),
    .Z(_1301_));
 MUX2_X1 _3421_ (.A(\mem[1][29] ),
    .B(\mem[5][29] ),
    .S(net201),
    .Z(_1302_));
 MUX2_X1 _3422_ (.A(_1301_),
    .B(_1302_),
    .S(net207),
    .Z(_1303_));
 AOI22_X1 _3423_ (.A1(net190),
    .A2(_1300_),
    .B1(_1303_),
    .B2(net198),
    .ZN(_1304_));
 BUF_X1 input11 (.A(wr_data[16]),
    .Z(net11));
 MUX2_X1 _3425_ (.A(\mem[10][29] ),
    .B(\mem[14][29] ),
    .S(net201),
    .Z(_1306_));
 MUX2_X1 _3426_ (.A(\mem[11][29] ),
    .B(\mem[15][29] ),
    .S(net201),
    .Z(_1307_));
 MUX2_X1 _3427_ (.A(_1306_),
    .B(_1307_),
    .S(net207),
    .Z(_1308_));
 MUX2_X1 _3428_ (.A(\mem[2][29] ),
    .B(\mem[6][29] ),
    .S(net201),
    .Z(_1309_));
 BUF_X1 input10 (.A(wr_data[15]),
    .Z(net10));
 MUX2_X1 _3430_ (.A(\mem[3][29] ),
    .B(\mem[7][29] ),
    .S(net201),
    .Z(_1311_));
 MUX2_X1 _3431_ (.A(_1309_),
    .B(_1311_),
    .S(net205),
    .Z(_1312_));
 AOI22_X1 _3432_ (.A1(_0894_),
    .A2(_1308_),
    .B1(_1312_),
    .B2(_0892_),
    .ZN(_1313_));
 NAND2_X1 _3433_ (.A1(_1304_),
    .A2(_1313_),
    .ZN(_1314_));
 NAND3_X1 _3434_ (.A1(net210),
    .A2(net174),
    .A3(_1314_),
    .ZN(_1315_));
 OAI21_X1 _3435_ (.A(\last_valid_data[29] ),
    .B1(net172),
    .B2(net209),
    .ZN(_1316_));
 AOI21_X1 _3436_ (.A(net208),
    .B1(_1315_),
    .B2(_1316_),
    .ZN(_0068_));
 MUX2_X1 _3437_ (.A(\mem[8][2] ),
    .B(\mem[12][2] ),
    .S(net201),
    .Z(_1317_));
 MUX2_X1 _3438_ (.A(\mem[9][2] ),
    .B(\mem[13][2] ),
    .S(net201),
    .Z(_1318_));
 MUX2_X1 _3439_ (.A(_1317_),
    .B(_1318_),
    .S(net205),
    .Z(_1319_));
 BUF_X1 input9 (.A(wr_data[14]),
    .Z(net9));
 MUX2_X1 _3441_ (.A(\mem[0][2] ),
    .B(\mem[4][2] ),
    .S(net201),
    .Z(_1321_));
 MUX2_X1 _3442_ (.A(\mem[1][2] ),
    .B(\mem[5][2] ),
    .S(net201),
    .Z(_1322_));
 MUX2_X1 _3443_ (.A(_1321_),
    .B(_1322_),
    .S(net205),
    .Z(_1323_));
 AOI22_X1 _3444_ (.A1(net190),
    .A2(_1319_),
    .B1(_1323_),
    .B2(net198),
    .ZN(_1324_));
 MUX2_X1 _3445_ (.A(\mem[10][2] ),
    .B(\mem[14][2] ),
    .S(net201),
    .Z(_1325_));
 MUX2_X1 _3446_ (.A(\mem[11][2] ),
    .B(\mem[15][2] ),
    .S(net201),
    .Z(_1326_));
 MUX2_X1 _3447_ (.A(_1325_),
    .B(_1326_),
    .S(net205),
    .Z(_1327_));
 MUX2_X1 _3448_ (.A(\mem[2][2] ),
    .B(\mem[6][2] ),
    .S(net201),
    .Z(_1328_));
 MUX2_X1 _3449_ (.A(\mem[3][2] ),
    .B(\mem[7][2] ),
    .S(net201),
    .Z(_1329_));
 MUX2_X1 _3450_ (.A(_1328_),
    .B(_1329_),
    .S(net205),
    .Z(_1330_));
 AOI22_X1 _3451_ (.A1(_0894_),
    .A2(_1327_),
    .B1(_1330_),
    .B2(_0892_),
    .ZN(_1331_));
 NAND2_X1 _3452_ (.A1(_1324_),
    .A2(_1331_),
    .ZN(_1332_));
 NAND3_X1 _3453_ (.A1(net210),
    .A2(net174),
    .A3(_1332_),
    .ZN(_1333_));
 OAI21_X1 _3454_ (.A(\last_valid_data[2] ),
    .B1(net172),
    .B2(net209),
    .ZN(_1334_));
 AOI21_X1 _3455_ (.A(net208),
    .B1(_1333_),
    .B2(_1334_),
    .ZN(_0069_));
 MUX2_X1 _3456_ (.A(\mem[8][30] ),
    .B(\mem[12][30] ),
    .S(net201),
    .Z(_1335_));
 MUX2_X1 _3457_ (.A(\mem[9][30] ),
    .B(\mem[13][30] ),
    .S(net201),
    .Z(_1336_));
 MUX2_X1 _3458_ (.A(_1335_),
    .B(_1336_),
    .S(net205),
    .Z(_1337_));
 MUX2_X1 _3459_ (.A(\mem[0][30] ),
    .B(\mem[4][30] ),
    .S(net201),
    .Z(_1338_));
 MUX2_X1 _3460_ (.A(\mem[1][30] ),
    .B(\mem[5][30] ),
    .S(net201),
    .Z(_1339_));
 MUX2_X1 _3461_ (.A(_1338_),
    .B(_1339_),
    .S(net205),
    .Z(_1340_));
 AOI22_X1 _3462_ (.A1(net190),
    .A2(_1337_),
    .B1(_1340_),
    .B2(net198),
    .ZN(_1341_));
 MUX2_X1 _3463_ (.A(\mem[10][30] ),
    .B(\mem[14][30] ),
    .S(net201),
    .Z(_1342_));
 MUX2_X1 _3464_ (.A(\mem[11][30] ),
    .B(\mem[15][30] ),
    .S(net201),
    .Z(_1343_));
 MUX2_X1 _3465_ (.A(_1342_),
    .B(_1343_),
    .S(net205),
    .Z(_1344_));
 MUX2_X1 _3466_ (.A(\mem[2][30] ),
    .B(\mem[6][30] ),
    .S(net201),
    .Z(_1345_));
 MUX2_X1 _3467_ (.A(\mem[3][30] ),
    .B(\mem[7][30] ),
    .S(net201),
    .Z(_1346_));
 MUX2_X1 _3468_ (.A(_1345_),
    .B(_1346_),
    .S(net205),
    .Z(_1347_));
 AOI22_X1 _3469_ (.A1(net188),
    .A2(_1344_),
    .B1(_1347_),
    .B2(_0892_),
    .ZN(_1348_));
 NAND2_X1 _3470_ (.A1(_1341_),
    .A2(_1348_),
    .ZN(_1349_));
 NAND3_X1 _3471_ (.A1(net210),
    .A2(net174),
    .A3(_1349_),
    .ZN(_1350_));
 OAI21_X1 _3472_ (.A(\last_valid_data[30] ),
    .B1(net172),
    .B2(net209),
    .ZN(_1351_));
 AOI21_X1 _3473_ (.A(net208),
    .B1(_1350_),
    .B2(_1351_),
    .ZN(_0070_));
 MUX2_X1 _3474_ (.A(\mem[8][31] ),
    .B(\mem[12][31] ),
    .S(net203),
    .Z(_1352_));
 MUX2_X1 _3475_ (.A(\mem[9][31] ),
    .B(\mem[13][31] ),
    .S(net203),
    .Z(_1353_));
 MUX2_X1 _3476_ (.A(_1352_),
    .B(_1353_),
    .S(net206),
    .Z(_1354_));
 MUX2_X1 _3477_ (.A(\mem[0][31] ),
    .B(\mem[4][31] ),
    .S(net201),
    .Z(_1355_));
 MUX2_X1 _3478_ (.A(\mem[1][31] ),
    .B(\mem[5][31] ),
    .S(net201),
    .Z(_1356_));
 MUX2_X1 _3479_ (.A(_1355_),
    .B(_1356_),
    .S(net205),
    .Z(_1357_));
 AOI22_X1 _3480_ (.A1(net190),
    .A2(_1354_),
    .B1(_1357_),
    .B2(net198),
    .ZN(_1358_));
 MUX2_X1 _3481_ (.A(\mem[10][31] ),
    .B(\mem[14][31] ),
    .S(net203),
    .Z(_1359_));
 MUX2_X1 _3482_ (.A(\mem[11][31] ),
    .B(\mem[15][31] ),
    .S(net203),
    .Z(_1360_));
 MUX2_X1 _3483_ (.A(_1359_),
    .B(_1360_),
    .S(net206),
    .Z(_1361_));
 MUX2_X1 _3484_ (.A(\mem[2][31] ),
    .B(\mem[6][31] ),
    .S(net201),
    .Z(_1362_));
 MUX2_X1 _3485_ (.A(\mem[3][31] ),
    .B(\mem[7][31] ),
    .S(net201),
    .Z(_1363_));
 MUX2_X1 _3486_ (.A(_1362_),
    .B(_1363_),
    .S(net206),
    .Z(_1364_));
 AOI22_X1 _3487_ (.A1(net188),
    .A2(_1361_),
    .B1(_1364_),
    .B2(net189),
    .ZN(_1365_));
 NAND2_X1 _3488_ (.A1(_1358_),
    .A2(_1365_),
    .ZN(_1366_));
 NAND3_X1 _3489_ (.A1(net210),
    .A2(net174),
    .A3(_1366_),
    .ZN(_1367_));
 OAI21_X1 _3490_ (.A(\last_valid_data[31] ),
    .B1(net172),
    .B2(net209),
    .ZN(_1368_));
 AOI21_X1 _3491_ (.A(net208),
    .B1(_1367_),
    .B2(_1368_),
    .ZN(_0071_));
 MUX2_X1 _3492_ (.A(\mem[8][3] ),
    .B(\mem[12][3] ),
    .S(net201),
    .Z(_1369_));
 MUX2_X1 _3493_ (.A(\mem[9][3] ),
    .B(\mem[13][3] ),
    .S(net201),
    .Z(_1370_));
 MUX2_X1 _3494_ (.A(_1369_),
    .B(_1370_),
    .S(net206),
    .Z(_1371_));
 MUX2_X1 _3495_ (.A(\mem[0][3] ),
    .B(\mem[4][3] ),
    .S(net201),
    .Z(_1372_));
 MUX2_X1 _3496_ (.A(\mem[1][3] ),
    .B(\mem[5][3] ),
    .S(net201),
    .Z(_1373_));
 MUX2_X1 _3497_ (.A(_1372_),
    .B(_1373_),
    .S(net205),
    .Z(_1374_));
 AOI22_X1 _3498_ (.A1(net190),
    .A2(_1371_),
    .B1(_1374_),
    .B2(net198),
    .ZN(_1375_));
 MUX2_X1 _3499_ (.A(\mem[10][3] ),
    .B(\mem[14][3] ),
    .S(net201),
    .Z(_1376_));
 MUX2_X1 _3500_ (.A(\mem[11][3] ),
    .B(\mem[15][3] ),
    .S(net201),
    .Z(_1377_));
 MUX2_X1 _3501_ (.A(_1376_),
    .B(_1377_),
    .S(net205),
    .Z(_1378_));
 MUX2_X1 _3502_ (.A(\mem[2][3] ),
    .B(\mem[6][3] ),
    .S(net201),
    .Z(_1379_));
 MUX2_X1 _3503_ (.A(\mem[3][3] ),
    .B(\mem[7][3] ),
    .S(net201),
    .Z(_1380_));
 MUX2_X1 _3504_ (.A(_1379_),
    .B(_1380_),
    .S(net205),
    .Z(_1381_));
 AOI22_X1 _3505_ (.A1(net188),
    .A2(_1378_),
    .B1(_1381_),
    .B2(net189),
    .ZN(_1382_));
 NAND2_X1 _3506_ (.A1(_1375_),
    .A2(_1382_),
    .ZN(_1383_));
 NAND3_X1 _3507_ (.A1(net210),
    .A2(net174),
    .A3(_1383_),
    .ZN(_1384_));
 OAI21_X1 _3508_ (.A(\last_valid_data[3] ),
    .B1(net172),
    .B2(net209),
    .ZN(_1385_));
 AOI21_X1 _3509_ (.A(net208),
    .B1(_1384_),
    .B2(_1385_),
    .ZN(_0072_));
 MUX2_X1 _3510_ (.A(\mem[8][4] ),
    .B(\mem[12][4] ),
    .S(net203),
    .Z(_1386_));
 MUX2_X1 _3511_ (.A(\mem[9][4] ),
    .B(\mem[13][4] ),
    .S(net203),
    .Z(_1387_));
 MUX2_X1 _3512_ (.A(_1386_),
    .B(_1387_),
    .S(net206),
    .Z(_1388_));
 MUX2_X1 _3513_ (.A(\mem[0][4] ),
    .B(\mem[4][4] ),
    .S(net201),
    .Z(_1389_));
 MUX2_X1 _3514_ (.A(\mem[1][4] ),
    .B(\mem[5][4] ),
    .S(net201),
    .Z(_1390_));
 MUX2_X1 _3515_ (.A(_1389_),
    .B(_1390_),
    .S(net206),
    .Z(_1391_));
 AOI22_X1 _3516_ (.A1(net190),
    .A2(_1388_),
    .B1(_1391_),
    .B2(net198),
    .ZN(_1392_));
 MUX2_X1 _3517_ (.A(\mem[10][4] ),
    .B(\mem[14][4] ),
    .S(net203),
    .Z(_1393_));
 MUX2_X1 _3518_ (.A(\mem[11][4] ),
    .B(\mem[15][4] ),
    .S(net203),
    .Z(_1394_));
 MUX2_X1 _3519_ (.A(_1393_),
    .B(_1394_),
    .S(net206),
    .Z(_1395_));
 MUX2_X1 _3520_ (.A(\mem[2][4] ),
    .B(\mem[6][4] ),
    .S(net201),
    .Z(_1396_));
 MUX2_X1 _3521_ (.A(\mem[3][4] ),
    .B(\mem[7][4] ),
    .S(net201),
    .Z(_1397_));
 MUX2_X1 _3522_ (.A(_1396_),
    .B(_1397_),
    .S(net206),
    .Z(_1398_));
 AOI22_X1 _3523_ (.A1(net188),
    .A2(_1395_),
    .B1(_1398_),
    .B2(net189),
    .ZN(_1399_));
 NAND2_X1 _3524_ (.A1(_1392_),
    .A2(_1399_),
    .ZN(_1400_));
 NAND3_X1 _3525_ (.A1(net210),
    .A2(net174),
    .A3(_1400_),
    .ZN(_1401_));
 OAI21_X1 _3526_ (.A(\last_valid_data[4] ),
    .B1(net172),
    .B2(net209),
    .ZN(_1402_));
 AOI21_X1 _3527_ (.A(net208),
    .B1(_1401_),
    .B2(_1402_),
    .ZN(_0073_));
 MUX2_X1 _3528_ (.A(\mem[8][5] ),
    .B(\mem[12][5] ),
    .S(net203),
    .Z(_1403_));
 MUX2_X1 _3529_ (.A(\mem[9][5] ),
    .B(\mem[13][5] ),
    .S(net203),
    .Z(_1404_));
 MUX2_X1 _3530_ (.A(_1403_),
    .B(_1404_),
    .S(net206),
    .Z(_1405_));
 MUX2_X1 _3531_ (.A(\mem[0][5] ),
    .B(\mem[4][5] ),
    .S(net203),
    .Z(_1406_));
 MUX2_X1 _3532_ (.A(\mem[1][5] ),
    .B(\mem[5][5] ),
    .S(net203),
    .Z(_1407_));
 MUX2_X1 _3533_ (.A(_1406_),
    .B(_1407_),
    .S(net206),
    .Z(_1408_));
 AOI22_X1 _3534_ (.A1(net190),
    .A2(_1405_),
    .B1(_1408_),
    .B2(net198),
    .ZN(_1409_));
 MUX2_X1 _3535_ (.A(\mem[10][5] ),
    .B(\mem[14][5] ),
    .S(net203),
    .Z(_1410_));
 MUX2_X1 _3536_ (.A(\mem[11][5] ),
    .B(\mem[15][5] ),
    .S(net203),
    .Z(_1411_));
 MUX2_X1 _3537_ (.A(_1410_),
    .B(_1411_),
    .S(net206),
    .Z(_1412_));
 MUX2_X1 _3538_ (.A(\mem[2][5] ),
    .B(\mem[6][5] ),
    .S(net203),
    .Z(_1413_));
 MUX2_X1 _3539_ (.A(\mem[3][5] ),
    .B(\mem[7][5] ),
    .S(net203),
    .Z(_1414_));
 MUX2_X1 _3540_ (.A(_1413_),
    .B(_1414_),
    .S(net206),
    .Z(_1415_));
 AOI22_X1 _3541_ (.A1(net188),
    .A2(_1412_),
    .B1(_1415_),
    .B2(net189),
    .ZN(_1416_));
 NAND2_X1 _3542_ (.A1(_1409_),
    .A2(_1416_),
    .ZN(_1417_));
 NAND3_X1 _3543_ (.A1(net210),
    .A2(net173),
    .A3(_1417_),
    .ZN(_1418_));
 OAI21_X1 _3544_ (.A(\last_valid_data[5] ),
    .B1(net172),
    .B2(net209),
    .ZN(_1419_));
 AOI21_X1 _3545_ (.A(net208),
    .B1(_1418_),
    .B2(_1419_),
    .ZN(_0074_));
 MUX2_X1 _3546_ (.A(\mem[8][6] ),
    .B(\mem[12][6] ),
    .S(net203),
    .Z(_1420_));
 MUX2_X1 _3547_ (.A(\mem[9][6] ),
    .B(\mem[13][6] ),
    .S(net203),
    .Z(_1421_));
 MUX2_X1 _3548_ (.A(_1420_),
    .B(_1421_),
    .S(net206),
    .Z(_1422_));
 MUX2_X1 _3549_ (.A(\mem[0][6] ),
    .B(\mem[4][6] ),
    .S(net203),
    .Z(_1423_));
 MUX2_X1 _3550_ (.A(\mem[1][6] ),
    .B(\mem[5][6] ),
    .S(net203),
    .Z(_1424_));
 MUX2_X1 _3551_ (.A(_1423_),
    .B(_1424_),
    .S(net206),
    .Z(_1425_));
 AOI22_X1 _3552_ (.A1(net190),
    .A2(_1422_),
    .B1(_1425_),
    .B2(net198),
    .ZN(_1426_));
 MUX2_X1 _3553_ (.A(\mem[10][6] ),
    .B(\mem[14][6] ),
    .S(net203),
    .Z(_1427_));
 MUX2_X1 _3554_ (.A(\mem[11][6] ),
    .B(\mem[15][6] ),
    .S(net203),
    .Z(_1428_));
 MUX2_X1 _3555_ (.A(_1427_),
    .B(_1428_),
    .S(net206),
    .Z(_1429_));
 MUX2_X1 _3556_ (.A(\mem[2][6] ),
    .B(\mem[6][6] ),
    .S(net203),
    .Z(_1430_));
 MUX2_X1 _3557_ (.A(\mem[3][6] ),
    .B(\mem[7][6] ),
    .S(net203),
    .Z(_1431_));
 MUX2_X1 _3558_ (.A(_1430_),
    .B(_1431_),
    .S(net206),
    .Z(_1432_));
 AOI22_X1 _3559_ (.A1(net188),
    .A2(_1429_),
    .B1(_1432_),
    .B2(net189),
    .ZN(_1433_));
 NAND2_X1 _3560_ (.A1(_1426_),
    .A2(_1433_),
    .ZN(_1434_));
 NAND3_X1 _3561_ (.A1(net210),
    .A2(net173),
    .A3(_1434_),
    .ZN(_1435_));
 OAI21_X1 _3562_ (.A(\last_valid_data[6] ),
    .B1(net172),
    .B2(net209),
    .ZN(_1436_));
 AOI21_X1 _3563_ (.A(net208),
    .B1(_1435_),
    .B2(_1436_),
    .ZN(_0075_));
 MUX2_X1 _3564_ (.A(\mem[8][7] ),
    .B(\mem[12][7] ),
    .S(net203),
    .Z(_1437_));
 MUX2_X1 _3565_ (.A(\mem[9][7] ),
    .B(\mem[13][7] ),
    .S(net203),
    .Z(_1438_));
 MUX2_X1 _3566_ (.A(_1437_),
    .B(_1438_),
    .S(net206),
    .Z(_1439_));
 MUX2_X1 _3567_ (.A(\mem[0][7] ),
    .B(\mem[4][7] ),
    .S(net203),
    .Z(_1440_));
 MUX2_X1 _3568_ (.A(\mem[1][7] ),
    .B(\mem[5][7] ),
    .S(net203),
    .Z(_1441_));
 MUX2_X1 _3569_ (.A(_1440_),
    .B(_1441_),
    .S(net206),
    .Z(_1442_));
 AOI22_X1 _3570_ (.A1(net190),
    .A2(_1439_),
    .B1(_1442_),
    .B2(net198),
    .ZN(_1443_));
 MUX2_X1 _3571_ (.A(\mem[10][7] ),
    .B(\mem[14][7] ),
    .S(net203),
    .Z(_1444_));
 MUX2_X1 _3572_ (.A(\mem[11][7] ),
    .B(\mem[15][7] ),
    .S(net203),
    .Z(_1445_));
 MUX2_X1 _3573_ (.A(_1444_),
    .B(_1445_),
    .S(net206),
    .Z(_1446_));
 MUX2_X1 _3574_ (.A(\mem[2][7] ),
    .B(\mem[6][7] ),
    .S(net203),
    .Z(_1447_));
 MUX2_X1 _3575_ (.A(\mem[3][7] ),
    .B(\mem[7][7] ),
    .S(net203),
    .Z(_1448_));
 MUX2_X1 _3576_ (.A(_1447_),
    .B(_1448_),
    .S(net206),
    .Z(_1449_));
 AOI22_X1 _3577_ (.A1(net188),
    .A2(_1446_),
    .B1(_1449_),
    .B2(net189),
    .ZN(_1450_));
 NAND2_X1 _3578_ (.A1(_1443_),
    .A2(_1450_),
    .ZN(_1451_));
 NAND3_X1 _3579_ (.A1(net210),
    .A2(net173),
    .A3(_1451_),
    .ZN(_1452_));
 OAI21_X1 _3580_ (.A(\last_valid_data[7] ),
    .B1(net44),
    .B2(net209),
    .ZN(_1453_));
 AOI21_X1 _3581_ (.A(net208),
    .B1(_1452_),
    .B2(_1453_),
    .ZN(_0076_));
 MUX2_X1 _3582_ (.A(\mem[8][8] ),
    .B(\mem[12][8] ),
    .S(net203),
    .Z(_1454_));
 MUX2_X1 _3583_ (.A(\mem[9][8] ),
    .B(\mem[13][8] ),
    .S(net203),
    .Z(_1455_));
 MUX2_X1 _3584_ (.A(_1454_),
    .B(_1455_),
    .S(net206),
    .Z(_1456_));
 MUX2_X1 _3585_ (.A(\mem[0][8] ),
    .B(\mem[4][8] ),
    .S(net203),
    .Z(_1457_));
 MUX2_X1 _3586_ (.A(\mem[1][8] ),
    .B(\mem[5][8] ),
    .S(net203),
    .Z(_1458_));
 MUX2_X1 _3587_ (.A(_1457_),
    .B(_1458_),
    .S(net206),
    .Z(_1459_));
 AOI22_X1 _3588_ (.A1(net190),
    .A2(_1456_),
    .B1(_1459_),
    .B2(net198),
    .ZN(_1460_));
 MUX2_X1 _3589_ (.A(\mem[10][8] ),
    .B(\mem[14][8] ),
    .S(net203),
    .Z(_1461_));
 MUX2_X1 _3590_ (.A(\mem[11][8] ),
    .B(\mem[15][8] ),
    .S(net203),
    .Z(_1462_));
 MUX2_X1 _3591_ (.A(_1461_),
    .B(_1462_),
    .S(net206),
    .Z(_1463_));
 MUX2_X1 _3592_ (.A(\mem[2][8] ),
    .B(\mem[6][8] ),
    .S(net203),
    .Z(_1464_));
 MUX2_X1 _3593_ (.A(\mem[3][8] ),
    .B(\mem[7][8] ),
    .S(net203),
    .Z(_1465_));
 MUX2_X1 _3594_ (.A(_1464_),
    .B(_1465_),
    .S(net206),
    .Z(_1466_));
 AOI22_X1 _3595_ (.A1(net188),
    .A2(_1463_),
    .B1(_1466_),
    .B2(net189),
    .ZN(_1467_));
 NAND2_X1 _3596_ (.A1(_1460_),
    .A2(_1467_),
    .ZN(_1468_));
 NAND3_X1 _3597_ (.A1(net210),
    .A2(net173),
    .A3(_1468_),
    .ZN(_1469_));
 OAI21_X1 _3598_ (.A(\last_valid_data[8] ),
    .B1(net44),
    .B2(net209),
    .ZN(_1470_));
 AOI21_X1 _3599_ (.A(net208),
    .B1(_1469_),
    .B2(_1470_),
    .ZN(_0077_));
 MUX2_X1 _3600_ (.A(\mem[8][9] ),
    .B(\mem[12][9] ),
    .S(net203),
    .Z(_1471_));
 MUX2_X1 _3601_ (.A(\mem[9][9] ),
    .B(\mem[13][9] ),
    .S(net203),
    .Z(_1472_));
 MUX2_X1 _3602_ (.A(_1471_),
    .B(_1472_),
    .S(net206),
    .Z(_1473_));
 MUX2_X1 _3603_ (.A(\mem[0][9] ),
    .B(\mem[4][9] ),
    .S(net203),
    .Z(_1474_));
 MUX2_X1 _3604_ (.A(\mem[1][9] ),
    .B(\mem[5][9] ),
    .S(net203),
    .Z(_1475_));
 MUX2_X1 _3605_ (.A(_1474_),
    .B(_1475_),
    .S(net206),
    .Z(_1476_));
 AOI22_X1 _3606_ (.A1(net190),
    .A2(_1473_),
    .B1(_1476_),
    .B2(net198),
    .ZN(_1477_));
 MUX2_X1 _3607_ (.A(\mem[10][9] ),
    .B(\mem[14][9] ),
    .S(net203),
    .Z(_1478_));
 MUX2_X1 _3608_ (.A(\mem[11][9] ),
    .B(\mem[15][9] ),
    .S(net203),
    .Z(_1479_));
 MUX2_X1 _3609_ (.A(_1478_),
    .B(_1479_),
    .S(net206),
    .Z(_1480_));
 MUX2_X1 _3610_ (.A(\mem[2][9] ),
    .B(\mem[6][9] ),
    .S(net203),
    .Z(_1481_));
 MUX2_X1 _3611_ (.A(\mem[3][9] ),
    .B(\mem[7][9] ),
    .S(net203),
    .Z(_1482_));
 MUX2_X1 _3612_ (.A(_1481_),
    .B(_1482_),
    .S(net206),
    .Z(_1483_));
 AOI22_X1 _3613_ (.A1(net188),
    .A2(_1480_),
    .B1(_1483_),
    .B2(net189),
    .ZN(_1484_));
 NAND2_X1 _3614_ (.A1(_1477_),
    .A2(_1484_),
    .ZN(_1485_));
 NAND3_X1 _3615_ (.A1(net210),
    .A2(net173),
    .A3(_1485_),
    .ZN(_1486_));
 OAI21_X1 _3616_ (.A(\last_valid_data[9] ),
    .B1(net44),
    .B2(net209),
    .ZN(_1487_));
 AOI21_X1 _3617_ (.A(net208),
    .B1(_1486_),
    .B2(_1487_),
    .ZN(_0078_));
 BUF_X1 input8 (.A(wr_data[13]),
    .Z(net8));
 INV_X1 _3619_ (.A(last_valid_data_available),
    .ZN(_1489_));
 AOI21_X1 _3620_ (.A(net208),
    .B1(_0787_),
    .B2(_1489_),
    .ZN(_0079_));
 NAND2_X1 _3621_ (.A1(_0004_),
    .A2(net3),
    .ZN(_1490_));
 OAI21_X1 _3622_ (.A(_0782_),
    .B1(_1490_),
    .B2(_0787_),
    .ZN(_0592_));
 AOI21_X1 _3623_ (.A(_0783_),
    .B1(_0790_),
    .B2(_0791_),
    .ZN(_0593_));
 MUX2_X1 _3624_ (.A(_0792_),
    .B(_0793_),
    .S(_0794_),
    .Z(_0594_));
 AOI21_X1 _3625_ (.A(net208),
    .B1(_0796_),
    .B2(_0797_),
    .ZN(_0595_));
 NAND4_X1 _3626_ (.A1(net210),
    .A2(_0014_),
    .A3(\rd_ptr[2] ),
    .A4(\rd_ptr[3] ),
    .ZN(_1491_));
 OAI21_X1 _3627_ (.A(\rd_ptr[4] ),
    .B1(net172),
    .B2(_1491_),
    .ZN(_1492_));
 OR3_X1 _3628_ (.A1(\rd_ptr[4] ),
    .A2(net172),
    .A3(_1491_),
    .ZN(_1493_));
 AOI21_X1 _3629_ (.A(net208),
    .B1(_1492_),
    .B2(_1493_),
    .ZN(_0596_));
 AND2_X1 _3630_ (.A1(\wr_ptr[0] ),
    .A2(net3),
    .ZN(_1494_));
 AND2_X1 _3631_ (.A1(_0018_),
    .A2(net3),
    .ZN(_1495_));
 AND2_X1 _3632_ (.A1(net36),
    .A2(net98),
    .ZN(_1496_));
 MUX2_X1 _3633_ (.A(_1494_),
    .B(_1495_),
    .S(_1496_),
    .Z(_0597_));
 AND2_X1 _3634_ (.A1(\wr_ptr[1] ),
    .A2(net3),
    .ZN(_1497_));
 AND2_X1 _3635_ (.A1(_0020_),
    .A2(net3),
    .ZN(_1498_));
 MUX2_X1 _3636_ (.A(_1497_),
    .B(_1498_),
    .S(_1496_),
    .Z(_0598_));
 NOR2_X1 _3637_ (.A1(\wr_ptr[2] ),
    .A2(_0783_),
    .ZN(_1499_));
 AND2_X1 _3638_ (.A1(\wr_ptr[2] ),
    .A2(net3),
    .ZN(_1500_));
 NAND3_X1 _3639_ (.A1(net36),
    .A2(_0023_),
    .A3(net98),
    .ZN(_1501_));
 MUX2_X1 _3640_ (.A(_1499_),
    .B(_1500_),
    .S(_1501_),
    .Z(_0599_));
 NOR2_X1 _3641_ (.A1(\wr_ptr[3] ),
    .A2(_0783_),
    .ZN(_1502_));
 NOR2_X1 _3642_ (.A1(_0704_),
    .A2(_0783_),
    .ZN(_1503_));
 NAND4_X1 _3643_ (.A1(\wr_ptr[1] ),
    .A2(\wr_ptr[0] ),
    .A3(net98),
    .A4(_0715_),
    .ZN(_1504_));
 MUX2_X1 _3644_ (.A(_1502_),
    .B(_1503_),
    .S(_1504_),
    .Z(_0600_));
 NOR2_X1 _3645_ (.A1(\wr_ptr[4] ),
    .A2(_0783_),
    .ZN(_1505_));
 AND2_X1 _3646_ (.A1(\wr_ptr[4] ),
    .A2(net3),
    .ZN(_1506_));
 NAND3_X1 _3647_ (.A1(_0023_),
    .A2(net98),
    .A3(_0716_),
    .ZN(_1507_));
 MUX2_X1 _3648_ (.A(_1505_),
    .B(_1506_),
    .S(_1507_),
    .Z(_0601_));
 XOR2_X1 _3649_ (.A(net40),
    .B(_0025_),
    .Z(_1508_));
 NOR4_X1 _3650_ (.A1(net41),
    .A2(net42),
    .A3(net43),
    .A4(_1508_),
    .ZN(net37));
 NAND2_X1 _3651_ (.A1(net40),
    .A2(net41),
    .ZN(_1509_));
 OAI21_X1 _3652_ (.A(_0617_),
    .B1(_1509_),
    .B2(_0612_),
    .ZN(net38));
 NOR2_X1 _3653_ (.A1(_0633_),
    .A2(net98),
    .ZN(net63));
 NAND2_X1 _3654_ (.A1(net173),
    .A2(_0899_),
    .ZN(_1510_));
 BUF_X1 input7 (.A(wr_data[12]),
    .Z(net7));
 NAND3_X1 _3656_ (.A1(last_valid_data_available),
    .A2(\last_valid_data[0] ),
    .A3(net44),
    .ZN(_1512_));
 NAND2_X1 _3657_ (.A1(_1510_),
    .A2(_1512_),
    .ZN(net64));
 NAND2_X1 _3658_ (.A1(net96),
    .A2(_0932_),
    .ZN(_1513_));
 NAND3_X1 _3659_ (.A1(last_valid_data_available),
    .A2(\last_valid_data[10] ),
    .A3(net44),
    .ZN(_1514_));
 NAND2_X1 _3660_ (.A1(_1513_),
    .A2(_1514_),
    .ZN(net65));
 NAND2_X1 _3661_ (.A1(net173),
    .A2(_0950_),
    .ZN(_1515_));
 NAND3_X1 _3662_ (.A1(last_valid_data_available),
    .A2(\last_valid_data[11] ),
    .A3(net44),
    .ZN(_1516_));
 NAND2_X1 _3663_ (.A1(_1515_),
    .A2(_1516_),
    .ZN(net66));
 NAND2_X1 _3664_ (.A1(net96),
    .A2(_0968_),
    .ZN(_1517_));
 NAND3_X1 _3665_ (.A1(last_valid_data_available),
    .A2(\last_valid_data[12] ),
    .A3(net44),
    .ZN(_1518_));
 NAND2_X1 _3666_ (.A1(_1517_),
    .A2(_1518_),
    .ZN(net67));
 NAND2_X1 _3667_ (.A1(net173),
    .A2(_0986_),
    .ZN(_1519_));
 NAND3_X1 _3668_ (.A1(last_valid_data_available),
    .A2(\last_valid_data[13] ),
    .A3(net44),
    .ZN(_1520_));
 NAND2_X1 _3669_ (.A1(_1519_),
    .A2(_1520_),
    .ZN(net68));
 NAND2_X1 _3670_ (.A1(net173),
    .A2(_1005_),
    .ZN(_1521_));
 NAND3_X1 _3671_ (.A1(last_valid_data_available),
    .A2(\last_valid_data[14] ),
    .A3(net44),
    .ZN(_1522_));
 NAND2_X1 _3672_ (.A1(_1521_),
    .A2(_1522_),
    .ZN(net69));
 NAND2_X1 _3673_ (.A1(net173),
    .A2(_1024_),
    .ZN(_1523_));
 NAND3_X1 _3674_ (.A1(last_valid_data_available),
    .A2(\last_valid_data[15] ),
    .A3(net44),
    .ZN(_1524_));
 NAND2_X1 _3675_ (.A1(_1523_),
    .A2(_1524_),
    .ZN(net70));
 NAND2_X1 _3676_ (.A1(net96),
    .A2(_1044_),
    .ZN(_1525_));
 NAND3_X1 _3677_ (.A1(last_valid_data_available),
    .A2(\last_valid_data[16] ),
    .A3(net44),
    .ZN(_1526_));
 NAND2_X1 _3678_ (.A1(_1525_),
    .A2(_1526_),
    .ZN(net71));
 NAND2_X1 _3679_ (.A1(net173),
    .A2(_1063_),
    .ZN(_1527_));
 NAND3_X1 _3680_ (.A1(last_valid_data_available),
    .A2(\last_valid_data[17] ),
    .A3(net44),
    .ZN(_1528_));
 NAND2_X1 _3681_ (.A1(_1527_),
    .A2(_1528_),
    .ZN(net72));
 BUF_X1 input6 (.A(wr_data[11]),
    .Z(net6));
 NAND2_X1 _3683_ (.A1(net173),
    .A2(_1082_),
    .ZN(_1530_));
 BUF_X1 input5 (.A(wr_data[10]),
    .Z(net5));
 NAND3_X1 _3685_ (.A1(last_valid_data_available),
    .A2(\last_valid_data[18] ),
    .A3(net44),
    .ZN(_1532_));
 NAND2_X1 _3686_ (.A1(_1530_),
    .A2(_1532_),
    .ZN(net73));
 NAND2_X1 _3687_ (.A1(net96),
    .A2(_1102_),
    .ZN(_1533_));
 BUF_X1 input4 (.A(wr_data[0]),
    .Z(net4));
 NAND3_X1 _3689_ (.A1(net199),
    .A2(\last_valid_data[19] ),
    .A3(net172),
    .ZN(_1535_));
 NAND2_X1 _3690_ (.A1(_1533_),
    .A2(_1535_),
    .ZN(net74));
 NAND2_X1 _3691_ (.A1(net96),
    .A2(_1123_),
    .ZN(_1536_));
 NAND3_X1 _3692_ (.A1(net199),
    .A2(\last_valid_data[1] ),
    .A3(net172),
    .ZN(_1537_));
 NAND2_X1 _3693_ (.A1(_1536_),
    .A2(_1537_),
    .ZN(net75));
 NAND2_X1 _3694_ (.A1(net96),
    .A2(_1141_),
    .ZN(_1538_));
 NAND3_X1 _3695_ (.A1(net199),
    .A2(\last_valid_data[20] ),
    .A3(net172),
    .ZN(_1539_));
 NAND2_X1 _3696_ (.A1(_1538_),
    .A2(_1539_),
    .ZN(net76));
 NAND2_X1 _3697_ (.A1(net96),
    .A2(_1159_),
    .ZN(_1540_));
 NAND3_X1 _3698_ (.A1(net199),
    .A2(\last_valid_data[21] ),
    .A3(net172),
    .ZN(_1541_));
 NAND2_X1 _3699_ (.A1(_1540_),
    .A2(_1541_),
    .ZN(net77));
 NAND2_X1 _3700_ (.A1(net174),
    .A2(_1177_),
    .ZN(_1542_));
 NAND3_X1 _3701_ (.A1(net199),
    .A2(\last_valid_data[22] ),
    .A3(net172),
    .ZN(_1543_));
 NAND2_X1 _3702_ (.A1(_1542_),
    .A2(_1543_),
    .ZN(net78));
 NAND2_X1 _3703_ (.A1(net174),
    .A2(_1196_),
    .ZN(_1544_));
 NAND3_X1 _3704_ (.A1(net199),
    .A2(\last_valid_data[23] ),
    .A3(net172),
    .ZN(_1545_));
 NAND2_X1 _3705_ (.A1(_1544_),
    .A2(_1545_),
    .ZN(net79));
 NAND2_X1 _3706_ (.A1(net174),
    .A2(_1215_),
    .ZN(_1546_));
 NAND3_X1 _3707_ (.A1(net199),
    .A2(\last_valid_data[24] ),
    .A3(net172),
    .ZN(_1547_));
 NAND2_X1 _3708_ (.A1(_1546_),
    .A2(_1547_),
    .ZN(net80));
 NAND2_X1 _3709_ (.A1(net96),
    .A2(_1235_),
    .ZN(_1548_));
 NAND3_X1 _3710_ (.A1(net199),
    .A2(\last_valid_data[25] ),
    .A3(net172),
    .ZN(_1549_));
 NAND2_X1 _3711_ (.A1(_1548_),
    .A2(_1549_),
    .ZN(net81));
 NAND2_X1 _3712_ (.A1(net96),
    .A2(_1254_),
    .ZN(_1550_));
 NAND3_X1 _3713_ (.A1(net199),
    .A2(\last_valid_data[26] ),
    .A3(net172),
    .ZN(_1551_));
 NAND2_X1 _3714_ (.A1(_1550_),
    .A2(_1551_),
    .ZN(net82));
 BUF_X1 input3 (.A(rst_n),
    .Z(net3));
 NAND2_X1 _3716_ (.A1(net174),
    .A2(_1273_),
    .ZN(_1553_));
 BUF_X1 input2 (.A(rd_en),
    .Z(net2));
 NAND3_X1 _3718_ (.A1(net199),
    .A2(\last_valid_data[27] ),
    .A3(net172),
    .ZN(_1555_));
 NAND2_X1 _3719_ (.A1(_1553_),
    .A2(_1555_),
    .ZN(net83));
 NAND2_X1 _3720_ (.A1(net174),
    .A2(_1293_),
    .ZN(_1556_));
 BUF_X1 input1 (.A(clear_errors),
    .Z(net1));
 NAND3_X1 _3722_ (.A1(net199),
    .A2(\last_valid_data[28] ),
    .A3(net172),
    .ZN(_1558_));
 NAND2_X1 _3723_ (.A1(_1556_),
    .A2(_1558_),
    .ZN(net84));
 NAND2_X1 _3724_ (.A1(net174),
    .A2(_1314_),
    .ZN(_1559_));
 NAND3_X1 _3725_ (.A1(net199),
    .A2(\last_valid_data[29] ),
    .A3(net172),
    .ZN(_1560_));
 NAND2_X1 _3726_ (.A1(_1559_),
    .A2(_1560_),
    .ZN(net85));
 NAND2_X1 _3727_ (.A1(net174),
    .A2(_1332_),
    .ZN(_1561_));
 NAND3_X1 _3728_ (.A1(net199),
    .A2(\last_valid_data[2] ),
    .A3(net172),
    .ZN(_1562_));
 NAND2_X1 _3729_ (.A1(_1561_),
    .A2(_1562_),
    .ZN(net86));
 NAND2_X1 _3730_ (.A1(net174),
    .A2(_1349_),
    .ZN(_1563_));
 NAND3_X1 _3731_ (.A1(net199),
    .A2(\last_valid_data[30] ),
    .A3(net172),
    .ZN(_1564_));
 NAND2_X1 _3732_ (.A1(_1563_),
    .A2(_1564_),
    .ZN(net87));
 NAND2_X1 _3733_ (.A1(net174),
    .A2(_1366_),
    .ZN(_1565_));
 NAND3_X1 _3734_ (.A1(net199),
    .A2(\last_valid_data[31] ),
    .A3(net172),
    .ZN(_1566_));
 NAND2_X1 _3735_ (.A1(_1565_),
    .A2(_1566_),
    .ZN(net88));
 NAND2_X1 _3736_ (.A1(net174),
    .A2(_1383_),
    .ZN(_1567_));
 NAND3_X1 _3737_ (.A1(net199),
    .A2(\last_valid_data[3] ),
    .A3(net172),
    .ZN(_1568_));
 NAND2_X1 _3738_ (.A1(_1567_),
    .A2(_1568_),
    .ZN(net89));
 NAND2_X1 _3739_ (.A1(net174),
    .A2(_1400_),
    .ZN(_1569_));
 NAND3_X1 _3740_ (.A1(net199),
    .A2(\last_valid_data[4] ),
    .A3(net172),
    .ZN(_1570_));
 NAND2_X1 _3741_ (.A1(_1569_),
    .A2(_1570_),
    .ZN(net90));
 NAND2_X1 _3742_ (.A1(net173),
    .A2(_1417_),
    .ZN(_1571_));
 NAND3_X1 _3743_ (.A1(net199),
    .A2(\last_valid_data[5] ),
    .A3(net172),
    .ZN(_1572_));
 NAND2_X1 _3744_ (.A1(_1571_),
    .A2(_1572_),
    .ZN(net91));
 NAND2_X1 _3745_ (.A1(net173),
    .A2(_1434_),
    .ZN(_1573_));
 NAND3_X1 _3746_ (.A1(net199),
    .A2(\last_valid_data[6] ),
    .A3(net172),
    .ZN(_1574_));
 NAND2_X1 _3747_ (.A1(_1573_),
    .A2(_1574_),
    .ZN(net92));
 NAND2_X1 _3748_ (.A1(net173),
    .A2(_1451_),
    .ZN(_1575_));
 NAND3_X1 _3749_ (.A1(last_valid_data_available),
    .A2(\last_valid_data[7] ),
    .A3(net44),
    .ZN(_1576_));
 NAND2_X1 _3750_ (.A1(_1575_),
    .A2(_1576_),
    .ZN(net93));
 NAND2_X1 _3751_ (.A1(net173),
    .A2(_1468_),
    .ZN(_1577_));
 NAND3_X1 _3752_ (.A1(last_valid_data_available),
    .A2(\last_valid_data[8] ),
    .A3(net44),
    .ZN(_1578_));
 NAND2_X1 _3753_ (.A1(_1577_),
    .A2(_1578_),
    .ZN(net94));
 NAND2_X1 _3754_ (.A1(net173),
    .A2(_1485_),
    .ZN(_1579_));
 NAND3_X1 _3755_ (.A1(last_valid_data_available),
    .A2(\last_valid_data[9] ),
    .A3(net44),
    .ZN(_1580_));
 NAND2_X1 _3756_ (.A1(_1579_),
    .A2(_1580_),
    .ZN(net95));
 FA_X1 _3757_ (.A(_2150_),
    .B(\wr_ptr[1] ),
    .CI(_0006_),
    .CO(_0007_),
    .S(net40));
 HA_X1 _3758_ (.A(_2151_),
    .B(\wr_ptr[2] ),
    .CO(_0008_),
    .S(_0009_));
 HA_X1 _3759_ (.A(_2150_),
    .B(\wr_ptr[1] ),
    .CO(_0010_),
    .S(_0011_));
 HA_X1 _3760_ (.A(_2152_),
    .B(\wr_ptr[3] ),
    .CO(_0012_),
    .S(_0013_));
 HA_X1 _3761_ (.A(\rd_ptr[0] ),
    .B(\rd_ptr[1] ),
    .CO(_0014_),
    .S(_0015_));
 HA_X1 _3762_ (.A(net45),
    .B(net52),
    .CO(_0016_),
    .S(_0017_));
 HA_X1 _3763_ (.A(_0018_),
    .B(_2153_),
    .CO(_0019_),
    .S(_0020_));
 HA_X1 _3764_ (.A(_0018_),
    .B(\wr_ptr[1] ),
    .CO(_0021_),
    .S(_2154_));
 HA_X1 _3765_ (.A(\wr_ptr[0] ),
    .B(_2153_),
    .CO(_0022_),
    .S(_2155_));
 HA_X1 _3766_ (.A(\wr_ptr[0] ),
    .B(\wr_ptr[1] ),
    .CO(_0023_),
    .S(_2156_));
 HA_X1 _3767_ (.A(\rd_ptr[0] ),
    .B(_0018_),
    .CO(_0024_),
    .S(_0025_));
 DFF_X2 _3768_ (.D(_0026_),
    .CK(clknet_leaf_41_clk),
    .Q(_0000_),
    .QN(_2149_));
 DFF_X1 _3769_ (.D(_0027_),
    .CK(clknet_leaf_41_clk),
    .Q(_0001_),
    .QN(_2148_));
 DFF_X2 _3770_ (.D(_0028_),
    .CK(clknet_leaf_48_clk),
    .Q(_0002_),
    .QN(_2147_));
 DFF_X1 _3771_ (.D(_0029_),
    .CK(clknet_leaf_43_clk),
    .Q(_0003_),
    .QN(_2146_));
 DFF_X1 \error_count[0]$_SDFFE_PN0P_  (.D(_0030_),
    .CK(clknet_leaf_48_clk),
    .Q(net45),
    .QN(_0005_));
 DFF_X1 \error_count[10]$_SDFFE_PN0P_  (.D(_0031_),
    .CK(clknet_leaf_49_clk),
    .Q(net46),
    .QN(_2145_));
 DFF_X1 \error_count[11]$_SDFFE_PN0P_  (.D(_0032_),
    .CK(clknet_leaf_49_clk),
    .Q(net47),
    .QN(_2144_));
 DFF_X1 \error_count[12]$_SDFFE_PN0P_  (.D(_0033_),
    .CK(clknet_leaf_41_clk),
    .Q(net48),
    .QN(_2143_));
 DFF_X1 \error_count[13]$_SDFFE_PN0P_  (.D(_0034_),
    .CK(clknet_leaf_40_clk),
    .Q(net49),
    .QN(_2142_));
 DFF_X1 \error_count[14]$_SDFFE_PN0P_  (.D(_0035_),
    .CK(clknet_leaf_40_clk),
    .Q(net50),
    .QN(_2141_));
 DFF_X1 \error_count[15]$_SDFFE_PN0P_  (.D(_0036_),
    .CK(clknet_leaf_40_clk),
    .Q(net51),
    .QN(_2140_));
 DFF_X1 \error_count[1]$_SDFFE_PN0P_  (.D(_0037_),
    .CK(clknet_leaf_49_clk),
    .Q(net52),
    .QN(_2139_));
 DFF_X1 \error_count[2]$_SDFFE_PN0P_  (.D(_0038_),
    .CK(clknet_leaf_49_clk),
    .Q(net53),
    .QN(_2138_));
 DFF_X1 \error_count[3]$_SDFFE_PN0P_  (.D(_0039_),
    .CK(clknet_leaf_50_clk),
    .Q(net54),
    .QN(_2137_));
 DFF_X1 \error_count[4]$_SDFFE_PN0P_  (.D(_0040_),
    .CK(clknet_leaf_50_clk),
    .Q(net55),
    .QN(_2136_));
 DFF_X1 \error_count[5]$_SDFFE_PN0P_  (.D(_0041_),
    .CK(clknet_leaf_49_clk),
    .Q(net56),
    .QN(_2135_));
 DFF_X1 \error_count[6]$_SDFFE_PN0P_  (.D(_0042_),
    .CK(clknet_leaf_50_clk),
    .Q(net57),
    .QN(_2134_));
 DFF_X1 \error_count[7]$_SDFFE_PN0P_  (.D(_0043_),
    .CK(clknet_leaf_50_clk),
    .Q(net58),
    .QN(_2133_));
 DFF_X1 \error_count[8]$_SDFFE_PN0P_  (.D(_0044_),
    .CK(clknet_leaf_49_clk),
    .Q(net59),
    .QN(_2132_));
 DFF_X1 \error_count[9]$_SDFFE_PN0P_  (.D(_0045_),
    .CK(clknet_leaf_49_clk),
    .Q(net60),
    .QN(_2131_));
 DFF_X1 \error_detected$_SDFF_PN0_  (.D(_0046_),
    .CK(clknet_leaf_50_clk),
    .Q(net61),
    .QN(_2130_));
 DFF_X1 \last_valid_data[0]$_SDFFE_PN0P_  (.D(_0047_),
    .CK(clknet_leaf_63_clk),
    .Q(\last_valid_data[0] ),
    .QN(_2129_));
 DFF_X1 \last_valid_data[10]$_SDFFE_PN0P_  (.D(_0048_),
    .CK(clknet_leaf_48_clk),
    .Q(\last_valid_data[10] ),
    .QN(_2128_));
 DFF_X1 \last_valid_data[11]$_SDFFE_PN0P_  (.D(_0049_),
    .CK(clknet_leaf_63_clk),
    .Q(\last_valid_data[11] ),
    .QN(_2127_));
 DFF_X1 \last_valid_data[12]$_SDFFE_PN0P_  (.D(_0050_),
    .CK(clknet_leaf_48_clk),
    .Q(\last_valid_data[12] ),
    .QN(_2126_));
 DFF_X1 \last_valid_data[13]$_SDFFE_PN0P_  (.D(_0051_),
    .CK(clknet_leaf_65_clk),
    .Q(\last_valid_data[13] ),
    .QN(_2125_));
 DFF_X1 \last_valid_data[14]$_SDFFE_PN0P_  (.D(_0052_),
    .CK(clknet_leaf_62_clk),
    .Q(\last_valid_data[14] ),
    .QN(_2124_));
 DFF_X1 \last_valid_data[15]$_SDFFE_PN0P_  (.D(_0053_),
    .CK(clknet_leaf_47_clk),
    .Q(\last_valid_data[15] ),
    .QN(_2123_));
 DFF_X1 \last_valid_data[16]$_SDFFE_PN0P_  (.D(_0054_),
    .CK(clknet_leaf_48_clk),
    .Q(\last_valid_data[16] ),
    .QN(_2122_));
 DFF_X1 \last_valid_data[17]$_SDFFE_PN0P_  (.D(_0055_),
    .CK(clknet_leaf_45_clk),
    .Q(\last_valid_data[17] ),
    .QN(_2121_));
 DFF_X1 \last_valid_data[18]$_SDFFE_PN0P_  (.D(_0056_),
    .CK(clknet_leaf_45_clk),
    .Q(\last_valid_data[18] ),
    .QN(_2120_));
 DFF_X1 \last_valid_data[19]$_SDFFE_PN0P_  (.D(_0057_),
    .CK(clknet_leaf_43_clk),
    .Q(\last_valid_data[19] ),
    .QN(_2119_));
 DFF_X1 \last_valid_data[1]$_SDFFE_PN0P_  (.D(_0058_),
    .CK(clknet_leaf_43_clk),
    .Q(\last_valid_data[1] ),
    .QN(_2118_));
 DFF_X1 \last_valid_data[20]$_SDFFE_PN0P_  (.D(_0059_),
    .CK(clknet_leaf_43_clk),
    .Q(\last_valid_data[20] ),
    .QN(_2117_));
 DFF_X1 \last_valid_data[21]$_SDFFE_PN0P_  (.D(_0060_),
    .CK(clknet_leaf_46_clk),
    .Q(\last_valid_data[21] ),
    .QN(_2116_));
 DFF_X1 \last_valid_data[22]$_SDFFE_PN0P_  (.D(_0061_),
    .CK(clknet_leaf_44_clk),
    .Q(\last_valid_data[22] ),
    .QN(_2115_));
 DFF_X1 \last_valid_data[23]$_SDFFE_PN0P_  (.D(_0062_),
    .CK(clknet_leaf_27_clk),
    .Q(\last_valid_data[23] ),
    .QN(_2114_));
 DFF_X1 \last_valid_data[24]$_SDFFE_PN0P_  (.D(_0063_),
    .CK(clknet_leaf_27_clk),
    .Q(\last_valid_data[24] ),
    .QN(_2113_));
 DFF_X1 \last_valid_data[25]$_SDFFE_PN0P_  (.D(_0064_),
    .CK(clknet_leaf_43_clk),
    .Q(\last_valid_data[25] ),
    .QN(_2112_));
 DFF_X1 \last_valid_data[26]$_SDFFE_PN0P_  (.D(_0065_),
    .CK(clknet_leaf_43_clk),
    .Q(\last_valid_data[26] ),
    .QN(_2111_));
 DFF_X1 \last_valid_data[27]$_SDFFE_PN0P_  (.D(_0066_),
    .CK(clknet_leaf_27_clk),
    .Q(\last_valid_data[27] ),
    .QN(_2110_));
 DFF_X1 \last_valid_data[28]$_SDFFE_PN0P_  (.D(_0067_),
    .CK(clknet_leaf_6_clk),
    .Q(\last_valid_data[28] ),
    .QN(_2109_));
 DFF_X1 \last_valid_data[29]$_SDFFE_PN0P_  (.D(_0068_),
    .CK(clknet_leaf_7_clk),
    .Q(\last_valid_data[29] ),
    .QN(_2108_));
 DFF_X1 \last_valid_data[2]$_SDFFE_PN0P_  (.D(_0069_),
    .CK(clknet_leaf_7_clk),
    .Q(\last_valid_data[2] ),
    .QN(_2107_));
 DFF_X1 \last_valid_data[30]$_SDFFE_PN0P_  (.D(_0070_),
    .CK(clknet_leaf_8_clk),
    .Q(\last_valid_data[30] ),
    .QN(_2106_));
 DFF_X1 \last_valid_data[31]$_SDFFE_PN0P_  (.D(_0071_),
    .CK(clknet_leaf_7_clk),
    .Q(\last_valid_data[31] ),
    .QN(_2105_));
 DFF_X1 \last_valid_data[3]$_SDFFE_PN0P_  (.D(_0072_),
    .CK(clknet_leaf_7_clk),
    .Q(\last_valid_data[3] ),
    .QN(_2104_));
 DFF_X1 \last_valid_data[4]$_SDFFE_PN0P_  (.D(_0073_),
    .CK(clknet_leaf_7_clk),
    .Q(\last_valid_data[4] ),
    .QN(_2103_));
 DFF_X1 \last_valid_data[5]$_SDFFE_PN0P_  (.D(_0074_),
    .CK(clknet_leaf_5_clk),
    .Q(\last_valid_data[5] ),
    .QN(_2102_));
 DFF_X1 \last_valid_data[6]$_SDFFE_PN0P_  (.D(_0075_),
    .CK(clknet_leaf_5_clk),
    .Q(\last_valid_data[6] ),
    .QN(_2101_));
 DFF_X1 \last_valid_data[7]$_SDFFE_PN0P_  (.D(_0076_),
    .CK(clknet_leaf_65_clk),
    .Q(\last_valid_data[7] ),
    .QN(_2100_));
 DFF_X1 \last_valid_data[8]$_SDFFE_PN0P_  (.D(_0077_),
    .CK(clknet_leaf_64_clk),
    .Q(\last_valid_data[8] ),
    .QN(_2099_));
 DFF_X1 \last_valid_data[9]$_SDFFE_PN0P_  (.D(_0078_),
    .CK(clknet_leaf_64_clk),
    .Q(\last_valid_data[9] ),
    .QN(_2098_));
 DFF_X1 \last_valid_data_available$_SDFFE_PN0P_  (.D(_0079_),
    .CK(clknet_leaf_48_clk),
    .Q(last_valid_data_available),
    .QN(_2097_));
 DFF_X1 \mem[0][0]$_DFFE_PP_  (.D(_0080_),
    .CK(clknet_leaf_65_clk),
    .Q(\mem[0][0] ),
    .QN(_2096_));
 DFF_X1 \mem[0][10]$_DFFE_PP_  (.D(_0081_),
    .CK(clknet_leaf_55_clk),
    .Q(\mem[0][10] ),
    .QN(_2095_));
 DFF_X1 \mem[0][11]$_DFFE_PP_  (.D(_0082_),
    .CK(clknet_leaf_58_clk),
    .Q(\mem[0][11] ),
    .QN(_2094_));
 DFF_X1 \mem[0][12]$_DFFE_PP_  (.D(_0083_),
    .CK(clknet_leaf_54_clk),
    .Q(\mem[0][12] ),
    .QN(_2093_));
 DFF_X1 \mem[0][13]$_DFFE_PP_  (.D(_0084_),
    .CK(clknet_leaf_70_clk),
    .Q(\mem[0][13] ),
    .QN(_2092_));
 DFF_X1 \mem[0][14]$_DFFE_PP_  (.D(_0085_),
    .CK(clknet_leaf_57_clk),
    .Q(\mem[0][14] ),
    .QN(_2091_));
 DFF_X1 \mem[0][15]$_DFFE_PP_  (.D(_0086_),
    .CK(clknet_leaf_57_clk),
    .Q(\mem[0][15] ),
    .QN(_2090_));
 DFF_X1 \mem[0][16]$_DFFE_PP_  (.D(_0087_),
    .CK(clknet_leaf_47_clk),
    .Q(\mem[0][16] ),
    .QN(_2089_));
 DFF_X1 \mem[0][17]$_DFFE_PP_  (.D(_0088_),
    .CK(clknet_leaf_44_clk),
    .Q(\mem[0][17] ),
    .QN(_2088_));
 DFF_X1 \mem[0][18]$_DFFE_PP_  (.D(_0089_),
    .CK(clknet_leaf_62_clk),
    .Q(\mem[0][18] ),
    .QN(_2087_));
 DFF_X1 \mem[0][19]$_DFFE_PP_  (.D(_0090_),
    .CK(clknet_leaf_6_clk),
    .Q(\mem[0][19] ),
    .QN(_2086_));
 DFF_X1 \mem[0][1]$_DFFE_PP_  (.D(_0091_),
    .CK(clknet_leaf_29_clk),
    .Q(\mem[0][1] ),
    .QN(_2085_));
 DFF_X1 \mem[0][20]$_DFFE_PP_  (.D(_0092_),
    .CK(clknet_leaf_30_clk),
    .Q(\mem[0][20] ),
    .QN(_2084_));
 DFF_X1 \mem[0][21]$_DFFE_PP_  (.D(_0093_),
    .CK(clknet_leaf_34_clk),
    .Q(\mem[0][21] ),
    .QN(_2083_));
 DFF_X1 \mem[0][22]$_DFFE_PP_  (.D(_0094_),
    .CK(clknet_leaf_30_clk),
    .Q(\mem[0][22] ),
    .QN(_2082_));
 DFF_X1 \mem[0][23]$_DFFE_PP_  (.D(_0095_),
    .CK(clknet_leaf_23_clk),
    .Q(\mem[0][23] ),
    .QN(_2081_));
 DFF_X1 \mem[0][24]$_DFFE_PP_  (.D(_0096_),
    .CK(clknet_leaf_22_clk),
    .Q(\mem[0][24] ),
    .QN(_2080_));
 DFF_X1 \mem[0][25]$_DFFE_PP_  (.D(_0097_),
    .CK(clknet_leaf_26_clk),
    .Q(\mem[0][25] ),
    .QN(_2079_));
 DFF_X1 \mem[0][26]$_DFFE_PP_  (.D(_0098_),
    .CK(clknet_leaf_23_clk),
    .Q(\mem[0][26] ),
    .QN(_2078_));
 DFF_X1 \mem[0][27]$_DFFE_PP_  (.D(_0099_),
    .CK(clknet_leaf_23_clk),
    .Q(\mem[0][27] ),
    .QN(_2077_));
 DFF_X1 \mem[0][28]$_DFFE_PP_  (.D(_0100_),
    .CK(clknet_leaf_19_clk),
    .Q(\mem[0][28] ),
    .QN(_2076_));
 DFF_X1 \mem[0][29]$_DFFE_PP_  (.D(_0101_),
    .CK(clknet_leaf_18_clk),
    .Q(\mem[0][29] ),
    .QN(_2075_));
 DFF_X1 \mem[0][2]$_DFFE_PP_  (.D(_0102_),
    .CK(clknet_leaf_19_clk),
    .Q(\mem[0][2] ),
    .QN(_2074_));
 DFF_X1 \mem[0][30]$_DFFE_PP_  (.D(_0103_),
    .CK(clknet_leaf_14_clk),
    .Q(\mem[0][30] ),
    .QN(_2073_));
 DFF_X1 \mem[0][31]$_DFFE_PP_  (.D(_0104_),
    .CK(clknet_leaf_9_clk),
    .Q(\mem[0][31] ),
    .QN(_2072_));
 DFF_X1 \mem[0][3]$_DFFE_PP_  (.D(_0105_),
    .CK(clknet_leaf_9_clk),
    .Q(\mem[0][3] ),
    .QN(_2071_));
 DFF_X1 \mem[0][4]$_DFFE_PP_  (.D(_0106_),
    .CK(clknet_leaf_9_clk),
    .Q(\mem[0][4] ),
    .QN(_2070_));
 DFF_X1 \mem[0][5]$_DFFE_PP_  (.D(_0107_),
    .CK(clknet_leaf_4_clk),
    .Q(\mem[0][5] ),
    .QN(_2069_));
 DFF_X1 \mem[0][6]$_DFFE_PP_  (.D(_0108_),
    .CK(clknet_leaf_66_clk),
    .Q(\mem[0][6] ),
    .QN(_2068_));
 DFF_X1 \mem[0][7]$_DFFE_PP_  (.D(_0109_),
    .CK(clknet_leaf_71_clk),
    .Q(\mem[0][7] ),
    .QN(_2067_));
 DFF_X1 \mem[0][8]$_DFFE_PP_  (.D(_0110_),
    .CK(clknet_leaf_66_clk),
    .Q(\mem[0][8] ),
    .QN(_2066_));
 DFF_X1 \mem[0][9]$_DFFE_PP_  (.D(_0111_),
    .CK(clknet_leaf_71_clk),
    .Q(\mem[0][9] ),
    .QN(_2065_));
 DFF_X1 \mem[10][0]$_DFFE_PP_  (.D(_0112_),
    .CK(clknet_leaf_66_clk),
    .Q(\mem[10][0] ),
    .QN(_2064_));
 DFF_X1 \mem[10][10]$_DFFE_PP_  (.D(_0113_),
    .CK(clknet_leaf_51_clk),
    .Q(\mem[10][10] ),
    .QN(_2063_));
 DFF_X1 \mem[10][11]$_DFFE_PP_  (.D(_0114_),
    .CK(clknet_leaf_69_clk),
    .Q(\mem[10][11] ),
    .QN(_2062_));
 DFF_X1 \mem[10][12]$_DFFE_PP_  (.D(_0115_),
    .CK(clknet_leaf_55_clk),
    .Q(\mem[10][12] ),
    .QN(_2061_));
 DFF_X1 \mem[10][13]$_DFFE_PP_  (.D(_0116_),
    .CK(clknet_leaf_69_clk),
    .Q(\mem[10][13] ),
    .QN(_2060_));
 DFF_X1 \mem[10][14]$_DFFE_PP_  (.D(_0117_),
    .CK(clknet_leaf_60_clk),
    .Q(\mem[10][14] ),
    .QN(_2059_));
 DFF_X1 \mem[10][15]$_DFFE_PP_  (.D(_0118_),
    .CK(clknet_leaf_60_clk),
    .Q(\mem[10][15] ),
    .QN(_2058_));
 DFF_X1 \mem[10][16]$_DFFE_PP_  (.D(_0119_),
    .CK(clknet_leaf_51_clk),
    .Q(\mem[10][16] ),
    .QN(_2057_));
 DFF_X1 \mem[10][17]$_DFFE_PP_  (.D(_0120_),
    .CK(clknet_leaf_46_clk),
    .Q(\mem[10][17] ),
    .QN(_2056_));
 DFF_X1 \mem[10][18]$_DFFE_PP_  (.D(_0121_),
    .CK(clknet_leaf_62_clk),
    .Q(\mem[10][18] ),
    .QN(_2055_));
 DFF_X1 \mem[10][19]$_DFFE_PP_  (.D(_0122_),
    .CK(clknet_leaf_5_clk),
    .Q(\mem[10][19] ),
    .QN(_2054_));
 DFF_X1 \mem[10][1]$_DFFE_PP_  (.D(_0123_),
    .CK(clknet_leaf_39_clk),
    .Q(\mem[10][1] ),
    .QN(_2053_));
 DFF_X1 \mem[10][20]$_DFFE_PP_  (.D(_0124_),
    .CK(clknet_leaf_36_clk),
    .Q(\mem[10][20] ),
    .QN(_2052_));
 DFF_X1 \mem[10][21]$_DFFE_PP_  (.D(_0125_),
    .CK(clknet_leaf_37_clk),
    .Q(\mem[10][21] ),
    .QN(_2051_));
 DFF_X1 \mem[10][22]$_DFFE_PP_  (.D(_0126_),
    .CK(clknet_leaf_34_clk),
    .Q(\mem[10][22] ),
    .QN(_2050_));
 DFF_X1 \mem[10][23]$_DFFE_PP_  (.D(_0127_),
    .CK(clknet_leaf_21_clk),
    .Q(\mem[10][23] ),
    .QN(_2049_));
 DFF_X1 \mem[10][24]$_DFFE_PP_  (.D(_0128_),
    .CK(clknet_leaf_32_clk),
    .Q(\mem[10][24] ),
    .QN(_2048_));
 DFF_X1 \mem[10][25]$_DFFE_PP_  (.D(_0129_),
    .CK(clknet_leaf_28_clk),
    .Q(\mem[10][25] ),
    .QN(_2047_));
 DFF_X1 \mem[10][26]$_DFFE_PP_  (.D(_0130_),
    .CK(clknet_leaf_31_clk),
    .Q(\mem[10][26] ),
    .QN(_2046_));
 DFF_X1 \mem[10][27]$_DFFE_PP_  (.D(_0131_),
    .CK(clknet_leaf_8_clk),
    .Q(\mem[10][27] ),
    .QN(_2045_));
 DFF_X1 \mem[10][28]$_DFFE_PP_  (.D(_0132_),
    .CK(clknet_leaf_18_clk),
    .Q(\mem[10][28] ),
    .QN(_2044_));
 DFF_X1 \mem[10][29]$_DFFE_PP_  (.D(_0133_),
    .CK(clknet_leaf_17_clk),
    .Q(\mem[10][29] ),
    .QN(_2043_));
 DFF_X1 \mem[10][2]$_DFFE_PP_  (.D(_0134_),
    .CK(clknet_leaf_16_clk),
    .Q(\mem[10][2] ),
    .QN(_2042_));
 DFF_X1 \mem[10][30]$_DFFE_PP_  (.D(_0135_),
    .CK(clknet_leaf_13_clk),
    .Q(\mem[10][30] ),
    .QN(_2041_));
 DFF_X1 \mem[10][31]$_DFFE_PP_  (.D(_0136_),
    .CK(clknet_leaf_1_clk),
    .Q(\mem[10][31] ),
    .QN(_2040_));
 DFF_X1 \mem[10][3]$_DFFE_PP_  (.D(_0137_),
    .CK(clknet_leaf_12_clk),
    .Q(\mem[10][3] ),
    .QN(_2039_));
 DFF_X1 \mem[10][4]$_DFFE_PP_  (.D(_0138_),
    .CK(clknet_leaf_11_clk),
    .Q(\mem[10][4] ),
    .QN(_2038_));
 DFF_X1 \mem[10][5]$_DFFE_PP_  (.D(_0139_),
    .CK(clknet_leaf_1_clk),
    .Q(\mem[10][5] ),
    .QN(_2037_));
 DFF_X1 \mem[10][6]$_DFFE_PP_  (.D(_0140_),
    .CK(clknet_leaf_75_clk),
    .Q(\mem[10][6] ),
    .QN(_2036_));
 DFF_X1 \mem[10][7]$_DFFE_PP_  (.D(_0141_),
    .CK(clknet_leaf_73_clk),
    .Q(\mem[10][7] ),
    .QN(_2035_));
 DFF_X1 \mem[10][8]$_DFFE_PP_  (.D(_0142_),
    .CK(clknet_leaf_0_clk),
    .Q(\mem[10][8] ),
    .QN(_2034_));
 DFF_X1 \mem[10][9]$_DFFE_PP_  (.D(_0143_),
    .CK(clknet_leaf_73_clk),
    .Q(\mem[10][9] ),
    .QN(_2033_));
 DFF_X1 \mem[11][0]$_DFFE_PP_  (.D(_0144_),
    .CK(clknet_leaf_66_clk),
    .Q(\mem[11][0] ),
    .QN(_2032_));
 DFF_X1 \mem[11][10]$_DFFE_PP_  (.D(_0145_),
    .CK(clknet_leaf_52_clk),
    .Q(\mem[11][10] ),
    .QN(_2031_));
 DFF_X1 \mem[11][11]$_DFFE_PP_  (.D(_0146_),
    .CK(clknet_leaf_59_clk),
    .Q(\mem[11][11] ),
    .QN(_2030_));
 DFF_X1 \mem[11][12]$_DFFE_PP_  (.D(_0147_),
    .CK(clknet_leaf_52_clk),
    .Q(\mem[11][12] ),
    .QN(_2029_));
 DFF_X1 \mem[11][13]$_DFFE_PP_  (.D(_0148_),
    .CK(clknet_leaf_68_clk),
    .Q(\mem[11][13] ),
    .QN(_2028_));
 DFF_X1 \mem[11][14]$_DFFE_PP_  (.D(_0149_),
    .CK(clknet_leaf_59_clk),
    .Q(\mem[11][14] ),
    .QN(_2027_));
 DFF_X1 \mem[11][15]$_DFFE_PP_  (.D(_0150_),
    .CK(clknet_leaf_61_clk),
    .Q(\mem[11][15] ),
    .QN(_2026_));
 DFF_X1 \mem[11][16]$_DFFE_PP_  (.D(_0151_),
    .CK(clknet_leaf_50_clk),
    .Q(\mem[11][16] ),
    .QN(_2025_));
 DFF_X1 \mem[11][17]$_DFFE_PP_  (.D(_0152_),
    .CK(clknet_leaf_46_clk),
    .Q(\mem[11][17] ),
    .QN(_2024_));
 DFF_X1 \mem[11][18]$_DFFE_PP_  (.D(_0153_),
    .CK(clknet_leaf_61_clk),
    .Q(\mem[11][18] ),
    .QN(_2023_));
 DFF_X1 \mem[11][19]$_DFFE_PP_  (.D(_0154_),
    .CK(clknet_leaf_6_clk),
    .Q(\mem[11][19] ),
    .QN(_2022_));
 DFF_X1 \mem[11][1]$_DFFE_PP_  (.D(_0155_),
    .CK(clknet_leaf_38_clk),
    .Q(\mem[11][1] ),
    .QN(_2021_));
 DFF_X1 \mem[11][20]$_DFFE_PP_  (.D(_0156_),
    .CK(clknet_leaf_38_clk),
    .Q(\mem[11][20] ),
    .QN(_2020_));
 DFF_X1 \mem[11][21]$_DFFE_PP_  (.D(_0157_),
    .CK(clknet_leaf_37_clk),
    .Q(\mem[11][21] ),
    .QN(_2019_));
 DFF_X1 \mem[11][22]$_DFFE_PP_  (.D(_0158_),
    .CK(clknet_leaf_34_clk),
    .Q(\mem[11][22] ),
    .QN(_2018_));
 DFF_X1 \mem[11][23]$_DFFE_PP_  (.D(_0159_),
    .CK(clknet_leaf_22_clk),
    .Q(\mem[11][23] ),
    .QN(_2017_));
 DFF_X1 \mem[11][24]$_DFFE_PP_  (.D(_0160_),
    .CK(clknet_leaf_33_clk),
    .Q(\mem[11][24] ),
    .QN(_2016_));
 DFF_X1 \mem[11][25]$_DFFE_PP_  (.D(_0161_),
    .CK(clknet_leaf_28_clk),
    .Q(\mem[11][25] ),
    .QN(_2015_));
 DFF_X1 \mem[11][26]$_DFFE_PP_  (.D(_0162_),
    .CK(clknet_leaf_31_clk),
    .Q(\mem[11][26] ),
    .QN(_2014_));
 DFF_X1 \mem[11][27]$_DFFE_PP_  (.D(_0163_),
    .CK(clknet_leaf_8_clk),
    .Q(\mem[11][27] ),
    .QN(_2013_));
 DFF_X1 \mem[11][28]$_DFFE_PP_  (.D(_0164_),
    .CK(clknet_leaf_21_clk),
    .Q(\mem[11][28] ),
    .QN(_2012_));
 DFF_X1 \mem[11][29]$_DFFE_PP_  (.D(_0165_),
    .CK(clknet_leaf_17_clk),
    .Q(\mem[11][29] ),
    .QN(_2011_));
 DFF_X1 \mem[11][2]$_DFFE_PP_  (.D(_0166_),
    .CK(clknet_leaf_16_clk),
    .Q(\mem[11][2] ),
    .QN(_2010_));
 DFF_X1 \mem[11][30]$_DFFE_PP_  (.D(_0167_),
    .CK(clknet_leaf_13_clk),
    .Q(\mem[11][30] ),
    .QN(_2009_));
 DFF_X1 \mem[11][31]$_DFFE_PP_  (.D(_0168_),
    .CK(clknet_leaf_2_clk),
    .Q(\mem[11][31] ),
    .QN(_2008_));
 DFF_X1 \mem[11][3]$_DFFE_PP_  (.D(_0169_),
    .CK(clknet_leaf_11_clk),
    .Q(\mem[11][3] ),
    .QN(_2007_));
 DFF_X1 \mem[11][4]$_DFFE_PP_  (.D(_0170_),
    .CK(clknet_leaf_1_clk),
    .Q(\mem[11][4] ),
    .QN(_2006_));
 DFF_X1 \mem[11][5]$_DFFE_PP_  (.D(_0171_),
    .CK(clknet_leaf_0_clk),
    .Q(\mem[11][5] ),
    .QN(_2005_));
 DFF_X1 \mem[11][6]$_DFFE_PP_  (.D(_0172_),
    .CK(clknet_leaf_0_clk),
    .Q(\mem[11][6] ),
    .QN(_2004_));
 DFF_X1 \mem[11][7]$_DFFE_PP_  (.D(_0173_),
    .CK(clknet_leaf_73_clk),
    .Q(\mem[11][7] ),
    .QN(_2003_));
 DFF_X1 \mem[11][8]$_DFFE_PP_  (.D(_0174_),
    .CK(clknet_leaf_0_clk),
    .Q(\mem[11][8] ),
    .QN(_2002_));
 DFF_X1 \mem[11][9]$_DFFE_PP_  (.D(_0175_),
    .CK(clknet_leaf_73_clk),
    .Q(\mem[11][9] ),
    .QN(_2001_));
 DFF_X1 \mem[12][0]$_DFFE_PP_  (.D(_0176_),
    .CK(clknet_leaf_63_clk),
    .Q(\mem[12][0] ),
    .QN(_2000_));
 DFF_X1 \mem[12][10]$_DFFE_PP_  (.D(_0177_),
    .CK(clknet_leaf_53_clk),
    .Q(\mem[12][10] ),
    .QN(_1999_));
 DFF_X1 \mem[12][11]$_DFFE_PP_  (.D(_0178_),
    .CK(clknet_leaf_69_clk),
    .Q(\mem[12][11] ),
    .QN(_1998_));
 DFF_X1 \mem[12][12]$_DFFE_PP_  (.D(_0179_),
    .CK(clknet_leaf_53_clk),
    .Q(\mem[12][12] ),
    .QN(_1997_));
 DFF_X1 \mem[12][13]$_DFFE_PP_  (.D(_0180_),
    .CK(clknet_leaf_70_clk),
    .Q(\mem[12][13] ),
    .QN(_1996_));
 DFF_X1 \mem[12][14]$_DFFE_PP_  (.D(_0181_),
    .CK(clknet_leaf_58_clk),
    .Q(\mem[12][14] ),
    .QN(_1995_));
 DFF_X1 \mem[12][15]$_DFFE_PP_  (.D(_0182_),
    .CK(clknet_leaf_53_clk),
    .Q(\mem[12][15] ),
    .QN(_1994_));
 DFF_X1 \mem[12][16]$_DFFE_PP_  (.D(_0183_),
    .CK(clknet_leaf_50_clk),
    .Q(\mem[12][16] ),
    .QN(_1993_));
 DFF_X1 \mem[12][17]$_DFFE_PP_  (.D(_0184_),
    .CK(clknet_leaf_63_clk),
    .Q(\mem[12][17] ),
    .QN(_1992_));
 DFF_X1 \mem[12][18]$_DFFE_PP_  (.D(_0185_),
    .CK(clknet_leaf_61_clk),
    .Q(\mem[12][18] ),
    .QN(_1991_));
 DFF_X1 \mem[12][19]$_DFFE_PP_  (.D(_0186_),
    .CK(clknet_leaf_64_clk),
    .Q(\mem[12][19] ),
    .QN(_1990_));
 DFF_X1 \mem[12][1]$_DFFE_PP_  (.D(_0187_),
    .CK(clknet_leaf_39_clk),
    .Q(\mem[12][1] ),
    .QN(_1989_));
 DFF_X1 \mem[12][20]$_DFFE_PP_  (.D(_0188_),
    .CK(clknet_leaf_38_clk),
    .Q(\mem[12][20] ),
    .QN(_1988_));
 DFF_X1 \mem[12][21]$_DFFE_PP_  (.D(_0189_),
    .CK(clknet_leaf_36_clk),
    .Q(\mem[12][21] ),
    .QN(_1987_));
 DFF_X1 \mem[12][22]$_DFFE_PP_  (.D(_0190_),
    .CK(clknet_leaf_33_clk),
    .Q(\mem[12][22] ),
    .QN(_1986_));
 DFF_X1 \mem[12][23]$_DFFE_PP_  (.D(_0191_),
    .CK(clknet_leaf_21_clk),
    .Q(\mem[12][23] ),
    .QN(_1985_));
 DFF_X1 \mem[12][24]$_DFFE_PP_  (.D(_0192_),
    .CK(clknet_leaf_32_clk),
    .Q(\mem[12][24] ),
    .QN(_1984_));
 DFF_X1 \mem[12][25]$_DFFE_PP_  (.D(_0193_),
    .CK(clknet_leaf_43_clk),
    .Q(\mem[12][25] ),
    .QN(_1983_));
 DFF_X1 \mem[12][26]$_DFFE_PP_  (.D(_0194_),
    .CK(clknet_leaf_29_clk),
    .Q(\mem[12][26] ),
    .QN(_1982_));
 DFF_X1 \mem[12][27]$_DFFE_PP_  (.D(_0195_),
    .CK(clknet_leaf_25_clk),
    .Q(\mem[12][27] ),
    .QN(_1981_));
 DFF_X1 \mem[12][28]$_DFFE_PP_  (.D(_0196_),
    .CK(clknet_leaf_20_clk),
    .Q(\mem[12][28] ),
    .QN(_1980_));
 DFF_X1 \mem[12][29]$_DFFE_PP_  (.D(_0197_),
    .CK(clknet_leaf_17_clk),
    .Q(\mem[12][29] ),
    .QN(_1979_));
 DFF_X1 \mem[12][2]$_DFFE_PP_  (.D(_0198_),
    .CK(clknet_leaf_18_clk),
    .Q(\mem[12][2] ),
    .QN(_1978_));
 DFF_X1 \mem[12][30]$_DFFE_PP_  (.D(_0199_),
    .CK(clknet_leaf_14_clk),
    .Q(\mem[12][30] ),
    .QN(_1977_));
 DFF_X1 \mem[12][31]$_DFFE_PP_  (.D(_0200_),
    .CK(clknet_leaf_5_clk),
    .Q(\mem[12][31] ),
    .QN(_1976_));
 DFF_X1 \mem[12][3]$_DFFE_PP_  (.D(_0201_),
    .CK(clknet_leaf_10_clk),
    .Q(\mem[12][3] ),
    .QN(_1975_));
 DFF_X1 \mem[12][4]$_DFFE_PP_  (.D(_0202_),
    .CK(clknet_leaf_2_clk),
    .Q(\mem[12][4] ),
    .QN(_1974_));
 DFF_X1 \mem[12][5]$_DFFE_PP_  (.D(_0203_),
    .CK(clknet_leaf_4_clk),
    .Q(\mem[12][5] ),
    .QN(_1973_));
 DFF_X1 \mem[12][6]$_DFFE_PP_  (.D(_0204_),
    .CK(clknet_leaf_67_clk),
    .Q(\mem[12][6] ),
    .QN(_1972_));
 DFF_X1 \mem[12][7]$_DFFE_PP_  (.D(_0205_),
    .CK(clknet_leaf_74_clk),
    .Q(\mem[12][7] ),
    .QN(_1971_));
 DFF_X1 \mem[12][8]$_DFFE_PP_  (.D(_0206_),
    .CK(clknet_leaf_3_clk),
    .Q(\mem[12][8] ),
    .QN(_1970_));
 DFF_X1 \mem[12][9]$_DFFE_PP_  (.D(_0207_),
    .CK(clknet_leaf_71_clk),
    .Q(\mem[12][9] ),
    .QN(_1969_));
 DFF_X1 \mem[13][0]$_DFFE_PP_  (.D(_0208_),
    .CK(clknet_leaf_64_clk),
    .Q(\mem[13][0] ),
    .QN(_1968_));
 DFF_X1 \mem[13][10]$_DFFE_PP_  (.D(_0209_),
    .CK(clknet_leaf_52_clk),
    .Q(\mem[13][10] ),
    .QN(_1967_));
 DFF_X1 \mem[13][11]$_DFFE_PP_  (.D(_0210_),
    .CK(clknet_leaf_58_clk),
    .Q(\mem[13][11] ),
    .QN(_1966_));
 DFF_X1 \mem[13][12]$_DFFE_PP_  (.D(_0211_),
    .CK(clknet_leaf_53_clk),
    .Q(\mem[13][12] ),
    .QN(_1965_));
 DFF_X1 \mem[13][13]$_DFFE_PP_  (.D(_0212_),
    .CK(clknet_leaf_69_clk),
    .Q(\mem[13][13] ),
    .QN(_1964_));
 DFF_X1 \mem[13][14]$_DFFE_PP_  (.D(_0213_),
    .CK(clknet_leaf_57_clk),
    .Q(\mem[13][14] ),
    .QN(_1963_));
 DFF_X1 \mem[13][15]$_DFFE_PP_  (.D(_0214_),
    .CK(clknet_leaf_58_clk),
    .Q(\mem[13][15] ),
    .QN(_1962_));
 DFF_X1 \mem[13][16]$_DFFE_PP_  (.D(_0215_),
    .CK(clknet_leaf_52_clk),
    .Q(\mem[13][16] ),
    .QN(_1961_));
 DFF_X1 \mem[13][17]$_DFFE_PP_  (.D(_0216_),
    .CK(clknet_leaf_45_clk),
    .Q(\mem[13][17] ),
    .QN(_1960_));
 DFF_X1 \mem[13][18]$_DFFE_PP_  (.D(_0217_),
    .CK(clknet_leaf_61_clk),
    .Q(\mem[13][18] ),
    .QN(_1959_));
 DFF_X1 \mem[13][19]$_DFFE_PP_  (.D(_0218_),
    .CK(clknet_leaf_45_clk),
    .Q(\mem[13][19] ),
    .QN(_1958_));
 DFF_X1 \mem[13][1]$_DFFE_PP_  (.D(_0219_),
    .CK(clknet_leaf_39_clk),
    .Q(\mem[13][1] ),
    .QN(_1957_));
 DFF_X1 \mem[13][20]$_DFFE_PP_  (.D(_0220_),
    .CK(clknet_leaf_38_clk),
    .Q(\mem[13][20] ),
    .QN(_1956_));
 DFF_X1 \mem[13][21]$_DFFE_PP_  (.D(_0221_),
    .CK(clknet_leaf_34_clk),
    .Q(\mem[13][21] ),
    .QN(_1955_));
 DFF_X1 \mem[13][22]$_DFFE_PP_  (.D(_0222_),
    .CK(clknet_leaf_33_clk),
    .Q(\mem[13][22] ),
    .QN(_1954_));
 DFF_X1 \mem[13][23]$_DFFE_PP_  (.D(_0223_),
    .CK(clknet_leaf_22_clk),
    .Q(\mem[13][23] ),
    .QN(_1953_));
 DFF_X1 \mem[13][24]$_DFFE_PP_  (.D(_0224_),
    .CK(clknet_leaf_32_clk),
    .Q(\mem[13][24] ),
    .QN(_1952_));
 DFF_X1 \mem[13][25]$_DFFE_PP_  (.D(_0225_),
    .CK(clknet_leaf_29_clk),
    .Q(\mem[13][25] ),
    .QN(_1951_));
 DFF_X1 \mem[13][26]$_DFFE_PP_  (.D(_0226_),
    .CK(clknet_leaf_30_clk),
    .Q(\mem[13][26] ),
    .QN(_1950_));
 DFF_X1 \mem[13][27]$_DFFE_PP_  (.D(_0227_),
    .CK(clknet_leaf_24_clk),
    .Q(\mem[13][27] ),
    .QN(_1949_));
 DFF_X1 \mem[13][28]$_DFFE_PP_  (.D(_0228_),
    .CK(clknet_leaf_21_clk),
    .Q(\mem[13][28] ),
    .QN(_1948_));
 DFF_X1 \mem[13][29]$_DFFE_PP_  (.D(_0229_),
    .CK(clknet_leaf_17_clk),
    .Q(\mem[13][29] ),
    .QN(_1947_));
 DFF_X1 \mem[13][2]$_DFFE_PP_  (.D(_0230_),
    .CK(clknet_leaf_15_clk),
    .Q(\mem[13][2] ),
    .QN(_1946_));
 DFF_X1 \mem[13][30]$_DFFE_PP_  (.D(_0231_),
    .CK(clknet_leaf_15_clk),
    .Q(\mem[13][30] ),
    .QN(_1945_));
 DFF_X1 \mem[13][31]$_DFFE_PP_  (.D(_0232_),
    .CK(clknet_leaf_4_clk),
    .Q(\mem[13][31] ),
    .QN(_1944_));
 DFF_X1 \mem[13][3]$_DFFE_PP_  (.D(_0233_),
    .CK(clknet_leaf_10_clk),
    .Q(\mem[13][3] ),
    .QN(_1943_));
 DFF_X1 \mem[13][4]$_DFFE_PP_  (.D(_0234_),
    .CK(clknet_leaf_2_clk),
    .Q(\mem[13][4] ),
    .QN(_1942_));
 DFF_X1 \mem[13][5]$_DFFE_PP_  (.D(_0235_),
    .CK(clknet_leaf_2_clk),
    .Q(\mem[13][5] ),
    .QN(_1941_));
 DFF_X1 \mem[13][6]$_DFFE_PP_  (.D(_0236_),
    .CK(clknet_leaf_72_clk),
    .Q(\mem[13][6] ),
    .QN(_1940_));
 DFF_X1 \mem[13][7]$_DFFE_PP_  (.D(_0237_),
    .CK(clknet_leaf_71_clk),
    .Q(\mem[13][7] ),
    .QN(_1939_));
 DFF_X1 \mem[13][8]$_DFFE_PP_  (.D(_0238_),
    .CK(clknet_leaf_3_clk),
    .Q(\mem[13][8] ),
    .QN(_1938_));
 DFF_X1 \mem[13][9]$_DFFE_PP_  (.D(_0239_),
    .CK(clknet_leaf_70_clk),
    .Q(\mem[13][9] ),
    .QN(_1937_));
 DFF_X1 \mem[14][0]$_DFFE_PP_  (.D(_0240_),
    .CK(clknet_leaf_65_clk),
    .Q(\mem[14][0] ),
    .QN(_1936_));
 DFF_X1 \mem[14][10]$_DFFE_PP_  (.D(_0241_),
    .CK(clknet_leaf_51_clk),
    .Q(\mem[14][10] ),
    .QN(_1935_));
 DFF_X1 \mem[14][11]$_DFFE_PP_  (.D(_0242_),
    .CK(clknet_leaf_69_clk),
    .Q(\mem[14][11] ),
    .QN(_1934_));
 DFF_X1 \mem[14][12]$_DFFE_PP_  (.D(_0243_),
    .CK(clknet_leaf_53_clk),
    .Q(\mem[14][12] ),
    .QN(_1933_));
 DFF_X1 \mem[14][13]$_DFFE_PP_  (.D(_0244_),
    .CK(clknet_leaf_67_clk),
    .Q(\mem[14][13] ),
    .QN(_1932_));
 DFF_X1 \mem[14][14]$_DFFE_PP_  (.D(_0245_),
    .CK(clknet_leaf_60_clk),
    .Q(\mem[14][14] ),
    .QN(_1931_));
 DFF_X1 \mem[14][15]$_DFFE_PP_  (.D(_0246_),
    .CK(clknet_leaf_60_clk),
    .Q(\mem[14][15] ),
    .QN(_1930_));
 DFF_X1 \mem[14][16]$_DFFE_PP_  (.D(_0247_),
    .CK(clknet_leaf_48_clk),
    .Q(\mem[14][16] ),
    .QN(_1929_));
 DFF_X1 \mem[14][17]$_DFFE_PP_  (.D(_0248_),
    .CK(clknet_leaf_46_clk),
    .Q(\mem[14][17] ),
    .QN(_1928_));
 DFF_X1 \mem[14][18]$_DFFE_PP_  (.D(_0249_),
    .CK(clknet_leaf_62_clk),
    .Q(\mem[14][18] ),
    .QN(_1927_));
 DFF_X1 \mem[14][19]$_DFFE_PP_  (.D(_0250_),
    .CK(clknet_leaf_5_clk),
    .Q(\mem[14][19] ),
    .QN(_1926_));
 DFF_X1 \mem[14][1]$_DFFE_PP_  (.D(_0251_),
    .CK(clknet_leaf_39_clk),
    .Q(\mem[14][1] ),
    .QN(_1925_));
 DFF_X1 \mem[14][20]$_DFFE_PP_  (.D(_0252_),
    .CK(clknet_leaf_36_clk),
    .Q(\mem[14][20] ),
    .QN(_1924_));
 DFF_X1 \mem[14][21]$_DFFE_PP_  (.D(_0253_),
    .CK(clknet_leaf_36_clk),
    .Q(\mem[14][21] ),
    .QN(_1923_));
 DFF_X1 \mem[14][22]$_DFFE_PP_  (.D(_0254_),
    .CK(clknet_leaf_33_clk),
    .Q(\mem[14][22] ),
    .QN(_1922_));
 DFF_X1 \mem[14][23]$_DFFE_PP_  (.D(_0255_),
    .CK(clknet_leaf_21_clk),
    .Q(\mem[14][23] ),
    .QN(_1921_));
 DFF_X1 \mem[14][24]$_DFFE_PP_  (.D(_0256_),
    .CK(clknet_leaf_32_clk),
    .Q(\mem[14][24] ),
    .QN(_1920_));
 DFF_X1 \mem[14][25]$_DFFE_PP_  (.D(_0257_),
    .CK(clknet_leaf_44_clk),
    .Q(\mem[14][25] ),
    .QN(_1919_));
 DFF_X1 \mem[14][26]$_DFFE_PP_  (.D(_0258_),
    .CK(clknet_leaf_31_clk),
    .Q(\mem[14][26] ),
    .QN(_1918_));
 DFF_X1 \mem[14][27]$_DFFE_PP_  (.D(_0259_),
    .CK(clknet_leaf_8_clk),
    .Q(\mem[14][27] ),
    .QN(_1917_));
 DFF_X1 \mem[14][28]$_DFFE_PP_  (.D(_0260_),
    .CK(clknet_leaf_20_clk),
    .Q(\mem[14][28] ),
    .QN(_1916_));
 DFF_X1 \mem[14][29]$_DFFE_PP_  (.D(_0261_),
    .CK(clknet_leaf_17_clk),
    .Q(\mem[14][29] ),
    .QN(_1915_));
 DFF_X1 \mem[14][2]$_DFFE_PP_  (.D(_0262_),
    .CK(clknet_leaf_16_clk),
    .Q(\mem[14][2] ),
    .QN(_1914_));
 DFF_X1 \mem[14][30]$_DFFE_PP_  (.D(_0263_),
    .CK(clknet_leaf_16_clk),
    .Q(\mem[14][30] ),
    .QN(_1913_));
 DFF_X1 \mem[14][31]$_DFFE_PP_  (.D(_0264_),
    .CK(clknet_leaf_1_clk),
    .Q(\mem[14][31] ),
    .QN(_1912_));
 DFF_X1 \mem[14][3]$_DFFE_PP_  (.D(_0265_),
    .CK(clknet_leaf_12_clk),
    .Q(\mem[14][3] ),
    .QN(_1911_));
 DFF_X1 \mem[14][4]$_DFFE_PP_  (.D(_0266_),
    .CK(clknet_leaf_2_clk),
    .Q(\mem[14][4] ),
    .QN(_1910_));
 DFF_X1 \mem[14][5]$_DFFE_PP_  (.D(_0267_),
    .CK(clknet_leaf_1_clk),
    .Q(\mem[14][5] ),
    .QN(_1909_));
 DFF_X1 \mem[14][6]$_DFFE_PP_  (.D(_0268_),
    .CK(clknet_leaf_75_clk),
    .Q(\mem[14][6] ),
    .QN(_1908_));
 DFF_X1 \mem[14][7]$_DFFE_PP_  (.D(_0269_),
    .CK(clknet_leaf_73_clk),
    .Q(\mem[14][7] ),
    .QN(_1907_));
 DFF_X1 \mem[14][8]$_DFFE_PP_  (.D(_0270_),
    .CK(clknet_leaf_0_clk),
    .Q(\mem[14][8] ),
    .QN(_1906_));
 DFF_X1 \mem[14][9]$_DFFE_PP_  (.D(_0271_),
    .CK(clknet_leaf_73_clk),
    .Q(\mem[14][9] ),
    .QN(_1905_));
 DFF_X1 \mem[15][0]$_DFFE_PP_  (.D(_0272_),
    .CK(clknet_leaf_65_clk),
    .Q(\mem[15][0] ),
    .QN(_1904_));
 DFF_X1 \mem[15][10]$_DFFE_PP_  (.D(_0273_),
    .CK(clknet_leaf_52_clk),
    .Q(\mem[15][10] ),
    .QN(_1903_));
 DFF_X1 \mem[15][11]$_DFFE_PP_  (.D(_0274_),
    .CK(clknet_leaf_59_clk),
    .Q(\mem[15][11] ),
    .QN(_1902_));
 DFF_X1 \mem[15][12]$_DFFE_PP_  (.D(_0275_),
    .CK(clknet_leaf_55_clk),
    .Q(\mem[15][12] ),
    .QN(_1901_));
 DFF_X1 \mem[15][13]$_DFFE_PP_  (.D(_0276_),
    .CK(clknet_leaf_68_clk),
    .Q(\mem[15][13] ),
    .QN(_1900_));
 DFF_X1 \mem[15][14]$_DFFE_PP_  (.D(_0277_),
    .CK(clknet_leaf_59_clk),
    .Q(\mem[15][14] ),
    .QN(_1899_));
 DFF_X1 \mem[15][15]$_DFFE_PP_  (.D(_0278_),
    .CK(clknet_leaf_60_clk),
    .Q(\mem[15][15] ),
    .QN(_1898_));
 DFF_X1 \mem[15][16]$_DFFE_PP_  (.D(_0279_),
    .CK(clknet_leaf_50_clk),
    .Q(\mem[15][16] ),
    .QN(_1897_));
 DFF_X1 \mem[15][17]$_DFFE_PP_  (.D(_0280_),
    .CK(clknet_leaf_46_clk),
    .Q(\mem[15][17] ),
    .QN(_1896_));
 DFF_X1 \mem[15][18]$_DFFE_PP_  (.D(_0281_),
    .CK(clknet_leaf_62_clk),
    .Q(\mem[15][18] ),
    .QN(_1895_));
 DFF_X1 \mem[15][19]$_DFFE_PP_  (.D(_0282_),
    .CK(clknet_leaf_6_clk),
    .Q(\mem[15][19] ),
    .QN(_1894_));
 DFF_X1 \mem[15][1]$_DFFE_PP_  (.D(_0283_),
    .CK(clknet_leaf_39_clk),
    .Q(\mem[15][1] ),
    .QN(_1893_));
 DFF_X1 \mem[15][20]$_DFFE_PP_  (.D(_0284_),
    .CK(clknet_leaf_37_clk),
    .Q(\mem[15][20] ),
    .QN(_1892_));
 DFF_X1 \mem[15][21]$_DFFE_PP_  (.D(_0285_),
    .CK(clknet_leaf_37_clk),
    .Q(\mem[15][21] ),
    .QN(_1891_));
 DFF_X1 \mem[15][22]$_DFFE_PP_  (.D(_0286_),
    .CK(clknet_leaf_34_clk),
    .Q(\mem[15][22] ),
    .QN(_1890_));
 DFF_X1 \mem[15][23]$_DFFE_PP_  (.D(_0287_),
    .CK(clknet_leaf_22_clk),
    .Q(\mem[15][23] ),
    .QN(_1889_));
 DFF_X1 \mem[15][24]$_DFFE_PP_  (.D(_0288_),
    .CK(clknet_leaf_33_clk),
    .Q(\mem[15][24] ),
    .QN(_1888_));
 DFF_X1 \mem[15][25]$_DFFE_PP_  (.D(_0289_),
    .CK(clknet_leaf_29_clk),
    .Q(\mem[15][25] ),
    .QN(_1887_));
 DFF_X1 \mem[15][26]$_DFFE_PP_  (.D(_0290_),
    .CK(clknet_leaf_31_clk),
    .Q(\mem[15][26] ),
    .QN(_1886_));
 DFF_X1 \mem[15][27]$_DFFE_PP_  (.D(_0291_),
    .CK(clknet_leaf_25_clk),
    .Q(\mem[15][27] ),
    .QN(_1885_));
 DFF_X1 \mem[15][28]$_DFFE_PP_  (.D(_0292_),
    .CK(clknet_leaf_20_clk),
    .Q(\mem[15][28] ),
    .QN(_1884_));
 DFF_X1 \mem[15][29]$_DFFE_PP_  (.D(_0293_),
    .CK(clknet_leaf_17_clk),
    .Q(\mem[15][29] ),
    .QN(_1883_));
 DFF_X1 \mem[15][2]$_DFFE_PP_  (.D(_0294_),
    .CK(clknet_leaf_16_clk),
    .Q(\mem[15][2] ),
    .QN(_1882_));
 DFF_X1 \mem[15][30]$_DFFE_PP_  (.D(_0295_),
    .CK(clknet_leaf_13_clk),
    .Q(\mem[15][30] ),
    .QN(_1881_));
 DFF_X1 \mem[15][31]$_DFFE_PP_  (.D(_0296_),
    .CK(clknet_leaf_2_clk),
    .Q(\mem[15][31] ),
    .QN(_1880_));
 DFF_X1 \mem[15][3]$_DFFE_PP_  (.D(_0297_),
    .CK(clknet_leaf_12_clk),
    .Q(\mem[15][3] ),
    .QN(_1879_));
 DFF_X1 \mem[15][4]$_DFFE_PP_  (.D(_0298_),
    .CK(clknet_leaf_1_clk),
    .Q(\mem[15][4] ),
    .QN(_1878_));
 DFF_X1 \mem[15][5]$_DFFE_PP_  (.D(_0299_),
    .CK(clknet_leaf_1_clk),
    .Q(\mem[15][5] ),
    .QN(_1877_));
 DFF_X1 \mem[15][6]$_DFFE_PP_  (.D(_0300_),
    .CK(clknet_leaf_0_clk),
    .Q(\mem[15][6] ),
    .QN(_1876_));
 DFF_X1 \mem[15][7]$_DFFE_PP_  (.D(_0301_),
    .CK(clknet_leaf_75_clk),
    .Q(\mem[15][7] ),
    .QN(_1875_));
 DFF_X1 \mem[15][8]$_DFFE_PP_  (.D(_0302_),
    .CK(clknet_leaf_0_clk),
    .Q(\mem[15][8] ),
    .QN(_1874_));
 DFF_X1 \mem[15][9]$_DFFE_PP_  (.D(_0303_),
    .CK(clknet_leaf_73_clk),
    .Q(\mem[15][9] ),
    .QN(_1873_));
 DFF_X1 \mem[1][0]$_DFFE_PP_  (.D(_0304_),
    .CK(clknet_leaf_64_clk),
    .Q(\mem[1][0] ),
    .QN(_1872_));
 DFF_X1 \mem[1][10]$_DFFE_PP_  (.D(_0305_),
    .CK(clknet_leaf_54_clk),
    .Q(\mem[1][10] ),
    .QN(_1871_));
 DFF_X1 \mem[1][11]$_DFFE_PP_  (.D(_0306_),
    .CK(clknet_leaf_69_clk),
    .Q(\mem[1][11] ),
    .QN(_1870_));
 DFF_X1 \mem[1][12]$_DFFE_PP_  (.D(_0307_),
    .CK(clknet_leaf_54_clk),
    .Q(\mem[1][12] ),
    .QN(_1869_));
 DFF_X1 \mem[1][13]$_DFFE_PP_  (.D(_0308_),
    .CK(clknet_leaf_70_clk),
    .Q(\mem[1][13] ),
    .QN(_1868_));
 DFF_X1 \mem[1][14]$_DFFE_PP_  (.D(_0309_),
    .CK(clknet_leaf_57_clk),
    .Q(\mem[1][14] ),
    .QN(_1867_));
 DFF_X1 \mem[1][15]$_DFFE_PP_  (.D(_0310_),
    .CK(clknet_leaf_56_clk),
    .Q(\mem[1][15] ),
    .QN(_1866_));
 DFF_X1 \mem[1][16]$_DFFE_PP_  (.D(_0311_),
    .CK(clknet_leaf_51_clk),
    .Q(\mem[1][16] ),
    .QN(_1865_));
 DFF_X1 \mem[1][17]$_DFFE_PP_  (.D(_0312_),
    .CK(clknet_leaf_45_clk),
    .Q(\mem[1][17] ),
    .QN(_1864_));
 DFF_X1 \mem[1][18]$_DFFE_PP_  (.D(_0313_),
    .CK(clknet_leaf_46_clk),
    .Q(\mem[1][18] ),
    .QN(_1863_));
 DFF_X1 \mem[1][19]$_DFFE_PP_  (.D(_0314_),
    .CK(clknet_leaf_27_clk),
    .Q(\mem[1][19] ),
    .QN(_1862_));
 DFF_X1 \mem[1][1]$_DFFE_PP_  (.D(_0315_),
    .CK(clknet_leaf_42_clk),
    .Q(\mem[1][1] ),
    .QN(_1861_));
 DFF_X1 \mem[1][20]$_DFFE_PP_  (.D(_0316_),
    .CK(clknet_leaf_30_clk),
    .Q(\mem[1][20] ),
    .QN(_1860_));
 DFF_X1 \mem[1][21]$_DFFE_PP_  (.D(_0317_),
    .CK(clknet_leaf_36_clk),
    .Q(\mem[1][21] ),
    .QN(_1859_));
 DFF_X1 \mem[1][22]$_DFFE_PP_  (.D(_0318_),
    .CK(clknet_leaf_34_clk),
    .Q(\mem[1][22] ),
    .QN(_1858_));
 DFF_X1 \mem[1][23]$_DFFE_PP_  (.D(_0319_),
    .CK(clknet_leaf_20_clk),
    .Q(\mem[1][23] ),
    .QN(_1857_));
 DFF_X1 \mem[1][24]$_DFFE_PP_  (.D(_0320_),
    .CK(clknet_leaf_32_clk),
    .Q(\mem[1][24] ),
    .QN(_1856_));
 DFF_X1 \mem[1][25]$_DFFE_PP_  (.D(_0321_),
    .CK(clknet_leaf_26_clk),
    .Q(\mem[1][25] ),
    .QN(_1855_));
 DFF_X1 \mem[1][26]$_DFFE_PP_  (.D(_0322_),
    .CK(clknet_leaf_28_clk),
    .Q(\mem[1][26] ),
    .QN(_1854_));
 DFF_X1 \mem[1][27]$_DFFE_PP_  (.D(_0323_),
    .CK(clknet_leaf_24_clk),
    .Q(\mem[1][27] ),
    .QN(_1853_));
 DFF_X1 \mem[1][28]$_DFFE_PP_  (.D(_0324_),
    .CK(clknet_leaf_20_clk),
    .Q(\mem[1][28] ),
    .QN(_1852_));
 DFF_X1 \mem[1][29]$_DFFE_PP_  (.D(_0325_),
    .CK(clknet_leaf_18_clk),
    .Q(\mem[1][29] ),
    .QN(_1851_));
 DFF_X1 \mem[1][2]$_DFFE_PP_  (.D(_0326_),
    .CK(clknet_leaf_15_clk),
    .Q(\mem[1][2] ),
    .QN(_1850_));
 DFF_X1 \mem[1][30]$_DFFE_PP_  (.D(_0327_),
    .CK(clknet_leaf_14_clk),
    .Q(\mem[1][30] ),
    .QN(_1849_));
 DFF_X1 \mem[1][31]$_DFFE_PP_  (.D(_0328_),
    .CK(clknet_leaf_10_clk),
    .Q(\mem[1][31] ),
    .QN(_1848_));
 DFF_X1 \mem[1][3]$_DFFE_PP_  (.D(_0329_),
    .CK(clknet_leaf_9_clk),
    .Q(\mem[1][3] ),
    .QN(_1847_));
 DFF_X1 \mem[1][4]$_DFFE_PP_  (.D(_0330_),
    .CK(clknet_leaf_10_clk),
    .Q(\mem[1][4] ),
    .QN(_1846_));
 DFF_X1 \mem[1][5]$_DFFE_PP_  (.D(_0331_),
    .CK(clknet_leaf_4_clk),
    .Q(\mem[1][5] ),
    .QN(_1845_));
 DFF_X1 \mem[1][6]$_DFFE_PP_  (.D(_0332_),
    .CK(clknet_leaf_67_clk),
    .Q(\mem[1][6] ),
    .QN(_1844_));
 DFF_X1 \mem[1][7]$_DFFE_PP_  (.D(_0333_),
    .CK(clknet_leaf_73_clk),
    .Q(\mem[1][7] ),
    .QN(_1843_));
 DFF_X1 \mem[1][8]$_DFFE_PP_  (.D(_0334_),
    .CK(clknet_leaf_4_clk),
    .Q(\mem[1][8] ),
    .QN(_1842_));
 DFF_X1 \mem[1][9]$_DFFE_PP_  (.D(_0335_),
    .CK(clknet_leaf_72_clk),
    .Q(\mem[1][9] ),
    .QN(_1841_));
 DFF_X1 \mem[2][0]$_DFFE_PP_  (.D(_0336_),
    .CK(clknet_leaf_68_clk),
    .Q(\mem[2][0] ),
    .QN(_1840_));
 DFF_X1 \mem[2][10]$_DFFE_PP_  (.D(_0337_),
    .CK(clknet_leaf_56_clk),
    .Q(\mem[2][10] ),
    .QN(_1839_));
 DFF_X1 \mem[2][11]$_DFFE_PP_  (.D(_0338_),
    .CK(clknet_leaf_68_clk),
    .Q(\mem[2][11] ),
    .QN(_1838_));
 DFF_X1 \mem[2][12]$_DFFE_PP_  (.D(_0339_),
    .CK(clknet_leaf_55_clk),
    .Q(\mem[2][12] ),
    .QN(_1837_));
 DFF_X1 \mem[2][13]$_DFFE_PP_  (.D(_0340_),
    .CK(clknet_leaf_67_clk),
    .Q(\mem[2][13] ),
    .QN(_1836_));
 DFF_X1 \mem[2][14]$_DFFE_PP_  (.D(_0341_),
    .CK(clknet_leaf_61_clk),
    .Q(\mem[2][14] ),
    .QN(_1835_));
 DFF_X1 \mem[2][15]$_DFFE_PP_  (.D(_0342_),
    .CK(clknet_leaf_61_clk),
    .Q(\mem[2][15] ),
    .QN(_1834_));
 DFF_X1 \mem[2][16]$_DFFE_PP_  (.D(_0343_),
    .CK(clknet_leaf_47_clk),
    .Q(\mem[2][16] ),
    .QN(_1833_));
 DFF_X1 \mem[2][17]$_DFFE_PP_  (.D(_0344_),
    .CK(clknet_leaf_44_clk),
    .Q(\mem[2][17] ),
    .QN(_1832_));
 DFF_X1 \mem[2][18]$_DFFE_PP_  (.D(_0345_),
    .CK(clknet_leaf_62_clk),
    .Q(\mem[2][18] ),
    .QN(_1831_));
 DFF_X1 \mem[2][19]$_DFFE_PP_  (.D(_0346_),
    .CK(clknet_leaf_6_clk),
    .Q(\mem[2][19] ),
    .QN(_1830_));
 DFF_X1 \mem[2][1]$_DFFE_PP_  (.D(_0347_),
    .CK(clknet_leaf_42_clk),
    .Q(\mem[2][1] ),
    .QN(_1829_));
 DFF_X1 \mem[2][20]$_DFFE_PP_  (.D(_0348_),
    .CK(clknet_leaf_35_clk),
    .Q(\mem[2][20] ),
    .QN(_1828_));
 DFF_X1 \mem[2][21]$_DFFE_PP_  (.D(_0349_),
    .CK(clknet_leaf_35_clk),
    .Q(\mem[2][21] ),
    .QN(_1827_));
 DFF_X1 \mem[2][22]$_DFFE_PP_  (.D(_0350_),
    .CK(clknet_leaf_30_clk),
    .Q(\mem[2][22] ),
    .QN(_1826_));
 DFF_X1 \mem[2][23]$_DFFE_PP_  (.D(_0351_),
    .CK(clknet_leaf_23_clk),
    .Q(\mem[2][23] ),
    .QN(_1825_));
 DFF_X1 \mem[2][24]$_DFFE_PP_  (.D(_0352_),
    .CK(clknet_leaf_23_clk),
    .Q(\mem[2][24] ),
    .QN(_1824_));
 DFF_X1 \mem[2][25]$_DFFE_PP_  (.D(_0353_),
    .CK(clknet_leaf_28_clk),
    .Q(\mem[2][25] ),
    .QN(_1823_));
 DFF_X1 \mem[2][26]$_DFFE_PP_  (.D(_0354_),
    .CK(clknet_leaf_26_clk),
    .Q(\mem[2][26] ),
    .QN(_1822_));
 DFF_X1 \mem[2][27]$_DFFE_PP_  (.D(_0355_),
    .CK(clknet_leaf_8_clk),
    .Q(\mem[2][27] ),
    .QN(_1821_));
 DFF_X1 \mem[2][28]$_DFFE_PP_  (.D(_0356_),
    .CK(clknet_leaf_24_clk),
    .Q(\mem[2][28] ),
    .QN(_1820_));
 DFF_X1 \mem[2][29]$_DFFE_PP_  (.D(_0357_),
    .CK(clknet_leaf_16_clk),
    .Q(\mem[2][29] ),
    .QN(_1819_));
 DFF_X1 \mem[2][2]$_DFFE_PP_  (.D(_0358_),
    .CK(clknet_leaf_16_clk),
    .Q(\mem[2][2] ),
    .QN(_1818_));
 DFF_X1 \mem[2][30]$_DFFE_PP_  (.D(_0359_),
    .CK(clknet_leaf_12_clk),
    .Q(\mem[2][30] ),
    .QN(_1817_));
 DFF_X1 \mem[2][31]$_DFFE_PP_  (.D(_0360_),
    .CK(clknet_leaf_11_clk),
    .Q(\mem[2][31] ),
    .QN(_1816_));
 DFF_X1 \mem[2][3]$_DFFE_PP_  (.D(_0361_),
    .CK(clknet_leaf_12_clk),
    .Q(\mem[2][3] ),
    .QN(_1815_));
 DFF_X1 \mem[2][4]$_DFFE_PP_  (.D(_0362_),
    .CK(clknet_leaf_11_clk),
    .Q(\mem[2][4] ),
    .QN(_1814_));
 DFF_X1 \mem[2][5]$_DFFE_PP_  (.D(_0363_),
    .CK(clknet_leaf_76_clk),
    .Q(\mem[2][5] ),
    .QN(_1813_));
 DFF_X1 \mem[2][6]$_DFFE_PP_  (.D(_0364_),
    .CK(clknet_leaf_75_clk),
    .Q(\mem[2][6] ),
    .QN(_1812_));
 DFF_X1 \mem[2][7]$_DFFE_PP_  (.D(_0365_),
    .CK(clknet_leaf_75_clk),
    .Q(\mem[2][7] ),
    .QN(_1811_));
 DFF_X1 \mem[2][8]$_DFFE_PP_  (.D(_0366_),
    .CK(clknet_leaf_76_clk),
    .Q(\mem[2][8] ),
    .QN(_1810_));
 DFF_X1 \mem[2][9]$_DFFE_PP_  (.D(_0367_),
    .CK(clknet_leaf_72_clk),
    .Q(\mem[2][9] ),
    .QN(_1809_));
 DFF_X1 \mem[3][0]$_DFFE_PP_  (.D(_0368_),
    .CK(clknet_leaf_65_clk),
    .Q(\mem[3][0] ),
    .QN(_1808_));
 DFF_X1 \mem[3][10]$_DFFE_PP_  (.D(_0369_),
    .CK(clknet_leaf_55_clk),
    .Q(\mem[3][10] ),
    .QN(_1807_));
 DFF_X1 \mem[3][11]$_DFFE_PP_  (.D(_0370_),
    .CK(clknet_leaf_60_clk),
    .Q(\mem[3][11] ),
    .QN(_1806_));
 DFF_X1 \mem[3][12]$_DFFE_PP_  (.D(_0371_),
    .CK(clknet_leaf_55_clk),
    .Q(\mem[3][12] ),
    .QN(_1805_));
 DFF_X1 \mem[3][13]$_DFFE_PP_  (.D(_0372_),
    .CK(clknet_leaf_68_clk),
    .Q(\mem[3][13] ),
    .QN(_1804_));
 DFF_X1 \mem[3][14]$_DFFE_PP_  (.D(_0373_),
    .CK(clknet_leaf_56_clk),
    .Q(\mem[3][14] ),
    .QN(_1803_));
 DFF_X1 \mem[3][15]$_DFFE_PP_  (.D(_0374_),
    .CK(clknet_leaf_56_clk),
    .Q(\mem[3][15] ),
    .QN(_1802_));
 DFF_X1 \mem[3][16]$_DFFE_PP_  (.D(_0375_),
    .CK(clknet_leaf_47_clk),
    .Q(\mem[3][16] ),
    .QN(_1801_));
 DFF_X1 \mem[3][17]$_DFFE_PP_  (.D(_0376_),
    .CK(clknet_leaf_27_clk),
    .Q(\mem[3][17] ),
    .QN(_1800_));
 DFF_X1 \mem[3][18]$_DFFE_PP_  (.D(_0377_),
    .CK(clknet_leaf_62_clk),
    .Q(\mem[3][18] ),
    .QN(_1799_));
 DFF_X1 \mem[3][19]$_DFFE_PP_  (.D(_0378_),
    .CK(clknet_leaf_7_clk),
    .Q(\mem[3][19] ),
    .QN(_1798_));
 DFF_X1 \mem[3][1]$_DFFE_PP_  (.D(_0379_),
    .CK(clknet_leaf_42_clk),
    .Q(\mem[3][1] ),
    .QN(_1797_));
 DFF_X1 \mem[3][20]$_DFFE_PP_  (.D(_0380_),
    .CK(clknet_leaf_35_clk),
    .Q(\mem[3][20] ),
    .QN(_1796_));
 DFF_X1 \mem[3][21]$_DFFE_PP_  (.D(_0381_),
    .CK(clknet_leaf_35_clk),
    .Q(\mem[3][21] ),
    .QN(_1795_));
 DFF_X1 \mem[3][22]$_DFFE_PP_  (.D(_0382_),
    .CK(clknet_leaf_30_clk),
    .Q(\mem[3][22] ),
    .QN(_1794_));
 DFF_X1 \mem[3][23]$_DFFE_PP_  (.D(_0383_),
    .CK(clknet_leaf_24_clk),
    .Q(\mem[3][23] ),
    .QN(_1793_));
 DFF_X1 \mem[3][24]$_DFFE_PP_  (.D(_0384_),
    .CK(clknet_leaf_31_clk),
    .Q(\mem[3][24] ),
    .QN(_1792_));
 DFF_X1 \mem[3][25]$_DFFE_PP_  (.D(_0385_),
    .CK(clknet_leaf_26_clk),
    .Q(\mem[3][25] ),
    .QN(_1791_));
 DFF_X1 \mem[3][26]$_DFFE_PP_  (.D(_0386_),
    .CK(clknet_leaf_26_clk),
    .Q(\mem[3][26] ),
    .QN(_1790_));
 DFF_X1 \mem[3][27]$_DFFE_PP_  (.D(_0387_),
    .CK(clknet_leaf_25_clk),
    .Q(\mem[3][27] ),
    .QN(_1789_));
 DFF_X1 \mem[3][28]$_DFFE_PP_  (.D(_0388_),
    .CK(clknet_leaf_19_clk),
    .Q(\mem[3][28] ),
    .QN(_1788_));
 DFF_X1 \mem[3][29]$_DFFE_PP_  (.D(_0389_),
    .CK(clknet_leaf_14_clk),
    .Q(\mem[3][29] ),
    .QN(_1787_));
 DFF_X1 \mem[3][2]$_DFFE_PP_  (.D(_0390_),
    .CK(clknet_leaf_13_clk),
    .Q(\mem[3][2] ),
    .QN(_1786_));
 DFF_X1 \mem[3][30]$_DFFE_PP_  (.D(_0391_),
    .CK(clknet_leaf_13_clk),
    .Q(\mem[3][30] ),
    .QN(_1785_));
 DFF_X1 \mem[3][31]$_DFFE_PP_  (.D(_0392_),
    .CK(clknet_leaf_11_clk),
    .Q(\mem[3][31] ),
    .QN(_1784_));
 DFF_X1 \mem[3][3]$_DFFE_PP_  (.D(_0393_),
    .CK(clknet_leaf_12_clk),
    .Q(\mem[3][3] ),
    .QN(_1783_));
 DFF_X1 \mem[3][4]$_DFFE_PP_  (.D(_0394_),
    .CK(clknet_leaf_12_clk),
    .Q(\mem[3][4] ),
    .QN(_1782_));
 DFF_X1 \mem[3][5]$_DFFE_PP_  (.D(_0395_),
    .CK(clknet_leaf_76_clk),
    .Q(\mem[3][5] ),
    .QN(_1781_));
 DFF_X1 \mem[3][6]$_DFFE_PP_  (.D(_0396_),
    .CK(clknet_leaf_76_clk),
    .Q(\mem[3][6] ),
    .QN(_1780_));
 DFF_X1 \mem[3][7]$_DFFE_PP_  (.D(_0397_),
    .CK(clknet_leaf_75_clk),
    .Q(\mem[3][7] ),
    .QN(_1779_));
 DFF_X1 \mem[3][8]$_DFFE_PP_  (.D(_0398_),
    .CK(clknet_leaf_76_clk),
    .Q(\mem[3][8] ),
    .QN(_1778_));
 DFF_X1 \mem[3][9]$_DFFE_PP_  (.D(_0399_),
    .CK(clknet_leaf_72_clk),
    .Q(\mem[3][9] ),
    .QN(_1777_));
 DFF_X1 \mem[4][0]$_DFFE_PP_  (.D(_0400_),
    .CK(clknet_leaf_63_clk),
    .Q(\mem[4][0] ),
    .QN(_1776_));
 DFF_X1 \mem[4][10]$_DFFE_PP_  (.D(_0401_),
    .CK(clknet_leaf_54_clk),
    .Q(\mem[4][10] ),
    .QN(_1775_));
 DFF_X1 \mem[4][11]$_DFFE_PP_  (.D(_0402_),
    .CK(clknet_leaf_59_clk),
    .Q(\mem[4][11] ),
    .QN(_1774_));
 DFF_X1 \mem[4][12]$_DFFE_PP_  (.D(_0403_),
    .CK(clknet_leaf_54_clk),
    .Q(\mem[4][12] ),
    .QN(_1773_));
 DFF_X1 \mem[4][13]$_DFFE_PP_  (.D(_0404_),
    .CK(clknet_leaf_70_clk),
    .Q(\mem[4][13] ),
    .QN(_1772_));
 DFF_X1 \mem[4][14]$_DFFE_PP_  (.D(_0405_),
    .CK(clknet_leaf_57_clk),
    .Q(\mem[4][14] ),
    .QN(_1771_));
 DFF_X1 \mem[4][15]$_DFFE_PP_  (.D(_0406_),
    .CK(clknet_leaf_57_clk),
    .Q(\mem[4][15] ),
    .QN(_1770_));
 DFF_X1 \mem[4][16]$_DFFE_PP_  (.D(_0407_),
    .CK(clknet_leaf_47_clk),
    .Q(\mem[4][16] ),
    .QN(_1769_));
 DFF_X1 \mem[4][17]$_DFFE_PP_  (.D(_0408_),
    .CK(clknet_leaf_44_clk),
    .Q(\mem[4][17] ),
    .QN(_1768_));
 DFF_X1 \mem[4][18]$_DFFE_PP_  (.D(_0409_),
    .CK(clknet_leaf_47_clk),
    .Q(\mem[4][18] ),
    .QN(_1767_));
 DFF_X1 \mem[4][19]$_DFFE_PP_  (.D(_0410_),
    .CK(clknet_leaf_6_clk),
    .Q(\mem[4][19] ),
    .QN(_1766_));
 DFF_X1 \mem[4][1]$_DFFE_PP_  (.D(_0411_),
    .CK(clknet_leaf_29_clk),
    .Q(\mem[4][1] ),
    .QN(_1765_));
 DFF_X1 \mem[4][20]$_DFFE_PP_  (.D(_0412_),
    .CK(clknet_leaf_30_clk),
    .Q(\mem[4][20] ),
    .QN(_1764_));
 DFF_X1 \mem[4][21]$_DFFE_PP_  (.D(_0413_),
    .CK(clknet_leaf_35_clk),
    .Q(\mem[4][21] ),
    .QN(_1763_));
 DFF_X1 \mem[4][22]$_DFFE_PP_  (.D(_0414_),
    .CK(clknet_leaf_33_clk),
    .Q(\mem[4][22] ),
    .QN(_1762_));
 DFF_X1 \mem[4][23]$_DFFE_PP_  (.D(_0415_),
    .CK(clknet_leaf_23_clk),
    .Q(\mem[4][23] ),
    .QN(_1761_));
 DFF_X1 \mem[4][24]$_DFFE_PP_  (.D(_0416_),
    .CK(clknet_leaf_31_clk),
    .Q(\mem[4][24] ),
    .QN(_1760_));
 DFF_X1 \mem[4][25]$_DFFE_PP_  (.D(_0417_),
    .CK(clknet_leaf_28_clk),
    .Q(\mem[4][25] ),
    .QN(_1759_));
 DFF_X1 \mem[4][26]$_DFFE_PP_  (.D(_0418_),
    .CK(clknet_leaf_28_clk),
    .Q(\mem[4][26] ),
    .QN(_1758_));
 DFF_X1 \mem[4][27]$_DFFE_PP_  (.D(_0419_),
    .CK(clknet_leaf_25_clk),
    .Q(\mem[4][27] ),
    .QN(_1757_));
 DFF_X1 \mem[4][28]$_DFFE_PP_  (.D(_0420_),
    .CK(clknet_leaf_19_clk),
    .Q(\mem[4][28] ),
    .QN(_1756_));
 DFF_X1 \mem[4][29]$_DFFE_PP_  (.D(_0421_),
    .CK(clknet_leaf_18_clk),
    .Q(\mem[4][29] ),
    .QN(_1755_));
 DFF_X1 \mem[4][2]$_DFFE_PP_  (.D(_0422_),
    .CK(clknet_leaf_19_clk),
    .Q(\mem[4][2] ),
    .QN(_1754_));
 DFF_X1 \mem[4][30]$_DFFE_PP_  (.D(_0423_),
    .CK(clknet_leaf_9_clk),
    .Q(\mem[4][30] ),
    .QN(_1753_));
 DFF_X1 \mem[4][31]$_DFFE_PP_  (.D(_0424_),
    .CK(clknet_leaf_8_clk),
    .Q(\mem[4][31] ),
    .QN(_1752_));
 DFF_X1 \mem[4][3]$_DFFE_PP_  (.D(_0425_),
    .CK(clknet_leaf_9_clk),
    .Q(\mem[4][3] ),
    .QN(_1751_));
 DFF_X1 \mem[4][4]$_DFFE_PP_  (.D(_0426_),
    .CK(clknet_leaf_10_clk),
    .Q(\mem[4][4] ),
    .QN(_1750_));
 DFF_X1 \mem[4][5]$_DFFE_PP_  (.D(_0427_),
    .CK(clknet_leaf_4_clk),
    .Q(\mem[4][5] ),
    .QN(_1749_));
 DFF_X1 \mem[4][6]$_DFFE_PP_  (.D(_0428_),
    .CK(clknet_leaf_67_clk),
    .Q(\mem[4][6] ),
    .QN(_1748_));
 DFF_X1 \mem[4][7]$_DFFE_PP_  (.D(_0429_),
    .CK(clknet_leaf_74_clk),
    .Q(\mem[4][7] ),
    .QN(_1747_));
 DFF_X1 \mem[4][8]$_DFFE_PP_  (.D(_0430_),
    .CK(clknet_leaf_66_clk),
    .Q(\mem[4][8] ),
    .QN(_1746_));
 DFF_X1 \mem[4][9]$_DFFE_PP_  (.D(_0431_),
    .CK(clknet_leaf_71_clk),
    .Q(\mem[4][9] ),
    .QN(_1745_));
 DFF_X1 \mem[5][0]$_DFFE_PP_  (.D(_0432_),
    .CK(clknet_leaf_64_clk),
    .Q(\mem[5][0] ),
    .QN(_1744_));
 DFF_X1 \mem[5][10]$_DFFE_PP_  (.D(_0433_),
    .CK(clknet_leaf_54_clk),
    .Q(\mem[5][10] ),
    .QN(_1743_));
 DFF_X1 \mem[5][11]$_DFFE_PP_  (.D(_0434_),
    .CK(clknet_leaf_59_clk),
    .Q(\mem[5][11] ),
    .QN(_1742_));
 DFF_X1 \mem[5][12]$_DFFE_PP_  (.D(_0435_),
    .CK(clknet_leaf_54_clk),
    .Q(\mem[5][12] ),
    .QN(_1741_));
 DFF_X1 \mem[5][13]$_DFFE_PP_  (.D(_0436_),
    .CK(clknet_leaf_69_clk),
    .Q(\mem[5][13] ),
    .QN(_1740_));
 DFF_X1 \mem[5][14]$_DFFE_PP_  (.D(_0437_),
    .CK(clknet_leaf_57_clk),
    .Q(\mem[5][14] ),
    .QN(_1739_));
 DFF_X1 \mem[5][15]$_DFFE_PP_  (.D(_0438_),
    .CK(clknet_leaf_57_clk),
    .Q(\mem[5][15] ),
    .QN(_1738_));
 DFF_X1 \mem[5][16]$_DFFE_PP_  (.D(_0439_),
    .CK(clknet_leaf_51_clk),
    .Q(\mem[5][16] ),
    .QN(_1737_));
 DFF_X1 \mem[5][17]$_DFFE_PP_  (.D(_0440_),
    .CK(clknet_leaf_45_clk),
    .Q(\mem[5][17] ),
    .QN(_1736_));
 DFF_X1 \mem[5][18]$_DFFE_PP_  (.D(_0441_),
    .CK(clknet_leaf_46_clk),
    .Q(\mem[5][18] ),
    .QN(_1735_));
 DFF_X1 \mem[5][19]$_DFFE_PP_  (.D(_0442_),
    .CK(clknet_leaf_26_clk),
    .Q(\mem[5][19] ),
    .QN(_1734_));
 DFF_X1 \mem[5][1]$_DFFE_PP_  (.D(_0443_),
    .CK(clknet_leaf_29_clk),
    .Q(\mem[5][1] ),
    .QN(_1733_));
 DFF_X1 \mem[5][20]$_DFFE_PP_  (.D(_0444_),
    .CK(clknet_leaf_30_clk),
    .Q(\mem[5][20] ),
    .QN(_1732_));
 DFF_X1 \mem[5][21]$_DFFE_PP_  (.D(_0445_),
    .CK(clknet_leaf_36_clk),
    .Q(\mem[5][21] ),
    .QN(_1731_));
 DFF_X1 \mem[5][22]$_DFFE_PP_  (.D(_0446_),
    .CK(clknet_leaf_34_clk),
    .Q(\mem[5][22] ),
    .QN(_1730_));
 DFF_X1 \mem[5][23]$_DFFE_PP_  (.D(_0447_),
    .CK(clknet_leaf_21_clk),
    .Q(\mem[5][23] ),
    .QN(_1729_));
 DFF_X1 \mem[5][24]$_DFFE_PP_  (.D(_0448_),
    .CK(clknet_leaf_32_clk),
    .Q(\mem[5][24] ),
    .QN(_1728_));
 DFF_X1 \mem[5][25]$_DFFE_PP_  (.D(_0449_),
    .CK(clknet_leaf_27_clk),
    .Q(\mem[5][25] ),
    .QN(_1727_));
 DFF_X1 \mem[5][26]$_DFFE_PP_  (.D(_0450_),
    .CK(clknet_leaf_28_clk),
    .Q(\mem[5][26] ),
    .QN(_1726_));
 DFF_X1 \mem[5][27]$_DFFE_PP_  (.D(_0451_),
    .CK(clknet_leaf_24_clk),
    .Q(\mem[5][27] ),
    .QN(_1725_));
 DFF_X1 \mem[5][28]$_DFFE_PP_  (.D(_0452_),
    .CK(clknet_leaf_20_clk),
    .Q(\mem[5][28] ),
    .QN(_1724_));
 DFF_X1 \mem[5][29]$_DFFE_PP_  (.D(_0453_),
    .CK(clknet_leaf_18_clk),
    .Q(\mem[5][29] ),
    .QN(_1723_));
 DFF_X1 \mem[5][2]$_DFFE_PP_  (.D(_0454_),
    .CK(clknet_leaf_15_clk),
    .Q(\mem[5][2] ),
    .QN(_1722_));
 DFF_X1 \mem[5][30]$_DFFE_PP_  (.D(_0455_),
    .CK(clknet_leaf_9_clk),
    .Q(\mem[5][30] ),
    .QN(_1721_));
 DFF_X1 \mem[5][31]$_DFFE_PP_  (.D(_0456_),
    .CK(clknet_leaf_8_clk),
    .Q(\mem[5][31] ),
    .QN(_1720_));
 DFF_X1 \mem[5][3]$_DFFE_PP_  (.D(_0457_),
    .CK(clknet_leaf_9_clk),
    .Q(\mem[5][3] ),
    .QN(_1719_));
 DFF_X1 \mem[5][4]$_DFFE_PP_  (.D(_0458_),
    .CK(clknet_leaf_10_clk),
    .Q(\mem[5][4] ),
    .QN(_1718_));
 DFF_X1 \mem[5][5]$_DFFE_PP_  (.D(_0459_),
    .CK(clknet_leaf_4_clk),
    .Q(\mem[5][5] ),
    .QN(_1717_));
 DFF_X1 \mem[5][6]$_DFFE_PP_  (.D(_0460_),
    .CK(clknet_leaf_67_clk),
    .Q(\mem[5][6] ),
    .QN(_1716_));
 DFF_X1 \mem[5][7]$_DFFE_PP_  (.D(_0461_),
    .CK(clknet_leaf_71_clk),
    .Q(\mem[5][7] ),
    .QN(_1715_));
 DFF_X1 \mem[5][8]$_DFFE_PP_  (.D(_0462_),
    .CK(clknet_leaf_66_clk),
    .Q(\mem[5][8] ),
    .QN(_1714_));
 DFF_X1 \mem[5][9]$_DFFE_PP_  (.D(_0463_),
    .CK(clknet_leaf_72_clk),
    .Q(\mem[5][9] ),
    .QN(_1713_));
 DFF_X1 \mem[6][0]$_DFFE_PP_  (.D(_0464_),
    .CK(clknet_leaf_68_clk),
    .Q(\mem[6][0] ),
    .QN(_1712_));
 DFF_X1 \mem[6][10]$_DFFE_PP_  (.D(_0465_),
    .CK(clknet_leaf_51_clk),
    .Q(\mem[6][10] ),
    .QN(_1711_));
 DFF_X1 \mem[6][11]$_DFFE_PP_  (.D(_0466_),
    .CK(clknet_leaf_68_clk),
    .Q(\mem[6][11] ),
    .QN(_1710_));
 DFF_X1 \mem[6][12]$_DFFE_PP_  (.D(_0467_),
    .CK(clknet_leaf_55_clk),
    .Q(\mem[6][12] ),
    .QN(_1709_));
 DFF_X1 \mem[6][13]$_DFFE_PP_  (.D(_0468_),
    .CK(clknet_leaf_67_clk),
    .Q(\mem[6][13] ),
    .QN(_1708_));
 DFF_X1 \mem[6][14]$_DFFE_PP_  (.D(_0469_),
    .CK(clknet_leaf_56_clk),
    .Q(\mem[6][14] ),
    .QN(_1707_));
 DFF_X1 \mem[6][15]$_DFFE_PP_  (.D(_0470_),
    .CK(clknet_leaf_61_clk),
    .Q(\mem[6][15] ),
    .QN(_1706_));
 DFF_X1 \mem[6][16]$_DFFE_PP_  (.D(_0471_),
    .CK(clknet_leaf_47_clk),
    .Q(\mem[6][16] ),
    .QN(_1705_));
 DFF_X1 \mem[6][17]$_DFFE_PP_  (.D(_0472_),
    .CK(clknet_leaf_44_clk),
    .Q(\mem[6][17] ),
    .QN(_1704_));
 DFF_X1 \mem[6][18]$_DFFE_PP_  (.D(_0473_),
    .CK(clknet_leaf_63_clk),
    .Q(\mem[6][18] ),
    .QN(_1703_));
 DFF_X1 \mem[6][19]$_DFFE_PP_  (.D(_0474_),
    .CK(clknet_leaf_5_clk),
    .Q(\mem[6][19] ),
    .QN(_1702_));
 DFF_X1 \mem[6][1]$_DFFE_PP_  (.D(_0475_),
    .CK(clknet_leaf_42_clk),
    .Q(\mem[6][1] ),
    .QN(_1701_));
 DFF_X1 \mem[6][20]$_DFFE_PP_  (.D(_0476_),
    .CK(clknet_leaf_35_clk),
    .Q(\mem[6][20] ),
    .QN(_1700_));
 DFF_X1 \mem[6][21]$_DFFE_PP_  (.D(_0477_),
    .CK(clknet_leaf_35_clk),
    .Q(\mem[6][21] ),
    .QN(_1699_));
 DFF_X1 \mem[6][22]$_DFFE_PP_  (.D(_0478_),
    .CK(clknet_leaf_32_clk),
    .Q(\mem[6][22] ),
    .QN(_1698_));
 DFF_X1 \mem[6][23]$_DFFE_PP_  (.D(_0479_),
    .CK(clknet_leaf_24_clk),
    .Q(\mem[6][23] ),
    .QN(_1697_));
 DFF_X1 \mem[6][24]$_DFFE_PP_  (.D(_0480_),
    .CK(clknet_leaf_23_clk),
    .Q(\mem[6][24] ),
    .QN(_1696_));
 DFF_X1 \mem[6][25]$_DFFE_PP_  (.D(_0481_),
    .CK(clknet_leaf_28_clk),
    .Q(\mem[6][25] ),
    .QN(_1695_));
 DFF_X1 \mem[6][26]$_DFFE_PP_  (.D(_0482_),
    .CK(clknet_leaf_26_clk),
    .Q(\mem[6][26] ),
    .QN(_1694_));
 DFF_X1 \mem[6][27]$_DFFE_PP_  (.D(_0483_),
    .CK(clknet_leaf_25_clk),
    .Q(\mem[6][27] ),
    .QN(_1693_));
 DFF_X1 \mem[6][28]$_DFFE_PP_  (.D(_0484_),
    .CK(clknet_leaf_19_clk),
    .Q(\mem[6][28] ),
    .QN(_1692_));
 DFF_X1 \mem[6][29]$_DFFE_PP_  (.D(_0485_),
    .CK(clknet_leaf_16_clk),
    .Q(\mem[6][29] ),
    .QN(_1691_));
 DFF_X1 \mem[6][2]$_DFFE_PP_  (.D(_0486_),
    .CK(clknet_leaf_16_clk),
    .Q(\mem[6][2] ),
    .QN(_1690_));
 DFF_X1 \mem[6][30]$_DFFE_PP_  (.D(_0487_),
    .CK(clknet_leaf_13_clk),
    .Q(\mem[6][30] ),
    .QN(_1689_));
 DFF_X1 \mem[6][31]$_DFFE_PP_  (.D(_0488_),
    .CK(clknet_leaf_11_clk),
    .Q(\mem[6][31] ),
    .QN(_1688_));
 DFF_X1 \mem[6][3]$_DFFE_PP_  (.D(_0489_),
    .CK(clknet_leaf_12_clk),
    .Q(\mem[6][3] ),
    .QN(_1687_));
 DFF_X1 \mem[6][4]$_DFFE_PP_  (.D(_0490_),
    .CK(clknet_leaf_11_clk),
    .Q(\mem[6][4] ),
    .QN(_1686_));
 DFF_X1 \mem[6][5]$_DFFE_PP_  (.D(_0491_),
    .CK(clknet_leaf_1_clk),
    .Q(\mem[6][5] ),
    .QN(_1685_));
 DFF_X1 \mem[6][6]$_DFFE_PP_  (.D(_0492_),
    .CK(clknet_leaf_75_clk),
    .Q(\mem[6][6] ),
    .QN(_1684_));
 DFF_X1 \mem[6][7]$_DFFE_PP_  (.D(_0493_),
    .CK(clknet_leaf_75_clk),
    .Q(\mem[6][7] ),
    .QN(_1683_));
 DFF_X1 \mem[6][8]$_DFFE_PP_  (.D(_0494_),
    .CK(clknet_leaf_0_clk),
    .Q(\mem[6][8] ),
    .QN(_1682_));
 DFF_X1 \mem[6][9]$_DFFE_PP_  (.D(_0495_),
    .CK(clknet_leaf_72_clk),
    .Q(\mem[6][9] ),
    .QN(_1681_));
 DFF_X1 \mem[7][0]$_DFFE_PP_  (.D(_0496_),
    .CK(clknet_leaf_65_clk),
    .Q(\mem[7][0] ),
    .QN(_1680_));
 DFF_X1 \mem[7][10]$_DFFE_PP_  (.D(_0497_),
    .CK(clknet_leaf_52_clk),
    .Q(\mem[7][10] ),
    .QN(_1679_));
 DFF_X1 \mem[7][11]$_DFFE_PP_  (.D(_0498_),
    .CK(clknet_leaf_60_clk),
    .Q(\mem[7][11] ),
    .QN(_1678_));
 DFF_X1 \mem[7][12]$_DFFE_PP_  (.D(_0499_),
    .CK(clknet_leaf_51_clk),
    .Q(\mem[7][12] ),
    .QN(_1677_));
 DFF_X1 \mem[7][13]$_DFFE_PP_  (.D(_0500_),
    .CK(clknet_leaf_68_clk),
    .Q(\mem[7][13] ),
    .QN(_1676_));
 DFF_X1 \mem[7][14]$_DFFE_PP_  (.D(_0501_),
    .CK(clknet_leaf_56_clk),
    .Q(\mem[7][14] ),
    .QN(_1675_));
 DFF_X1 \mem[7][15]$_DFFE_PP_  (.D(_0502_),
    .CK(clknet_leaf_56_clk),
    .Q(\mem[7][15] ),
    .QN(_1674_));
 DFF_X1 \mem[7][16]$_DFFE_PP_  (.D(_0503_),
    .CK(clknet_leaf_48_clk),
    .Q(\mem[7][16] ),
    .QN(_1673_));
 DFF_X1 \mem[7][17]$_DFFE_PP_  (.D(_0504_),
    .CK(clknet_leaf_27_clk),
    .Q(\mem[7][17] ),
    .QN(_1672_));
 DFF_X1 \mem[7][18]$_DFFE_PP_  (.D(_0505_),
    .CK(clknet_leaf_62_clk),
    .Q(\mem[7][18] ),
    .QN(_1671_));
 DFF_X1 \mem[7][19]$_DFFE_PP_  (.D(_0506_),
    .CK(clknet_leaf_6_clk),
    .Q(\mem[7][19] ),
    .QN(_1670_));
 DFF_X1 \mem[7][1]$_DFFE_PP_  (.D(_0507_),
    .CK(clknet_leaf_42_clk),
    .Q(\mem[7][1] ),
    .QN(_1669_));
 DFF_X1 \mem[7][20]$_DFFE_PP_  (.D(_0508_),
    .CK(clknet_leaf_38_clk),
    .Q(\mem[7][20] ),
    .QN(_1668_));
 DFF_X1 \mem[7][21]$_DFFE_PP_  (.D(_0509_),
    .CK(clknet_leaf_36_clk),
    .Q(\mem[7][21] ),
    .QN(_1667_));
 DFF_X1 \mem[7][22]$_DFFE_PP_  (.D(_0510_),
    .CK(clknet_leaf_35_clk),
    .Q(\mem[7][22] ),
    .QN(_1666_));
 DFF_X1 \mem[7][23]$_DFFE_PP_  (.D(_0511_),
    .CK(clknet_leaf_24_clk),
    .Q(\mem[7][23] ),
    .QN(_1665_));
 DFF_X1 \mem[7][24]$_DFFE_PP_  (.D(_0512_),
    .CK(clknet_leaf_31_clk),
    .Q(\mem[7][24] ),
    .QN(_1664_));
 DFF_X1 \mem[7][25]$_DFFE_PP_  (.D(_0513_),
    .CK(clknet_leaf_28_clk),
    .Q(\mem[7][25] ),
    .QN(_1663_));
 DFF_X1 \mem[7][26]$_DFFE_PP_  (.D(_0514_),
    .CK(clknet_leaf_23_clk),
    .Q(\mem[7][26] ),
    .QN(_1662_));
 DFF_X1 \mem[7][27]$_DFFE_PP_  (.D(_0515_),
    .CK(clknet_leaf_26_clk),
    .Q(\mem[7][27] ),
    .QN(_1661_));
 DFF_X1 \mem[7][28]$_DFFE_PP_  (.D(_0516_),
    .CK(clknet_leaf_19_clk),
    .Q(\mem[7][28] ),
    .QN(_1660_));
 DFF_X1 \mem[7][29]$_DFFE_PP_  (.D(_0517_),
    .CK(clknet_leaf_15_clk),
    .Q(\mem[7][29] ),
    .QN(_1659_));
 DFF_X1 \mem[7][2]$_DFFE_PP_  (.D(_0518_),
    .CK(clknet_leaf_13_clk),
    .Q(\mem[7][2] ),
    .QN(_1658_));
 DFF_X1 \mem[7][30]$_DFFE_PP_  (.D(_0519_),
    .CK(clknet_leaf_14_clk),
    .Q(\mem[7][30] ),
    .QN(_1657_));
 DFF_X1 \mem[7][31]$_DFFE_PP_  (.D(_0520_),
    .CK(clknet_leaf_11_clk),
    .Q(\mem[7][31] ),
    .QN(_1656_));
 DFF_X1 \mem[7][3]$_DFFE_PP_  (.D(_0521_),
    .CK(clknet_leaf_12_clk),
    .Q(\mem[7][3] ),
    .QN(_1655_));
 DFF_X1 \mem[7][4]$_DFFE_PP_  (.D(_0522_),
    .CK(clknet_leaf_11_clk),
    .Q(\mem[7][4] ),
    .QN(_1654_));
 DFF_X1 \mem[7][5]$_DFFE_PP_  (.D(_0523_),
    .CK(clknet_leaf_3_clk),
    .Q(\mem[7][5] ),
    .QN(_1653_));
 DFF_X1 \mem[7][6]$_DFFE_PP_  (.D(_0524_),
    .CK(clknet_leaf_76_clk),
    .Q(\mem[7][6] ),
    .QN(_1652_));
 DFF_X1 \mem[7][7]$_DFFE_PP_  (.D(_0525_),
    .CK(clknet_leaf_76_clk),
    .Q(\mem[7][7] ),
    .QN(_1651_));
 DFF_X1 \mem[7][8]$_DFFE_PP_  (.D(_0526_),
    .CK(clknet_leaf_3_clk),
    .Q(\mem[7][8] ),
    .QN(_1650_));
 DFF_X1 \mem[7][9]$_DFFE_PP_  (.D(_0527_),
    .CK(clknet_leaf_72_clk),
    .Q(\mem[7][9] ),
    .QN(_1649_));
 DFF_X1 \mem[8][0]$_DFFE_PP_  (.D(_0528_),
    .CK(clknet_leaf_63_clk),
    .Q(\mem[8][0] ),
    .QN(_1648_));
 DFF_X1 \mem[8][10]$_DFFE_PP_  (.D(_0529_),
    .CK(clknet_leaf_53_clk),
    .Q(\mem[8][10] ),
    .QN(_1647_));
 DFF_X1 \mem[8][11]$_DFFE_PP_  (.D(_0530_),
    .CK(clknet_leaf_70_clk),
    .Q(\mem[8][11] ),
    .QN(_1646_));
 DFF_X1 \mem[8][12]$_DFFE_PP_  (.D(_0531_),
    .CK(clknet_leaf_54_clk),
    .Q(\mem[8][12] ),
    .QN(_1645_));
 DFF_X1 \mem[8][13]$_DFFE_PP_  (.D(_0532_),
    .CK(clknet_leaf_70_clk),
    .Q(\mem[8][13] ),
    .QN(_1644_));
 DFF_X1 \mem[8][14]$_DFFE_PP_  (.D(_0533_),
    .CK(clknet_leaf_58_clk),
    .Q(\mem[8][14] ),
    .QN(_1643_));
 DFF_X1 \mem[8][15]$_DFFE_PP_  (.D(_0534_),
    .CK(clknet_leaf_53_clk),
    .Q(\mem[8][15] ),
    .QN(_1642_));
 DFF_X1 \mem[8][16]$_DFFE_PP_  (.D(_0535_),
    .CK(clknet_leaf_50_clk),
    .Q(\mem[8][16] ),
    .QN(_1641_));
 DFF_X1 \mem[8][17]$_DFFE_PP_  (.D(_0536_),
    .CK(clknet_leaf_45_clk),
    .Q(\mem[8][17] ),
    .QN(_1640_));
 DFF_X1 \mem[8][18]$_DFFE_PP_  (.D(_0537_),
    .CK(clknet_leaf_61_clk),
    .Q(\mem[8][18] ),
    .QN(_1639_));
 DFF_X1 \mem[8][19]$_DFFE_PP_  (.D(_0538_),
    .CK(clknet_leaf_64_clk),
    .Q(\mem[8][19] ),
    .QN(_1638_));
 DFF_X1 \mem[8][1]$_DFFE_PP_  (.D(_0539_),
    .CK(clknet_leaf_39_clk),
    .Q(\mem[8][1] ),
    .QN(_1637_));
 DFF_X1 \mem[8][20]$_DFFE_PP_  (.D(_0540_),
    .CK(clknet_leaf_38_clk),
    .Q(\mem[8][20] ),
    .QN(_1636_));
 DFF_X1 \mem[8][21]$_DFFE_PP_  (.D(_0541_),
    .CK(clknet_leaf_37_clk),
    .Q(\mem[8][21] ),
    .QN(_1635_));
 DFF_X1 \mem[8][22]$_DFFE_PP_  (.D(_0542_),
    .CK(clknet_leaf_33_clk),
    .Q(\mem[8][22] ),
    .QN(_1634_));
 DFF_X1 \mem[8][23]$_DFFE_PP_  (.D(_0543_),
    .CK(clknet_leaf_21_clk),
    .Q(\mem[8][23] ),
    .QN(_1633_));
 DFF_X1 \mem[8][24]$_DFFE_PP_  (.D(_0544_),
    .CK(clknet_leaf_22_clk),
    .Q(\mem[8][24] ),
    .QN(_1632_));
 DFF_X1 \mem[8][25]$_DFFE_PP_  (.D(_0545_),
    .CK(clknet_leaf_42_clk),
    .Q(\mem[8][25] ),
    .QN(_1631_));
 DFF_X1 \mem[8][26]$_DFFE_PP_  (.D(_0546_),
    .CK(clknet_leaf_29_clk),
    .Q(\mem[8][26] ),
    .QN(_1630_));
 DFF_X1 \mem[8][27]$_DFFE_PP_  (.D(_0547_),
    .CK(clknet_leaf_25_clk),
    .Q(\mem[8][27] ),
    .QN(_1629_));
 DFF_X1 \mem[8][28]$_DFFE_PP_  (.D(_0548_),
    .CK(clknet_leaf_20_clk),
    .Q(\mem[8][28] ),
    .QN(_1628_));
 DFF_X1 \mem[8][29]$_DFFE_PP_  (.D(_0549_),
    .CK(clknet_leaf_17_clk),
    .Q(\mem[8][29] ),
    .QN(_1627_));
 DFF_X1 \mem[8][2]$_DFFE_PP_  (.D(_0550_),
    .CK(clknet_leaf_15_clk),
    .Q(\mem[8][2] ),
    .QN(_1626_));
 DFF_X1 \mem[8][30]$_DFFE_PP_  (.D(_0551_),
    .CK(clknet_leaf_14_clk),
    .Q(\mem[8][30] ),
    .QN(_1625_));
 DFF_X1 \mem[8][31]$_DFFE_PP_  (.D(_0552_),
    .CK(clknet_leaf_5_clk),
    .Q(\mem[8][31] ),
    .QN(_1624_));
 DFF_X1 \mem[8][3]$_DFFE_PP_  (.D(_0553_),
    .CK(clknet_leaf_10_clk),
    .Q(\mem[8][3] ),
    .QN(_1623_));
 DFF_X1 \mem[8][4]$_DFFE_PP_  (.D(_0554_),
    .CK(clknet_leaf_2_clk),
    .Q(\mem[8][4] ),
    .QN(_1622_));
 DFF_X1 \mem[8][5]$_DFFE_PP_  (.D(_0555_),
    .CK(clknet_leaf_3_clk),
    .Q(\mem[8][5] ),
    .QN(_1621_));
 DFF_X1 \mem[8][6]$_DFFE_PP_  (.D(_0556_),
    .CK(clknet_leaf_66_clk),
    .Q(\mem[8][6] ),
    .QN(_1620_));
 DFF_X1 \mem[8][7]$_DFFE_PP_  (.D(_0557_),
    .CK(clknet_leaf_74_clk),
    .Q(\mem[8][7] ),
    .QN(_1619_));
 DFF_X1 \mem[8][8]$_DFFE_PP_  (.D(_0558_),
    .CK(clknet_leaf_3_clk),
    .Q(\mem[8][8] ),
    .QN(_1618_));
 DFF_X1 \mem[8][9]$_DFFE_PP_  (.D(_0559_),
    .CK(clknet_leaf_74_clk),
    .Q(\mem[8][9] ),
    .QN(_1617_));
 DFF_X1 \mem[9][0]$_DFFE_PP_  (.D(_0560_),
    .CK(clknet_leaf_64_clk),
    .Q(\mem[9][0] ),
    .QN(_1616_));
 DFF_X1 \mem[9][10]$_DFFE_PP_  (.D(_0561_),
    .CK(clknet_leaf_52_clk),
    .Q(\mem[9][10] ),
    .QN(_1615_));
 DFF_X1 \mem[9][11]$_DFFE_PP_  (.D(_0562_),
    .CK(clknet_leaf_58_clk),
    .Q(\mem[9][11] ),
    .QN(_1614_));
 DFF_X1 \mem[9][12]$_DFFE_PP_  (.D(_0563_),
    .CK(clknet_leaf_53_clk),
    .Q(\mem[9][12] ),
    .QN(_1613_));
 DFF_X1 \mem[9][13]$_DFFE_PP_  (.D(_0564_),
    .CK(clknet_leaf_69_clk),
    .Q(\mem[9][13] ),
    .QN(_1612_));
 DFF_X1 \mem[9][14]$_DFFE_PP_  (.D(_0565_),
    .CK(clknet_leaf_58_clk),
    .Q(\mem[9][14] ),
    .QN(_1611_));
 DFF_X1 \mem[9][15]$_DFFE_PP_  (.D(_0566_),
    .CK(clknet_leaf_59_clk),
    .Q(\mem[9][15] ),
    .QN(_1610_));
 DFF_X1 \mem[9][16]$_DFFE_PP_  (.D(_0567_),
    .CK(clknet_leaf_52_clk),
    .Q(\mem[9][16] ),
    .QN(_1609_));
 DFF_X1 \mem[9][17]$_DFFE_PP_  (.D(_0568_),
    .CK(clknet_leaf_44_clk),
    .Q(\mem[9][17] ),
    .QN(_1608_));
 DFF_X1 \mem[9][18]$_DFFE_PP_  (.D(_0569_),
    .CK(clknet_leaf_47_clk),
    .Q(\mem[9][18] ),
    .QN(_1607_));
 DFF_X1 \mem[9][19]$_DFFE_PP_  (.D(_0570_),
    .CK(clknet_leaf_44_clk),
    .Q(\mem[9][19] ),
    .QN(_1606_));
 DFF_X1 \mem[9][1]$_DFFE_PP_  (.D(_0571_),
    .CK(clknet_leaf_39_clk),
    .Q(\mem[9][1] ),
    .QN(_1605_));
 DFF_X1 \mem[9][20]$_DFFE_PP_  (.D(_0572_),
    .CK(clknet_leaf_38_clk),
    .Q(\mem[9][20] ),
    .QN(_1604_));
 DFF_X1 \mem[9][21]$_DFFE_PP_  (.D(_0573_),
    .CK(clknet_leaf_34_clk),
    .Q(\mem[9][21] ),
    .QN(_1603_));
 DFF_X1 \mem[9][22]$_DFFE_PP_  (.D(_0574_),
    .CK(clknet_leaf_33_clk),
    .Q(\mem[9][22] ),
    .QN(_1602_));
 DFF_X1 \mem[9][23]$_DFFE_PP_  (.D(_0575_),
    .CK(clknet_leaf_22_clk),
    .Q(\mem[9][23] ),
    .QN(_1601_));
 DFF_X1 \mem[9][24]$_DFFE_PP_  (.D(_0576_),
    .CK(clknet_leaf_32_clk),
    .Q(\mem[9][24] ),
    .QN(_1600_));
 DFF_X1 \mem[9][25]$_DFFE_PP_  (.D(_0577_),
    .CK(clknet_leaf_42_clk),
    .Q(\mem[9][25] ),
    .QN(_1599_));
 DFF_X1 \mem[9][26]$_DFFE_PP_  (.D(_0578_),
    .CK(clknet_leaf_31_clk),
    .Q(\mem[9][26] ),
    .QN(_1598_));
 DFF_X1 \mem[9][27]$_DFFE_PP_  (.D(_0579_),
    .CK(clknet_leaf_25_clk),
    .Q(\mem[9][27] ),
    .QN(_1597_));
 DFF_X1 \mem[9][28]$_DFFE_PP_  (.D(_0580_),
    .CK(clknet_leaf_21_clk),
    .Q(\mem[9][28] ),
    .QN(_1596_));
 DFF_X1 \mem[9][29]$_DFFE_PP_  (.D(_0581_),
    .CK(clknet_leaf_18_clk),
    .Q(\mem[9][29] ),
    .QN(_1595_));
 DFF_X1 \mem[9][2]$_DFFE_PP_  (.D(_0582_),
    .CK(clknet_leaf_15_clk),
    .Q(\mem[9][2] ),
    .QN(_1594_));
 DFF_X1 \mem[9][30]$_DFFE_PP_  (.D(_0583_),
    .CK(clknet_leaf_14_clk),
    .Q(\mem[9][30] ),
    .QN(_1593_));
 DFF_X1 \mem[9][31]$_DFFE_PP_  (.D(_0584_),
    .CK(clknet_leaf_4_clk),
    .Q(\mem[9][31] ),
    .QN(_1592_));
 DFF_X1 \mem[9][3]$_DFFE_PP_  (.D(_0585_),
    .CK(clknet_leaf_7_clk),
    .Q(\mem[9][3] ),
    .QN(_1591_));
 DFF_X1 \mem[9][4]$_DFFE_PP_  (.D(_0586_),
    .CK(clknet_leaf_2_clk),
    .Q(\mem[9][4] ),
    .QN(_1590_));
 DFF_X1 \mem[9][5]$_DFFE_PP_  (.D(_0587_),
    .CK(clknet_leaf_3_clk),
    .Q(\mem[9][5] ),
    .QN(_1589_));
 DFF_X1 \mem[9][6]$_DFFE_PP_  (.D(_0588_),
    .CK(clknet_leaf_72_clk),
    .Q(\mem[9][6] ),
    .QN(_1588_));
 DFF_X1 \mem[9][7]$_DFFE_PP_  (.D(_0589_),
    .CK(clknet_leaf_71_clk),
    .Q(\mem[9][7] ),
    .QN(_1587_));
 DFF_X1 \mem[9][8]$_DFFE_PP_  (.D(_0590_),
    .CK(clknet_leaf_3_clk),
    .Q(\mem[9][8] ),
    .QN(_1586_));
 DFF_X1 \mem[9][9]$_DFFE_PP_  (.D(_0591_),
    .CK(clknet_leaf_70_clk),
    .Q(\mem[9][9] ),
    .QN(_1585_));
 DFF_X1 \rd_ptr[0]$_SDFFE_PN0P_  (.D(_0592_),
    .CK(clknet_leaf_41_clk),
    .Q(\rd_ptr[0] ),
    .QN(_0004_));
 DFF_X1 \rd_ptr[1]$_SDFFE_PN0P_  (.D(_0593_),
    .CK(clknet_leaf_41_clk),
    .Q(\rd_ptr[1] ),
    .QN(_2150_));
 DFF_X1 \rd_ptr[2]$_SDFFE_PN0P_  (.D(_0594_),
    .CK(clknet_leaf_40_clk),
    .Q(\rd_ptr[2] ),
    .QN(_2151_));
 DFF_X1 \rd_ptr[3]$_SDFFE_PN0P_  (.D(_0595_),
    .CK(clknet_leaf_43_clk),
    .Q(\rd_ptr[3] ),
    .QN(_2152_));
 DFF_X1 \rd_ptr[4]$_SDFFE_PN0P_  (.D(_0596_),
    .CK(clknet_leaf_41_clk),
    .Q(\rd_ptr[4] ),
    .QN(_1584_));
 DFF_X1 \wr_ptr[0]$_SDFFE_PN0P_  (.D(_0597_),
    .CK(clknet_leaf_41_clk),
    .Q(\wr_ptr[0] ),
    .QN(_0018_));
 DFF_X1 \wr_ptr[1]$_SDFFE_PN0P_  (.D(_0598_),
    .CK(clknet_leaf_41_clk),
    .Q(\wr_ptr[1] ),
    .QN(_2153_));
 DFF_X1 \wr_ptr[2]$_SDFFE_PN0P_  (.D(_0599_),
    .CK(clknet_leaf_42_clk),
    .Q(\wr_ptr[2] ),
    .QN(_1583_));
 DFF_X1 \wr_ptr[3]$_SDFFE_PN0P_  (.D(_0600_),
    .CK(clknet_leaf_40_clk),
    .Q(\wr_ptr[3] ),
    .QN(_1582_));
 DFF_X1 \wr_ptr[4]$_SDFFE_PN0P_  (.D(_0601_),
    .CK(clknet_leaf_40_clk),
    .Q(\wr_ptr[4] ),
    .QN(_1581_));
 CLKBUF_X3 clkload4 (.A(clknet_3_5__leaf_clk));
 INV_X2 clkload5 (.A(clknet_3_6__leaf_clk));
 INV_X2 clkload6 (.A(clknet_3_7__leaf_clk));
 CLKBUF_X1 clkload7 (.A(clknet_leaf_67_clk));
 CLKBUF_X1 clkload8 (.A(clknet_leaf_71_clk));
 INV_X2 clkload9 (.A(clknet_leaf_74_clk));
 CLKBUF_X1 clkload10 (.A(clknet_leaf_5_clk));
 CLKBUF_X1 clkload11 (.A(clknet_leaf_65_clk));
 CLKBUF_X1 clkload12 (.A(clknet_leaf_66_clk));
 CLKBUF_X1 clkload13 (.A(clknet_leaf_76_clk));
 CLKBUF_X1 clkload14 (.A(clknet_leaf_55_clk));
 CLKBUF_X1 clkload15 (.A(clknet_leaf_56_clk));
 CLKBUF_X1 clkload16 (.A(clknet_leaf_58_clk));
 CLKBUF_X1 clkload17 (.A(clknet_leaf_59_clk));
 CLKBUF_X1 clkload18 (.A(clknet_leaf_60_clk));
 INV_X1 clkload19 (.A(clknet_leaf_45_clk));
 INV_X1 clkload20 (.A(clknet_leaf_46_clk));
 CLKBUF_X1 clkload21 (.A(clknet_leaf_47_clk));
 CLKBUF_X1 clkload22 (.A(clknet_leaf_48_clk));
 INV_X1 clkload23 (.A(clknet_leaf_49_clk));
 INV_X1 clkload24 (.A(clknet_leaf_51_clk));
 CLKBUF_X1 clkload25 (.A(clknet_leaf_61_clk));
 CLKBUF_X1 clkload26 (.A(clknet_leaf_62_clk));
 INV_X1 clkload27 (.A(clknet_leaf_63_clk));
 INV_X1 clkload28 (.A(clknet_leaf_6_clk));
 INV_X1 clkload29 (.A(clknet_leaf_7_clk));
 INV_X1 clkload30 (.A(clknet_leaf_8_clk));
 CLKBUF_X1 clkload31 (.A(clknet_leaf_9_clk));
 INV_X1 clkload32 (.A(clknet_leaf_10_clk));
 INV_X1 clkload33 (.A(clknet_leaf_13_clk));
 INV_X1 clkload34 (.A(clknet_leaf_14_clk));
 INV_X1 clkload35 (.A(clknet_leaf_25_clk));
 CLKBUF_X1 clkload36 (.A(clknet_leaf_26_clk));
 INV_X1 clkload37 (.A(clknet_leaf_15_clk));
 INV_X1 clkload38 (.A(clknet_leaf_17_clk));
 INV_X1 clkload39 (.A(clknet_leaf_18_clk));
 INV_X1 clkload40 (.A(clknet_leaf_19_clk));
 INV_X1 clkload41 (.A(clknet_leaf_20_clk));
 CLKBUF_X1 clkload42 (.A(clknet_leaf_21_clk));
 INV_X2 clkload43 (.A(clknet_leaf_22_clk));
 CLKBUF_X1 clkload44 (.A(clknet_leaf_23_clk));
 INV_X1 clkload45 (.A(clknet_leaf_24_clk));
 INV_X1 clkload46 (.A(clknet_leaf_27_clk));
 INV_X1 clkload47 (.A(clknet_leaf_29_clk));
 INV_X1 clkload48 (.A(clknet_leaf_39_clk));
 INV_X2 clkload49 (.A(clknet_leaf_40_clk));
 CLKBUF_X1 clkload50 (.A(clknet_leaf_41_clk));
 CLKBUF_X1 clkload51 (.A(clknet_leaf_42_clk));
 CLKBUF_X1 clkload52 (.A(clknet_leaf_43_clk));
 CLKBUF_X1 clkload53 (.A(clknet_leaf_44_clk));
 CLKBUF_X1 clkload54 (.A(clknet_leaf_36_clk));
 INV_X2 clkload55 (.A(clknet_leaf_37_clk));
 CLKBUF_X1 clkload56 (.A(clknet_leaf_38_clk));
endmodule
