module parameterized_i2c_master (ack_error,
    busy,
    clk,
    done,
    read,
    rst_n,
    scl,
    scl_internal_debug,
    sda,
    sda_internal_debug,
    start,
    stop,
    write,
    addr,
    bit_counter_debug,
    data_in,
    data_out,
    phase,
    shift_reg_debug,
    state);
 output ack_error;
 output busy;
 input clk;
 output done;
 input read;
 input rst_n;
 output scl;
 output scl_internal_debug;
 inout sda;
 output sda_internal_debug;
 input start;
 input stop;
 input write;
 input [6:0] addr;
 output [2:0] bit_counter_debug;
 input [7:0] data_in;
 output [7:0] data_out;
 output [1:0] phase;
 output [7:0] shift_reg_debug;
 output [3:0] state;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire clknet_0_clk;
 wire cmd_read;
 wire cmd_write;
 wire \divider_counter[0] ;
 wire \divider_counter[1] ;
 wire \divider_counter[2] ;
 wire \divider_counter[3] ;
 wire \divider_counter[4] ;
 wire \divider_counter[5] ;
 wire \divider_counter[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 CLKBUF_X2 _352_ (.A(_346_),
    .Z(_041_));
 CLKBUF_X3 _353_ (.A(_041_),
    .Z(_042_));
 BUF_X1 _354_ (.A(\divider_counter[3] ),
    .Z(_043_));
 BUF_X2 _355_ (.A(\divider_counter[2] ),
    .Z(_044_));
 OR4_X4 _356_ (.A1(\divider_counter[5] ),
    .A2(\divider_counter[4] ),
    .A3(_043_),
    .A4(_044_),
    .ZN(_045_));
 OR3_X2 _357_ (.A1(\divider_counter[6] ),
    .A2(\divider_counter[1] ),
    .A3(\divider_counter[0] ),
    .ZN(_046_));
 NOR2_X4 _358_ (.A1(_045_),
    .A2(_046_),
    .ZN(_047_));
 CLKBUF_X3 _359_ (.A(net46),
    .Z(_048_));
 BUF_X4 _360_ (.A(_048_),
    .Z(_049_));
 BUF_X4 _361_ (.A(net45),
    .Z(_050_));
 CLKBUF_X3 _362_ (.A(net47),
    .Z(_051_));
 BUF_X4 _363_ (.A(_051_),
    .Z(_052_));
 NOR3_X4 _364_ (.A1(_049_),
    .A2(_050_),
    .A3(_052_),
    .ZN(_053_));
 CLKBUF_X3 _365_ (.A(net48),
    .Z(_054_));
 INV_X2 _366_ (.A(_054_),
    .ZN(_055_));
 BUF_X4 _367_ (.A(_055_),
    .Z(_056_));
 BUF_X2 _368_ (.A(rst_n),
    .Z(_057_));
 INV_X2 _369_ (.A(_057_),
    .ZN(_058_));
 NOR2_X1 _370_ (.A1(_056_),
    .A2(_058_),
    .ZN(_059_));
 AND4_X1 _371_ (.A1(_042_),
    .A2(_047_),
    .A3(_053_),
    .A4(_059_),
    .ZN(_024_));
 BUF_X2 _372_ (.A(_057_),
    .Z(_060_));
 NAND2_X1 _373_ (.A1(net19),
    .A2(_060_),
    .ZN(_061_));
 CLKBUF_X3 _374_ (.A(_049_),
    .Z(_062_));
 INV_X2 _375_ (.A(_050_),
    .ZN(_063_));
 INV_X2 _376_ (.A(_051_),
    .ZN(_064_));
 NAND2_X1 _377_ (.A1(_063_),
    .A2(_064_),
    .ZN(_065_));
 BUF_X4 _378_ (.A(_050_),
    .Z(_066_));
 CLKBUF_X3 _379_ (.A(_052_),
    .Z(_067_));
 BUF_X2 _380_ (.A(_342_),
    .Z(_068_));
 NAND3_X1 _381_ (.A1(_066_),
    .A2(_067_),
    .A3(_068_),
    .ZN(_069_));
 AOI21_X1 _382_ (.A(_062_),
    .B1(_065_),
    .B2(_069_),
    .ZN(_070_));
 NOR4_X4 _383_ (.A1(_048_),
    .A2(net45),
    .A3(_051_),
    .A4(net17),
    .ZN(_071_));
 NOR4_X2 _384_ (.A1(_054_),
    .A2(_045_),
    .A3(_046_),
    .A4(_071_),
    .ZN(_072_));
 AOI21_X1 _385_ (.A(_061_),
    .B1(_070_),
    .B2(_072_),
    .ZN(_002_));
 CLKBUF_X3 _386_ (.A(_058_),
    .Z(_073_));
 CLKBUF_X2 _387_ (.A(net20),
    .Z(_074_));
 NAND2_X1 _388_ (.A1(_050_),
    .A2(_064_),
    .ZN(_075_));
 MUX2_X1 _389_ (.A(_068_),
    .B(_041_),
    .S(_048_),
    .Z(_076_));
 INV_X2 _390_ (.A(_048_),
    .ZN(_077_));
 NAND4_X2 _391_ (.A1(_077_),
    .A2(_050_),
    .A3(_055_),
    .A4(_052_),
    .ZN(_078_));
 INV_X1 _392_ (.A(_041_),
    .ZN(_079_));
 INV_X1 _393_ (.A(cmd_write),
    .ZN(_080_));
 BUF_X1 _394_ (.A(stop),
    .Z(_081_));
 NOR3_X1 _395_ (.A1(_079_),
    .A2(_080_),
    .A3(_081_),
    .ZN(_082_));
 OAI221_X2 _396_ (.A(_072_),
    .B1(_075_),
    .B2(_076_),
    .C1(_078_),
    .C2(_082_),
    .ZN(_083_));
 AND2_X1 _397_ (.A1(_048_),
    .A2(net45),
    .ZN(_084_));
 NOR2_X4 _398_ (.A1(_054_),
    .A2(_051_),
    .ZN(_085_));
 NAND4_X2 _399_ (.A1(_041_),
    .A2(net19),
    .A3(_084_),
    .A4(_085_),
    .ZN(_086_));
 NAND3_X2 _400_ (.A1(_055_),
    .A2(_052_),
    .A3(_084_),
    .ZN(_087_));
 INV_X1 _401_ (.A(_081_),
    .ZN(_088_));
 CLKBUF_X2 _402_ (.A(cmd_read),
    .Z(_089_));
 AND2_X1 _403_ (.A1(_088_),
    .A2(_089_),
    .ZN(_090_));
 NOR2_X1 _404_ (.A1(_050_),
    .A2(_054_),
    .ZN(_091_));
 OAI21_X2 _405_ (.A(_091_),
    .B1(_052_),
    .B2(_049_),
    .ZN(_092_));
 CLKBUF_X2 _406_ (.A(net21),
    .Z(_093_));
 BUF_X1 _407_ (.A(net22),
    .Z(_094_));
 NOR2_X2 _408_ (.A1(_093_),
    .A2(_094_),
    .ZN(_095_));
 NAND2_X2 _409_ (.A1(_330_),
    .A2(_095_),
    .ZN(_096_));
 OAI221_X2 _410_ (.A(_086_),
    .B1(_087_),
    .B2(_090_),
    .C1(_092_),
    .C2(_096_),
    .ZN(_097_));
 CLKBUF_X3 _411_ (.A(_054_),
    .Z(_098_));
 NAND2_X1 _412_ (.A1(_063_),
    .A2(_067_),
    .ZN(_099_));
 OAI21_X1 _413_ (.A(_049_),
    .B1(_063_),
    .B2(_067_),
    .ZN(_100_));
 AOI21_X2 _414_ (.A(_098_),
    .B1(_099_),
    .B2(_100_),
    .ZN(_101_));
 BUF_X4 _415_ (.A(_079_),
    .Z(_102_));
 AOI211_X2 _416_ (.A(_083_),
    .B(_097_),
    .C1(_101_),
    .C2(_102_),
    .ZN(_103_));
 NOR3_X1 _417_ (.A1(_073_),
    .A2(_074_),
    .A3(_103_),
    .ZN(_104_));
 NOR3_X1 _418_ (.A1(_330_),
    .A2(_073_),
    .A3(_092_),
    .ZN(_105_));
 AOI21_X1 _419_ (.A(_104_),
    .B1(_105_),
    .B2(_103_),
    .ZN(_003_));
 BUF_X2 _420_ (.A(_057_),
    .Z(_106_));
 NOR2_X1 _421_ (.A1(_093_),
    .A2(_103_),
    .ZN(_107_));
 NOR2_X1 _422_ (.A1(_049_),
    .A2(_052_),
    .ZN(_108_));
 NOR3_X1 _423_ (.A1(_066_),
    .A2(_098_),
    .A3(_108_),
    .ZN(_109_));
 AND3_X1 _424_ (.A1(_333_),
    .A2(_109_),
    .A3(_103_),
    .ZN(_110_));
 OAI21_X1 _425_ (.A(_106_),
    .B1(_107_),
    .B2(_110_),
    .ZN(_004_));
 OR2_X1 _426_ (.A1(_332_),
    .A2(_092_),
    .ZN(_111_));
 AOI21_X1 _427_ (.A(_094_),
    .B1(_103_),
    .B2(_111_),
    .ZN(_112_));
 AND4_X1 _428_ (.A1(_094_),
    .A2(_332_),
    .A3(_109_),
    .A4(_103_),
    .ZN(_113_));
 OAI21_X1 _429_ (.A(_106_),
    .B1(_112_),
    .B2(_113_),
    .ZN(_005_));
 OAI21_X1 _430_ (.A(_057_),
    .B1(net23),
    .B2(_047_),
    .ZN(_114_));
 NOR2_X1 _431_ (.A1(_098_),
    .A2(_071_),
    .ZN(_115_));
 NOR2_X1 _432_ (.A1(_056_),
    .A2(_042_),
    .ZN(_116_));
 AOI21_X1 _433_ (.A(_115_),
    .B1(_116_),
    .B2(_053_),
    .ZN(_117_));
 AOI21_X1 _434_ (.A(_114_),
    .B1(_117_),
    .B2(_047_),
    .ZN(_006_));
 NOR2_X2 _435_ (.A1(_062_),
    .A2(_066_),
    .ZN(_118_));
 NAND4_X2 _436_ (.A1(net17),
    .A2(_047_),
    .A3(_118_),
    .A4(_085_),
    .ZN(_119_));
 MUX2_X1 _437_ (.A(net16),
    .B(_089_),
    .S(_119_),
    .Z(_120_));
 AND2_X1 _438_ (.A1(_106_),
    .A2(_120_),
    .ZN(_007_));
 MUX2_X1 _439_ (.A(net18),
    .B(cmd_write),
    .S(_119_),
    .Z(_121_));
 AND2_X1 _440_ (.A1(_106_),
    .A2(_121_),
    .ZN(_008_));
 OR2_X1 _441_ (.A1(_045_),
    .A2(_046_),
    .ZN(_122_));
 CLKBUF_X3 _442_ (.A(_122_),
    .Z(_123_));
 NAND4_X4 _443_ (.A1(_049_),
    .A2(_063_),
    .A3(_055_),
    .A4(_052_),
    .ZN(_124_));
 NOR4_X4 _444_ (.A1(_102_),
    .A2(_123_),
    .A3(_096_),
    .A4(_124_),
    .ZN(_125_));
 MUX2_X1 _445_ (.A(net24),
    .B(net37),
    .S(_125_),
    .Z(_126_));
 AND2_X1 _446_ (.A1(_060_),
    .A2(_126_),
    .ZN(_009_));
 BUF_X2 _447_ (.A(net38),
    .Z(_127_));
 MUX2_X1 _448_ (.A(net25),
    .B(_127_),
    .S(_125_),
    .Z(_128_));
 AND2_X1 _449_ (.A1(_060_),
    .A2(_128_),
    .ZN(_010_));
 MUX2_X1 _450_ (.A(net26),
    .B(net39),
    .S(_125_),
    .Z(_129_));
 AND2_X1 _451_ (.A1(_060_),
    .A2(_129_),
    .ZN(_011_));
 BUF_X2 _452_ (.A(net40),
    .Z(_130_));
 MUX2_X1 _453_ (.A(net27),
    .B(_130_),
    .S(_125_),
    .Z(_131_));
 AND2_X1 _454_ (.A1(_060_),
    .A2(_131_),
    .ZN(_012_));
 MUX2_X1 _455_ (.A(net28),
    .B(net41),
    .S(_125_),
    .Z(_132_));
 AND2_X1 _456_ (.A1(_060_),
    .A2(_132_),
    .ZN(_013_));
 BUF_X2 _457_ (.A(net42),
    .Z(_133_));
 MUX2_X1 _458_ (.A(net29),
    .B(_133_),
    .S(_125_),
    .Z(_134_));
 AND2_X1 _459_ (.A1(_060_),
    .A2(_134_),
    .ZN(_014_));
 MUX2_X1 _460_ (.A(net30),
    .B(net43),
    .S(_125_),
    .Z(_135_));
 AND2_X1 _461_ (.A1(_060_),
    .A2(_135_),
    .ZN(_015_));
 BUF_X2 _462_ (.A(net44),
    .Z(_136_));
 MUX2_X1 _463_ (.A(net31),
    .B(_136_),
    .S(_125_),
    .Z(_137_));
 AND2_X1 _464_ (.A1(_060_),
    .A2(_137_),
    .ZN(_016_));
 AND3_X1 _465_ (.A1(_060_),
    .A2(_001_),
    .A3(_123_),
    .ZN(_017_));
 NOR3_X1 _466_ (.A1(_073_),
    .A2(_350_),
    .A3(_047_),
    .ZN(_018_));
 XNOR2_X1 _467_ (.A(_044_),
    .B(_349_),
    .ZN(_138_));
 NAND3_X1 _468_ (.A1(_106_),
    .A2(_123_),
    .A3(_138_),
    .ZN(_019_));
 OR2_X1 _469_ (.A1(\divider_counter[1] ),
    .A2(\divider_counter[0] ),
    .ZN(_139_));
 NOR2_X1 _470_ (.A1(_044_),
    .A2(_139_),
    .ZN(_140_));
 XNOR2_X1 _471_ (.A(_043_),
    .B(_140_),
    .ZN(_141_));
 NAND2_X1 _472_ (.A1(_106_),
    .A2(_141_),
    .ZN(_020_));
 INV_X1 _473_ (.A(_349_),
    .ZN(_142_));
 NOR3_X1 _474_ (.A1(_043_),
    .A2(_044_),
    .A3(_142_),
    .ZN(_143_));
 XNOR2_X1 _475_ (.A(\divider_counter[4] ),
    .B(_143_),
    .ZN(_144_));
 NAND3_X1 _476_ (.A1(_106_),
    .A2(_123_),
    .A3(_144_),
    .ZN(_021_));
 NOR4_X1 _477_ (.A1(\divider_counter[4] ),
    .A2(_043_),
    .A3(_044_),
    .A4(_139_),
    .ZN(_145_));
 XNOR2_X1 _478_ (.A(\divider_counter[5] ),
    .B(_145_),
    .ZN(_146_));
 NAND2_X1 _479_ (.A1(_106_),
    .A2(_146_),
    .ZN(_022_));
 AOI21_X1 _480_ (.A(_045_),
    .B1(_139_),
    .B2(_142_),
    .ZN(_147_));
 NAND2_X1 _481_ (.A1(\divider_counter[6] ),
    .A2(_349_),
    .ZN(_148_));
 OAI22_X1 _482_ (.A1(\divider_counter[6] ),
    .A2(_147_),
    .B1(_148_),
    .B2(_045_),
    .ZN(_149_));
 NAND2_X1 _483_ (.A1(_106_),
    .A2(_149_),
    .ZN(_023_));
 NOR2_X1 _484_ (.A1(net33),
    .A2(_047_),
    .ZN(_150_));
 NOR3_X1 _485_ (.A1(_340_),
    .A2(_068_),
    .A3(_123_),
    .ZN(_151_));
 NOR3_X1 _486_ (.A1(_073_),
    .A2(_150_),
    .A3(_151_),
    .ZN(_025_));
 NAND2_X1 _487_ (.A1(_341_),
    .A2(_047_),
    .ZN(_152_));
 NAND2_X1 _488_ (.A1(net34),
    .A2(_123_),
    .ZN(_153_));
 AOI21_X1 _489_ (.A(_073_),
    .B1(_152_),
    .B2(_153_),
    .ZN(_026_));
 NAND2_X1 _490_ (.A1(net35),
    .A2(_123_),
    .ZN(_154_));
 NAND3_X1 _491_ (.A1(_098_),
    .A2(_340_),
    .A3(_053_),
    .ZN(_155_));
 OR3_X1 _492_ (.A1(_098_),
    .A2(_341_),
    .A3(_053_),
    .ZN(_156_));
 NAND3_X1 _493_ (.A1(_047_),
    .A2(_155_),
    .A3(_156_),
    .ZN(_157_));
 NAND3_X1 _494_ (.A1(_106_),
    .A2(_154_),
    .A3(_157_),
    .ZN(_027_));
 INV_X1 _495_ (.A(net36),
    .ZN(_158_));
 NAND2_X1 _496_ (.A1(_057_),
    .A2(_158_),
    .ZN(_159_));
 NAND4_X1 _497_ (.A1(_062_),
    .A2(_056_),
    .A3(_067_),
    .A4(_081_),
    .ZN(_160_));
 AOI21_X1 _498_ (.A(_160_),
    .B1(_042_),
    .B2(_066_),
    .ZN(_161_));
 XNOR2_X2 _499_ (.A(_048_),
    .B(_052_),
    .ZN(_162_));
 OR4_X1 _500_ (.A1(_050_),
    .A2(_098_),
    .A3(_102_),
    .A4(_162_),
    .ZN(_163_));
 AOI21_X1 _501_ (.A(_163_),
    .B1(_096_),
    .B2(_158_),
    .ZN(_164_));
 NOR2_X1 _502_ (.A1(_042_),
    .A2(_068_),
    .ZN(_165_));
 NAND4_X1 _503_ (.A1(_077_),
    .A2(_066_),
    .A3(_085_),
    .A4(_165_),
    .ZN(_166_));
 NOR2_X1 _504_ (.A1(_089_),
    .A2(_136_),
    .ZN(_167_));
 NAND2_X1 _505_ (.A1(_084_),
    .A2(_085_),
    .ZN(_168_));
 NAND3_X1 _506_ (.A1(cmd_write),
    .A2(_088_),
    .A3(net15),
    .ZN(_169_));
 OAI221_X1 _507_ (.A(_166_),
    .B1(_167_),
    .B2(_168_),
    .C1(_169_),
    .C2(_078_),
    .ZN(_170_));
 NOR4_X1 _508_ (.A1(_058_),
    .A2(_161_),
    .A3(_164_),
    .A4(_170_),
    .ZN(_171_));
 NAND2_X1 _509_ (.A1(_088_),
    .A2(_089_),
    .ZN(_172_));
 OAI21_X1 _510_ (.A(_042_),
    .B1(_172_),
    .B2(_087_),
    .ZN(_173_));
 CLKBUF_X3 _511_ (.A(_124_),
    .Z(_174_));
 NAND3_X1 _512_ (.A1(_102_),
    .A2(_168_),
    .A3(_174_),
    .ZN(_175_));
 NAND2_X1 _513_ (.A1(_173_),
    .A2(_175_),
    .ZN(_176_));
 INV_X1 _514_ (.A(_136_),
    .ZN(_177_));
 XOR2_X1 _515_ (.A(_066_),
    .B(_067_),
    .Z(_178_));
 OAI221_X1 _516_ (.A(_056_),
    .B1(_177_),
    .B2(_065_),
    .C1(_178_),
    .C2(_062_),
    .ZN(_179_));
 NOR3_X1 _517_ (.A1(_098_),
    .A2(_102_),
    .A3(_053_),
    .ZN(_180_));
 NOR3_X1 _518_ (.A1(_056_),
    .A2(_042_),
    .A3(_068_),
    .ZN(_181_));
 AOI21_X1 _519_ (.A(_180_),
    .B1(_181_),
    .B2(_053_),
    .ZN(_182_));
 AND4_X1 _520_ (.A1(_056_),
    .A2(_067_),
    .A3(_102_),
    .A4(_118_),
    .ZN(_183_));
 MUX2_X1 _521_ (.A(net37),
    .B(_127_),
    .S(_074_),
    .Z(_184_));
 MUX2_X1 _522_ (.A(net39),
    .B(_130_),
    .S(_074_),
    .Z(_185_));
 MUX2_X1 _523_ (.A(_184_),
    .B(_185_),
    .S(_093_),
    .Z(_186_));
 MUX2_X1 _524_ (.A(net41),
    .B(_133_),
    .S(_074_),
    .Z(_187_));
 MUX2_X1 _525_ (.A(net43),
    .B(_136_),
    .S(_074_),
    .Z(_188_));
 MUX2_X1 _526_ (.A(_187_),
    .B(_188_),
    .S(_093_),
    .Z(_189_));
 MUX2_X1 _527_ (.A(_186_),
    .B(_189_),
    .S(_094_),
    .Z(_190_));
 AOI22_X1 _528_ (.A1(_179_),
    .A2(_182_),
    .B1(_183_),
    .B2(_190_),
    .ZN(_191_));
 NAND3_X1 _529_ (.A1(_171_),
    .A2(_176_),
    .A3(_191_),
    .ZN(_192_));
 INV_X1 _530_ (.A(_330_),
    .ZN(_193_));
 OR2_X1 _531_ (.A1(_093_),
    .A2(_094_),
    .ZN(_194_));
 OAI21_X1 _532_ (.A(_042_),
    .B1(_193_),
    .B2(_194_),
    .ZN(_195_));
 OAI21_X1 _533_ (.A(_086_),
    .B1(_124_),
    .B2(_195_),
    .ZN(_196_));
 OR2_X2 _534_ (.A1(_123_),
    .A2(_196_),
    .ZN(_197_));
 NOR2_X1 _535_ (.A1(_042_),
    .A2(_340_),
    .ZN(_198_));
 OAI21_X1 _536_ (.A(_078_),
    .B1(_168_),
    .B2(_344_),
    .ZN(_199_));
 AOI221_X2 _537_ (.A(_197_),
    .B1(_198_),
    .B2(_199_),
    .C1(_101_),
    .C2(_341_),
    .ZN(_200_));
 MUX2_X1 _538_ (.A(_159_),
    .B(_192_),
    .S(_200_),
    .Z(_028_));
 NAND2_X1 _539_ (.A1(_049_),
    .A2(_050_),
    .ZN(_201_));
 OR2_X2 _540_ (.A1(_054_),
    .A2(_051_),
    .ZN(_202_));
 OAI21_X1 _541_ (.A(_041_),
    .B1(net19),
    .B2(_089_),
    .ZN(_203_));
 OR3_X1 _542_ (.A1(_201_),
    .A2(_202_),
    .A3(_203_),
    .ZN(_204_));
 AND3_X1 _543_ (.A1(_049_),
    .A2(_063_),
    .A3(_068_),
    .ZN(_205_));
 OAI21_X1 _544_ (.A(_052_),
    .B1(_063_),
    .B2(_049_),
    .ZN(_206_));
 NAND3_X1 _545_ (.A1(_062_),
    .A2(_063_),
    .A3(_085_),
    .ZN(_207_));
 AOI21_X1 _546_ (.A(_102_),
    .B1(_330_),
    .B2(_095_),
    .ZN(_208_));
 OAI221_X2 _547_ (.A(_204_),
    .B1(_205_),
    .B2(_206_),
    .C1(_207_),
    .C2(_208_),
    .ZN(_209_));
 NOR2_X2 _548_ (.A1(_083_),
    .A2(_209_),
    .ZN(_210_));
 OAI21_X1 _549_ (.A(net16),
    .B1(_118_),
    .B2(_098_),
    .ZN(_211_));
 AOI221_X1 _550_ (.A(_077_),
    .B1(_067_),
    .B2(net16),
    .C1(_085_),
    .C2(net8),
    .ZN(_212_));
 OR2_X1 _551_ (.A1(_063_),
    .A2(_212_),
    .ZN(_213_));
 MUX2_X1 _552_ (.A(_089_),
    .B(net8),
    .S(_067_),
    .Z(_214_));
 AOI21_X1 _553_ (.A(_062_),
    .B1(_056_),
    .B2(_214_),
    .ZN(_215_));
 OAI21_X1 _554_ (.A(_211_),
    .B1(_213_),
    .B2(_215_),
    .ZN(_216_));
 NAND2_X1 _555_ (.A1(_210_),
    .A2(_216_),
    .ZN(_217_));
 OR2_X1 _556_ (.A1(_083_),
    .A2(_209_),
    .ZN(_218_));
 BUF_X2 _557_ (.A(_218_),
    .Z(_219_));
 XOR2_X2 _558_ (.A(_332_),
    .B(_000_),
    .Z(_220_));
 NOR3_X1 _559_ (.A1(_333_),
    .A2(_096_),
    .A3(_220_),
    .ZN(_221_));
 NOR2_X1 _560_ (.A1(_174_),
    .A2(_221_),
    .ZN(_222_));
 OAI21_X1 _561_ (.A(net37),
    .B1(_219_),
    .B2(_222_),
    .ZN(_223_));
 AOI21_X1 _562_ (.A(_073_),
    .B1(_217_),
    .B2(_223_),
    .ZN(_029_));
 NAND2_X1 _563_ (.A1(_050_),
    .A2(_067_),
    .ZN(_224_));
 XNOR2_X2 _564_ (.A(_062_),
    .B(_224_),
    .ZN(_225_));
 NAND2_X4 _565_ (.A1(_056_),
    .A2(_225_),
    .ZN(_226_));
 NAND2_X1 _566_ (.A1(net1),
    .A2(_226_),
    .ZN(_227_));
 NOR3_X4 _567_ (.A1(_077_),
    .A2(_066_),
    .A3(_202_),
    .ZN(_228_));
 AOI21_X1 _568_ (.A(_174_),
    .B1(_220_),
    .B2(_334_),
    .ZN(_229_));
 NAND2_X2 _569_ (.A1(_050_),
    .A2(_056_),
    .ZN(_230_));
 NOR2_X4 _570_ (.A1(_162_),
    .A2(_230_),
    .ZN(_231_));
 AOI222_X2 _571_ (.A1(net37),
    .A2(_228_),
    .B1(_229_),
    .B2(_127_),
    .C1(_231_),
    .C2(net9),
    .ZN(_232_));
 NAND3_X1 _572_ (.A1(_210_),
    .A2(_227_),
    .A3(_232_),
    .ZN(_233_));
 INV_X1 _573_ (.A(_127_),
    .ZN(_234_));
 AOI21_X1 _574_ (.A(_073_),
    .B1(_234_),
    .B2(_219_),
    .ZN(_235_));
 AND2_X1 _575_ (.A1(_233_),
    .A2(_235_),
    .ZN(_030_));
 AOI222_X2 _576_ (.A1(_127_),
    .A2(_228_),
    .B1(_226_),
    .B2(net2),
    .C1(_231_),
    .C2(net10),
    .ZN(_236_));
 OR2_X1 _577_ (.A1(_219_),
    .A2(_236_),
    .ZN(_237_));
 NOR2_X1 _578_ (.A1(_193_),
    .A2(_095_),
    .ZN(_238_));
 AND2_X1 _579_ (.A1(_333_),
    .A2(_238_),
    .ZN(_239_));
 AOI21_X1 _580_ (.A(_174_),
    .B1(_220_),
    .B2(_239_),
    .ZN(_240_));
 OAI21_X1 _581_ (.A(net39),
    .B1(_219_),
    .B2(_240_),
    .ZN(_241_));
 AOI21_X1 _582_ (.A(_073_),
    .B1(_237_),
    .B2(_241_),
    .ZN(_031_));
 NAND2_X1 _583_ (.A1(net3),
    .A2(_226_),
    .ZN(_242_));
 AOI21_X1 _584_ (.A(_174_),
    .B1(_220_),
    .B2(_336_),
    .ZN(_243_));
 AOI222_X2 _585_ (.A1(net39),
    .A2(_228_),
    .B1(_231_),
    .B2(net11),
    .C1(_243_),
    .C2(_130_),
    .ZN(_244_));
 NAND3_X1 _586_ (.A1(_210_),
    .A2(_242_),
    .A3(_244_),
    .ZN(_245_));
 INV_X1 _587_ (.A(_130_),
    .ZN(_246_));
 AOI21_X1 _588_ (.A(_058_),
    .B1(_246_),
    .B2(_219_),
    .ZN(_247_));
 AND2_X1 _589_ (.A1(_245_),
    .A2(_247_),
    .ZN(_032_));
 AOI222_X2 _590_ (.A1(_130_),
    .A2(_228_),
    .B1(_226_),
    .B2(net4),
    .C1(_231_),
    .C2(net12),
    .ZN(_248_));
 OR2_X1 _591_ (.A1(_219_),
    .A2(_248_),
    .ZN(_249_));
 XNOR2_X2 _592_ (.A(_332_),
    .B(_000_),
    .ZN(_250_));
 NOR2_X1 _593_ (.A1(_333_),
    .A2(_250_),
    .ZN(_251_));
 AOI21_X1 _594_ (.A(_174_),
    .B1(_238_),
    .B2(_251_),
    .ZN(_252_));
 OAI21_X1 _595_ (.A(net41),
    .B1(_219_),
    .B2(_252_),
    .ZN(_253_));
 AOI21_X1 _596_ (.A(_073_),
    .B1(_249_),
    .B2(_253_),
    .ZN(_033_));
 NAND2_X1 _597_ (.A1(net5),
    .A2(_226_),
    .ZN(_254_));
 AOI21_X1 _598_ (.A(_174_),
    .B1(_250_),
    .B2(_334_),
    .ZN(_255_));
 AOI222_X2 _599_ (.A1(net41),
    .A2(_228_),
    .B1(_231_),
    .B2(net13),
    .C1(_255_),
    .C2(_133_),
    .ZN(_256_));
 NAND3_X1 _600_ (.A1(_210_),
    .A2(_254_),
    .A3(_256_),
    .ZN(_257_));
 INV_X1 _601_ (.A(_133_),
    .ZN(_258_));
 AOI21_X1 _602_ (.A(_058_),
    .B1(_258_),
    .B2(_219_),
    .ZN(_259_));
 AND2_X1 _603_ (.A1(_257_),
    .A2(_259_),
    .ZN(_034_));
 AOI222_X2 _604_ (.A1(_133_),
    .A2(_228_),
    .B1(_226_),
    .B2(net6),
    .C1(_231_),
    .C2(net14),
    .ZN(_260_));
 OR2_X1 _605_ (.A1(_218_),
    .A2(_260_),
    .ZN(_261_));
 AOI21_X1 _606_ (.A(_174_),
    .B1(_250_),
    .B2(_239_),
    .ZN(_262_));
 OAI21_X1 _607_ (.A(net43),
    .B1(_219_),
    .B2(_262_),
    .ZN(_263_));
 AOI21_X1 _608_ (.A(_073_),
    .B1(_261_),
    .B2(_263_),
    .ZN(_035_));
 NAND2_X1 _609_ (.A1(net7),
    .A2(_226_),
    .ZN(_264_));
 AOI21_X1 _610_ (.A(_174_),
    .B1(_250_),
    .B2(_336_),
    .ZN(_265_));
 AOI222_X2 _611_ (.A1(net43),
    .A2(_228_),
    .B1(_231_),
    .B2(net15),
    .C1(_265_),
    .C2(_136_),
    .ZN(_266_));
 NAND3_X1 _612_ (.A1(_210_),
    .A2(_264_),
    .A3(_266_),
    .ZN(_267_));
 AOI21_X1 _613_ (.A(_058_),
    .B1(_177_),
    .B2(_219_),
    .ZN(_268_));
 AND2_X1 _614_ (.A1(_267_),
    .A2(_268_),
    .ZN(_036_));
 NOR2_X1 _615_ (.A1(_063_),
    .A2(_058_),
    .ZN(_269_));
 AND2_X1 _616_ (.A1(_057_),
    .A2(_091_),
    .ZN(_270_));
 NAND2_X1 _617_ (.A1(_108_),
    .A2(_116_),
    .ZN(_271_));
 AND3_X1 _618_ (.A1(_049_),
    .A2(_052_),
    .A3(_041_),
    .ZN(_272_));
 NOR3_X1 _619_ (.A1(_098_),
    .A2(_108_),
    .A3(_272_),
    .ZN(_273_));
 OAI21_X1 _620_ (.A(_273_),
    .B1(_096_),
    .B2(_102_),
    .ZN(_274_));
 AOI21_X2 _621_ (.A(_066_),
    .B1(_271_),
    .B2(_274_),
    .ZN(_275_));
 NAND3_X1 _622_ (.A1(_062_),
    .A2(_064_),
    .A3(_068_),
    .ZN(_276_));
 AOI21_X2 _623_ (.A(_230_),
    .B1(_276_),
    .B2(_042_),
    .ZN(_277_));
 NOR4_X2 _624_ (.A1(_062_),
    .A2(_066_),
    .A3(net17),
    .A4(_202_),
    .ZN(_278_));
 NOR4_X4 _625_ (.A1(_197_),
    .A2(_275_),
    .A3(_277_),
    .A4(_278_),
    .ZN(_279_));
 MUX2_X1 _626_ (.A(_269_),
    .B(_270_),
    .S(_279_),
    .Z(_037_));
 NOR2_X1 _627_ (.A1(_077_),
    .A2(_058_),
    .ZN(_280_));
 OAI21_X1 _628_ (.A(_084_),
    .B1(_172_),
    .B2(_064_),
    .ZN(_281_));
 NAND2_X1 _629_ (.A1(_077_),
    .A2(_075_),
    .ZN(_282_));
 NAND3_X1 _630_ (.A1(_056_),
    .A2(_281_),
    .A3(_282_),
    .ZN(_283_));
 NOR2_X1 _631_ (.A1(_201_),
    .A2(_202_),
    .ZN(_284_));
 NAND3_X1 _632_ (.A1(_042_),
    .A2(_089_),
    .A3(_284_),
    .ZN(_285_));
 AOI21_X1 _633_ (.A(_058_),
    .B1(_283_),
    .B2(_285_),
    .ZN(_286_));
 MUX2_X1 _634_ (.A(_280_),
    .B(_286_),
    .S(_279_),
    .Z(_038_));
 NOR2_X1 _635_ (.A1(_064_),
    .A2(_058_),
    .ZN(_287_));
 NOR3_X1 _636_ (.A1(_067_),
    .A2(_102_),
    .A3(_201_),
    .ZN(_288_));
 OAI21_X1 _637_ (.A(_066_),
    .B1(_080_),
    .B2(_081_),
    .ZN(_289_));
 NOR2_X1 _638_ (.A1(_062_),
    .A2(_064_),
    .ZN(_290_));
 AOI21_X1 _639_ (.A(_288_),
    .B1(_289_),
    .B2(_290_),
    .ZN(_291_));
 OAI221_X1 _640_ (.A(_174_),
    .B1(_291_),
    .B2(_098_),
    .C1(_172_),
    .C2(_087_),
    .ZN(_292_));
 AND2_X1 _641_ (.A1(_057_),
    .A2(_292_),
    .ZN(_293_));
 MUX2_X1 _642_ (.A(_287_),
    .B(_293_),
    .S(_279_),
    .Z(_039_));
 NAND2_X1 _643_ (.A1(_102_),
    .A2(_284_),
    .ZN(_294_));
 NOR2_X1 _644_ (.A1(_080_),
    .A2(_081_),
    .ZN(_295_));
 OAI221_X1 _645_ (.A(_294_),
    .B1(_087_),
    .B2(_090_),
    .C1(_078_),
    .C2(_295_),
    .ZN(_296_));
 AND2_X1 _646_ (.A1(_057_),
    .A2(_296_),
    .ZN(_297_));
 MUX2_X1 _647_ (.A(_059_),
    .B(_297_),
    .S(_279_),
    .Z(_040_));
 HA_X1 _648_ (.A(_330_),
    .B(_331_),
    .CO(_332_),
    .S(_333_));
 HA_X1 _649_ (.A(net20),
    .B(_331_),
    .CO(_334_),
    .S(_335_));
 HA_X1 _650_ (.A(net20),
    .B(net21),
    .CO(_336_),
    .S(_337_));
 HA_X1 _651_ (.A(_338_),
    .B(_339_),
    .CO(_340_),
    .S(_341_));
 HA_X1 _652_ (.A(_338_),
    .B(net34),
    .CO(_342_),
    .S(_343_));
 HA_X1 _653_ (.A(net33),
    .B(_339_),
    .CO(_344_),
    .S(_345_));
 HA_X1 _654_ (.A(net33),
    .B(net34),
    .CO(_346_),
    .S(_347_));
 HA_X1 _655_ (.A(_001_),
    .B(_348_),
    .CO(_349_),
    .S(_350_));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 BUF_X1 _657_ (.A(net49),
    .Z(scl));
 BUF_X1 _658_ (.A(net50),
    .Z(sda));
 DFF_X2 \ack_error$_SDFFE_PN0P_  (.D(_002_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net19),
    .QN(_329_));
 DFF_X2 \bit_counter_debug[0]$_SDFFE_PN1P_  (.D(_003_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net20),
    .QN(_330_));
 DFF_X1 \bit_counter_debug[1]$_SDFFE_PN1P_  (.D(_004_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net21),
    .QN(_331_));
 DFF_X2 \bit_counter_debug[2]$_SDFFE_PN1P_  (.D(_005_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net22),
    .QN(_000_));
 DFF_X1 \busy$_SDFFE_PN0N_  (.D(_006_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net23),
    .QN(_328_));
 DFF_X1 \cmd_read$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_2_0__leaf_clk),
    .Q(cmd_read),
    .QN(_327_));
 DFF_X1 \cmd_write$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_2_0__leaf_clk),
    .Q(cmd_write),
    .QN(_326_));
 DFF_X1 \data_out[0]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net24),
    .QN(_325_));
 DFF_X1 \data_out[1]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net25),
    .QN(_324_));
 DFF_X1 \data_out[2]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net26),
    .QN(_323_));
 DFF_X1 \data_out[3]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net27),
    .QN(_322_));
 DFF_X1 \data_out[4]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net28),
    .QN(_321_));
 DFF_X1 \data_out[5]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net29),
    .QN(_320_));
 DFF_X1 \data_out[6]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net30),
    .QN(_319_));
 DFF_X1 \data_out[7]$_SDFFE_PN0P_  (.D(_016_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net31),
    .QN(_318_));
 DFF_X1 \divider_counter[0]$_SDFF_PN0_  (.D(_017_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\divider_counter[0] ),
    .QN(_001_));
 DFF_X1 \divider_counter[1]$_SDFF_PN0_  (.D(_018_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\divider_counter[1] ),
    .QN(_348_));
 DFF_X1 \divider_counter[2]$_SDFF_PN1_  (.D(_019_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\divider_counter[2] ),
    .QN(_317_));
 DFF_X1 \divider_counter[3]$_SDFF_PN1_  (.D(_020_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\divider_counter[3] ),
    .QN(_316_));
 DFF_X1 \divider_counter[4]$_SDFF_PN1_  (.D(_021_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\divider_counter[4] ),
    .QN(_315_));
 DFF_X1 \divider_counter[5]$_SDFF_PN1_  (.D(_022_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\divider_counter[5] ),
    .QN(_314_));
 DFF_X1 \divider_counter[6]$_SDFF_PN1_  (.D(_023_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\divider_counter[6] ),
    .QN(_313_));
 DFF_X1 \done$_SDFF_PP0_  (.D(_024_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net32),
    .QN(_312_));
 DFF_X2 \phase[0]$_SDFFE_PN0N_  (.D(_025_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net33),
    .QN(_338_));
 DFF_X2 \phase[1]$_SDFFE_PN0N_  (.D(_026_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net34),
    .QN(_339_));
 DFF_X1 \scl_internal$_SDFFE_PN1N_  (.D(_027_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net35),
    .QN(_311_));
 DFF_X1 \sda_internal$_SDFFE_PN1P_  (.D(_028_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net36),
    .QN(_310_));
 DFF_X2 \shift_reg_debug[0]$_SDFFE_PN0P_  (.D(_029_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net37),
    .QN(_309_));
 DFF_X1 \shift_reg_debug[1]$_SDFFE_PN0P_  (.D(_030_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net38),
    .QN(_308_));
 DFF_X2 \shift_reg_debug[2]$_SDFFE_PN0P_  (.D(_031_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net39),
    .QN(_307_));
 DFF_X1 \shift_reg_debug[3]$_SDFFE_PN0P_  (.D(_032_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net40),
    .QN(_306_));
 DFF_X2 \shift_reg_debug[4]$_SDFFE_PN0P_  (.D(_033_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net41),
    .QN(_305_));
 DFF_X1 \shift_reg_debug[5]$_SDFFE_PN0P_  (.D(_034_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net42),
    .QN(_304_));
 DFF_X2 \shift_reg_debug[6]$_SDFFE_PN0P_  (.D(_035_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net43),
    .QN(_303_));
 DFF_X1 \shift_reg_debug[7]$_SDFFE_PN0P_  (.D(_036_),
    .CK(clknet_2_3__leaf_clk),
    .Q(net44),
    .QN(_302_));
 DFF_X2 \state[0]$_SDFFE_PN0P_  (.D(_037_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net45),
    .QN(_301_));
 DFF_X1 \state[1]$_SDFFE_PN0P_  (.D(_038_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net46),
    .QN(_300_));
 DFF_X1 \state[2]$_SDFFE_PN0P_  (.D(_039_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net47),
    .QN(_299_));
 DFF_X1 \state[3]$_SDFFE_PN0P_  (.D(_040_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net48),
    .QN(_298_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_63 ();
 BUF_X1 input1 (.A(addr[0]),
    .Z(net1));
 BUF_X1 input2 (.A(addr[1]),
    .Z(net2));
 BUF_X1 input3 (.A(addr[2]),
    .Z(net3));
 BUF_X1 input4 (.A(addr[3]),
    .Z(net4));
 BUF_X1 input5 (.A(addr[4]),
    .Z(net5));
 BUF_X1 input6 (.A(addr[5]),
    .Z(net6));
 BUF_X1 input7 (.A(addr[6]),
    .Z(net7));
 BUF_X1 input8 (.A(data_in[0]),
    .Z(net8));
 BUF_X1 input9 (.A(data_in[1]),
    .Z(net9));
 BUF_X1 input10 (.A(data_in[2]),
    .Z(net10));
 BUF_X1 input11 (.A(data_in[3]),
    .Z(net11));
 BUF_X1 input12 (.A(data_in[4]),
    .Z(net12));
 BUF_X1 input13 (.A(data_in[5]),
    .Z(net13));
 BUF_X1 input14 (.A(data_in[6]),
    .Z(net14));
 BUF_X1 input15 (.A(data_in[7]),
    .Z(net15));
 BUF_X1 input16 (.A(read),
    .Z(net16));
 BUF_X2 input17 (.A(start),
    .Z(net17));
 BUF_X1 input18 (.A(write),
    .Z(net18));
 BUF_X1 output19 (.A(net19),
    .Z(ack_error));
 BUF_X1 output20 (.A(net20),
    .Z(bit_counter_debug[0]));
 BUF_X1 output21 (.A(net21),
    .Z(bit_counter_debug[1]));
 BUF_X1 output22 (.A(net22),
    .Z(bit_counter_debug[2]));
 BUF_X1 output23 (.A(net23),
    .Z(busy));
 BUF_X1 output24 (.A(net24),
    .Z(data_out[0]));
 BUF_X1 output25 (.A(net25),
    .Z(data_out[1]));
 BUF_X1 output26 (.A(net26),
    .Z(data_out[2]));
 BUF_X1 output27 (.A(net27),
    .Z(data_out[3]));
 BUF_X1 output28 (.A(net28),
    .Z(data_out[4]));
 BUF_X1 output29 (.A(net29),
    .Z(data_out[5]));
 BUF_X1 output30 (.A(net30),
    .Z(data_out[6]));
 BUF_X1 output31 (.A(net31),
    .Z(data_out[7]));
 BUF_X1 output32 (.A(net32),
    .Z(done));
 BUF_X1 output33 (.A(net33),
    .Z(phase[0]));
 BUF_X1 output34 (.A(net34),
    .Z(phase[1]));
 BUF_X1 output35 (.A(net35),
    .Z(scl_internal_debug));
 BUF_X1 output36 (.A(net36),
    .Z(sda_internal_debug));
 BUF_X1 output37 (.A(net37),
    .Z(shift_reg_debug[0]));
 BUF_X1 output38 (.A(net38),
    .Z(shift_reg_debug[1]));
 BUF_X1 output39 (.A(net39),
    .Z(shift_reg_debug[2]));
 BUF_X1 output40 (.A(net40),
    .Z(shift_reg_debug[3]));
 BUF_X1 output41 (.A(net41),
    .Z(shift_reg_debug[4]));
 BUF_X1 output42 (.A(net42),
    .Z(shift_reg_debug[5]));
 BUF_X1 output43 (.A(net43),
    .Z(shift_reg_debug[6]));
 BUF_X1 output44 (.A(net44),
    .Z(shift_reg_debug[7]));
 BUF_X1 output45 (.A(net45),
    .Z(state[0]));
 BUF_X1 output46 (.A(net46),
    .Z(state[1]));
 BUF_X1 output47 (.A(net47),
    .Z(state[2]));
 BUF_X1 output48 (.A(net48),
    .Z(state[3]));
 LOGIC0_X1 _657__49 (.Z(net49));
 LOGIC0_X1 _658__50 (.Z(net50));
 CLKBUF_X3 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 CLKBUF_X3 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 CLKBUF_X3 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 INV_X2 clkload0 (.A(clknet_2_1__leaf_clk));
 CLKBUF_X1 clkload1 (.A(clknet_2_2__leaf_clk));
 INV_X2 clkload2 (.A(clknet_2_3__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X8 FILLER_0_97 ();
 FILLCELL_X4 FILLER_0_105 ();
 FILLCELL_X8 FILLER_0_112 ();
 FILLCELL_X4 FILLER_0_120 ();
 FILLCELL_X1 FILLER_0_127 ();
 FILLCELL_X32 FILLER_0_131 ();
 FILLCELL_X8 FILLER_0_163 ();
 FILLCELL_X1 FILLER_0_171 ();
 FILLCELL_X32 FILLER_0_175 ();
 FILLCELL_X32 FILLER_0_207 ();
 FILLCELL_X4 FILLER_0_239 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X8 FILLER_1_97 ();
 FILLCELL_X2 FILLER_1_105 ();
 FILLCELL_X1 FILLER_1_107 ();
 FILLCELL_X32 FILLER_1_111 ();
 FILLCELL_X32 FILLER_1_143 ();
 FILLCELL_X32 FILLER_1_175 ();
 FILLCELL_X32 FILLER_1_207 ();
 FILLCELL_X4 FILLER_1_239 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X16 FILLER_2_225 ();
 FILLCELL_X2 FILLER_2_241 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X16 FILLER_3_225 ();
 FILLCELL_X2 FILLER_3_241 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X16 FILLER_4_225 ();
 FILLCELL_X2 FILLER_4_241 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X16 FILLER_5_225 ();
 FILLCELL_X2 FILLER_5_241 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X8 FILLER_6_33 ();
 FILLCELL_X4 FILLER_6_41 ();
 FILLCELL_X2 FILLER_6_45 ();
 FILLCELL_X16 FILLER_6_82 ();
 FILLCELL_X2 FILLER_6_98 ();
 FILLCELL_X1 FILLER_6_100 ();
 FILLCELL_X1 FILLER_6_118 ();
 FILLCELL_X2 FILLER_6_126 ();
 FILLCELL_X1 FILLER_6_128 ();
 FILLCELL_X32 FILLER_6_158 ();
 FILLCELL_X32 FILLER_6_190 ();
 FILLCELL_X16 FILLER_6_222 ();
 FILLCELL_X4 FILLER_6_238 ();
 FILLCELL_X1 FILLER_6_242 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X16 FILLER_7_33 ();
 FILLCELL_X8 FILLER_7_49 ();
 FILLCELL_X2 FILLER_7_57 ();
 FILLCELL_X8 FILLER_7_94 ();
 FILLCELL_X2 FILLER_7_109 ();
 FILLCELL_X4 FILLER_7_140 ();
 FILLCELL_X1 FILLER_7_144 ();
 FILLCELL_X1 FILLER_7_155 ();
 FILLCELL_X1 FILLER_7_160 ();
 FILLCELL_X8 FILLER_7_178 ();
 FILLCELL_X2 FILLER_7_203 ();
 FILLCELL_X1 FILLER_7_205 ();
 FILLCELL_X32 FILLER_7_209 ();
 FILLCELL_X2 FILLER_7_241 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X8 FILLER_8_33 ();
 FILLCELL_X4 FILLER_8_41 ();
 FILLCELL_X32 FILLER_8_82 ();
 FILLCELL_X8 FILLER_8_114 ();
 FILLCELL_X8 FILLER_8_146 ();
 FILLCELL_X4 FILLER_8_158 ();
 FILLCELL_X2 FILLER_8_162 ();
 FILLCELL_X1 FILLER_8_164 ();
 FILLCELL_X16 FILLER_8_173 ();
 FILLCELL_X8 FILLER_8_189 ();
 FILLCELL_X4 FILLER_8_197 ();
 FILLCELL_X32 FILLER_8_205 ();
 FILLCELL_X4 FILLER_8_237 ();
 FILLCELL_X2 FILLER_8_241 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X4 FILLER_9_33 ();
 FILLCELL_X2 FILLER_9_37 ();
 FILLCELL_X1 FILLER_9_39 ();
 FILLCELL_X1 FILLER_9_57 ();
 FILLCELL_X1 FILLER_9_62 ();
 FILLCELL_X1 FILLER_9_67 ();
 FILLCELL_X2 FILLER_9_74 ();
 FILLCELL_X16 FILLER_9_78 ();
 FILLCELL_X4 FILLER_9_94 ();
 FILLCELL_X2 FILLER_9_98 ();
 FILLCELL_X8 FILLER_9_104 ();
 FILLCELL_X4 FILLER_9_112 ();
 FILLCELL_X1 FILLER_9_116 ();
 FILLCELL_X8 FILLER_9_120 ();
 FILLCELL_X4 FILLER_9_128 ();
 FILLCELL_X2 FILLER_9_132 ();
 FILLCELL_X1 FILLER_9_134 ();
 FILLCELL_X16 FILLER_9_144 ();
 FILLCELL_X8 FILLER_9_160 ();
 FILLCELL_X32 FILLER_9_174 ();
 FILLCELL_X32 FILLER_9_206 ();
 FILLCELL_X4 FILLER_9_238 ();
 FILLCELL_X1 FILLER_9_242 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X2 FILLER_10_68 ();
 FILLCELL_X1 FILLER_10_70 ();
 FILLCELL_X8 FILLER_10_83 ();
 FILLCELL_X2 FILLER_10_91 ();
 FILLCELL_X2 FILLER_10_97 ();
 FILLCELL_X1 FILLER_10_99 ();
 FILLCELL_X2 FILLER_10_114 ();
 FILLCELL_X8 FILLER_10_125 ();
 FILLCELL_X2 FILLER_10_133 ();
 FILLCELL_X1 FILLER_10_135 ();
 FILLCELL_X16 FILLER_10_143 ();
 FILLCELL_X4 FILLER_10_171 ();
 FILLCELL_X8 FILLER_10_222 ();
 FILLCELL_X8 FILLER_10_233 ();
 FILLCELL_X2 FILLER_10_241 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X16 FILLER_11_33 ();
 FILLCELL_X2 FILLER_11_49 ();
 FILLCELL_X1 FILLER_11_51 ();
 FILLCELL_X4 FILLER_11_69 ();
 FILLCELL_X1 FILLER_11_73 ();
 FILLCELL_X8 FILLER_11_84 ();
 FILLCELL_X1 FILLER_11_92 ();
 FILLCELL_X4 FILLER_11_112 ();
 FILLCELL_X2 FILLER_11_116 ();
 FILLCELL_X1 FILLER_11_118 ();
 FILLCELL_X4 FILLER_11_121 ();
 FILLCELL_X2 FILLER_11_125 ();
 FILLCELL_X1 FILLER_11_127 ();
 FILLCELL_X1 FILLER_11_143 ();
 FILLCELL_X1 FILLER_11_150 ();
 FILLCELL_X1 FILLER_11_158 ();
 FILLCELL_X1 FILLER_11_163 ();
 FILLCELL_X1 FILLER_11_180 ();
 FILLCELL_X32 FILLER_11_196 ();
 FILLCELL_X8 FILLER_11_228 ();
 FILLCELL_X4 FILLER_11_236 ();
 FILLCELL_X2 FILLER_11_240 ();
 FILLCELL_X1 FILLER_11_242 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X8 FILLER_12_33 ();
 FILLCELL_X4 FILLER_12_41 ();
 FILLCELL_X2 FILLER_12_45 ();
 FILLCELL_X4 FILLER_12_69 ();
 FILLCELL_X16 FILLER_12_83 ();
 FILLCELL_X1 FILLER_12_104 ();
 FILLCELL_X2 FILLER_12_112 ();
 FILLCELL_X1 FILLER_12_114 ();
 FILLCELL_X2 FILLER_12_188 ();
 FILLCELL_X1 FILLER_12_190 ();
 FILLCELL_X4 FILLER_12_198 ();
 FILLCELL_X2 FILLER_12_202 ();
 FILLCELL_X32 FILLER_12_208 ();
 FILLCELL_X2 FILLER_12_240 ();
 FILLCELL_X1 FILLER_12_242 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X1 FILLER_13_65 ();
 FILLCELL_X16 FILLER_13_87 ();
 FILLCELL_X8 FILLER_13_103 ();
 FILLCELL_X2 FILLER_13_111 ();
 FILLCELL_X1 FILLER_13_113 ();
 FILLCELL_X1 FILLER_13_130 ();
 FILLCELL_X2 FILLER_13_134 ();
 FILLCELL_X8 FILLER_13_192 ();
 FILLCELL_X8 FILLER_13_219 ();
 FILLCELL_X1 FILLER_13_227 ();
 FILLCELL_X8 FILLER_13_231 ();
 FILLCELL_X4 FILLER_13_239 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X16 FILLER_14_97 ();
 FILLCELL_X1 FILLER_14_134 ();
 FILLCELL_X1 FILLER_14_142 ();
 FILLCELL_X1 FILLER_14_146 ();
 FILLCELL_X2 FILLER_14_156 ();
 FILLCELL_X2 FILLER_14_163 ();
 FILLCELL_X4 FILLER_14_193 ();
 FILLCELL_X2 FILLER_14_197 ();
 FILLCELL_X1 FILLER_14_199 ();
 FILLCELL_X2 FILLER_14_217 ();
 FILLCELL_X2 FILLER_14_224 ();
 FILLCELL_X1 FILLER_14_226 ();
 FILLCELL_X8 FILLER_14_230 ();
 FILLCELL_X4 FILLER_14_238 ();
 FILLCELL_X1 FILLER_14_242 ();
 FILLCELL_X4 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_8 ();
 FILLCELL_X16 FILLER_15_40 ();
 FILLCELL_X2 FILLER_15_56 ();
 FILLCELL_X1 FILLER_15_58 ();
 FILLCELL_X16 FILLER_15_66 ();
 FILLCELL_X4 FILLER_15_82 ();
 FILLCELL_X8 FILLER_15_93 ();
 FILLCELL_X2 FILLER_15_101 ();
 FILLCELL_X4 FILLER_15_107 ();
 FILLCELL_X2 FILLER_15_111 ();
 FILLCELL_X1 FILLER_15_113 ();
 FILLCELL_X1 FILLER_15_133 ();
 FILLCELL_X2 FILLER_15_152 ();
 FILLCELL_X2 FILLER_15_161 ();
 FILLCELL_X2 FILLER_15_167 ();
 FILLCELL_X1 FILLER_15_169 ();
 FILLCELL_X2 FILLER_15_177 ();
 FILLCELL_X1 FILLER_15_179 ();
 FILLCELL_X32 FILLER_15_194 ();
 FILLCELL_X16 FILLER_15_226 ();
 FILLCELL_X1 FILLER_15_242 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X16 FILLER_16_33 ();
 FILLCELL_X4 FILLER_16_49 ();
 FILLCELL_X1 FILLER_16_95 ();
 FILLCELL_X4 FILLER_16_153 ();
 FILLCELL_X2 FILLER_16_157 ();
 FILLCELL_X1 FILLER_16_170 ();
 FILLCELL_X4 FILLER_16_178 ();
 FILLCELL_X2 FILLER_16_186 ();
 FILLCELL_X1 FILLER_16_188 ();
 FILLCELL_X32 FILLER_16_192 ();
 FILLCELL_X16 FILLER_16_224 ();
 FILLCELL_X2 FILLER_16_240 ();
 FILLCELL_X1 FILLER_16_242 ();
 FILLCELL_X1 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_5 ();
 FILLCELL_X16 FILLER_17_37 ();
 FILLCELL_X8 FILLER_17_53 ();
 FILLCELL_X2 FILLER_17_61 ();
 FILLCELL_X1 FILLER_17_63 ();
 FILLCELL_X1 FILLER_17_72 ();
 FILLCELL_X32 FILLER_17_80 ();
 FILLCELL_X1 FILLER_17_112 ();
 FILLCELL_X1 FILLER_17_122 ();
 FILLCELL_X1 FILLER_17_126 ();
 FILLCELL_X1 FILLER_17_133 ();
 FILLCELL_X1 FILLER_17_138 ();
 FILLCELL_X2 FILLER_17_142 ();
 FILLCELL_X2 FILLER_17_147 ();
 FILLCELL_X1 FILLER_17_153 ();
 FILLCELL_X2 FILLER_17_168 ();
 FILLCELL_X2 FILLER_17_175 ();
 FILLCELL_X1 FILLER_17_177 ();
 FILLCELL_X2 FILLER_17_188 ();
 FILLCELL_X32 FILLER_17_197 ();
 FILLCELL_X8 FILLER_17_229 ();
 FILLCELL_X4 FILLER_17_237 ();
 FILLCELL_X2 FILLER_17_241 ();
 FILLCELL_X32 FILLER_18_4 ();
 FILLCELL_X16 FILLER_18_36 ();
 FILLCELL_X8 FILLER_18_52 ();
 FILLCELL_X1 FILLER_18_60 ();
 FILLCELL_X8 FILLER_18_78 ();
 FILLCELL_X2 FILLER_18_86 ();
 FILLCELL_X4 FILLER_18_91 ();
 FILLCELL_X8 FILLER_18_103 ();
 FILLCELL_X4 FILLER_18_111 ();
 FILLCELL_X2 FILLER_18_115 ();
 FILLCELL_X1 FILLER_18_117 ();
 FILLCELL_X1 FILLER_18_127 ();
 FILLCELL_X4 FILLER_18_144 ();
 FILLCELL_X1 FILLER_18_148 ();
 FILLCELL_X2 FILLER_18_158 ();
 FILLCELL_X2 FILLER_18_165 ();
 FILLCELL_X1 FILLER_18_167 ();
 FILLCELL_X4 FILLER_18_187 ();
 FILLCELL_X2 FILLER_18_191 ();
 FILLCELL_X1 FILLER_18_193 ();
 FILLCELL_X1 FILLER_18_213 ();
 FILLCELL_X16 FILLER_18_217 ();
 FILLCELL_X8 FILLER_18_233 ();
 FILLCELL_X2 FILLER_18_241 ();
 FILLCELL_X8 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_12 ();
 FILLCELL_X32 FILLER_19_44 ();
 FILLCELL_X1 FILLER_19_76 ();
 FILLCELL_X2 FILLER_19_80 ();
 FILLCELL_X4 FILLER_19_105 ();
 FILLCELL_X1 FILLER_19_109 ();
 FILLCELL_X8 FILLER_19_114 ();
 FILLCELL_X2 FILLER_19_122 ();
 FILLCELL_X1 FILLER_19_124 ();
 FILLCELL_X2 FILLER_19_145 ();
 FILLCELL_X1 FILLER_19_147 ();
 FILLCELL_X2 FILLER_19_174 ();
 FILLCELL_X32 FILLER_19_180 ();
 FILLCELL_X16 FILLER_19_212 ();
 FILLCELL_X8 FILLER_19_228 ();
 FILLCELL_X4 FILLER_19_236 ();
 FILLCELL_X2 FILLER_19_240 ();
 FILLCELL_X1 FILLER_19_242 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X16 FILLER_20_33 ();
 FILLCELL_X4 FILLER_20_49 ();
 FILLCELL_X1 FILLER_20_53 ();
 FILLCELL_X2 FILLER_20_73 ();
 FILLCELL_X1 FILLER_20_79 ();
 FILLCELL_X4 FILLER_20_103 ();
 FILLCELL_X1 FILLER_20_107 ();
 FILLCELL_X2 FILLER_20_110 ();
 FILLCELL_X4 FILLER_20_116 ();
 FILLCELL_X2 FILLER_20_120 ();
 FILLCELL_X1 FILLER_20_122 ();
 FILLCELL_X1 FILLER_20_160 ();
 FILLCELL_X2 FILLER_20_166 ();
 FILLCELL_X1 FILLER_20_175 ();
 FILLCELL_X32 FILLER_20_183 ();
 FILLCELL_X16 FILLER_20_215 ();
 FILLCELL_X8 FILLER_20_231 ();
 FILLCELL_X4 FILLER_20_239 ();
 FILLCELL_X8 FILLER_21_1 ();
 FILLCELL_X2 FILLER_21_9 ();
 FILLCELL_X16 FILLER_21_14 ();
 FILLCELL_X1 FILLER_21_30 ();
 FILLCELL_X16 FILLER_21_34 ();
 FILLCELL_X4 FILLER_21_50 ();
 FILLCELL_X1 FILLER_21_54 ();
 FILLCELL_X8 FILLER_21_72 ();
 FILLCELL_X4 FILLER_21_80 ();
 FILLCELL_X1 FILLER_21_88 ();
 FILLCELL_X1 FILLER_21_94 ();
 FILLCELL_X1 FILLER_21_105 ();
 FILLCELL_X2 FILLER_21_109 ();
 FILLCELL_X8 FILLER_21_116 ();
 FILLCELL_X4 FILLER_21_124 ();
 FILLCELL_X2 FILLER_21_128 ();
 FILLCELL_X4 FILLER_21_134 ();
 FILLCELL_X1 FILLER_21_153 ();
 FILLCELL_X2 FILLER_21_170 ();
 FILLCELL_X32 FILLER_21_181 ();
 FILLCELL_X16 FILLER_21_213 ();
 FILLCELL_X8 FILLER_21_229 ();
 FILLCELL_X4 FILLER_21_237 ();
 FILLCELL_X2 FILLER_21_241 ();
 FILLCELL_X16 FILLER_22_1 ();
 FILLCELL_X4 FILLER_22_17 ();
 FILLCELL_X16 FILLER_22_24 ();
 FILLCELL_X8 FILLER_22_40 ();
 FILLCELL_X4 FILLER_22_48 ();
 FILLCELL_X8 FILLER_22_59 ();
 FILLCELL_X4 FILLER_22_67 ();
 FILLCELL_X2 FILLER_22_71 ();
 FILLCELL_X4 FILLER_22_77 ();
 FILLCELL_X2 FILLER_22_95 ();
 FILLCELL_X4 FILLER_22_106 ();
 FILLCELL_X1 FILLER_22_110 ();
 FILLCELL_X8 FILLER_22_115 ();
 FILLCELL_X1 FILLER_22_123 ();
 FILLCELL_X8 FILLER_22_133 ();
 FILLCELL_X4 FILLER_22_141 ();
 FILLCELL_X1 FILLER_22_145 ();
 FILLCELL_X8 FILLER_22_150 ();
 FILLCELL_X4 FILLER_22_158 ();
 FILLCELL_X32 FILLER_22_172 ();
 FILLCELL_X32 FILLER_22_204 ();
 FILLCELL_X4 FILLER_22_236 ();
 FILLCELL_X2 FILLER_22_240 ();
 FILLCELL_X1 FILLER_22_242 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X4 FILLER_23_33 ();
 FILLCELL_X2 FILLER_23_37 ();
 FILLCELL_X1 FILLER_23_39 ();
 FILLCELL_X8 FILLER_23_61 ();
 FILLCELL_X2 FILLER_23_69 ();
 FILLCELL_X8 FILLER_23_91 ();
 FILLCELL_X8 FILLER_23_118 ();
 FILLCELL_X4 FILLER_23_126 ();
 FILLCELL_X2 FILLER_23_130 ();
 FILLCELL_X1 FILLER_23_132 ();
 FILLCELL_X2 FILLER_23_136 ();
 FILLCELL_X4 FILLER_23_141 ();
 FILLCELL_X1 FILLER_23_145 ();
 FILLCELL_X8 FILLER_23_149 ();
 FILLCELL_X4 FILLER_23_157 ();
 FILLCELL_X1 FILLER_23_161 ();
 FILLCELL_X4 FILLER_23_173 ();
 FILLCELL_X1 FILLER_23_177 ();
 FILLCELL_X16 FILLER_23_182 ();
 FILLCELL_X4 FILLER_23_198 ();
 FILLCELL_X2 FILLER_23_202 ();
 FILLCELL_X32 FILLER_23_207 ();
 FILLCELL_X4 FILLER_23_239 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X8 FILLER_24_65 ();
 FILLCELL_X4 FILLER_24_73 ();
 FILLCELL_X1 FILLER_24_77 ();
 FILLCELL_X4 FILLER_24_85 ();
 FILLCELL_X2 FILLER_24_89 ();
 FILLCELL_X1 FILLER_24_91 ();
 FILLCELL_X2 FILLER_24_107 ();
 FILLCELL_X1 FILLER_24_109 ();
 FILLCELL_X2 FILLER_24_136 ();
 FILLCELL_X4 FILLER_24_155 ();
 FILLCELL_X32 FILLER_24_184 ();
 FILLCELL_X16 FILLER_24_216 ();
 FILLCELL_X8 FILLER_24_232 ();
 FILLCELL_X2 FILLER_24_240 ();
 FILLCELL_X1 FILLER_24_242 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X16 FILLER_25_33 ();
 FILLCELL_X8 FILLER_25_49 ();
 FILLCELL_X4 FILLER_25_57 ();
 FILLCELL_X2 FILLER_25_61 ();
 FILLCELL_X1 FILLER_25_63 ();
 FILLCELL_X8 FILLER_25_68 ();
 FILLCELL_X4 FILLER_25_76 ();
 FILLCELL_X2 FILLER_25_80 ();
 FILLCELL_X1 FILLER_25_82 ();
 FILLCELL_X1 FILLER_25_97 ();
 FILLCELL_X2 FILLER_25_110 ();
 FILLCELL_X1 FILLER_25_112 ();
 FILLCELL_X2 FILLER_25_136 ();
 FILLCELL_X2 FILLER_25_142 ();
 FILLCELL_X1 FILLER_25_144 ();
 FILLCELL_X32 FILLER_25_164 ();
 FILLCELL_X32 FILLER_25_196 ();
 FILLCELL_X8 FILLER_25_228 ();
 FILLCELL_X4 FILLER_25_236 ();
 FILLCELL_X2 FILLER_25_240 ();
 FILLCELL_X1 FILLER_25_242 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X16 FILLER_26_33 ();
 FILLCELL_X1 FILLER_26_49 ();
 FILLCELL_X2 FILLER_26_74 ();
 FILLCELL_X1 FILLER_26_76 ();
 FILLCELL_X8 FILLER_26_98 ();
 FILLCELL_X2 FILLER_26_106 ();
 FILLCELL_X1 FILLER_26_108 ();
 FILLCELL_X1 FILLER_26_113 ();
 FILLCELL_X16 FILLER_26_118 ();
 FILLCELL_X8 FILLER_26_134 ();
 FILLCELL_X4 FILLER_26_142 ();
 FILLCELL_X32 FILLER_26_151 ();
 FILLCELL_X32 FILLER_26_183 ();
 FILLCELL_X16 FILLER_26_215 ();
 FILLCELL_X8 FILLER_26_231 ();
 FILLCELL_X4 FILLER_26_239 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X16 FILLER_27_65 ();
 FILLCELL_X8 FILLER_27_81 ();
 FILLCELL_X2 FILLER_27_89 ();
 FILLCELL_X1 FILLER_27_114 ();
 FILLCELL_X4 FILLER_27_119 ();
 FILLCELL_X2 FILLER_27_123 ();
 FILLCELL_X1 FILLER_27_125 ();
 FILLCELL_X2 FILLER_27_130 ();
 FILLCELL_X8 FILLER_27_138 ();
 FILLCELL_X2 FILLER_27_146 ();
 FILLCELL_X4 FILLER_27_151 ();
 FILLCELL_X1 FILLER_27_155 ();
 FILLCELL_X4 FILLER_27_158 ();
 FILLCELL_X1 FILLER_27_162 ();
 FILLCELL_X32 FILLER_27_165 ();
 FILLCELL_X32 FILLER_27_197 ();
 FILLCELL_X8 FILLER_27_229 ();
 FILLCELL_X4 FILLER_27_237 ();
 FILLCELL_X2 FILLER_27_241 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X8 FILLER_28_33 ();
 FILLCELL_X4 FILLER_28_41 ();
 FILLCELL_X1 FILLER_28_45 ();
 FILLCELL_X4 FILLER_28_74 ();
 FILLCELL_X4 FILLER_28_82 ();
 FILLCELL_X2 FILLER_28_86 ();
 FILLCELL_X8 FILLER_28_95 ();
 FILLCELL_X1 FILLER_28_103 ();
 FILLCELL_X8 FILLER_28_127 ();
 FILLCELL_X2 FILLER_28_160 ();
 FILLCELL_X1 FILLER_28_162 ();
 FILLCELL_X32 FILLER_28_167 ();
 FILLCELL_X32 FILLER_28_199 ();
 FILLCELL_X8 FILLER_28_231 ();
 FILLCELL_X4 FILLER_28_239 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X16 FILLER_29_33 ();
 FILLCELL_X4 FILLER_29_49 ();
 FILLCELL_X2 FILLER_29_53 ();
 FILLCELL_X2 FILLER_29_66 ();
 FILLCELL_X1 FILLER_29_68 ();
 FILLCELL_X2 FILLER_29_73 ();
 FILLCELL_X1 FILLER_29_75 ();
 FILLCELL_X8 FILLER_29_93 ();
 FILLCELL_X4 FILLER_29_101 ();
 FILLCELL_X2 FILLER_29_105 ();
 FILLCELL_X1 FILLER_29_107 ();
 FILLCELL_X1 FILLER_29_122 ();
 FILLCELL_X2 FILLER_29_141 ();
 FILLCELL_X4 FILLER_29_147 ();
 FILLCELL_X2 FILLER_29_155 ();
 FILLCELL_X1 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_183 ();
 FILLCELL_X16 FILLER_29_215 ();
 FILLCELL_X8 FILLER_29_231 ();
 FILLCELL_X4 FILLER_29_239 ();
 FILLCELL_X1 FILLER_30_1 ();
 FILLCELL_X16 FILLER_30_12 ();
 FILLCELL_X8 FILLER_30_28 ();
 FILLCELL_X4 FILLER_30_36 ();
 FILLCELL_X1 FILLER_30_121 ();
 FILLCELL_X1 FILLER_30_173 ();
 FILLCELL_X32 FILLER_30_181 ();
 FILLCELL_X16 FILLER_30_213 ();
 FILLCELL_X8 FILLER_30_229 ();
 FILLCELL_X4 FILLER_30_237 ();
 FILLCELL_X2 FILLER_30_241 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X16 FILLER_31_33 ();
 FILLCELL_X4 FILLER_31_49 ();
 FILLCELL_X2 FILLER_31_53 ();
 FILLCELL_X1 FILLER_31_55 ();
 FILLCELL_X2 FILLER_31_59 ();
 FILLCELL_X1 FILLER_31_61 ();
 FILLCELL_X4 FILLER_31_68 ();
 FILLCELL_X2 FILLER_31_72 ();
 FILLCELL_X4 FILLER_31_77 ();
 FILLCELL_X1 FILLER_31_81 ();
 FILLCELL_X1 FILLER_31_99 ();
 FILLCELL_X2 FILLER_31_176 ();
 FILLCELL_X32 FILLER_31_181 ();
 FILLCELL_X16 FILLER_31_213 ();
 FILLCELL_X8 FILLER_31_229 ();
 FILLCELL_X4 FILLER_31_237 ();
 FILLCELL_X2 FILLER_31_241 ();
endmodule
