module lfsr (bit_out,
    clk,
    enable,
    load,
    rst_n,
    lfsr_out,
    seed);
 output bit_out;
 input clk;
 input enable;
 input load;
 input rst_n;
 output [7:0] lfsr_out;
 input [7:0] seed;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire _34_;
 wire _35_;
 wire _36_;
 wire _37_;
 wire _38_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 CLKBUF_X2 _39_ (.A(rst_n),
    .Z(_08_));
 BUF_X4 _40_ (.A(enable),
    .Z(_09_));
 MUX2_X1 _41_ (.A(net10),
    .B(net12),
    .S(_09_),
    .Z(_10_));
 INV_X2 _42_ (.A(net1),
    .ZN(_11_));
 MUX2_X1 _43_ (.A(net2),
    .B(_10_),
    .S(_11_),
    .Z(_12_));
 AND2_X1 _44_ (.A1(_08_),
    .A2(_12_),
    .ZN(_00_));
 MUX2_X1 _45_ (.A(net12),
    .B(net13),
    .S(_09_),
    .Z(_13_));
 MUX2_X1 _46_ (.A(net3),
    .B(_13_),
    .S(_11_),
    .Z(_14_));
 AND2_X1 _47_ (.A1(_08_),
    .A2(_14_),
    .ZN(_01_));
 MUX2_X1 _48_ (.A(net13),
    .B(net14),
    .S(_09_),
    .Z(_15_));
 MUX2_X1 _49_ (.A(net4),
    .B(_15_),
    .S(_11_),
    .Z(_16_));
 AND2_X1 _50_ (.A1(_08_),
    .A2(_16_),
    .ZN(_02_));
 MUX2_X1 _51_ (.A(net14),
    .B(net15),
    .S(_09_),
    .Z(_17_));
 MUX2_X1 _52_ (.A(net5),
    .B(_17_),
    .S(_11_),
    .Z(_18_));
 AND2_X1 _53_ (.A1(_08_),
    .A2(_18_),
    .ZN(_03_));
 MUX2_X1 _54_ (.A(net15),
    .B(net16),
    .S(_09_),
    .Z(_19_));
 MUX2_X1 _55_ (.A(net6),
    .B(_19_),
    .S(_11_),
    .Z(_20_));
 AND2_X1 _56_ (.A1(_08_),
    .A2(_20_),
    .ZN(_04_));
 MUX2_X1 _57_ (.A(net16),
    .B(net17),
    .S(_09_),
    .Z(_21_));
 MUX2_X1 _58_ (.A(net7),
    .B(_21_),
    .S(_11_),
    .Z(_22_));
 AND2_X1 _59_ (.A1(_08_),
    .A2(_22_),
    .ZN(_05_));
 MUX2_X1 _60_ (.A(net17),
    .B(net18),
    .S(_09_),
    .Z(_23_));
 MUX2_X1 _61_ (.A(net8),
    .B(_23_),
    .S(_11_),
    .Z(_24_));
 AND2_X1 _62_ (.A1(_08_),
    .A2(_24_),
    .ZN(_06_));
 OR2_X1 _63_ (.A1(net1),
    .A2(net18),
    .ZN(_25_));
 XNOR2_X1 _64_ (.A(net15),
    .B(net16),
    .ZN(_26_));
 XNOR2_X1 _65_ (.A(net14),
    .B(_26_),
    .ZN(_27_));
 AOI21_X1 _66_ (.A(_25_),
    .B1(_27_),
    .B2(_09_),
    .ZN(_28_));
 AND4_X1 _67_ (.A1(_11_),
    .A2(_09_),
    .A3(net18),
    .A4(_27_),
    .ZN(_29_));
 OAI21_X1 _68_ (.A(_08_),
    .B1(net9),
    .B2(_11_),
    .ZN(_30_));
 NOR3_X1 _69_ (.A1(_28_),
    .A2(_29_),
    .A3(_30_),
    .ZN(_07_));
 BUF_X1 _70_ (.A(net10),
    .Z(net11));
 DFF_X1 \lfsr_reg[0]$_SDFFE_PN0P_  (.D(_00_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net10),
    .QN(_38_));
 DFF_X1 \lfsr_reg[1]$_SDFFE_PN0P_  (.D(_01_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net12),
    .QN(_37_));
 DFF_X1 \lfsr_reg[2]$_SDFFE_PN0P_  (.D(_02_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net13),
    .QN(_36_));
 DFF_X1 \lfsr_reg[3]$_SDFFE_PN0P_  (.D(_03_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net14),
    .QN(_35_));
 DFF_X1 \lfsr_reg[4]$_SDFFE_PN0P_  (.D(_04_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net15),
    .QN(_34_));
 DFF_X1 \lfsr_reg[5]$_SDFFE_PN0P_  (.D(_05_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net16),
    .QN(_33_));
 DFF_X1 \lfsr_reg[6]$_SDFFE_PN0P_  (.D(_06_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net17),
    .QN(_32_));
 DFF_X1 \lfsr_reg[7]$_SDFFE_PN0P_  (.D(_07_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net18),
    .QN(_31_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_59 ();
 BUF_X1 input1 (.A(load),
    .Z(net1));
 BUF_X1 input2 (.A(seed[0]),
    .Z(net2));
 BUF_X1 input3 (.A(seed[1]),
    .Z(net3));
 BUF_X1 input4 (.A(seed[2]),
    .Z(net4));
 BUF_X1 input5 (.A(seed[3]),
    .Z(net5));
 BUF_X1 input6 (.A(seed[4]),
    .Z(net6));
 BUF_X1 input7 (.A(seed[5]),
    .Z(net7));
 BUF_X1 input8 (.A(seed[6]),
    .Z(net8));
 BUF_X1 input9 (.A(seed[7]),
    .Z(net9));
 BUF_X1 output10 (.A(net10),
    .Z(bit_out));
 BUF_X1 output11 (.A(net11),
    .Z(lfsr_out[0]));
 BUF_X1 output12 (.A(net12),
    .Z(lfsr_out[1]));
 BUF_X1 output13 (.A(net13),
    .Z(lfsr_out[2]));
 BUF_X1 output14 (.A(net14),
    .Z(lfsr_out[3]));
 BUF_X1 output15 (.A(net15),
    .Z(lfsr_out[4]));
 BUF_X1 output16 (.A(net16),
    .Z(lfsr_out[5]));
 BUF_X1 output17 (.A(net17),
    .Z(lfsr_out[6]));
 BUF_X1 output18 (.A(net18),
    .Z(lfsr_out[7]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X8 FILLER_0_97 ();
 FILLCELL_X2 FILLER_0_105 ();
 FILLCELL_X8 FILLER_0_113 ();
 FILLCELL_X8 FILLER_0_127 ();
 FILLCELL_X1 FILLER_0_135 ();
 FILLCELL_X32 FILLER_0_139 ();
 FILLCELL_X32 FILLER_0_171 ();
 FILLCELL_X16 FILLER_0_203 ();
 FILLCELL_X8 FILLER_0_219 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X4 FILLER_1_97 ();
 FILLCELL_X1 FILLER_1_101 ();
 FILLCELL_X4 FILLER_1_106 ();
 FILLCELL_X8 FILLER_1_113 ();
 FILLCELL_X1 FILLER_1_121 ();
 FILLCELL_X8 FILLER_1_129 ();
 FILLCELL_X1 FILLER_1_137 ();
 FILLCELL_X32 FILLER_1_145 ();
 FILLCELL_X32 FILLER_1_177 ();
 FILLCELL_X16 FILLER_1_209 ();
 FILLCELL_X2 FILLER_1_225 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X8 FILLER_2_97 ();
 FILLCELL_X2 FILLER_2_105 ();
 FILLCELL_X1 FILLER_2_107 ();
 FILLCELL_X8 FILLER_2_129 ();
 FILLCELL_X4 FILLER_2_137 ();
 FILLCELL_X8 FILLER_2_148 ();
 FILLCELL_X2 FILLER_2_156 ();
 FILLCELL_X1 FILLER_2_158 ();
 FILLCELL_X32 FILLER_2_163 ();
 FILLCELL_X32 FILLER_2_195 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X16 FILLER_3_97 ();
 FILLCELL_X1 FILLER_3_113 ();
 FILLCELL_X8 FILLER_3_118 ();
 FILLCELL_X1 FILLER_3_126 ();
 FILLCELL_X8 FILLER_3_131 ();
 FILLCELL_X2 FILLER_3_139 ();
 FILLCELL_X32 FILLER_3_148 ();
 FILLCELL_X32 FILLER_3_180 ();
 FILLCELL_X8 FILLER_3_212 ();
 FILLCELL_X4 FILLER_3_220 ();
 FILLCELL_X2 FILLER_3_224 ();
 FILLCELL_X1 FILLER_3_226 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X16 FILLER_4_97 ();
 FILLCELL_X4 FILLER_4_113 ();
 FILLCELL_X1 FILLER_4_134 ();
 FILLCELL_X8 FILLER_4_152 ();
 FILLCELL_X1 FILLER_4_160 ();
 FILLCELL_X32 FILLER_4_178 ();
 FILLCELL_X16 FILLER_4_210 ();
 FILLCELL_X1 FILLER_4_226 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X2 FILLER_5_225 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X16 FILLER_6_129 ();
 FILLCELL_X8 FILLER_6_145 ();
 FILLCELL_X32 FILLER_6_158 ();
 FILLCELL_X32 FILLER_6_190 ();
 FILLCELL_X4 FILLER_6_222 ();
 FILLCELL_X1 FILLER_6_226 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X2 FILLER_7_225 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X2 FILLER_8_225 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X2 FILLER_9_225 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X16 FILLER_10_129 ();
 FILLCELL_X4 FILLER_10_145 ();
 FILLCELL_X4 FILLER_10_154 ();
 FILLCELL_X2 FILLER_10_158 ();
 FILLCELL_X8 FILLER_10_184 ();
 FILLCELL_X2 FILLER_10_192 ();
 FILLCELL_X1 FILLER_10_194 ();
 FILLCELL_X16 FILLER_10_198 ();
 FILLCELL_X4 FILLER_10_214 ();
 FILLCELL_X2 FILLER_10_218 ();
 FILLCELL_X1 FILLER_10_223 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X16 FILLER_11_172 ();
 FILLCELL_X4 FILLER_11_188 ();
 FILLCELL_X1 FILLER_11_192 ();
 FILLCELL_X16 FILLER_11_196 ();
 FILLCELL_X8 FILLER_11_212 ();
 FILLCELL_X4 FILLER_11_220 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X2 FILLER_12_225 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X2 FILLER_13_225 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X8 FILLER_14_97 ();
 FILLCELL_X4 FILLER_14_105 ();
 FILLCELL_X32 FILLER_14_142 ();
 FILLCELL_X32 FILLER_14_174 ();
 FILLCELL_X16 FILLER_14_206 ();
 FILLCELL_X4 FILLER_14_222 ();
 FILLCELL_X1 FILLER_14_226 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X4 FILLER_15_97 ();
 FILLCELL_X2 FILLER_15_101 ();
 FILLCELL_X4 FILLER_15_117 ();
 FILLCELL_X2 FILLER_15_121 ();
 FILLCELL_X1 FILLER_15_123 ();
 FILLCELL_X2 FILLER_15_131 ();
 FILLCELL_X32 FILLER_15_180 ();
 FILLCELL_X8 FILLER_15_212 ();
 FILLCELL_X4 FILLER_15_220 ();
 FILLCELL_X2 FILLER_15_224 ();
 FILLCELL_X1 FILLER_15_226 ();
 FILLCELL_X8 FILLER_16_1 ();
 FILLCELL_X4 FILLER_16_9 ();
 FILLCELL_X2 FILLER_16_13 ();
 FILLCELL_X32 FILLER_16_18 ();
 FILLCELL_X32 FILLER_16_50 ();
 FILLCELL_X16 FILLER_16_82 ();
 FILLCELL_X8 FILLER_16_98 ();
 FILLCELL_X4 FILLER_16_151 ();
 FILLCELL_X2 FILLER_16_155 ();
 FILLCELL_X1 FILLER_16_157 ();
 FILLCELL_X32 FILLER_16_166 ();
 FILLCELL_X16 FILLER_16_198 ();
 FILLCELL_X8 FILLER_16_214 ();
 FILLCELL_X4 FILLER_16_222 ();
 FILLCELL_X1 FILLER_16_226 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X8 FILLER_17_129 ();
 FILLCELL_X2 FILLER_17_137 ();
 FILLCELL_X1 FILLER_17_139 ();
 FILLCELL_X8 FILLER_17_147 ();
 FILLCELL_X4 FILLER_17_155 ();
 FILLCELL_X2 FILLER_17_159 ();
 FILLCELL_X16 FILLER_17_164 ();
 FILLCELL_X8 FILLER_17_180 ();
 FILLCELL_X4 FILLER_17_188 ();
 FILLCELL_X2 FILLER_17_192 ();
 FILLCELL_X1 FILLER_17_194 ();
 FILLCELL_X8 FILLER_17_198 ();
 FILLCELL_X1 FILLER_17_206 ();
 FILLCELL_X16 FILLER_17_210 ();
 FILLCELL_X1 FILLER_17_226 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X16 FILLER_18_161 ();
 FILLCELL_X8 FILLER_18_177 ();
 FILLCELL_X4 FILLER_18_185 ();
 FILLCELL_X2 FILLER_18_189 ();
 FILLCELL_X32 FILLER_18_194 ();
 FILLCELL_X1 FILLER_18_226 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X2 FILLER_19_225 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X2 FILLER_20_225 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X2 FILLER_21_225 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X2 FILLER_22_225 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X2 FILLER_23_225 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X2 FILLER_24_225 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X2 FILLER_25_225 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X2 FILLER_26_225 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X2 FILLER_27_225 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X8 FILLER_28_97 ();
 FILLCELL_X16 FILLER_28_108 ();
 FILLCELL_X8 FILLER_28_124 ();
 FILLCELL_X4 FILLER_28_132 ();
 FILLCELL_X2 FILLER_28_136 ();
 FILLCELL_X1 FILLER_28_138 ();
 FILLCELL_X32 FILLER_28_142 ();
 FILLCELL_X32 FILLER_28_174 ();
 FILLCELL_X16 FILLER_28_206 ();
 FILLCELL_X4 FILLER_28_222 ();
 FILLCELL_X1 FILLER_28_226 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X16 FILLER_29_97 ();
 FILLCELL_X16 FILLER_29_116 ();
 FILLCELL_X8 FILLER_29_132 ();
 FILLCELL_X4 FILLER_29_140 ();
 FILLCELL_X1 FILLER_29_144 ();
 FILLCELL_X32 FILLER_29_148 ();
 FILLCELL_X32 FILLER_29_180 ();
 FILLCELL_X8 FILLER_29_212 ();
 FILLCELL_X4 FILLER_29_220 ();
 FILLCELL_X2 FILLER_29_224 ();
 FILLCELL_X1 FILLER_29_226 ();
endmodule
