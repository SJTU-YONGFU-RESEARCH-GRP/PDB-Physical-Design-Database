module memory_mapped_fifo (clk,
    ext_empty,
    ext_full,
    ext_rd_en,
    ext_wr_en,
    mem_ready,
    mem_valid,
    mem_write,
    rst_n,
    ext_rd_data,
    ext_wr_data,
    mem_addr,
    mem_rdata,
    mem_wdata);
 input clk;
 output ext_empty;
 output ext_full;
 input ext_rd_en;
 input ext_wr_en;
 output mem_ready;
 input mem_valid;
 input mem_write;
 input rst_n;
 output [31:0] ext_rd_data;
 input [31:0] ext_wr_data;
 input [3:0] mem_addr;
 output [31:0] mem_rdata;
 input [31:0] mem_wdata;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire \mem[0][0] ;
 wire \mem[0][10] ;
 wire \mem[0][11] ;
 wire \mem[0][12] ;
 wire \mem[0][13] ;
 wire \mem[0][14] ;
 wire \mem[0][15] ;
 wire \mem[0][16] ;
 wire \mem[0][17] ;
 wire \mem[0][18] ;
 wire \mem[0][19] ;
 wire \mem[0][1] ;
 wire \mem[0][20] ;
 wire \mem[0][21] ;
 wire \mem[0][22] ;
 wire \mem[0][23] ;
 wire \mem[0][24] ;
 wire \mem[0][25] ;
 wire \mem[0][26] ;
 wire \mem[0][27] ;
 wire \mem[0][28] ;
 wire \mem[0][29] ;
 wire \mem[0][2] ;
 wire \mem[0][30] ;
 wire \mem[0][31] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[0][8] ;
 wire \mem[0][9] ;
 wire \mem[10][0] ;
 wire \mem[10][10] ;
 wire \mem[10][11] ;
 wire \mem[10][12] ;
 wire \mem[10][13] ;
 wire \mem[10][14] ;
 wire \mem[10][15] ;
 wire \mem[10][16] ;
 wire \mem[10][17] ;
 wire \mem[10][18] ;
 wire \mem[10][19] ;
 wire \mem[10][1] ;
 wire \mem[10][20] ;
 wire \mem[10][21] ;
 wire \mem[10][22] ;
 wire \mem[10][23] ;
 wire \mem[10][24] ;
 wire \mem[10][25] ;
 wire \mem[10][26] ;
 wire \mem[10][27] ;
 wire \mem[10][28] ;
 wire \mem[10][29] ;
 wire \mem[10][2] ;
 wire \mem[10][30] ;
 wire \mem[10][31] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[10][8] ;
 wire \mem[10][9] ;
 wire \mem[11][0] ;
 wire \mem[11][10] ;
 wire \mem[11][11] ;
 wire \mem[11][12] ;
 wire \mem[11][13] ;
 wire \mem[11][14] ;
 wire \mem[11][15] ;
 wire \mem[11][16] ;
 wire \mem[11][17] ;
 wire \mem[11][18] ;
 wire \mem[11][19] ;
 wire \mem[11][1] ;
 wire \mem[11][20] ;
 wire \mem[11][21] ;
 wire \mem[11][22] ;
 wire \mem[11][23] ;
 wire \mem[11][24] ;
 wire \mem[11][25] ;
 wire \mem[11][26] ;
 wire \mem[11][27] ;
 wire \mem[11][28] ;
 wire \mem[11][29] ;
 wire \mem[11][2] ;
 wire \mem[11][30] ;
 wire \mem[11][31] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[11][8] ;
 wire \mem[11][9] ;
 wire \mem[12][0] ;
 wire \mem[12][10] ;
 wire \mem[12][11] ;
 wire \mem[12][12] ;
 wire \mem[12][13] ;
 wire \mem[12][14] ;
 wire \mem[12][15] ;
 wire \mem[12][16] ;
 wire \mem[12][17] ;
 wire \mem[12][18] ;
 wire \mem[12][19] ;
 wire \mem[12][1] ;
 wire \mem[12][20] ;
 wire \mem[12][21] ;
 wire \mem[12][22] ;
 wire \mem[12][23] ;
 wire \mem[12][24] ;
 wire \mem[12][25] ;
 wire \mem[12][26] ;
 wire \mem[12][27] ;
 wire \mem[12][28] ;
 wire \mem[12][29] ;
 wire \mem[12][2] ;
 wire \mem[12][30] ;
 wire \mem[12][31] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[12][8] ;
 wire \mem[12][9] ;
 wire \mem[13][0] ;
 wire \mem[13][10] ;
 wire \mem[13][11] ;
 wire \mem[13][12] ;
 wire \mem[13][13] ;
 wire \mem[13][14] ;
 wire \mem[13][15] ;
 wire \mem[13][16] ;
 wire \mem[13][17] ;
 wire \mem[13][18] ;
 wire \mem[13][19] ;
 wire \mem[13][1] ;
 wire \mem[13][20] ;
 wire \mem[13][21] ;
 wire \mem[13][22] ;
 wire \mem[13][23] ;
 wire \mem[13][24] ;
 wire \mem[13][25] ;
 wire \mem[13][26] ;
 wire \mem[13][27] ;
 wire \mem[13][28] ;
 wire \mem[13][29] ;
 wire \mem[13][2] ;
 wire \mem[13][30] ;
 wire \mem[13][31] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[13][8] ;
 wire \mem[13][9] ;
 wire \mem[14][0] ;
 wire \mem[14][10] ;
 wire \mem[14][11] ;
 wire \mem[14][12] ;
 wire \mem[14][13] ;
 wire \mem[14][14] ;
 wire \mem[14][15] ;
 wire \mem[14][16] ;
 wire \mem[14][17] ;
 wire \mem[14][18] ;
 wire \mem[14][19] ;
 wire \mem[14][1] ;
 wire \mem[14][20] ;
 wire \mem[14][21] ;
 wire \mem[14][22] ;
 wire \mem[14][23] ;
 wire \mem[14][24] ;
 wire \mem[14][25] ;
 wire \mem[14][26] ;
 wire \mem[14][27] ;
 wire \mem[14][28] ;
 wire \mem[14][29] ;
 wire \mem[14][2] ;
 wire \mem[14][30] ;
 wire \mem[14][31] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[14][8] ;
 wire \mem[14][9] ;
 wire \mem[15][0] ;
 wire \mem[15][10] ;
 wire \mem[15][11] ;
 wire \mem[15][12] ;
 wire \mem[15][13] ;
 wire \mem[15][14] ;
 wire \mem[15][15] ;
 wire \mem[15][16] ;
 wire \mem[15][17] ;
 wire \mem[15][18] ;
 wire \mem[15][19] ;
 wire \mem[15][1] ;
 wire \mem[15][20] ;
 wire \mem[15][21] ;
 wire \mem[15][22] ;
 wire \mem[15][23] ;
 wire \mem[15][24] ;
 wire \mem[15][25] ;
 wire \mem[15][26] ;
 wire \mem[15][27] ;
 wire \mem[15][28] ;
 wire \mem[15][29] ;
 wire \mem[15][2] ;
 wire \mem[15][30] ;
 wire \mem[15][31] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[15][8] ;
 wire \mem[15][9] ;
 wire \mem[1][0] ;
 wire \mem[1][10] ;
 wire \mem[1][11] ;
 wire \mem[1][12] ;
 wire \mem[1][13] ;
 wire \mem[1][14] ;
 wire \mem[1][15] ;
 wire \mem[1][16] ;
 wire \mem[1][17] ;
 wire \mem[1][18] ;
 wire \mem[1][19] ;
 wire \mem[1][1] ;
 wire \mem[1][20] ;
 wire \mem[1][21] ;
 wire \mem[1][22] ;
 wire \mem[1][23] ;
 wire \mem[1][24] ;
 wire \mem[1][25] ;
 wire \mem[1][26] ;
 wire \mem[1][27] ;
 wire \mem[1][28] ;
 wire \mem[1][29] ;
 wire \mem[1][2] ;
 wire \mem[1][30] ;
 wire \mem[1][31] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[1][8] ;
 wire \mem[1][9] ;
 wire \mem[2][0] ;
 wire \mem[2][10] ;
 wire \mem[2][11] ;
 wire \mem[2][12] ;
 wire \mem[2][13] ;
 wire \mem[2][14] ;
 wire \mem[2][15] ;
 wire \mem[2][16] ;
 wire \mem[2][17] ;
 wire \mem[2][18] ;
 wire \mem[2][19] ;
 wire \mem[2][1] ;
 wire \mem[2][20] ;
 wire \mem[2][21] ;
 wire \mem[2][22] ;
 wire \mem[2][23] ;
 wire \mem[2][24] ;
 wire \mem[2][25] ;
 wire \mem[2][26] ;
 wire \mem[2][27] ;
 wire \mem[2][28] ;
 wire \mem[2][29] ;
 wire \mem[2][2] ;
 wire \mem[2][30] ;
 wire \mem[2][31] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[2][8] ;
 wire \mem[2][9] ;
 wire \mem[3][0] ;
 wire \mem[3][10] ;
 wire \mem[3][11] ;
 wire \mem[3][12] ;
 wire \mem[3][13] ;
 wire \mem[3][14] ;
 wire \mem[3][15] ;
 wire \mem[3][16] ;
 wire \mem[3][17] ;
 wire \mem[3][18] ;
 wire \mem[3][19] ;
 wire \mem[3][1] ;
 wire \mem[3][20] ;
 wire \mem[3][21] ;
 wire \mem[3][22] ;
 wire \mem[3][23] ;
 wire \mem[3][24] ;
 wire \mem[3][25] ;
 wire \mem[3][26] ;
 wire \mem[3][27] ;
 wire \mem[3][28] ;
 wire \mem[3][29] ;
 wire \mem[3][2] ;
 wire \mem[3][30] ;
 wire \mem[3][31] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[3][8] ;
 wire \mem[3][9] ;
 wire \mem[4][0] ;
 wire \mem[4][10] ;
 wire \mem[4][11] ;
 wire \mem[4][12] ;
 wire \mem[4][13] ;
 wire \mem[4][14] ;
 wire \mem[4][15] ;
 wire \mem[4][16] ;
 wire \mem[4][17] ;
 wire \mem[4][18] ;
 wire \mem[4][19] ;
 wire \mem[4][1] ;
 wire \mem[4][20] ;
 wire \mem[4][21] ;
 wire \mem[4][22] ;
 wire \mem[4][23] ;
 wire \mem[4][24] ;
 wire \mem[4][25] ;
 wire \mem[4][26] ;
 wire \mem[4][27] ;
 wire \mem[4][28] ;
 wire \mem[4][29] ;
 wire \mem[4][2] ;
 wire \mem[4][30] ;
 wire \mem[4][31] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[4][8] ;
 wire \mem[4][9] ;
 wire \mem[5][0] ;
 wire \mem[5][10] ;
 wire \mem[5][11] ;
 wire \mem[5][12] ;
 wire \mem[5][13] ;
 wire \mem[5][14] ;
 wire \mem[5][15] ;
 wire \mem[5][16] ;
 wire \mem[5][17] ;
 wire \mem[5][18] ;
 wire \mem[5][19] ;
 wire \mem[5][1] ;
 wire \mem[5][20] ;
 wire \mem[5][21] ;
 wire \mem[5][22] ;
 wire \mem[5][23] ;
 wire \mem[5][24] ;
 wire \mem[5][25] ;
 wire \mem[5][26] ;
 wire \mem[5][27] ;
 wire \mem[5][28] ;
 wire \mem[5][29] ;
 wire \mem[5][2] ;
 wire \mem[5][30] ;
 wire \mem[5][31] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[5][8] ;
 wire \mem[5][9] ;
 wire \mem[6][0] ;
 wire \mem[6][10] ;
 wire \mem[6][11] ;
 wire \mem[6][12] ;
 wire \mem[6][13] ;
 wire \mem[6][14] ;
 wire \mem[6][15] ;
 wire \mem[6][16] ;
 wire \mem[6][17] ;
 wire \mem[6][18] ;
 wire \mem[6][19] ;
 wire \mem[6][1] ;
 wire \mem[6][20] ;
 wire \mem[6][21] ;
 wire \mem[6][22] ;
 wire \mem[6][23] ;
 wire \mem[6][24] ;
 wire \mem[6][25] ;
 wire \mem[6][26] ;
 wire \mem[6][27] ;
 wire \mem[6][28] ;
 wire \mem[6][29] ;
 wire \mem[6][2] ;
 wire \mem[6][30] ;
 wire \mem[6][31] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[6][8] ;
 wire \mem[6][9] ;
 wire \mem[7][0] ;
 wire \mem[7][10] ;
 wire \mem[7][11] ;
 wire \mem[7][12] ;
 wire \mem[7][13] ;
 wire \mem[7][14] ;
 wire \mem[7][15] ;
 wire \mem[7][16] ;
 wire \mem[7][17] ;
 wire \mem[7][18] ;
 wire \mem[7][19] ;
 wire \mem[7][1] ;
 wire \mem[7][20] ;
 wire \mem[7][21] ;
 wire \mem[7][22] ;
 wire \mem[7][23] ;
 wire \mem[7][24] ;
 wire \mem[7][25] ;
 wire \mem[7][26] ;
 wire \mem[7][27] ;
 wire \mem[7][28] ;
 wire \mem[7][29] ;
 wire \mem[7][2] ;
 wire \mem[7][30] ;
 wire \mem[7][31] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[7][8] ;
 wire \mem[7][9] ;
 wire \mem[8][0] ;
 wire \mem[8][10] ;
 wire \mem[8][11] ;
 wire \mem[8][12] ;
 wire \mem[8][13] ;
 wire \mem[8][14] ;
 wire \mem[8][15] ;
 wire \mem[8][16] ;
 wire \mem[8][17] ;
 wire \mem[8][18] ;
 wire \mem[8][19] ;
 wire \mem[8][1] ;
 wire \mem[8][20] ;
 wire \mem[8][21] ;
 wire \mem[8][22] ;
 wire \mem[8][23] ;
 wire \mem[8][24] ;
 wire \mem[8][25] ;
 wire \mem[8][26] ;
 wire \mem[8][27] ;
 wire \mem[8][28] ;
 wire \mem[8][29] ;
 wire \mem[8][2] ;
 wire \mem[8][30] ;
 wire \mem[8][31] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[8][8] ;
 wire \mem[8][9] ;
 wire \mem[9][0] ;
 wire \mem[9][10] ;
 wire \mem[9][11] ;
 wire \mem[9][12] ;
 wire \mem[9][13] ;
 wire \mem[9][14] ;
 wire \mem[9][15] ;
 wire \mem[9][16] ;
 wire \mem[9][17] ;
 wire \mem[9][18] ;
 wire \mem[9][19] ;
 wire \mem[9][1] ;
 wire \mem[9][20] ;
 wire \mem[9][21] ;
 wire \mem[9][22] ;
 wire \mem[9][23] ;
 wire \mem[9][24] ;
 wire \mem[9][25] ;
 wire \mem[9][26] ;
 wire \mem[9][27] ;
 wire \mem[9][28] ;
 wire \mem[9][29] ;
 wire \mem[9][2] ;
 wire \mem[9][30] ;
 wire \mem[9][31] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \mem[9][8] ;
 wire \mem[9][9] ;
 wire \rd_ptr[0] ;
 wire \rd_ptr[1] ;
 wire \rd_ptr[2] ;
 wire \rd_ptr[3] ;
 wire \rd_ptr[4] ;
 wire \wr_ptr[0] ;
 wire \wr_ptr[1] ;
 wire \wr_ptr[2] ;
 wire \wr_ptr[3] ;
 wire \wr_ptr[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net165;
 wire net166;

 sky130_fd_sc_hd__a21o_1 _0905_ (.A1(_0886_),
    .A2(_0874_),
    .B1(_0885_),
    .X(_0741_));
 sky130_fd_sc_hd__a21oi_2 _0906_ (.A1(_0883_),
    .A2(_0741_),
    .B1(_0882_),
    .Y(_0742_));
 sky130_fd_sc_hd__xor2_2 _0907_ (.A(\wr_ptr[4] ),
    .B(\rd_ptr[4] ),
    .X(_0743_));
 sky130_fd_sc_hd__xnor2_4 _0908_ (.A(_0742_),
    .B(_0743_),
    .Y(_0744_));
 sky130_fd_sc_hd__xnor2_1 _0909_ (.A(_0886_),
    .B(_0874_),
    .Y(_0745_));
 sky130_fd_sc_hd__nand3b_1 _0910_ (.A_N(_0875_),
    .B(_0745_),
    .C(_0878_),
    .Y(_0746_));
 sky130_fd_sc_hd__nand2b_1 _0911_ (.A_N(_0877_),
    .B(_0880_),
    .Y(_0747_));
 sky130_fd_sc_hd__nor2_1 _0912_ (.A(_0879_),
    .B(_0885_),
    .Y(_0748_));
 sky130_fd_sc_hd__nor2_1 _0913_ (.A(_0886_),
    .B(_0885_),
    .Y(_0749_));
 sky130_fd_sc_hd__a21oi_4 _0914_ (.A1(_0747_),
    .A2(_0748_),
    .B1(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__xor2_2 _0915_ (.A(_0883_),
    .B(_0750_),
    .X(_0751_));
 sky130_fd_sc_hd__nor3_1 _0916_ (.A(_0744_),
    .B(_0746_),
    .C(_0751_),
    .Y(net75));
 sky130_fd_sc_hd__buf_16 _0917_ (.A(net39),
    .X(_0752_));
 sky130_fd_sc_hd__buf_2 _0918_ (.A(mem_addr[3]),
    .X(_0753_));
 sky130_fd_sc_hd__nor4_4 _0919_ (.A(net37),
    .B(net36),
    .C(net38),
    .D(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__and3_1 _0920_ (.A(_0752_),
    .B(net72),
    .C(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__o32ai_4 _0921_ (.A1(_0744_),
    .A2(_0746_),
    .A3(_0751_),
    .B1(_0755_),
    .B2(net35),
    .Y(_0756_));
 sky130_fd_sc_hd__buf_6 _0922_ (.A(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__nor2b_1 _0923_ (.A(net38),
    .B_N(_0753_),
    .Y(_0758_));
 sky130_fd_sc_hd__nor2_1 _0924_ (.A(net37),
    .B(net36),
    .Y(_0759_));
 sky130_fd_sc_hd__o21a_1 _0925_ (.A1(net40),
    .A2(net51),
    .B1(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__and4_1 _0926_ (.A(_0752_),
    .B(net72),
    .C(_0758_),
    .D(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__buf_2 _0927_ (.A(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__clkbuf_8 _0928_ (.A(_0762_),
    .X(_0763_));
 sky130_fd_sc_hd__buf_4 _0929_ (.A(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__nand2b_4 _0930_ (.A_N(\wr_ptr[2] ),
    .B(net73),
    .Y(_0765_));
 sky130_fd_sc_hd__buf_2 _0931_ (.A(\wr_ptr[3] ),
    .X(_0766_));
 sky130_fd_sc_hd__nand2_2 _0932_ (.A(_0766_),
    .B(_0897_),
    .Y(_0767_));
 sky130_fd_sc_hd__nor4_4 _0933_ (.A(_0757_),
    .B(_0764_),
    .C(_0765_),
    .D(_0767_),
    .Y(_0007_));
 sky130_fd_sc_hd__nand2_4 _0934_ (.A(net73),
    .B(\wr_ptr[2] ),
    .Y(_0768_));
 sky130_fd_sc_hd__nor4_4 _0935_ (.A(_0757_),
    .B(_0764_),
    .C(_0767_),
    .D(_0768_),
    .Y(_0003_));
 sky130_fd_sc_hd__nor4_2 _0936_ (.A(_0766_),
    .B(_0756_),
    .C(_0762_),
    .D(_0765_),
    .Y(_0769_));
 sky130_fd_sc_hd__and2_4 _0937_ (.A(_0903_),
    .B(_0769_),
    .X(_0012_));
 sky130_fd_sc_hd__nand2_2 _0938_ (.A(_0766_),
    .B(_0903_),
    .Y(_0770_));
 sky130_fd_sc_hd__nor4_4 _0939_ (.A(_0757_),
    .B(_0763_),
    .C(_0765_),
    .D(_0770_),
    .Y(_0004_));
 sky130_fd_sc_hd__nor4_2 _0940_ (.A(_0766_),
    .B(_0756_),
    .C(_0762_),
    .D(_0768_),
    .Y(_0771_));
 sky130_fd_sc_hd__and2_4 _0941_ (.A(_0897_),
    .B(_0771_),
    .X(_0011_));
 sky130_fd_sc_hd__nand2_1 _0942_ (.A(_0766_),
    .B(_0899_),
    .Y(_0772_));
 sky130_fd_sc_hd__nor4_4 _0943_ (.A(_0757_),
    .B(_0763_),
    .C(_0765_),
    .D(_0772_),
    .Y(_0005_));
 sky130_fd_sc_hd__and2_4 _0944_ (.A(_0901_),
    .B(_0771_),
    .X(_0010_));
 sky130_fd_sc_hd__nand2_2 _0945_ (.A(_0766_),
    .B(_0901_),
    .Y(_0773_));
 sky130_fd_sc_hd__nor4_4 _0946_ (.A(_0757_),
    .B(_0763_),
    .C(_0765_),
    .D(_0773_),
    .Y(_0006_));
 sky130_fd_sc_hd__and2_4 _0947_ (.A(_0899_),
    .B(_0771_),
    .X(_0009_));
 sky130_fd_sc_hd__nor4_4 _0948_ (.A(_0757_),
    .B(_0763_),
    .C(_0768_),
    .D(_0773_),
    .Y(_0002_));
 sky130_fd_sc_hd__and2_4 _0949_ (.A(_0903_),
    .B(_0771_),
    .X(_0008_));
 sky130_fd_sc_hd__xor2_2 _0950_ (.A(_0886_),
    .B(_0874_),
    .X(_0774_));
 sky130_fd_sc_hd__nor3b_4 _0951_ (.A(_0875_),
    .B(_0774_),
    .C_N(_0878_),
    .Y(_0775_));
 sky130_fd_sc_hd__xnor2_4 _0952_ (.A(_0883_),
    .B(_0750_),
    .Y(_0776_));
 sky130_fd_sc_hd__nand3_2 _0953_ (.A(_0744_),
    .B(_0775_),
    .C(_0776_),
    .Y(_0777_));
 sky130_fd_sc_hd__inv_1 _0954_ (.A(_0777_),
    .Y(net74));
 sky130_fd_sc_hd__and2_4 _0955_ (.A(_0897_),
    .B(_0769_),
    .X(_0015_));
 sky130_fd_sc_hd__nor4_4 _0956_ (.A(_0757_),
    .B(_0763_),
    .C(_0768_),
    .D(_0770_),
    .Y(_0000_));
 sky130_fd_sc_hd__nor4_2 _0957_ (.A(_0757_),
    .B(_0763_),
    .C(_0768_),
    .D(_0772_),
    .Y(_0001_));
 sky130_fd_sc_hd__and2_4 _0958_ (.A(_0901_),
    .B(_0769_),
    .X(_0014_));
 sky130_fd_sc_hd__and2_4 _0959_ (.A(_0899_),
    .B(_0769_),
    .X(_0013_));
 sky130_fd_sc_hd__buf_8 _0960_ (.A(_0752_),
    .X(_0778_));
 sky130_fd_sc_hd__mux2_4 _0961_ (.A0(net33),
    .A1(net70),
    .S(_0778_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_4 _0962_ (.A0(net34),
    .A1(net71),
    .S(_0778_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_4 _0963_ (.A0(net4),
    .A1(net41),
    .S(_0778_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_4 _0964_ (.A0(net5),
    .A1(net42),
    .S(_0778_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_8 _0965_ (.A0(net6),
    .A1(net43),
    .S(_0778_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_8 _0966_ (.A0(net7),
    .A1(net44),
    .S(_0778_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_4 _0967_ (.A0(net8),
    .A1(net45),
    .S(_0778_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_8 _0968_ (.A0(net9),
    .A1(net46),
    .S(_0778_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_4 _0969_ (.A0(net10),
    .A1(net47),
    .S(_0778_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_4 _0970_ (.A0(net11),
    .A1(net48),
    .S(_0778_),
    .X(_0024_));
 sky130_fd_sc_hd__buf_16 _0971_ (.A(_0752_),
    .X(_0779_));
 sky130_fd_sc_hd__mux2_4 _0972_ (.A0(net12),
    .A1(net49),
    .S(_0779_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_4 _0973_ (.A0(net13),
    .A1(net50),
    .S(_0779_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_8 _0974_ (.A0(net15),
    .A1(net52),
    .S(_0779_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_4 _0975_ (.A0(net16),
    .A1(net53),
    .S(_0779_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_8 _0976_ (.A0(net17),
    .A1(net54),
    .S(_0779_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_4 _0977_ (.A0(net18),
    .A1(net55),
    .S(_0779_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_8 _0978_ (.A0(net19),
    .A1(net56),
    .S(_0779_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_4 _0979_ (.A0(net20),
    .A1(net57),
    .S(_0779_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_4 _0980_ (.A0(net21),
    .A1(net58),
    .S(_0779_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_8 _0981_ (.A0(net22),
    .A1(net59),
    .S(_0779_),
    .X(_0035_));
 sky130_fd_sc_hd__buf_16 _0982_ (.A(_0752_),
    .X(_0780_));
 sky130_fd_sc_hd__mux2_4 _0983_ (.A0(net23),
    .A1(net60),
    .S(_0780_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_4 _0984_ (.A0(net24),
    .A1(net61),
    .S(_0780_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_4 _0985_ (.A0(net26),
    .A1(net63),
    .S(_0780_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_8 _0986_ (.A0(net27),
    .A1(net64),
    .S(_0780_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_8 _0987_ (.A0(net3),
    .A1(net40),
    .S(_0780_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_8 _0988_ (.A0(net14),
    .A1(net51),
    .S(_0780_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_8 _0989_ (.A0(net25),
    .A1(net62),
    .S(_0780_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_4 _0990_ (.A0(net28),
    .A1(net65),
    .S(_0780_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_4 _0991_ (.A0(net29),
    .A1(net66),
    .S(_0780_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_8 _0992_ (.A0(net30),
    .A1(net67),
    .S(_0780_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_4 _0993_ (.A0(net31),
    .A1(net68),
    .S(_0752_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_4 _0994_ (.A0(net32),
    .A1(net69),
    .S(_0752_),
    .X(_0045_));
 sky130_fd_sc_hd__inv_1 _0995_ (.A(_0877_),
    .Y(_0873_));
 sky130_fd_sc_hd__buf_4 _0996_ (.A(\rd_ptr[3] ),
    .X(_0781_));
 sky130_fd_sc_hd__inv_1 _0997_ (.A(_0781_),
    .Y(_0782_));
 sky130_fd_sc_hd__buf_6 _0998_ (.A(_0782_),
    .X(_0783_));
 sky130_fd_sc_hd__buf_6 _0999_ (.A(_0783_),
    .X(_0881_));
 sky130_fd_sc_hd__buf_6 _1000_ (.A(\rd_ptr[2] ),
    .X(_0784_));
 sky130_fd_sc_hd__clkinv_4 _1001_ (.A(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__buf_6 _1002_ (.A(_0785_),
    .X(_0884_));
 sky130_fd_sc_hd__inv_1 _1003_ (.A(\rd_ptr[0] ),
    .Y(_0887_));
 sky130_fd_sc_hd__inv_1 _1004_ (.A(\wr_ptr[0] ),
    .Y(_0876_));
 sky130_fd_sc_hd__clkinvlp_4 _1005_ (.A(\rd_ptr[1] ),
    .Y(_0872_));
 sky130_fd_sc_hd__inv_1 _1006_ (.A(\wr_ptr[1] ),
    .Y(_0896_));
 sky130_fd_sc_hd__nor2b_2 _1007_ (.A(net72),
    .B_N(_0752_),
    .Y(_0786_));
 sky130_fd_sc_hd__a21oi_1 _1008_ (.A1(_0754_),
    .A2(_0786_),
    .B1(net2),
    .Y(_0787_));
 sky130_fd_sc_hd__a31oi_4 _1009_ (.A1(_0744_),
    .A2(_0775_),
    .A3(_0776_),
    .B1(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__nor2_4 _1010_ (.A(_0762_),
    .B(_0788_),
    .Y(_0789_));
 sky130_fd_sc_hd__buf_4 _1011_ (.A(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__nand4_4 _1012_ (.A(_0752_),
    .B(net72),
    .C(_0758_),
    .D(_0760_),
    .Y(_0791_));
 sky130_fd_sc_hd__and2_0 _1013_ (.A(_0791_),
    .B(_0788_),
    .X(_0792_));
 sky130_fd_sc_hd__clkbuf_4 _1014_ (.A(_0792_),
    .X(_0793_));
 sky130_fd_sc_hd__buf_6 _1015_ (.A(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__buf_4 _1016_ (.A(_0894_),
    .X(_0795_));
 sky130_fd_sc_hd__buf_6 _1017_ (.A(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__buf_2 _1018_ (.A(_0892_),
    .X(_0797_));
 sky130_fd_sc_hd__buf_4 _1019_ (.A(_0797_),
    .X(_0798_));
 sky130_fd_sc_hd__nand2b_1 _1020_ (.A_N(_0781_),
    .B(\rd_ptr[2] ),
    .Y(_0799_));
 sky130_fd_sc_hd__a221oi_1 _1021_ (.A1(_0796_),
    .A2(\mem[7][0] ),
    .B1(\mem[5][0] ),
    .B2(_0798_),
    .C1(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__buf_6 _1022_ (.A(_0888_),
    .X(_0801_));
 sky130_fd_sc_hd__buf_6 _1023_ (.A(_0801_),
    .X(_0802_));
 sky130_fd_sc_hd__buf_4 _1024_ (.A(_0890_),
    .X(_0803_));
 sky130_fd_sc_hd__buf_6 _1025_ (.A(_0803_),
    .X(_0804_));
 sky130_fd_sc_hd__a22oi_1 _1026_ (.A1(\mem[4][0] ),
    .A2(_0802_),
    .B1(_0804_),
    .B2(\mem[6][0] ),
    .Y(_0805_));
 sky130_fd_sc_hd__buf_6 _1027_ (.A(_0781_),
    .X(_0806_));
 sky130_fd_sc_hd__a222oi_1 _1028_ (.A1(_0894_),
    .A2(\mem[11][0] ),
    .B1(\mem[10][0] ),
    .B2(_0890_),
    .C1(_0797_),
    .C2(\mem[9][0] ),
    .Y(_0807_));
 sky130_fd_sc_hd__a21oi_1 _1029_ (.A1(\mem[8][0] ),
    .A2(_0801_),
    .B1(_0784_),
    .Y(_0808_));
 sky130_fd_sc_hd__and3_1 _1030_ (.A(_0806_),
    .B(_0807_),
    .C(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__a21oi_1 _1031_ (.A1(_0800_),
    .A2(_0805_),
    .B1(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__and2_0 _1032_ (.A(\rd_ptr[3] ),
    .B(\rd_ptr[2] ),
    .X(_0811_));
 sky130_fd_sc_hd__buf_4 _1033_ (.A(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__a22oi_1 _1034_ (.A1(_0796_),
    .A2(\mem[15][0] ),
    .B1(\mem[14][0] ),
    .B2(_0804_),
    .Y(_0813_));
 sky130_fd_sc_hd__buf_6 _1035_ (.A(_0797_),
    .X(_0814_));
 sky130_fd_sc_hd__a22oi_1 _1036_ (.A1(\mem[12][0] ),
    .A2(_0802_),
    .B1(_0814_),
    .B2(\mem[13][0] ),
    .Y(_0815_));
 sky130_fd_sc_hd__nand3_1 _1037_ (.A(_0812_),
    .B(_0813_),
    .C(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__buf_4 _1038_ (.A(_0803_),
    .X(_0817_));
 sky130_fd_sc_hd__a22oi_1 _1039_ (.A1(_0796_),
    .A2(\mem[3][0] ),
    .B1(\mem[2][0] ),
    .B2(_0817_),
    .Y(_0818_));
 sky130_fd_sc_hd__nor2_2 _1040_ (.A(_0781_),
    .B(_0784_),
    .Y(_0819_));
 sky130_fd_sc_hd__buf_4 _1041_ (.A(_0797_),
    .X(_0820_));
 sky130_fd_sc_hd__nand2_1 _1042_ (.A(\mem[1][0] ),
    .B(_0820_),
    .Y(_0821_));
 sky130_fd_sc_hd__nand3_1 _1043_ (.A(_0818_),
    .B(_0819_),
    .C(_0821_),
    .Y(_0822_));
 sky130_fd_sc_hd__or2_4 _1044_ (.A(\rd_ptr[3] ),
    .B(\rd_ptr[2] ),
    .X(_0823_));
 sky130_fd_sc_hd__a2111oi_4 _1045_ (.A1(_0888_),
    .A2(_0823_),
    .B1(_0890_),
    .C1(_0894_),
    .D1(_0797_),
    .Y(_0824_));
 sky130_fd_sc_hd__a32o_1 _1046_ (.A1(_0810_),
    .A2(_0816_),
    .A3(_0822_),
    .B1(_0824_),
    .B2(\mem[0][0] ),
    .X(_0825_));
 sky130_fd_sc_hd__a22o_1 _1047_ (.A1(net76),
    .A2(_0790_),
    .B1(_0794_),
    .B2(_0825_),
    .X(_0048_));
 sky130_fd_sc_hd__buf_4 _1048_ (.A(_0791_),
    .X(_0826_));
 sky130_fd_sc_hd__buf_6 _1049_ (.A(_0788_),
    .X(_0827_));
 sky130_fd_sc_hd__nand2_1 _1050_ (.A(_0826_),
    .B(_0827_),
    .Y(_0828_));
 sky130_fd_sc_hd__a2111o_4 _1051_ (.A1(_0888_),
    .A2(_0823_),
    .B1(_0803_),
    .C1(_0795_),
    .D1(_0797_),
    .X(_0829_));
 sky130_fd_sc_hd__buf_8 _1052_ (.A(_0829_),
    .X(_0830_));
 sky130_fd_sc_hd__buf_8 _1053_ (.A(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__buf_4 _1054_ (.A(_0806_),
    .X(_0832_));
 sky130_fd_sc_hd__buf_6 _1055_ (.A(_0832_),
    .X(_0833_));
 sky130_fd_sc_hd__buf_4 _1056_ (.A(\rd_ptr[2] ),
    .X(_0834_));
 sky130_fd_sc_hd__buf_8 _1057_ (.A(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__buf_6 _1058_ (.A(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__buf_6 _1059_ (.A(_0801_),
    .X(_0837_));
 sky130_fd_sc_hd__buf_8 _1060_ (.A(_0837_),
    .X(_0838_));
 sky130_fd_sc_hd__buf_8 _1061_ (.A(_0784_),
    .X(_0839_));
 sky130_fd_sc_hd__buf_6 _1062_ (.A(_0839_),
    .X(_0840_));
 sky130_fd_sc_hd__buf_8 _1063_ (.A(_0795_),
    .X(_0841_));
 sky130_fd_sc_hd__buf_6 _1064_ (.A(_0801_),
    .X(_0842_));
 sky130_fd_sc_hd__a22oi_1 _1065_ (.A1(_0841_),
    .A2(\mem[11][10] ),
    .B1(\mem[8][10] ),
    .B2(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hd__nor2_1 _1066_ (.A(_0840_),
    .B(_0843_),
    .Y(_0844_));
 sky130_fd_sc_hd__a31oi_1 _1067_ (.A1(_0836_),
    .A2(\mem[12][10] ),
    .A3(_0838_),
    .B1(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__nor2b_1 _1068_ (.A(\rd_ptr[2] ),
    .B_N(_0894_),
    .Y(_0846_));
 sky130_fd_sc_hd__buf_4 _1069_ (.A(_0846_),
    .X(_0847_));
 sky130_fd_sc_hd__buf_4 _1070_ (.A(_0785_),
    .X(_0848_));
 sky130_fd_sc_hd__buf_6 _1071_ (.A(_0795_),
    .X(_0849_));
 sky130_fd_sc_hd__buf_8 _1072_ (.A(_0801_),
    .X(_0850_));
 sky130_fd_sc_hd__buf_6 _1073_ (.A(_0803_),
    .X(_0851_));
 sky130_fd_sc_hd__a222oi_1 _1074_ (.A1(_0849_),
    .A2(\mem[7][10] ),
    .B1(\mem[4][10] ),
    .B2(_0850_),
    .C1(_0851_),
    .C2(\mem[6][10] ),
    .Y(_0852_));
 sky130_fd_sc_hd__nor2_1 _1075_ (.A(_0848_),
    .B(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__a211oi_1 _1076_ (.A1(\mem[3][10] ),
    .A2(_0847_),
    .B1(_0853_),
    .C1(_0833_),
    .Y(_0854_));
 sky130_fd_sc_hd__a21oi_1 _1077_ (.A1(_0833_),
    .A2(_0845_),
    .B1(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__nand2_1 _1078_ (.A(_0781_),
    .B(_0784_),
    .Y(_0856_));
 sky130_fd_sc_hd__buf_8 _1079_ (.A(_0856_),
    .X(_0857_));
 sky130_fd_sc_hd__buf_4 _1080_ (.A(_0849_),
    .X(_0858_));
 sky130_fd_sc_hd__buf_6 _1081_ (.A(_0803_),
    .X(_0859_));
 sky130_fd_sc_hd__buf_6 _1082_ (.A(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__a22oi_1 _1083_ (.A1(_0858_),
    .A2(\mem[15][10] ),
    .B1(\mem[14][10] ),
    .B2(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hd__buf_6 _1084_ (.A(_0798_),
    .X(_0862_));
 sky130_fd_sc_hd__buf_8 _1085_ (.A(_0862_),
    .X(_0863_));
 sky130_fd_sc_hd__nor2b_1 _1086_ (.A(\rd_ptr[3] ),
    .B_N(\rd_ptr[2] ),
    .Y(_0864_));
 sky130_fd_sc_hd__buf_8 _1087_ (.A(_0864_),
    .X(_0865_));
 sky130_fd_sc_hd__buf_8 _1088_ (.A(_0865_),
    .X(_0866_));
 sky130_fd_sc_hd__buf_8 _1089_ (.A(_0834_),
    .X(_0867_));
 sky130_fd_sc_hd__mux2i_1 _1090_ (.A0(\mem[9][10] ),
    .A1(\mem[13][10] ),
    .S(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__buf_6 _1091_ (.A(_0782_),
    .X(_0869_));
 sky130_fd_sc_hd__o2bb2ai_1 _1092_ (.A1_N(\mem[5][10] ),
    .A2_N(_0866_),
    .B1(_0868_),
    .B2(_0869_),
    .Y(_0870_));
 sky130_fd_sc_hd__nand2_1 _1093_ (.A(_0863_),
    .B(_0870_),
    .Y(_0871_));
 sky130_fd_sc_hd__buf_6 _1094_ (.A(_0781_),
    .X(_0122_));
 sky130_fd_sc_hd__buf_6 _1095_ (.A(_0122_),
    .X(_0123_));
 sky130_fd_sc_hd__buf_6 _1096_ (.A(_0804_),
    .X(_0124_));
 sky130_fd_sc_hd__a22oi_1 _1097_ (.A1(\mem[2][10] ),
    .A2(_0124_),
    .B1(_0862_),
    .B2(\mem[1][10] ),
    .Y(_0125_));
 sky130_fd_sc_hd__nand3_1 _1098_ (.A(_0123_),
    .B(\mem[10][10] ),
    .C(_0860_),
    .Y(_0126_));
 sky130_fd_sc_hd__o21ai_0 _1099_ (.A1(_0123_),
    .A2(_0125_),
    .B1(_0126_),
    .Y(_0127_));
 sky130_fd_sc_hd__nand2_1 _1100_ (.A(_0884_),
    .B(_0127_),
    .Y(_0128_));
 sky130_fd_sc_hd__buf_8 _1101_ (.A(_0830_),
    .X(_0129_));
 sky130_fd_sc_hd__o2111ai_2 _1102_ (.A1(_0857_),
    .A2(_0861_),
    .B1(_0871_),
    .C1(_0128_),
    .D1(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hd__o22ai_4 _1103_ (.A1(\mem[0][10] ),
    .A2(_0831_),
    .B1(_0855_),
    .B2(_0130_),
    .Y(_0131_));
 sky130_fd_sc_hd__o2bb2ai_1 _1104_ (.A1_N(net77),
    .A2_N(_0790_),
    .B1(_0828_),
    .B2(_0131_),
    .Y(_0049_));
 sky130_fd_sc_hd__buf_8 _1105_ (.A(_0824_),
    .X(_0132_));
 sky130_fd_sc_hd__buf_8 _1106_ (.A(_0806_),
    .X(_0133_));
 sky130_fd_sc_hd__buf_6 _1107_ (.A(_0801_),
    .X(_0134_));
 sky130_fd_sc_hd__a32oi_1 _1108_ (.A1(_0867_),
    .A2(\mem[4][11] ),
    .A3(_0134_),
    .B1(_0847_),
    .B2(\mem[3][11] ),
    .Y(_0135_));
 sky130_fd_sc_hd__buf_8 _1109_ (.A(_0795_),
    .X(_0136_));
 sky130_fd_sc_hd__buf_6 _1110_ (.A(_0798_),
    .X(_0137_));
 sky130_fd_sc_hd__a222oi_1 _1111_ (.A1(_0136_),
    .A2(\mem[15][11] ),
    .B1(\mem[12][11] ),
    .B2(_0850_),
    .C1(_0137_),
    .C2(\mem[13][11] ),
    .Y(_0138_));
 sky130_fd_sc_hd__o22ai_1 _1112_ (.A1(_0133_),
    .A2(_0135_),
    .B1(_0138_),
    .B2(_0857_),
    .Y(_0139_));
 sky130_fd_sc_hd__buf_6 _1113_ (.A(_0798_),
    .X(_0140_));
 sky130_fd_sc_hd__and3_1 _1114_ (.A(_0781_),
    .B(\mem[14][11] ),
    .C(_0803_),
    .X(_0141_));
 sky130_fd_sc_hd__a31oi_2 _1115_ (.A1(_0782_),
    .A2(\mem[5][11] ),
    .A3(_0140_),
    .B1(_0141_),
    .Y(_0142_));
 sky130_fd_sc_hd__buf_6 _1116_ (.A(_0803_),
    .X(_0143_));
 sky130_fd_sc_hd__nand2b_1 _1117_ (.A_N(\rd_ptr[2] ),
    .B(\rd_ptr[3] ),
    .Y(_0144_));
 sky130_fd_sc_hd__buf_8 _1118_ (.A(_0144_),
    .X(_0145_));
 sky130_fd_sc_hd__a221oi_1 _1119_ (.A1(\mem[8][11] ),
    .A2(_0850_),
    .B1(_0143_),
    .B2(\mem[10][11] ),
    .C1(_0145_),
    .Y(_0146_));
 sky130_fd_sc_hd__a221oi_1 _1120_ (.A1(\mem[2][11] ),
    .A2(_0143_),
    .B1(_0137_),
    .B2(\mem[1][11] ),
    .C1(_0823_),
    .Y(_0147_));
 sky130_fd_sc_hd__a211oi_1 _1121_ (.A1(_0840_),
    .A2(_0142_),
    .B1(_0146_),
    .C1(_0147_),
    .Y(_0148_));
 sky130_fd_sc_hd__buf_6 _1122_ (.A(_0796_),
    .X(_0149_));
 sky130_fd_sc_hd__buf_6 _1123_ (.A(_0798_),
    .X(_0150_));
 sky130_fd_sc_hd__a22oi_1 _1124_ (.A1(_0149_),
    .A2(\mem[11][11] ),
    .B1(\mem[9][11] ),
    .B2(_0150_),
    .Y(_0151_));
 sky130_fd_sc_hd__buf_4 _1125_ (.A(_0817_),
    .X(_0152_));
 sky130_fd_sc_hd__a22oi_1 _1126_ (.A1(_0858_),
    .A2(\mem[7][11] ),
    .B1(\mem[6][11] ),
    .B2(_0152_),
    .Y(_0153_));
 sky130_fd_sc_hd__buf_8 _1127_ (.A(_0799_),
    .X(_0154_));
 sky130_fd_sc_hd__o22ai_1 _1128_ (.A1(_0145_),
    .A2(_0151_),
    .B1(_0153_),
    .B2(_0154_),
    .Y(_0155_));
 sky130_fd_sc_hd__nor4_1 _1129_ (.A(_0132_),
    .B(_0139_),
    .C(_0148_),
    .D(_0155_),
    .Y(_0156_));
 sky130_fd_sc_hd__buf_16 _1130_ (.A(_0830_),
    .X(_0157_));
 sky130_fd_sc_hd__nor2_1 _1131_ (.A(\mem[0][11] ),
    .B(_0157_),
    .Y(_0158_));
 sky130_fd_sc_hd__nor2_2 _1132_ (.A(_0156_),
    .B(_0158_),
    .Y(_0159_));
 sky130_fd_sc_hd__a22o_1 _1133_ (.A1(net78),
    .A2(_0790_),
    .B1(_0794_),
    .B2(_0159_),
    .X(_0050_));
 sky130_fd_sc_hd__nor2b_4 _1134_ (.A(_0784_),
    .B_N(_0781_),
    .Y(_0160_));
 sky130_fd_sc_hd__a22o_1 _1135_ (.A1(\mem[9][12] ),
    .A2(_0160_),
    .B1(_0866_),
    .B2(\mem[5][12] ),
    .X(_0161_));
 sky130_fd_sc_hd__buf_6 _1136_ (.A(_0122_),
    .X(_0162_));
 sky130_fd_sc_hd__buf_8 _1137_ (.A(_0804_),
    .X(_0163_));
 sky130_fd_sc_hd__a32oi_1 _1138_ (.A1(_0835_),
    .A2(\mem[6][12] ),
    .A3(_0163_),
    .B1(_0847_),
    .B2(\mem[3][12] ),
    .Y(_0164_));
 sky130_fd_sc_hd__nand2_8 _1139_ (.A(_0785_),
    .B(_0851_),
    .Y(_0165_));
 sky130_fd_sc_hd__buf_8 _1140_ (.A(_0806_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2i_1 _1141_ (.A0(\mem[2][12] ),
    .A1(\mem[10][12] ),
    .S(_0166_),
    .Y(_0167_));
 sky130_fd_sc_hd__nand3_1 _1142_ (.A(\mem[4][12] ),
    .B(_0838_),
    .C(_0866_),
    .Y(_0168_));
 sky130_fd_sc_hd__o221ai_2 _1143_ (.A1(_0162_),
    .A2(_0164_),
    .B1(_0165_),
    .B2(_0167_),
    .C1(_0168_),
    .Y(_0169_));
 sky130_fd_sc_hd__a21oi_1 _1144_ (.A1(_0863_),
    .A2(_0161_),
    .B1(_0169_),
    .Y(_0170_));
 sky130_fd_sc_hd__buf_6 _1145_ (.A(_0819_),
    .X(_0171_));
 sky130_fd_sc_hd__nand3_1 _1146_ (.A(\mem[1][12] ),
    .B(_0150_),
    .C(_0171_),
    .Y(_0172_));
 sky130_fd_sc_hd__buf_4 _1147_ (.A(_0802_),
    .X(_0173_));
 sky130_fd_sc_hd__buf_6 _1148_ (.A(_0160_),
    .X(_0174_));
 sky130_fd_sc_hd__nand3_1 _1149_ (.A(\mem[8][12] ),
    .B(_0173_),
    .C(_0174_),
    .Y(_0175_));
 sky130_fd_sc_hd__nand2_1 _1150_ (.A(_0172_),
    .B(_0175_),
    .Y(_0176_));
 sky130_fd_sc_hd__nand3_1 _1151_ (.A(_0858_),
    .B(\mem[7][12] ),
    .C(_0866_),
    .Y(_0177_));
 sky130_fd_sc_hd__buf_6 _1152_ (.A(_0812_),
    .X(_0178_));
 sky130_fd_sc_hd__nand3_1 _1153_ (.A(\mem[13][12] ),
    .B(_0150_),
    .C(_0178_),
    .Y(_0179_));
 sky130_fd_sc_hd__nand2_1 _1154_ (.A(_0177_),
    .B(_0179_),
    .Y(_0180_));
 sky130_fd_sc_hd__buf_8 _1155_ (.A(_0801_),
    .X(_0181_));
 sky130_fd_sc_hd__buf_6 _1156_ (.A(_0804_),
    .X(_0182_));
 sky130_fd_sc_hd__a22oi_1 _1157_ (.A1(\mem[12][12] ),
    .A2(_0181_),
    .B1(_0182_),
    .B2(\mem[14][12] ),
    .Y(_0183_));
 sky130_fd_sc_hd__nand2_1 _1158_ (.A(_0133_),
    .B(_0858_),
    .Y(_0184_));
 sky130_fd_sc_hd__mux2i_1 _1159_ (.A0(\mem[11][12] ),
    .A1(\mem[15][12] ),
    .S(_0835_),
    .Y(_0185_));
 sky130_fd_sc_hd__o22ai_1 _1160_ (.A1(_0857_),
    .A2(_0183_),
    .B1(_0184_),
    .B2(_0185_),
    .Y(_0186_));
 sky130_fd_sc_hd__nor4_1 _1161_ (.A(_0132_),
    .B(_0176_),
    .C(_0180_),
    .D(_0186_),
    .Y(_0187_));
 sky130_fd_sc_hd__nor2_1 _1162_ (.A(\mem[0][12] ),
    .B(_0129_),
    .Y(_0188_));
 sky130_fd_sc_hd__a21oi_1 _1163_ (.A1(_0170_),
    .A2(_0187_),
    .B1(_0188_),
    .Y(_0189_));
 sky130_fd_sc_hd__a22o_1 _1164_ (.A1(net79),
    .A2(_0790_),
    .B1(_0794_),
    .B2(_0189_),
    .X(_0051_));
 sky130_fd_sc_hd__a222oi_1 _1165_ (.A1(\mem[14][13] ),
    .A2(_0859_),
    .B1(_0137_),
    .B2(\mem[13][13] ),
    .C1(\mem[12][13] ),
    .C2(_0181_),
    .Y(_0190_));
 sky130_fd_sc_hd__nand3_1 _1166_ (.A(_0848_),
    .B(\mem[8][13] ),
    .C(_0173_),
    .Y(_0191_));
 sky130_fd_sc_hd__o21ai_0 _1167_ (.A1(_0848_),
    .A2(_0190_),
    .B1(_0191_),
    .Y(_0192_));
 sky130_fd_sc_hd__buf_8 _1168_ (.A(_0814_),
    .X(_0193_));
 sky130_fd_sc_hd__a22oi_1 _1169_ (.A1(\mem[6][13] ),
    .A2(_0182_),
    .B1(_0193_),
    .B2(\mem[5][13] ),
    .Y(_0194_));
 sky130_fd_sc_hd__o21ai_0 _1170_ (.A1(_0154_),
    .A2(_0194_),
    .B1(_0830_),
    .Y(_0195_));
 sky130_fd_sc_hd__a21oi_1 _1171_ (.A1(_0833_),
    .A2(_0192_),
    .B1(_0195_),
    .Y(_0196_));
 sky130_fd_sc_hd__buf_6 _1172_ (.A(_0839_),
    .X(_0197_));
 sky130_fd_sc_hd__clkbuf_8 _1173_ (.A(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__buf_6 _1174_ (.A(_0781_),
    .X(_0199_));
 sky130_fd_sc_hd__clkbuf_8 _1175_ (.A(_0199_),
    .X(_0200_));
 sky130_fd_sc_hd__nand2_1 _1176_ (.A(_0858_),
    .B(\mem[15][13] ),
    .Y(_0201_));
 sky130_fd_sc_hd__a221oi_1 _1177_ (.A1(_0841_),
    .A2(\mem[7][13] ),
    .B1(\mem[4][13] ),
    .B2(_0181_),
    .C1(_0832_),
    .Y(_0202_));
 sky130_fd_sc_hd__a21oi_1 _1178_ (.A1(_0200_),
    .A2(_0201_),
    .B1(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__a222oi_1 _1179_ (.A1(_0796_),
    .A2(\mem[11][13] ),
    .B1(\mem[10][13] ),
    .B2(_0804_),
    .C1(_0820_),
    .C2(\mem[9][13] ),
    .Y(_0204_));
 sky130_fd_sc_hd__a22oi_2 _1180_ (.A1(_0841_),
    .A2(\mem[3][13] ),
    .B1(\mem[2][13] ),
    .B2(_0124_),
    .Y(_0205_));
 sky130_fd_sc_hd__a21oi_1 _1181_ (.A1(\mem[1][13] ),
    .A2(_0137_),
    .B1(_0166_),
    .Y(_0206_));
 sky130_fd_sc_hd__buf_16 _1182_ (.A(_0834_),
    .X(_0207_));
 sky130_fd_sc_hd__buf_6 _1183_ (.A(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__a221oi_4 _1184_ (.A1(_0133_),
    .A2(_0204_),
    .B1(_0205_),
    .B2(_0206_),
    .C1(_0208_),
    .Y(_0209_));
 sky130_fd_sc_hd__a21oi_1 _1185_ (.A1(_0198_),
    .A2(_0203_),
    .B1(_0209_),
    .Y(_0210_));
 sky130_fd_sc_hd__nor2_1 _1186_ (.A(\mem[0][13] ),
    .B(_0129_),
    .Y(_0211_));
 sky130_fd_sc_hd__a21oi_4 _1187_ (.A1(_0196_),
    .A2(_0210_),
    .B1(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__a22o_1 _1188_ (.A1(net80),
    .A2(_0790_),
    .B1(_0794_),
    .B2(_0212_),
    .X(_0052_));
 sky130_fd_sc_hd__nor2_1 _1189_ (.A(\mem[0][14] ),
    .B(_0830_),
    .Y(_0213_));
 sky130_fd_sc_hd__mux2i_1 _1190_ (.A0(\mem[9][14] ),
    .A1(\mem[13][14] ),
    .S(_0839_),
    .Y(_0214_));
 sky130_fd_sc_hd__nand2_1 _1191_ (.A(\mem[5][14] ),
    .B(_0865_),
    .Y(_0215_));
 sky130_fd_sc_hd__o21ai_0 _1192_ (.A1(_0783_),
    .A2(_0214_),
    .B1(_0215_),
    .Y(_0216_));
 sky130_fd_sc_hd__a22o_1 _1193_ (.A1(\mem[15][14] ),
    .A2(_0812_),
    .B1(_0171_),
    .B2(\mem[3][14] ),
    .X(_0217_));
 sky130_fd_sc_hd__buf_6 _1194_ (.A(_0841_),
    .X(_0218_));
 sky130_fd_sc_hd__a221oi_1 _1195_ (.A1(_0193_),
    .A2(_0216_),
    .B1(_0217_),
    .B2(_0218_),
    .C1(_0132_),
    .Y(_0219_));
 sky130_fd_sc_hd__a221o_1 _1196_ (.A1(\mem[12][14] ),
    .A2(_0842_),
    .B1(_0152_),
    .B2(\mem[14][14] ),
    .C1(_0783_),
    .X(_0220_));
 sky130_fd_sc_hd__a21oi_1 _1197_ (.A1(\mem[4][14] ),
    .A2(_0173_),
    .B1(_0123_),
    .Y(_0221_));
 sky130_fd_sc_hd__a22oi_1 _1198_ (.A1(_0858_),
    .A2(\mem[7][14] ),
    .B1(\mem[6][14] ),
    .B2(_0152_),
    .Y(_0222_));
 sky130_fd_sc_hd__a21oi_1 _1199_ (.A1(_0221_),
    .A2(_0222_),
    .B1(_0884_),
    .Y(_0223_));
 sky130_fd_sc_hd__buf_4 _1200_ (.A(_0795_),
    .X(_0224_));
 sky130_fd_sc_hd__a222oi_1 _1201_ (.A1(_0224_),
    .A2(\mem[11][14] ),
    .B1(\mem[8][14] ),
    .B2(_0837_),
    .C1(_0182_),
    .C2(\mem[10][14] ),
    .Y(_0225_));
 sky130_fd_sc_hd__buf_6 _1202_ (.A(_0798_),
    .X(_0226_));
 sky130_fd_sc_hd__a221oi_1 _1203_ (.A1(\mem[2][14] ),
    .A2(_0163_),
    .B1(_0226_),
    .B2(\mem[1][14] ),
    .C1(_0832_),
    .Y(_0227_));
 sky130_fd_sc_hd__a211oi_1 _1204_ (.A1(_0200_),
    .A2(_0225_),
    .B1(_0227_),
    .C1(_0198_),
    .Y(_0228_));
 sky130_fd_sc_hd__a21oi_1 _1205_ (.A1(_0220_),
    .A2(_0223_),
    .B1(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__o21ai_2 _1206_ (.A1(_0213_),
    .A2(_0219_),
    .B1(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__a22o_1 _1207_ (.A1(net81),
    .A2(_0790_),
    .B1(_0794_),
    .B2(_0230_),
    .X(_0053_));
 sky130_fd_sc_hd__clkbuf_4 _1208_ (.A(_0827_),
    .X(_0231_));
 sky130_fd_sc_hd__nand2_1 _1209_ (.A(net82),
    .B(_0826_),
    .Y(_0232_));
 sky130_fd_sc_hd__a22oi_1 _1210_ (.A1(\mem[14][15] ),
    .A2(_0124_),
    .B1(_0862_),
    .B2(\mem[13][15] ),
    .Y(_0233_));
 sky130_fd_sc_hd__buf_6 _1211_ (.A(_0839_),
    .X(_0234_));
 sky130_fd_sc_hd__a21oi_1 _1212_ (.A1(_0858_),
    .A2(\mem[11][15] ),
    .B1(_0234_),
    .Y(_0235_));
 sky130_fd_sc_hd__a211oi_1 _1213_ (.A1(_0836_),
    .A2(_0233_),
    .B1(_0235_),
    .C1(_0881_),
    .Y(_0236_));
 sky130_fd_sc_hd__nor2_1 _1214_ (.A(_0132_),
    .B(_0236_),
    .Y(_0237_));
 sky130_fd_sc_hd__nand2_1 _1215_ (.A(\mem[2][15] ),
    .B(_0152_),
    .Y(_0238_));
 sky130_fd_sc_hd__nand3_1 _1216_ (.A(_0133_),
    .B(\mem[8][15] ),
    .C(_0173_),
    .Y(_0239_));
 sky130_fd_sc_hd__o21ai_0 _1217_ (.A1(_0123_),
    .A2(_0238_),
    .B1(_0239_),
    .Y(_0240_));
 sky130_fd_sc_hd__a32oi_1 _1218_ (.A1(_0218_),
    .A2(\mem[7][15] ),
    .A3(_0866_),
    .B1(_0240_),
    .B2(_0884_),
    .Y(_0241_));
 sky130_fd_sc_hd__nor2b_1 _1219_ (.A(\rd_ptr[3] ),
    .B_N(_0894_),
    .Y(_0242_));
 sky130_fd_sc_hd__buf_6 _1220_ (.A(_0242_),
    .X(_0243_));
 sky130_fd_sc_hd__a32oi_1 _1221_ (.A1(_0122_),
    .A2(\mem[10][15] ),
    .A3(_0143_),
    .B1(_0243_),
    .B2(\mem[3][15] ),
    .Y(_0244_));
 sky130_fd_sc_hd__buf_6 _1222_ (.A(_0801_),
    .X(_0245_));
 sky130_fd_sc_hd__a221oi_1 _1223_ (.A1(\mem[4][15] ),
    .A2(_0245_),
    .B1(_0851_),
    .B2(\mem[6][15] ),
    .C1(_0154_),
    .Y(_0246_));
 sky130_fd_sc_hd__buf_6 _1224_ (.A(_0795_),
    .X(_0247_));
 sky130_fd_sc_hd__a221oi_1 _1225_ (.A1(_0247_),
    .A2(\mem[15][15] ),
    .B1(\mem[12][15] ),
    .B2(_0134_),
    .C1(_0857_),
    .Y(_0248_));
 sky130_fd_sc_hd__a211o_1 _1226_ (.A1(_0848_),
    .A2(_0244_),
    .B1(_0246_),
    .C1(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2i_1 _1227_ (.A0(\mem[1][15] ),
    .A1(\mem[5][15] ),
    .S(_0835_),
    .Y(_0250_));
 sky130_fd_sc_hd__nor2_1 _1228_ (.A(_0162_),
    .B(_0250_),
    .Y(_0251_));
 sky130_fd_sc_hd__and2_0 _1229_ (.A(\mem[9][15] ),
    .B(_0174_),
    .X(_0252_));
 sky130_fd_sc_hd__o21ai_0 _1230_ (.A1(_0251_),
    .A2(_0252_),
    .B1(_0863_),
    .Y(_0253_));
 sky130_fd_sc_hd__nand4_1 _1231_ (.A(_0237_),
    .B(_0241_),
    .C(_0249_),
    .D(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hd__o2111ai_1 _1232_ (.A1(\mem[0][15] ),
    .A2(_0831_),
    .B1(_0254_),
    .C1(_0826_),
    .D1(_0231_),
    .Y(_0255_));
 sky130_fd_sc_hd__o21ai_0 _1233_ (.A1(_0231_),
    .A2(_0232_),
    .B1(_0255_),
    .Y(_0054_));
 sky130_fd_sc_hd__a222oi_1 _1234_ (.A1(_0136_),
    .A2(\mem[15][16] ),
    .B1(\mem[12][16] ),
    .B2(_0850_),
    .C1(_0851_),
    .C2(\mem[14][16] ),
    .Y(_0256_));
 sky130_fd_sc_hd__nand2_1 _1235_ (.A(_0208_),
    .B(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__a22oi_1 _1236_ (.A1(_0224_),
    .A2(\mem[11][16] ),
    .B1(\mem[8][16] ),
    .B2(_0837_),
    .Y(_0258_));
 sky130_fd_sc_hd__a21oi_1 _1237_ (.A1(\mem[10][16] ),
    .A2(_0143_),
    .B1(_0867_),
    .Y(_0259_));
 sky130_fd_sc_hd__a21oi_1 _1238_ (.A1(_0258_),
    .A2(_0259_),
    .B1(_0783_),
    .Y(_0260_));
 sky130_fd_sc_hd__mux2i_1 _1239_ (.A0(\mem[9][16] ),
    .A1(\mem[13][16] ),
    .S(_0839_),
    .Y(_0261_));
 sky130_fd_sc_hd__nand2_1 _1240_ (.A(\mem[5][16] ),
    .B(_0865_),
    .Y(_0262_));
 sky130_fd_sc_hd__o21ai_0 _1241_ (.A1(_0783_),
    .A2(_0261_),
    .B1(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__a222oi_1 _1242_ (.A1(_0796_),
    .A2(\mem[7][16] ),
    .B1(\mem[4][16] ),
    .B2(_0801_),
    .C1(_0817_),
    .C2(\mem[6][16] ),
    .Y(_0264_));
 sky130_fd_sc_hd__a22oi_1 _1243_ (.A1(_0136_),
    .A2(\mem[3][16] ),
    .B1(\mem[1][16] ),
    .B2(_0820_),
    .Y(_0265_));
 sky130_fd_sc_hd__a21oi_1 _1244_ (.A1(\mem[2][16] ),
    .A2(_0143_),
    .B1(_0207_),
    .Y(_0266_));
 sky130_fd_sc_hd__a221oi_2 _1245_ (.A1(_0197_),
    .A2(_0264_),
    .B1(_0265_),
    .B2(_0266_),
    .C1(_0133_),
    .Y(_0267_));
 sky130_fd_sc_hd__a221oi_2 _1246_ (.A1(_0257_),
    .A2(_0260_),
    .B1(_0263_),
    .B2(_0193_),
    .C1(_0267_),
    .Y(_0268_));
 sky130_fd_sc_hd__nor2_1 _1247_ (.A(\mem[0][16] ),
    .B(_0129_),
    .Y(_0269_));
 sky130_fd_sc_hd__a21oi_4 _1248_ (.A1(_0831_),
    .A2(_0268_),
    .B1(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__a22o_1 _1249_ (.A1(net83),
    .A2(_0790_),
    .B1(_0794_),
    .B2(_0270_),
    .X(_0055_));
 sky130_fd_sc_hd__a22oi_1 _1250_ (.A1(\mem[8][17] ),
    .A2(_0134_),
    .B1(_0124_),
    .B2(\mem[10][17] ),
    .Y(_0271_));
 sky130_fd_sc_hd__and2_2 _1251_ (.A(_0834_),
    .B(_0795_),
    .X(_0272_));
 sky130_fd_sc_hd__nand2_1 _1252_ (.A(\mem[15][17] ),
    .B(_0272_),
    .Y(_0273_));
 sky130_fd_sc_hd__o21ai_0 _1253_ (.A1(_0234_),
    .A2(_0271_),
    .B1(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__nand3_1 _1254_ (.A(_0234_),
    .B(\mem[5][17] ),
    .C(_0150_),
    .Y(_0275_));
 sky130_fd_sc_hd__buf_4 _1255_ (.A(_0785_),
    .X(_0276_));
 sky130_fd_sc_hd__nand3_1 _1256_ (.A(_0276_),
    .B(\mem[2][17] ),
    .C(_0182_),
    .Y(_0277_));
 sky130_fd_sc_hd__a21oi_1 _1257_ (.A1(_0275_),
    .A2(_0277_),
    .B1(_0200_),
    .Y(_0278_));
 sky130_fd_sc_hd__nand2_1 _1258_ (.A(_0276_),
    .B(_0150_),
    .Y(_0279_));
 sky130_fd_sc_hd__mux2i_1 _1259_ (.A0(\mem[1][17] ),
    .A1(\mem[9][17] ),
    .S(_0199_),
    .Y(_0280_));
 sky130_fd_sc_hd__mux2i_1 _1260_ (.A0(\mem[3][17] ),
    .A1(\mem[11][17] ),
    .S(_0199_),
    .Y(_0281_));
 sky130_fd_sc_hd__nand2_1 _1261_ (.A(_0276_),
    .B(_0149_),
    .Y(_0282_));
 sky130_fd_sc_hd__o22ai_1 _1262_ (.A1(_0279_),
    .A2(_0280_),
    .B1(_0281_),
    .B2(_0282_),
    .Y(_0283_));
 sky130_fd_sc_hd__a211oi_2 _1263_ (.A1(_0833_),
    .A2(_0274_),
    .B1(_0278_),
    .C1(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__a222oi_1 _1264_ (.A1(\mem[14][17] ),
    .A2(_0163_),
    .B1(_0226_),
    .B2(\mem[13][17] ),
    .C1(\mem[12][17] ),
    .C2(_0842_),
    .Y(_0285_));
 sky130_fd_sc_hd__nand2_1 _1265_ (.A(_0833_),
    .B(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__a222oi_1 _1266_ (.A1(_0136_),
    .A2(\mem[7][17] ),
    .B1(\mem[4][17] ),
    .B2(_0245_),
    .C1(_0124_),
    .C2(\mem[6][17] ),
    .Y(_0287_));
 sky130_fd_sc_hd__a21oi_1 _1267_ (.A1(_0869_),
    .A2(_0287_),
    .B1(_0884_),
    .Y(_0288_));
 sky130_fd_sc_hd__a21oi_1 _1268_ (.A1(_0286_),
    .A2(_0288_),
    .B1(_0132_),
    .Y(_0289_));
 sky130_fd_sc_hd__nor2_1 _1269_ (.A(\mem[0][17] ),
    .B(_0129_),
    .Y(_0290_));
 sky130_fd_sc_hd__a21oi_4 _1270_ (.A1(_0284_),
    .A2(_0289_),
    .B1(_0290_),
    .Y(_0291_));
 sky130_fd_sc_hd__a22o_1 _1271_ (.A1(net84),
    .A2(_0790_),
    .B1(_0794_),
    .B2(_0291_),
    .X(_0056_));
 sky130_fd_sc_hd__a22oi_2 _1272_ (.A1(\mem[8][18] ),
    .A2(_0134_),
    .B1(_0163_),
    .B2(\mem[10][18] ),
    .Y(_0292_));
 sky130_fd_sc_hd__a21oi_1 _1273_ (.A1(_0149_),
    .A2(\mem[3][18] ),
    .B1(_0832_),
    .Y(_0293_));
 sky130_fd_sc_hd__a211oi_1 _1274_ (.A1(_0123_),
    .A2(_0292_),
    .B1(_0293_),
    .C1(_0208_),
    .Y(_0294_));
 sky130_fd_sc_hd__a22oi_1 _1275_ (.A1(\mem[12][18] ),
    .A2(_0134_),
    .B1(_0226_),
    .B2(\mem[13][18] ),
    .Y(_0295_));
 sky130_fd_sc_hd__a21oi_1 _1276_ (.A1(_0149_),
    .A2(\mem[11][18] ),
    .B1(_0197_),
    .Y(_0296_));
 sky130_fd_sc_hd__a211oi_1 _1277_ (.A1(_0208_),
    .A2(_0295_),
    .B1(_0296_),
    .C1(_0869_),
    .Y(_0297_));
 sky130_fd_sc_hd__nor2_1 _1278_ (.A(_0294_),
    .B(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__mux2i_2 _1279_ (.A0(\mem[2][18] ),
    .A1(\mem[6][18] ),
    .S(_0207_),
    .Y(_0299_));
 sky130_fd_sc_hd__nand2_1 _1280_ (.A(\mem[14][18] ),
    .B(_0178_),
    .Y(_0300_));
 sky130_fd_sc_hd__o21ai_0 _1281_ (.A1(_0133_),
    .A2(_0299_),
    .B1(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__a222oi_1 _1282_ (.A1(_0224_),
    .A2(\mem[7][18] ),
    .B1(\mem[4][18] ),
    .B2(_0245_),
    .C1(_0226_),
    .C2(\mem[5][18] ),
    .Y(_0302_));
 sky130_fd_sc_hd__and3_2 _1283_ (.A(_0806_),
    .B(_0834_),
    .C(_0796_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _1284_ (.A0(\mem[1][18] ),
    .A1(\mem[9][18] ),
    .S(_0781_),
    .X(_0304_));
 sky130_fd_sc_hd__nor2b_2 _1285_ (.A(_0834_),
    .B_N(_0798_),
    .Y(_0305_));
 sky130_fd_sc_hd__a22oi_1 _1286_ (.A1(\mem[15][18] ),
    .A2(_0303_),
    .B1(_0304_),
    .B2(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__o21ai_0 _1287_ (.A1(_0154_),
    .A2(_0302_),
    .B1(_0306_),
    .Y(_0307_));
 sky130_fd_sc_hd__a21oi_1 _1288_ (.A1(_0860_),
    .A2(_0301_),
    .B1(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__buf_6 _1289_ (.A(_0829_),
    .X(_0309_));
 sky130_fd_sc_hd__nor2_1 _1290_ (.A(\mem[0][18] ),
    .B(_0309_),
    .Y(_0310_));
 sky130_fd_sc_hd__a31oi_4 _1291_ (.A1(_0157_),
    .A2(_0298_),
    .A3(_0308_),
    .B1(_0310_),
    .Y(_0311_));
 sky130_fd_sc_hd__a22o_1 _1292_ (.A1(net85),
    .A2(_0790_),
    .B1(_0794_),
    .B2(_0311_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2i_1 _1293_ (.A0(\mem[9][19] ),
    .A1(\mem[13][19] ),
    .S(_0867_),
    .Y(_0312_));
 sky130_fd_sc_hd__nand2_1 _1294_ (.A(\mem[5][19] ),
    .B(_0866_),
    .Y(_0313_));
 sky130_fd_sc_hd__o21ai_1 _1295_ (.A1(_0869_),
    .A2(_0312_),
    .B1(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__a22oi_1 _1296_ (.A1(\mem[4][19] ),
    .A2(_0842_),
    .B1(_0152_),
    .B2(\mem[6][19] ),
    .Y(_0315_));
 sky130_fd_sc_hd__nand3_1 _1297_ (.A(_0162_),
    .B(\mem[12][19] ),
    .C(_0173_),
    .Y(_0316_));
 sky130_fd_sc_hd__o21ai_0 _1298_ (.A1(_0162_),
    .A2(_0315_),
    .B1(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__a22oi_1 _1299_ (.A1(_0863_),
    .A2(_0314_),
    .B1(_0317_),
    .B2(_0198_),
    .Y(_0318_));
 sky130_fd_sc_hd__a22o_1 _1300_ (.A1(\mem[15][19] ),
    .A2(_0812_),
    .B1(_0171_),
    .B2(\mem[3][19] ),
    .X(_0319_));
 sky130_fd_sc_hd__clkinv_4 _1301_ (.A(_0851_),
    .Y(_0320_));
 sky130_fd_sc_hd__a22oi_1 _1302_ (.A1(\mem[10][19] ),
    .A2(_0160_),
    .B1(_0812_),
    .B2(\mem[14][19] ),
    .Y(_0321_));
 sky130_fd_sc_hd__nand3_1 _1303_ (.A(_0858_),
    .B(\mem[7][19] ),
    .C(_0865_),
    .Y(_0322_));
 sky130_fd_sc_hd__o21ai_0 _1304_ (.A1(_0320_),
    .A2(_0321_),
    .B1(_0322_),
    .Y(_0323_));
 sky130_fd_sc_hd__a22oi_1 _1305_ (.A1(\mem[2][19] ),
    .A2(_0851_),
    .B1(_0137_),
    .B2(\mem[1][19] ),
    .Y(_0324_));
 sky130_fd_sc_hd__a22oi_1 _1306_ (.A1(_0247_),
    .A2(\mem[11][19] ),
    .B1(\mem[8][19] ),
    .B2(_0181_),
    .Y(_0325_));
 sky130_fd_sc_hd__o221ai_2 _1307_ (.A1(_0823_),
    .A2(_0324_),
    .B1(_0325_),
    .B2(_0145_),
    .C1(_0829_),
    .Y(_0326_));
 sky130_fd_sc_hd__a211oi_1 _1308_ (.A1(_0218_),
    .A2(_0319_),
    .B1(_0323_),
    .C1(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__nor2_1 _1309_ (.A(\mem[0][19] ),
    .B(_0129_),
    .Y(_0328_));
 sky130_fd_sc_hd__a21oi_1 _1310_ (.A1(_0318_),
    .A2(_0327_),
    .B1(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__a22o_1 _1311_ (.A1(net86),
    .A2(_0790_),
    .B1(_0794_),
    .B2(_0329_),
    .X(_0058_));
 sky130_fd_sc_hd__buf_4 _1312_ (.A(_0789_),
    .X(_0330_));
 sky130_fd_sc_hd__buf_6 _1313_ (.A(_0806_),
    .X(_0331_));
 sky130_fd_sc_hd__a22oi_2 _1314_ (.A1(\mem[10][1] ),
    .A2(_0859_),
    .B1(_0140_),
    .B2(\mem[9][1] ),
    .Y(_0332_));
 sky130_fd_sc_hd__a21oi_1 _1315_ (.A1(\mem[2][1] ),
    .A2(_0163_),
    .B1(_0166_),
    .Y(_0333_));
 sky130_fd_sc_hd__a21oi_1 _1316_ (.A1(_0331_),
    .A2(_0332_),
    .B1(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__a32oi_1 _1317_ (.A1(_0166_),
    .A2(\mem[14][1] ),
    .A3(_0124_),
    .B1(_0243_),
    .B2(\mem[7][1] ),
    .Y(_0335_));
 sky130_fd_sc_hd__nand2_1 _1318_ (.A(_0836_),
    .B(_0335_),
    .Y(_0336_));
 sky130_fd_sc_hd__o21ai_2 _1319_ (.A1(_0836_),
    .A2(_0334_),
    .B1(_0336_),
    .Y(_0337_));
 sky130_fd_sc_hd__mux2i_1 _1320_ (.A0(\mem[1][1] ),
    .A1(\mem[5][1] ),
    .S(_0839_),
    .Y(_0338_));
 sky130_fd_sc_hd__nand2_1 _1321_ (.A(\mem[13][1] ),
    .B(_0178_),
    .Y(_0339_));
 sky130_fd_sc_hd__o21ai_0 _1322_ (.A1(_0166_),
    .A2(_0338_),
    .B1(_0339_),
    .Y(_0340_));
 sky130_fd_sc_hd__a22oi_2 _1323_ (.A1(_0849_),
    .A2(\mem[11][1] ),
    .B1(\mem[8][1] ),
    .B2(_0850_),
    .Y(_0341_));
 sky130_fd_sc_hd__a22oi_2 _1324_ (.A1(\mem[4][1] ),
    .A2(_0802_),
    .B1(_0859_),
    .B2(\mem[6][1] ),
    .Y(_0342_));
 sky130_fd_sc_hd__nand3_1 _1325_ (.A(\mem[12][1] ),
    .B(_0181_),
    .C(_0812_),
    .Y(_0343_));
 sky130_fd_sc_hd__o221ai_4 _1326_ (.A1(_0145_),
    .A2(_0341_),
    .B1(_0342_),
    .B2(_0154_),
    .C1(_0343_),
    .Y(_0344_));
 sky130_fd_sc_hd__a21oi_1 _1327_ (.A1(_0193_),
    .A2(_0340_),
    .B1(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__a22o_1 _1328_ (.A1(\mem[15][1] ),
    .A2(_0812_),
    .B1(_0819_),
    .B2(\mem[3][1] ),
    .X(_0346_));
 sky130_fd_sc_hd__a21oi_1 _1329_ (.A1(_0218_),
    .A2(_0346_),
    .B1(_0824_),
    .Y(_0347_));
 sky130_fd_sc_hd__nor2_1 _1330_ (.A(\mem[0][1] ),
    .B(_0830_),
    .Y(_0348_));
 sky130_fd_sc_hd__a31oi_4 _1331_ (.A1(_0337_),
    .A2(_0345_),
    .A3(_0347_),
    .B1(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__a22o_1 _1332_ (.A1(net87),
    .A2(_0330_),
    .B1(_0794_),
    .B2(_0349_),
    .X(_0059_));
 sky130_fd_sc_hd__buf_6 _1333_ (.A(_0793_),
    .X(_0350_));
 sky130_fd_sc_hd__a22o_1 _1334_ (.A1(_0149_),
    .A2(\mem[15][20] ),
    .B1(\mem[12][20] ),
    .B2(_0842_),
    .X(_0351_));
 sky130_fd_sc_hd__a22oi_1 _1335_ (.A1(\mem[4][20] ),
    .A2(_0181_),
    .B1(_0182_),
    .B2(\mem[6][20] ),
    .Y(_0352_));
 sky130_fd_sc_hd__a22oi_1 _1336_ (.A1(_0841_),
    .A2(\mem[3][20] ),
    .B1(\mem[2][20] ),
    .B2(_0182_),
    .Y(_0353_));
 sky130_fd_sc_hd__o22ai_1 _1337_ (.A1(_0154_),
    .A2(_0352_),
    .B1(_0353_),
    .B2(_0823_),
    .Y(_0354_));
 sky130_fd_sc_hd__a21oi_1 _1338_ (.A1(_0178_),
    .A2(_0351_),
    .B1(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__a32o_1 _1339_ (.A1(_0122_),
    .A2(\mem[14][20] ),
    .A3(_0859_),
    .B1(_0243_),
    .B2(\mem[7][20] ),
    .X(_0356_));
 sky130_fd_sc_hd__a22o_1 _1340_ (.A1(\mem[13][20] ),
    .A2(_0812_),
    .B1(_0171_),
    .B2(\mem[1][20] ),
    .X(_0357_));
 sky130_fd_sc_hd__a222oi_1 _1341_ (.A1(_0796_),
    .A2(\mem[11][20] ),
    .B1(\mem[8][20] ),
    .B2(_0802_),
    .C1(_0814_),
    .C2(\mem[9][20] ),
    .Y(_0358_));
 sky130_fd_sc_hd__nand2_1 _1342_ (.A(_0199_),
    .B(\mem[10][20] ),
    .Y(_0359_));
 sky130_fd_sc_hd__nand4_1 _1343_ (.A(_0783_),
    .B(_0197_),
    .C(\mem[5][20] ),
    .D(_0226_),
    .Y(_0360_));
 sky130_fd_sc_hd__o221ai_1 _1344_ (.A1(_0145_),
    .A2(_0358_),
    .B1(_0359_),
    .B2(_0165_),
    .C1(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__a221oi_2 _1345_ (.A1(_0836_),
    .A2(_0356_),
    .B1(_0357_),
    .B2(_0193_),
    .C1(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__nor2_1 _1346_ (.A(\mem[0][20] ),
    .B(_0309_),
    .Y(_0363_));
 sky130_fd_sc_hd__a31oi_2 _1347_ (.A1(_0157_),
    .A2(_0355_),
    .A3(_0362_),
    .B1(_0363_),
    .Y(_0364_));
 sky130_fd_sc_hd__a22o_1 _1348_ (.A1(net88),
    .A2(_0330_),
    .B1(_0350_),
    .B2(_0364_),
    .X(_0060_));
 sky130_fd_sc_hd__a22oi_1 _1349_ (.A1(\mem[6][21] ),
    .A2(_0804_),
    .B1(_0814_),
    .B2(\mem[5][21] ),
    .Y(_0365_));
 sky130_fd_sc_hd__nand2_1 _1350_ (.A(_0836_),
    .B(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__a22o_1 _1351_ (.A1(\mem[13][21] ),
    .A2(_0178_),
    .B1(_0171_),
    .B2(\mem[1][21] ),
    .X(_0367_));
 sky130_fd_sc_hd__a32oi_4 _1352_ (.A1(\mem[3][21] ),
    .A2(_0243_),
    .A3(_0366_),
    .B1(_0367_),
    .B2(_0863_),
    .Y(_0368_));
 sky130_fd_sc_hd__nand2_1 _1353_ (.A(\mem[14][21] ),
    .B(_0851_),
    .Y(_0369_));
 sky130_fd_sc_hd__a21oi_1 _1354_ (.A1(\mem[4][21] ),
    .A2(_0245_),
    .B1(_0122_),
    .Y(_0370_));
 sky130_fd_sc_hd__a221oi_1 _1355_ (.A1(_0832_),
    .A2(_0369_),
    .B1(_0370_),
    .B2(_0365_),
    .C1(_0276_),
    .Y(_0371_));
 sky130_fd_sc_hd__a311oi_2 _1356_ (.A1(\mem[8][21] ),
    .A2(_0838_),
    .A3(_0174_),
    .B1(_0824_),
    .C1(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__a32o_1 _1357_ (.A1(_0276_),
    .A2(\mem[2][21] ),
    .A3(_0124_),
    .B1(_0272_),
    .B2(\mem[7][21] ),
    .X(_0373_));
 sky130_fd_sc_hd__a222oi_1 _1358_ (.A1(_0849_),
    .A2(\mem[11][21] ),
    .B1(\mem[10][21] ),
    .B2(_0817_),
    .C1(_0140_),
    .C2(\mem[9][21] ),
    .Y(_0374_));
 sky130_fd_sc_hd__a221oi_1 _1359_ (.A1(_0224_),
    .A2(\mem[15][21] ),
    .B1(\mem[12][21] ),
    .B2(_0245_),
    .C1(_0785_),
    .Y(_0375_));
 sky130_fd_sc_hd__a211oi_1 _1360_ (.A1(_0848_),
    .A2(_0374_),
    .B1(_0375_),
    .C1(_0869_),
    .Y(_0376_));
 sky130_fd_sc_hd__a21oi_1 _1361_ (.A1(_0881_),
    .A2(_0373_),
    .B1(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__nor2_1 _1362_ (.A(\mem[0][21] ),
    .B(_0309_),
    .Y(_0378_));
 sky130_fd_sc_hd__a31oi_4 _1363_ (.A1(_0368_),
    .A2(_0372_),
    .A3(_0377_),
    .B1(_0378_),
    .Y(_0379_));
 sky130_fd_sc_hd__a22o_1 _1364_ (.A1(net89),
    .A2(_0330_),
    .B1(_0350_),
    .B2(_0379_),
    .X(_0061_));
 sky130_fd_sc_hd__nand2_1 _1365_ (.A(\mem[10][22] ),
    .B(_0152_),
    .Y(_0380_));
 sky130_fd_sc_hd__a221oi_1 _1366_ (.A1(_0247_),
    .A2(\mem[3][22] ),
    .B1(\mem[2][22] ),
    .B2(_0851_),
    .C1(_0166_),
    .Y(_0381_));
 sky130_fd_sc_hd__a21oi_1 _1367_ (.A1(_0162_),
    .A2(_0380_),
    .B1(_0381_),
    .Y(_0382_));
 sky130_fd_sc_hd__a32oi_1 _1368_ (.A1(_0331_),
    .A2(\mem[12][22] ),
    .A3(_0173_),
    .B1(_0243_),
    .B2(\mem[7][22] ),
    .Y(_0383_));
 sky130_fd_sc_hd__nand2_1 _1369_ (.A(_0198_),
    .B(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__o21ai_1 _1370_ (.A1(_0198_),
    .A2(_0382_),
    .B1(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__a32o_1 _1371_ (.A1(_0207_),
    .A2(\mem[13][22] ),
    .A3(_0814_),
    .B1(_0847_),
    .B2(\mem[11][22] ),
    .X(_0386_));
 sky130_fd_sc_hd__a22o_1 _1372_ (.A1(\mem[4][22] ),
    .A2(_0837_),
    .B1(_0226_),
    .B2(\mem[5][22] ),
    .X(_0387_));
 sky130_fd_sc_hd__a221oi_1 _1373_ (.A1(\mem[8][22] ),
    .A2(_0802_),
    .B1(_0814_),
    .B2(\mem[9][22] ),
    .C1(_0145_),
    .Y(_0388_));
 sky130_fd_sc_hd__a221oi_1 _1374_ (.A1(_0849_),
    .A2(\mem[15][22] ),
    .B1(\mem[14][22] ),
    .B2(_0859_),
    .C1(_0856_),
    .Y(_0389_));
 sky130_fd_sc_hd__and3_1 _1375_ (.A(_0834_),
    .B(\mem[6][22] ),
    .C(_0803_),
    .X(_0390_));
 sky130_fd_sc_hd__a311oi_1 _1376_ (.A1(_0785_),
    .A2(\mem[1][22] ),
    .A3(_0820_),
    .B1(_0390_),
    .C1(_0122_),
    .Y(_0391_));
 sky130_fd_sc_hd__nor3_1 _1377_ (.A(_0388_),
    .B(_0389_),
    .C(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__a221oi_2 _1378_ (.A1(_0200_),
    .A2(_0386_),
    .B1(_0387_),
    .B2(_0866_),
    .C1(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__nor2_1 _1379_ (.A(\mem[0][22] ),
    .B(_0309_),
    .Y(_0394_));
 sky130_fd_sc_hd__a31oi_4 _1380_ (.A1(_0157_),
    .A2(_0385_),
    .A3(_0393_),
    .B1(_0394_),
    .Y(_0395_));
 sky130_fd_sc_hd__a22o_1 _1381_ (.A1(net90),
    .A2(_0330_),
    .B1(_0350_),
    .B2(_0395_),
    .X(_0062_));
 sky130_fd_sc_hd__a32oi_1 _1382_ (.A1(_0234_),
    .A2(\mem[14][23] ),
    .A3(_0152_),
    .B1(_0847_),
    .B2(\mem[11][23] ),
    .Y(_0396_));
 sky130_fd_sc_hd__a222oi_1 _1383_ (.A1(_0849_),
    .A2(\mem[15][23] ),
    .B1(\mem[12][23] ),
    .B2(_0802_),
    .C1(_0820_),
    .C2(\mem[13][23] ),
    .Y(_0397_));
 sky130_fd_sc_hd__nand2_1 _1384_ (.A(_0840_),
    .B(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__a222oi_1 _1385_ (.A1(\mem[10][23] ),
    .A2(_0804_),
    .B1(_0814_),
    .B2(\mem[9][23] ),
    .C1(\mem[8][23] ),
    .C2(_0850_),
    .Y(_0399_));
 sky130_fd_sc_hd__nand2_1 _1386_ (.A(_0848_),
    .B(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__nand2_1 _1387_ (.A(_0398_),
    .B(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__and3_1 _1388_ (.A(_0785_),
    .B(\mem[1][23] ),
    .C(_0798_),
    .X(_0402_));
 sky130_fd_sc_hd__nand2_1 _1389_ (.A(\mem[5][23] ),
    .B(_0798_),
    .Y(_0403_));
 sky130_fd_sc_hd__a22oi_1 _1390_ (.A1(\mem[4][23] ),
    .A2(_0801_),
    .B1(_0804_),
    .B2(\mem[6][23] ),
    .Y(_0404_));
 sky130_fd_sc_hd__a221oi_1 _1391_ (.A1(_0795_),
    .A2(\mem[3][23] ),
    .B1(\mem[2][23] ),
    .B2(_0803_),
    .C1(_0834_),
    .Y(_0405_));
 sky130_fd_sc_hd__a31oi_1 _1392_ (.A1(_0839_),
    .A2(_0403_),
    .A3(_0404_),
    .B1(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__a2111oi_0 _1393_ (.A1(\mem[7][23] ),
    .A2(_0272_),
    .B1(_0402_),
    .C1(_0406_),
    .D1(_0331_),
    .Y(_0407_));
 sky130_fd_sc_hd__a31oi_1 _1394_ (.A1(_0833_),
    .A2(_0396_),
    .A3(_0401_),
    .B1(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__a21o_1 _1395_ (.A1(\mem[0][23] ),
    .A2(_0132_),
    .B1(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__a22o_1 _1396_ (.A1(net91),
    .A2(_0330_),
    .B1(_0350_),
    .B2(_0409_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2i_1 _1397_ (.A0(\mem[11][24] ),
    .A1(\mem[15][24] ),
    .S(_0839_),
    .Y(_0410_));
 sky130_fd_sc_hd__nand2_1 _1398_ (.A(\mem[7][24] ),
    .B(_0865_),
    .Y(_0411_));
 sky130_fd_sc_hd__o21ai_1 _1399_ (.A1(_0783_),
    .A2(_0410_),
    .B1(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__a22oi_1 _1400_ (.A1(_0247_),
    .A2(\mem[3][24] ),
    .B1(\mem[2][24] ),
    .B2(_0163_),
    .Y(_0413_));
 sky130_fd_sc_hd__a21oi_1 _1401_ (.A1(\mem[1][24] ),
    .A2(_0137_),
    .B1(_0166_),
    .Y(_0414_));
 sky130_fd_sc_hd__a21oi_2 _1402_ (.A1(_0413_),
    .A2(_0414_),
    .B1(_0840_),
    .Y(_0415_));
 sky130_fd_sc_hd__a222oi_1 _1403_ (.A1(\mem[10][24] ),
    .A2(_0817_),
    .B1(_0820_),
    .B2(\mem[9][24] ),
    .C1(\mem[8][24] ),
    .C2(_0837_),
    .Y(_0416_));
 sky130_fd_sc_hd__nand2_1 _1404_ (.A(_0162_),
    .B(_0416_),
    .Y(_0417_));
 sky130_fd_sc_hd__a222oi_1 _1405_ (.A1(\mem[6][24] ),
    .A2(_0817_),
    .B1(_0820_),
    .B2(\mem[5][24] ),
    .C1(\mem[4][24] ),
    .C2(_0837_),
    .Y(_0418_));
 sky130_fd_sc_hd__a222oi_1 _1406_ (.A1(\mem[14][24] ),
    .A2(_0817_),
    .B1(_0820_),
    .B2(\mem[13][24] ),
    .C1(\mem[12][24] ),
    .C2(_0837_),
    .Y(_0419_));
 sky130_fd_sc_hd__o22ai_2 _1407_ (.A1(_0154_),
    .A2(_0418_),
    .B1(_0419_),
    .B2(_0857_),
    .Y(_0420_));
 sky130_fd_sc_hd__a221oi_4 _1408_ (.A1(_0218_),
    .A2(_0412_),
    .B1(_0415_),
    .B2(_0417_),
    .C1(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__nor2_1 _1409_ (.A(\mem[0][24] ),
    .B(_0129_),
    .Y(_0422_));
 sky130_fd_sc_hd__a21oi_4 _1410_ (.A1(_0831_),
    .A2(_0421_),
    .B1(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__a22o_1 _1411_ (.A1(net92),
    .A2(_0330_),
    .B1(_0350_),
    .B2(_0423_),
    .X(_0064_));
 sky130_fd_sc_hd__nand2_1 _1412_ (.A(\mem[14][25] ),
    .B(_0182_),
    .Y(_0424_));
 sky130_fd_sc_hd__a22oi_1 _1413_ (.A1(\mem[12][25] ),
    .A2(_0134_),
    .B1(_0137_),
    .B2(\mem[13][25] ),
    .Y(_0425_));
 sky130_fd_sc_hd__a221oi_1 _1414_ (.A1(\mem[4][25] ),
    .A2(_0245_),
    .B1(_0851_),
    .B2(\mem[6][25] ),
    .C1(_0199_),
    .Y(_0426_));
 sky130_fd_sc_hd__a31oi_1 _1415_ (.A1(_0123_),
    .A2(_0424_),
    .A3(_0425_),
    .B1(_0426_),
    .Y(_0427_));
 sky130_fd_sc_hd__mux2i_1 _1416_ (.A0(\mem[3][25] ),
    .A1(\mem[11][25] ),
    .S(_0122_),
    .Y(_0428_));
 sky130_fd_sc_hd__mux2i_1 _1417_ (.A0(\mem[2][25] ),
    .A1(\mem[10][25] ),
    .S(_0199_),
    .Y(_0429_));
 sky130_fd_sc_hd__o22ai_1 _1418_ (.A1(_0282_),
    .A2(_0428_),
    .B1(_0429_),
    .B2(_0165_),
    .Y(_0430_));
 sky130_fd_sc_hd__a21oi_1 _1419_ (.A1(_0198_),
    .A2(_0427_),
    .B1(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__a22oi_1 _1420_ (.A1(\mem[8][25] ),
    .A2(_0181_),
    .B1(_0226_),
    .B2(\mem[9][25] ),
    .Y(_0432_));
 sky130_fd_sc_hd__nand2_1 _1421_ (.A(\mem[15][25] ),
    .B(_0272_),
    .Y(_0433_));
 sky130_fd_sc_hd__o21ai_0 _1422_ (.A1(_0840_),
    .A2(_0432_),
    .B1(_0433_),
    .Y(_0434_));
 sky130_fd_sc_hd__a22oi_1 _1423_ (.A1(_0149_),
    .A2(\mem[7][25] ),
    .B1(\mem[5][25] ),
    .B2(_0862_),
    .Y(_0435_));
 sky130_fd_sc_hd__a21oi_1 _1424_ (.A1(\mem[1][25] ),
    .A2(_0305_),
    .B1(_0123_),
    .Y(_0436_));
 sky130_fd_sc_hd__o21ai_0 _1425_ (.A1(_0848_),
    .A2(_0435_),
    .B1(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__o21ai_1 _1426_ (.A1(_0881_),
    .A2(_0434_),
    .B1(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__nor2_1 _1427_ (.A(\mem[0][25] ),
    .B(_0309_),
    .Y(_0439_));
 sky130_fd_sc_hd__a31oi_4 _1428_ (.A1(_0157_),
    .A2(_0431_),
    .A3(_0438_),
    .B1(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__a22o_1 _1429_ (.A1(net93),
    .A2(_0330_),
    .B1(_0350_),
    .B2(_0440_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2i_1 _1430_ (.A0(\mem[3][26] ),
    .A1(\mem[7][26] ),
    .S(_0197_),
    .Y(_0441_));
 sky130_fd_sc_hd__nand3_1 _1431_ (.A(_0200_),
    .B(_0208_),
    .C(\mem[15][26] ),
    .Y(_0442_));
 sky130_fd_sc_hd__o21ai_0 _1432_ (.A1(_0200_),
    .A2(_0441_),
    .B1(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__nand2_1 _1433_ (.A(_0218_),
    .B(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__mux2i_1 _1434_ (.A0(\mem[10][26] ),
    .A1(\mem[14][26] ),
    .S(_0207_),
    .Y(_0445_));
 sky130_fd_sc_hd__o31ai_1 _1435_ (.A1(_0783_),
    .A2(_0320_),
    .A3(_0445_),
    .B1(_0830_),
    .Y(_0446_));
 sky130_fd_sc_hd__a31oi_2 _1436_ (.A1(\mem[8][26] ),
    .A2(_0838_),
    .A3(_0174_),
    .B1(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__nand2_1 _1437_ (.A(\mem[5][26] ),
    .B(_0862_),
    .Y(_0448_));
 sky130_fd_sc_hd__a22oi_1 _1438_ (.A1(\mem[4][26] ),
    .A2(_0134_),
    .B1(_0124_),
    .B2(\mem[6][26] ),
    .Y(_0449_));
 sky130_fd_sc_hd__a221oi_1 _1439_ (.A1(\mem[2][26] ),
    .A2(_0143_),
    .B1(_0140_),
    .B2(\mem[1][26] ),
    .C1(_0835_),
    .Y(_0450_));
 sky130_fd_sc_hd__a31oi_1 _1440_ (.A1(_0208_),
    .A2(_0448_),
    .A3(_0449_),
    .B1(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__a221oi_1 _1441_ (.A1(_0247_),
    .A2(\mem[11][26] ),
    .B1(\mem[9][26] ),
    .B2(_0140_),
    .C1(_0835_),
    .Y(_0452_));
 sky130_fd_sc_hd__a221oi_1 _1442_ (.A1(\mem[12][26] ),
    .A2(_0134_),
    .B1(_0226_),
    .B2(\mem[13][26] ),
    .C1(_0276_),
    .Y(_0453_));
 sky130_fd_sc_hd__o21ai_0 _1443_ (.A1(_0452_),
    .A2(_0453_),
    .B1(_0200_),
    .Y(_0454_));
 sky130_fd_sc_hd__o21ai_1 _1444_ (.A1(_0833_),
    .A2(_0451_),
    .B1(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__nor2_1 _1445_ (.A(\mem[0][26] ),
    .B(_0309_),
    .Y(_0456_));
 sky130_fd_sc_hd__a31oi_4 _1446_ (.A1(_0444_),
    .A2(_0447_),
    .A3(_0455_),
    .B1(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__a22o_1 _1447_ (.A1(net94),
    .A2(_0330_),
    .B1(_0350_),
    .B2(_0457_),
    .X(_0066_));
 sky130_fd_sc_hd__nand2_1 _1448_ (.A(net95),
    .B(_0826_),
    .Y(_0458_));
 sky130_fd_sc_hd__a22oi_1 _1449_ (.A1(\mem[14][27] ),
    .A2(_0163_),
    .B1(_0862_),
    .B2(\mem[13][27] ),
    .Y(_0459_));
 sky130_fd_sc_hd__a221oi_1 _1450_ (.A1(_0247_),
    .A2(\mem[11][27] ),
    .B1(\mem[8][27] ),
    .B2(_0134_),
    .C1(_0197_),
    .Y(_0460_));
 sky130_fd_sc_hd__a21oi_1 _1451_ (.A1(_0208_),
    .A2(_0459_),
    .B1(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__a22oi_1 _1452_ (.A1(_0247_),
    .A2(\mem[7][27] ),
    .B1(\mem[4][27] ),
    .B2(_0181_),
    .Y(_0462_));
 sky130_fd_sc_hd__a221oi_1 _1453_ (.A1(\mem[2][27] ),
    .A2(_0859_),
    .B1(_0140_),
    .B2(\mem[1][27] ),
    .C1(_0835_),
    .Y(_0463_));
 sky130_fd_sc_hd__a211oi_1 _1454_ (.A1(_0208_),
    .A2(_0462_),
    .B1(_0463_),
    .C1(_0200_),
    .Y(_0464_));
 sky130_fd_sc_hd__a21oi_2 _1455_ (.A1(_0833_),
    .A2(_0461_),
    .B1(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__a22o_1 _1456_ (.A1(\mem[9][27] ),
    .A2(_0160_),
    .B1(_0865_),
    .B2(\mem[5][27] ),
    .X(_0466_));
 sky130_fd_sc_hd__a22o_1 _1457_ (.A1(\mem[15][27] ),
    .A2(_0178_),
    .B1(_0171_),
    .B2(\mem[3][27] ),
    .X(_0467_));
 sky130_fd_sc_hd__a22oi_1 _1458_ (.A1(_0863_),
    .A2(_0466_),
    .B1(_0467_),
    .B2(_0218_),
    .Y(_0468_));
 sky130_fd_sc_hd__a22o_1 _1459_ (.A1(\mem[10][27] ),
    .A2(_0160_),
    .B1(_0865_),
    .B2(\mem[6][27] ),
    .X(_0469_));
 sky130_fd_sc_hd__a32oi_1 _1460_ (.A1(\mem[12][27] ),
    .A2(_0838_),
    .A3(_0178_),
    .B1(_0469_),
    .B2(_0860_),
    .Y(_0470_));
 sky130_fd_sc_hd__nand4_1 _1461_ (.A(_0157_),
    .B(_0465_),
    .C(_0468_),
    .D(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__o2111ai_1 _1462_ (.A1(\mem[0][27] ),
    .A2(_0831_),
    .B1(_0471_),
    .C1(_0826_),
    .D1(_0231_),
    .Y(_0472_));
 sky130_fd_sc_hd__o21ai_0 _1463_ (.A1(_0231_),
    .A2(_0458_),
    .B1(_0472_),
    .Y(_0067_));
 sky130_fd_sc_hd__a22oi_1 _1464_ (.A1(_0136_),
    .A2(\mem[15][28] ),
    .B1(\mem[12][28] ),
    .B2(_0850_),
    .Y(_0473_));
 sky130_fd_sc_hd__a222oi_1 _1465_ (.A1(_0849_),
    .A2(\mem[7][28] ),
    .B1(\mem[4][28] ),
    .B2(_0802_),
    .C1(_0140_),
    .C2(\mem[5][28] ),
    .Y(_0474_));
 sky130_fd_sc_hd__a21oi_1 _1466_ (.A1(_0331_),
    .A2(_0473_),
    .B1(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__a221o_1 _1467_ (.A1(_0224_),
    .A2(\mem[3][28] ),
    .B1(\mem[2][28] ),
    .B2(_0143_),
    .C1(_0199_),
    .X(_0476_));
 sky130_fd_sc_hd__nand2_1 _1468_ (.A(\mem[8][28] ),
    .B(_0842_),
    .Y(_0477_));
 sky130_fd_sc_hd__a21oi_1 _1469_ (.A1(_0133_),
    .A2(_0477_),
    .B1(_0840_),
    .Y(_0478_));
 sky130_fd_sc_hd__mux2i_1 _1470_ (.A0(\mem[6][28] ),
    .A1(\mem[14][28] ),
    .S(_0806_),
    .Y(_0479_));
 sky130_fd_sc_hd__mux2i_1 _1471_ (.A0(\mem[1][28] ),
    .A1(\mem[9][28] ),
    .S(_0122_),
    .Y(_0480_));
 sky130_fd_sc_hd__o32ai_1 _1472_ (.A1(_0276_),
    .A2(_0320_),
    .A3(_0479_),
    .B1(_0480_),
    .B2(_0279_),
    .Y(_0481_));
 sky130_fd_sc_hd__a221oi_2 _1473_ (.A1(_0836_),
    .A2(_0475_),
    .B1(_0476_),
    .B2(_0478_),
    .C1(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__nand2_1 _1474_ (.A(\mem[13][28] ),
    .B(_0150_),
    .Y(_0483_));
 sky130_fd_sc_hd__a221oi_1 _1475_ (.A1(_0841_),
    .A2(\mem[11][28] ),
    .B1(\mem[10][28] ),
    .B2(_0163_),
    .C1(_0197_),
    .Y(_0484_));
 sky130_fd_sc_hd__a31oi_1 _1476_ (.A1(_0208_),
    .A2(_0473_),
    .A3(_0483_),
    .B1(_0484_),
    .Y(_0485_));
 sky130_fd_sc_hd__a21oi_1 _1477_ (.A1(_0833_),
    .A2(_0485_),
    .B1(_0132_),
    .Y(_0486_));
 sky130_fd_sc_hd__nor2_1 _1478_ (.A(\mem[0][28] ),
    .B(_0129_),
    .Y(_0487_));
 sky130_fd_sc_hd__a21oi_4 _1479_ (.A1(_0482_),
    .A2(_0486_),
    .B1(_0487_),
    .Y(_0488_));
 sky130_fd_sc_hd__a22o_1 _1480_ (.A1(net96),
    .A2(_0330_),
    .B1(_0350_),
    .B2(_0488_),
    .X(_0068_));
 sky130_fd_sc_hd__nand2_1 _1481_ (.A(\mem[2][29] ),
    .B(_0152_),
    .Y(_0489_));
 sky130_fd_sc_hd__nand3_1 _1482_ (.A(_0133_),
    .B(\mem[8][29] ),
    .C(_0173_),
    .Y(_0490_));
 sky130_fd_sc_hd__o21ai_0 _1483_ (.A1(_0123_),
    .A2(_0489_),
    .B1(_0490_),
    .Y(_0491_));
 sky130_fd_sc_hd__a22oi_1 _1484_ (.A1(_0149_),
    .A2(\mem[15][29] ),
    .B1(\mem[14][29] ),
    .B2(_0152_),
    .Y(_0492_));
 sky130_fd_sc_hd__a21oi_1 _1485_ (.A1(\mem[13][29] ),
    .A2(_0862_),
    .B1(_0857_),
    .Y(_0493_));
 sky130_fd_sc_hd__a221oi_1 _1486_ (.A1(\mem[4][29] ),
    .A2(_0181_),
    .B1(_0182_),
    .B2(\mem[6][29] ),
    .C1(_0154_),
    .Y(_0494_));
 sky130_fd_sc_hd__a21oi_1 _1487_ (.A1(_0492_),
    .A2(_0493_),
    .B1(_0494_),
    .Y(_0495_));
 sky130_fd_sc_hd__o21ai_0 _1488_ (.A1(_0198_),
    .A2(_0491_),
    .B1(_0495_),
    .Y(_0496_));
 sky130_fd_sc_hd__mux2i_1 _1489_ (.A0(\mem[1][29] ),
    .A1(\mem[5][29] ),
    .S(_0207_),
    .Y(_0497_));
 sky130_fd_sc_hd__nand2_1 _1490_ (.A(\mem[9][29] ),
    .B(_0174_),
    .Y(_0498_));
 sky130_fd_sc_hd__o21ai_0 _1491_ (.A1(_0133_),
    .A2(_0497_),
    .B1(_0498_),
    .Y(_0499_));
 sky130_fd_sc_hd__nand2_1 _1492_ (.A(_0832_),
    .B(_0842_),
    .Y(_0500_));
 sky130_fd_sc_hd__nand2_1 _1493_ (.A(_0234_),
    .B(\mem[12][29] ),
    .Y(_0501_));
 sky130_fd_sc_hd__mux2_1 _1494_ (.A0(\mem[3][29] ),
    .A1(\mem[7][29] ),
    .S(_0784_),
    .X(_0502_));
 sky130_fd_sc_hd__a22o_1 _1495_ (.A1(_0849_),
    .A2(\mem[11][29] ),
    .B1(\mem[10][29] ),
    .B2(_0817_),
    .X(_0503_));
 sky130_fd_sc_hd__a22oi_1 _1496_ (.A1(_0243_),
    .A2(_0502_),
    .B1(_0503_),
    .B2(_0174_),
    .Y(_0504_));
 sky130_fd_sc_hd__o21ai_1 _1497_ (.A1(_0500_),
    .A2(_0501_),
    .B1(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__a21oi_1 _1498_ (.A1(_0863_),
    .A2(_0499_),
    .B1(_0505_),
    .Y(_0506_));
 sky130_fd_sc_hd__nor2_1 _1499_ (.A(\mem[0][29] ),
    .B(_0309_),
    .Y(_0507_));
 sky130_fd_sc_hd__a31oi_1 _1500_ (.A1(_0157_),
    .A2(_0496_),
    .A3(_0506_),
    .B1(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__a22o_1 _1501_ (.A1(net97),
    .A2(_0330_),
    .B1(_0350_),
    .B2(_0508_),
    .X(_0069_));
 sky130_fd_sc_hd__nand2_1 _1502_ (.A(net98),
    .B(_0826_),
    .Y(_0509_));
 sky130_fd_sc_hd__mux2i_1 _1503_ (.A0(\mem[2][2] ),
    .A1(\mem[6][2] ),
    .S(_0867_),
    .Y(_0510_));
 sky130_fd_sc_hd__nor2_1 _1504_ (.A(_0162_),
    .B(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__a21oi_1 _1505_ (.A1(\mem[10][2] ),
    .A2(_0174_),
    .B1(_0511_),
    .Y(_0512_));
 sky130_fd_sc_hd__nor2_1 _1506_ (.A(\mem[0][2] ),
    .B(_0830_),
    .Y(_0513_));
 sky130_fd_sc_hd__a22oi_2 _1507_ (.A1(_0136_),
    .A2(\mem[7][2] ),
    .B1(\mem[4][2] ),
    .B2(_0837_),
    .Y(_0514_));
 sky130_fd_sc_hd__mux2i_2 _1508_ (.A0(\mem[8][2] ),
    .A1(\mem[12][2] ),
    .S(_0839_),
    .Y(_0515_));
 sky130_fd_sc_hd__o22ai_4 _1509_ (.A1(_0154_),
    .A2(_0514_),
    .B1(_0515_),
    .B2(_0500_),
    .Y(_0516_));
 sky130_fd_sc_hd__a311oi_4 _1510_ (.A1(\mem[1][2] ),
    .A2(_0193_),
    .A3(_0171_),
    .B1(_0824_),
    .C1(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__a221o_1 _1511_ (.A1(_0149_),
    .A2(\mem[11][2] ),
    .B1(\mem[9][2] ),
    .B2(_0862_),
    .C1(_0145_),
    .X(_0518_));
 sky130_fd_sc_hd__a22oi_1 _1512_ (.A1(_0858_),
    .A2(\mem[15][2] ),
    .B1(\mem[13][2] ),
    .B2(_0193_),
    .Y(_0519_));
 sky130_fd_sc_hd__nand2_1 _1513_ (.A(\mem[14][2] ),
    .B(_0860_),
    .Y(_0520_));
 sky130_fd_sc_hd__nand3_1 _1514_ (.A(_0178_),
    .B(_0519_),
    .C(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__nand2_1 _1515_ (.A(\mem[5][2] ),
    .B(_0150_),
    .Y(_0522_));
 sky130_fd_sc_hd__nand2_1 _1516_ (.A(_0858_),
    .B(\mem[3][2] ),
    .Y(_0523_));
 sky130_fd_sc_hd__a22oi_1 _1517_ (.A1(_0866_),
    .A2(_0522_),
    .B1(_0523_),
    .B2(_0171_),
    .Y(_0524_));
 sky130_fd_sc_hd__nand3_1 _1518_ (.A(_0518_),
    .B(_0521_),
    .C(_0524_),
    .Y(_0525_));
 sky130_fd_sc_hd__o221ai_4 _1519_ (.A1(_0320_),
    .A2(_0512_),
    .B1(_0513_),
    .B2(_0517_),
    .C1(_0525_),
    .Y(_0526_));
 sky130_fd_sc_hd__nand3_1 _1520_ (.A(_0826_),
    .B(_0231_),
    .C(_0526_),
    .Y(_0527_));
 sky130_fd_sc_hd__o21ai_0 _1521_ (.A1(_0231_),
    .A2(_0509_),
    .B1(_0527_),
    .Y(_0070_));
 sky130_fd_sc_hd__a22o_1 _1522_ (.A1(_0841_),
    .A2(\mem[15][30] ),
    .B1(\mem[12][30] ),
    .B2(_0181_),
    .X(_0528_));
 sky130_fd_sc_hd__a221o_1 _1523_ (.A1(_0247_),
    .A2(\mem[11][30] ),
    .B1(\mem[8][30] ),
    .B2(_0134_),
    .C1(_0835_),
    .X(_0529_));
 sky130_fd_sc_hd__o21ai_0 _1524_ (.A1(_0884_),
    .A2(_0528_),
    .B1(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__mux2_1 _1525_ (.A0(\mem[10][30] ),
    .A1(\mem[14][30] ),
    .S(_0834_),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _1526_ (.A0(\mem[9][30] ),
    .A1(\mem[13][30] ),
    .S(_0834_),
    .X(_0532_));
 sky130_fd_sc_hd__a221oi_1 _1527_ (.A1(_0860_),
    .A2(_0531_),
    .B1(_0532_),
    .B2(_0193_),
    .C1(_0869_),
    .Y(_0533_));
 sky130_fd_sc_hd__a22oi_1 _1528_ (.A1(_0136_),
    .A2(\mem[7][30] ),
    .B1(\mem[5][30] ),
    .B2(_0820_),
    .Y(_0534_));
 sky130_fd_sc_hd__a22oi_1 _1529_ (.A1(\mem[4][30] ),
    .A2(_0850_),
    .B1(_0143_),
    .B2(\mem[6][30] ),
    .Y(_0535_));
 sky130_fd_sc_hd__a221oi_1 _1530_ (.A1(_0849_),
    .A2(\mem[3][30] ),
    .B1(\mem[2][30] ),
    .B2(_0817_),
    .C1(_0207_),
    .Y(_0536_));
 sky130_fd_sc_hd__a31oi_1 _1531_ (.A1(_0234_),
    .A2(_0534_),
    .A3(_0535_),
    .B1(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__a211oi_1 _1532_ (.A1(\mem[1][30] ),
    .A2(_0305_),
    .B1(_0537_),
    .C1(_0200_),
    .Y(_0538_));
 sky130_fd_sc_hd__a21oi_1 _1533_ (.A1(_0530_),
    .A2(_0533_),
    .B1(_0538_),
    .Y(_0539_));
 sky130_fd_sc_hd__a21oi_4 _1534_ (.A1(\mem[0][30] ),
    .A2(_0132_),
    .B1(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__nor2_1 _1535_ (.A(net99),
    .B(_0827_),
    .Y(_0541_));
 sky130_fd_sc_hd__a211oi_1 _1536_ (.A1(_0231_),
    .A2(_0540_),
    .B1(_0541_),
    .C1(_0764_),
    .Y(_0071_));
 sky130_fd_sc_hd__mux2i_2 _1537_ (.A0(\mem[8][31] ),
    .A1(\mem[12][31] ),
    .S(_0207_),
    .Y(_0542_));
 sky130_fd_sc_hd__nand2_1 _1538_ (.A(_0162_),
    .B(_0542_),
    .Y(_0543_));
 sky130_fd_sc_hd__nand2_1 _1539_ (.A(_0234_),
    .B(\mem[4][31] ),
    .Y(_0544_));
 sky130_fd_sc_hd__nand2_1 _1540_ (.A(_0869_),
    .B(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__a32oi_2 _1541_ (.A1(_0122_),
    .A2(\mem[14][31] ),
    .A3(_0143_),
    .B1(_0243_),
    .B2(\mem[7][31] ),
    .Y(_0546_));
 sky130_fd_sc_hd__a22o_1 _1542_ (.A1(\mem[10][31] ),
    .A2(_0803_),
    .B1(_0797_),
    .B2(\mem[9][31] ),
    .X(_0547_));
 sky130_fd_sc_hd__a221oi_1 _1543_ (.A1(\mem[3][31] ),
    .A2(_0242_),
    .B1(_0547_),
    .B2(_0806_),
    .C1(_0867_),
    .Y(_0548_));
 sky130_fd_sc_hd__a21oi_1 _1544_ (.A1(_0840_),
    .A2(_0546_),
    .B1(_0548_),
    .Y(_0549_));
 sky130_fd_sc_hd__mux2_1 _1545_ (.A0(\mem[2][31] ),
    .A1(\mem[6][31] ),
    .S(_0784_),
    .X(_0550_));
 sky130_fd_sc_hd__mux2_1 _1546_ (.A0(\mem[1][31] ),
    .A1(\mem[5][31] ),
    .S(_0784_),
    .X(_0551_));
 sky130_fd_sc_hd__a221oi_1 _1547_ (.A1(_0163_),
    .A2(_0550_),
    .B1(_0551_),
    .B2(_0137_),
    .C1(_0166_),
    .Y(_0552_));
 sky130_fd_sc_hd__a22o_1 _1548_ (.A1(_0795_),
    .A2(\mem[15][31] ),
    .B1(\mem[13][31] ),
    .B2(_0798_),
    .X(_0553_));
 sky130_fd_sc_hd__a221oi_1 _1549_ (.A1(\mem[11][31] ),
    .A2(_0847_),
    .B1(_0553_),
    .B2(_0867_),
    .C1(_0783_),
    .Y(_0554_));
 sky130_fd_sc_hd__nor2_1 _1550_ (.A(_0552_),
    .B(_0554_),
    .Y(_0555_));
 sky130_fd_sc_hd__a311oi_1 _1551_ (.A1(_0838_),
    .A2(_0543_),
    .A3(_0545_),
    .B1(_0549_),
    .C1(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__nor2_1 _1552_ (.A(\mem[0][31] ),
    .B(_0129_),
    .Y(_0557_));
 sky130_fd_sc_hd__a21oi_1 _1553_ (.A1(_0831_),
    .A2(_0556_),
    .B1(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__a22o_1 _1554_ (.A1(net100),
    .A2(_0789_),
    .B1(_0350_),
    .B2(_0558_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2i_1 _1555_ (.A0(\mem[10][3] ),
    .A1(\mem[14][3] ),
    .S(_0839_),
    .Y(_0559_));
 sky130_fd_sc_hd__o2bb2ai_1 _1556_ (.A1_N(\mem[6][3] ),
    .A2_N(_0865_),
    .B1(_0559_),
    .B2(_0783_),
    .Y(_0560_));
 sky130_fd_sc_hd__a22oi_1 _1557_ (.A1(\mem[4][3] ),
    .A2(_0850_),
    .B1(_0140_),
    .B2(\mem[5][3] ),
    .Y(_0561_));
 sky130_fd_sc_hd__nand2_1 _1558_ (.A(_0841_),
    .B(\mem[7][3] ),
    .Y(_0562_));
 sky130_fd_sc_hd__nand3_1 _1559_ (.A(_0234_),
    .B(_0561_),
    .C(_0562_),
    .Y(_0563_));
 sky130_fd_sc_hd__a22oi_1 _1560_ (.A1(_0136_),
    .A2(\mem[3][3] ),
    .B1(\mem[2][3] ),
    .B2(_0859_),
    .Y(_0564_));
 sky130_fd_sc_hd__a21oi_1 _1561_ (.A1(\mem[1][3] ),
    .A2(_0814_),
    .B1(_0207_),
    .Y(_0565_));
 sky130_fd_sc_hd__a21oi_1 _1562_ (.A1(_0564_),
    .A2(_0565_),
    .B1(_0832_),
    .Y(_0566_));
 sky130_fd_sc_hd__a222oi_1 _1563_ (.A1(_0796_),
    .A2(\mem[15][3] ),
    .B1(\mem[12][3] ),
    .B2(_0802_),
    .C1(_0814_),
    .C2(\mem[13][3] ),
    .Y(_0567_));
 sky130_fd_sc_hd__a222oi_1 _1564_ (.A1(_0796_),
    .A2(\mem[11][3] ),
    .B1(\mem[8][3] ),
    .B2(_0802_),
    .C1(_0820_),
    .C2(\mem[9][3] ),
    .Y(_0568_));
 sky130_fd_sc_hd__o22ai_2 _1565_ (.A1(_0857_),
    .A2(_0567_),
    .B1(_0568_),
    .B2(_0145_),
    .Y(_0569_));
 sky130_fd_sc_hd__a221oi_2 _1566_ (.A1(_0860_),
    .A2(_0560_),
    .B1(_0563_),
    .B2(_0566_),
    .C1(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__nor2_1 _1567_ (.A(\mem[0][3] ),
    .B(_0830_),
    .Y(_0571_));
 sky130_fd_sc_hd__a21oi_4 _1568_ (.A1(_0157_),
    .A2(_0570_),
    .B1(_0571_),
    .Y(_0572_));
 sky130_fd_sc_hd__a22o_1 _1569_ (.A1(net101),
    .A2(_0789_),
    .B1(_0793_),
    .B2(_0572_),
    .X(_0073_));
 sky130_fd_sc_hd__mux4_1 _1570_ (.A0(\mem[2][4] ),
    .A1(\mem[6][4] ),
    .A2(\mem[10][4] ),
    .A3(\mem[14][4] ),
    .S0(_0784_),
    .S1(_0199_),
    .X(_0573_));
 sky130_fd_sc_hd__nand2_1 _1571_ (.A(_0860_),
    .B(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__mux2i_1 _1572_ (.A0(\mem[9][4] ),
    .A1(\mem[13][4] ),
    .S(_0835_),
    .Y(_0575_));
 sky130_fd_sc_hd__nand2_1 _1573_ (.A(_0200_),
    .B(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__nand2_1 _1574_ (.A(_0234_),
    .B(\mem[5][4] ),
    .Y(_0577_));
 sky130_fd_sc_hd__nand2_1 _1575_ (.A(_0869_),
    .B(_0577_),
    .Y(_0578_));
 sky130_fd_sc_hd__nand3_1 _1576_ (.A(_0863_),
    .B(_0576_),
    .C(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__a221o_1 _1577_ (.A1(_0224_),
    .A2(\mem[11][4] ),
    .B1(\mem[8][4] ),
    .B2(_0837_),
    .C1(_0145_),
    .X(_0580_));
 sky130_fd_sc_hd__a221o_1 _1578_ (.A1(_0224_),
    .A2(\mem[15][4] ),
    .B1(\mem[12][4] ),
    .B2(_0245_),
    .C1(_0857_),
    .X(_0581_));
 sky130_fd_sc_hd__a22oi_1 _1579_ (.A1(_0136_),
    .A2(\mem[7][4] ),
    .B1(\mem[4][4] ),
    .B2(_0837_),
    .Y(_0582_));
 sky130_fd_sc_hd__a22oi_1 _1580_ (.A1(_0247_),
    .A2(\mem[3][4] ),
    .B1(\mem[1][4] ),
    .B2(_0137_),
    .Y(_0583_));
 sky130_fd_sc_hd__a22oi_1 _1581_ (.A1(_0866_),
    .A2(_0582_),
    .B1(_0583_),
    .B2(_0171_),
    .Y(_0584_));
 sky130_fd_sc_hd__nand3_1 _1582_ (.A(_0580_),
    .B(_0581_),
    .C(_0584_),
    .Y(_0585_));
 sky130_fd_sc_hd__nor2_1 _1583_ (.A(\mem[0][4] ),
    .B(_0830_),
    .Y(_0586_));
 sky130_fd_sc_hd__a41oi_4 _1584_ (.A1(_0157_),
    .A2(_0574_),
    .A3(_0579_),
    .A4(_0585_),
    .B1(_0586_),
    .Y(_0587_));
 sky130_fd_sc_hd__a22o_1 _1585_ (.A1(net102),
    .A2(_0789_),
    .B1(_0793_),
    .B2(_0587_),
    .X(_0074_));
 sky130_fd_sc_hd__a22oi_1 _1586_ (.A1(\mem[6][5] ),
    .A2(_0124_),
    .B1(_0862_),
    .B2(\mem[5][5] ),
    .Y(_0588_));
 sky130_fd_sc_hd__a21oi_1 _1587_ (.A1(\mem[2][5] ),
    .A2(_0152_),
    .B1(_0234_),
    .Y(_0589_));
 sky130_fd_sc_hd__a21oi_1 _1588_ (.A1(_0836_),
    .A2(_0588_),
    .B1(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__a222oi_1 _1589_ (.A1(_0136_),
    .A2(\mem[11][5] ),
    .B1(\mem[10][5] ),
    .B2(_0859_),
    .C1(_0137_),
    .C2(\mem[9][5] ),
    .Y(_0591_));
 sky130_fd_sc_hd__a221oi_1 _1590_ (.A1(_0224_),
    .A2(\mem[15][5] ),
    .B1(\mem[14][5] ),
    .B2(_0851_),
    .C1(_0785_),
    .Y(_0592_));
 sky130_fd_sc_hd__a211oi_1 _1591_ (.A1(_0848_),
    .A2(_0591_),
    .B1(_0592_),
    .C1(_0881_),
    .Y(_0593_));
 sky130_fd_sc_hd__a21oi_1 _1592_ (.A1(_0881_),
    .A2(_0590_),
    .B1(_0593_),
    .Y(_0594_));
 sky130_fd_sc_hd__nand2_1 _1593_ (.A(\mem[1][5] ),
    .B(_0150_),
    .Y(_0595_));
 sky130_fd_sc_hd__nand3_1 _1594_ (.A(_0331_),
    .B(\mem[8][5] ),
    .C(_0173_),
    .Y(_0596_));
 sky130_fd_sc_hd__o21ai_0 _1595_ (.A1(_0123_),
    .A2(_0595_),
    .B1(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__a32oi_1 _1596_ (.A1(_0331_),
    .A2(\mem[12][5] ),
    .A3(_0173_),
    .B1(_0243_),
    .B2(\mem[7][5] ),
    .Y(_0598_));
 sky130_fd_sc_hd__nand2_1 _1597_ (.A(_0198_),
    .B(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__o21ai_0 _1598_ (.A1(_0198_),
    .A2(_0597_),
    .B1(_0599_),
    .Y(_0600_));
 sky130_fd_sc_hd__nand2_1 _1599_ (.A(\mem[3][5] ),
    .B(_0847_),
    .Y(_0601_));
 sky130_fd_sc_hd__nand4_1 _1600_ (.A(_0331_),
    .B(_0197_),
    .C(\mem[13][5] ),
    .D(_0862_),
    .Y(_0602_));
 sky130_fd_sc_hd__o21ai_0 _1601_ (.A1(_0331_),
    .A2(_0601_),
    .B1(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__a311oi_1 _1602_ (.A1(\mem[4][5] ),
    .A2(_0838_),
    .A3(_0866_),
    .B1(_0824_),
    .C1(_0603_),
    .Y(_0604_));
 sky130_fd_sc_hd__nor2_1 _1603_ (.A(\mem[0][5] ),
    .B(_0309_),
    .Y(_0605_));
 sky130_fd_sc_hd__a31oi_1 _1604_ (.A1(_0594_),
    .A2(_0600_),
    .A3(_0604_),
    .B1(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__a22o_1 _1605_ (.A1(net103),
    .A2(_0789_),
    .B1(_0793_),
    .B2(_0606_),
    .X(_0075_));
 sky130_fd_sc_hd__nand2_1 _1606_ (.A(net104),
    .B(_0791_),
    .Y(_0607_));
 sky130_fd_sc_hd__a22o_1 _1607_ (.A1(\mem[14][6] ),
    .A2(_0182_),
    .B1(_0150_),
    .B2(\mem[13][6] ),
    .X(_0608_));
 sky130_fd_sc_hd__a22oi_1 _1608_ (.A1(\mem[8][6] ),
    .A2(_0173_),
    .B1(_0860_),
    .B2(\mem[10][6] ),
    .Y(_0609_));
 sky130_fd_sc_hd__a21oi_1 _1609_ (.A1(\mem[9][6] ),
    .A2(_0150_),
    .B1(_0840_),
    .Y(_0610_));
 sky130_fd_sc_hd__a21oi_1 _1610_ (.A1(_0609_),
    .A2(_0610_),
    .B1(_0881_),
    .Y(_0611_));
 sky130_fd_sc_hd__o21ai_0 _1611_ (.A1(_0884_),
    .A2(_0608_),
    .B1(_0611_),
    .Y(_0612_));
 sky130_fd_sc_hd__mux2i_1 _1612_ (.A0(\mem[3][6] ),
    .A1(\mem[7][6] ),
    .S(_0835_),
    .Y(_0613_));
 sky130_fd_sc_hd__nor2_1 _1613_ (.A(_0162_),
    .B(_0613_),
    .Y(_0614_));
 sky130_fd_sc_hd__and3_1 _1614_ (.A(_0331_),
    .B(_0197_),
    .C(\mem[15][6] ),
    .X(_0615_));
 sky130_fd_sc_hd__o21ai_0 _1615_ (.A1(_0614_),
    .A2(_0615_),
    .B1(_0218_),
    .Y(_0616_));
 sky130_fd_sc_hd__mux2i_1 _1616_ (.A0(\mem[2][6] ),
    .A1(\mem[6][6] ),
    .S(_0197_),
    .Y(_0617_));
 sky130_fd_sc_hd__nand3_1 _1617_ (.A(_0208_),
    .B(\mem[5][6] ),
    .C(_0193_),
    .Y(_0618_));
 sky130_fd_sc_hd__o21ai_0 _1618_ (.A1(_0320_),
    .A2(_0617_),
    .B1(_0618_),
    .Y(_0619_));
 sky130_fd_sc_hd__nand2_1 _1619_ (.A(_0881_),
    .B(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__mux2_1 _1620_ (.A0(\mem[4][6] ),
    .A1(\mem[12][6] ),
    .S(_0806_),
    .X(_0621_));
 sky130_fd_sc_hd__nand3_1 _1621_ (.A(_0166_),
    .B(_0841_),
    .C(\mem[11][6] ),
    .Y(_0622_));
 sky130_fd_sc_hd__nand3b_1 _1622_ (.A_N(_0806_),
    .B(\mem[1][6] ),
    .C(_0226_),
    .Y(_0623_));
 sky130_fd_sc_hd__a21oi_1 _1623_ (.A1(_0622_),
    .A2(_0623_),
    .B1(_0840_),
    .Y(_0624_));
 sky130_fd_sc_hd__a311oi_2 _1624_ (.A1(_0836_),
    .A2(_0838_),
    .A3(_0621_),
    .B1(_0624_),
    .C1(_0132_),
    .Y(_0625_));
 sky130_fd_sc_hd__nand4_2 _1625_ (.A(_0612_),
    .B(_0616_),
    .C(_0620_),
    .D(_0625_),
    .Y(_0626_));
 sky130_fd_sc_hd__o2111ai_2 _1626_ (.A1(\mem[0][6] ),
    .A2(_0831_),
    .B1(_0626_),
    .C1(_0826_),
    .D1(_0827_),
    .Y(_0627_));
 sky130_fd_sc_hd__o21ai_0 _1627_ (.A1(_0231_),
    .A2(_0607_),
    .B1(_0627_),
    .Y(_0076_));
 sky130_fd_sc_hd__a22oi_2 _1628_ (.A1(\mem[6][7] ),
    .A2(_0804_),
    .B1(_0814_),
    .B2(\mem[5][7] ),
    .Y(_0628_));
 sky130_fd_sc_hd__nand2_1 _1629_ (.A(_0836_),
    .B(_0628_),
    .Y(_0629_));
 sky130_fd_sc_hd__a22o_1 _1630_ (.A1(\mem[13][7] ),
    .A2(_0178_),
    .B1(_0171_),
    .B2(\mem[1][7] ),
    .X(_0630_));
 sky130_fd_sc_hd__a32oi_2 _1631_ (.A1(\mem[3][7] ),
    .A2(_0243_),
    .A3(_0629_),
    .B1(_0630_),
    .B2(_0863_),
    .Y(_0631_));
 sky130_fd_sc_hd__nand2_1 _1632_ (.A(\mem[14][7] ),
    .B(_0143_),
    .Y(_0632_));
 sky130_fd_sc_hd__a21oi_1 _1633_ (.A1(\mem[4][7] ),
    .A2(_0245_),
    .B1(_0122_),
    .Y(_0633_));
 sky130_fd_sc_hd__a221oi_1 _1634_ (.A1(_0832_),
    .A2(_0632_),
    .B1(_0633_),
    .B2(_0628_),
    .C1(_0276_),
    .Y(_0634_));
 sky130_fd_sc_hd__a311oi_2 _1635_ (.A1(\mem[8][7] ),
    .A2(_0838_),
    .A3(_0174_),
    .B1(_0824_),
    .C1(_0634_),
    .Y(_0635_));
 sky130_fd_sc_hd__a32o_1 _1636_ (.A1(_0276_),
    .A2(\mem[2][7] ),
    .A3(_0124_),
    .B1(_0272_),
    .B2(\mem[7][7] ),
    .X(_0636_));
 sky130_fd_sc_hd__a222oi_1 _1637_ (.A1(_0849_),
    .A2(\mem[11][7] ),
    .B1(\mem[10][7] ),
    .B2(_0817_),
    .C1(_0140_),
    .C2(\mem[9][7] ),
    .Y(_0637_));
 sky130_fd_sc_hd__a221oi_1 _1638_ (.A1(_0224_),
    .A2(\mem[15][7] ),
    .B1(\mem[12][7] ),
    .B2(_0245_),
    .C1(_0785_),
    .Y(_0638_));
 sky130_fd_sc_hd__a211oi_1 _1639_ (.A1(_0848_),
    .A2(_0637_),
    .B1(_0638_),
    .C1(_0869_),
    .Y(_0639_));
 sky130_fd_sc_hd__a21oi_1 _1640_ (.A1(_0881_),
    .A2(_0636_),
    .B1(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__nor2_1 _1641_ (.A(\mem[0][7] ),
    .B(_0309_),
    .Y(_0641_));
 sky130_fd_sc_hd__a31oi_4 _1642_ (.A1(_0631_),
    .A2(_0635_),
    .A3(_0640_),
    .B1(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__a22o_1 _1643_ (.A1(net105),
    .A2(_0789_),
    .B1(_0793_),
    .B2(_0642_),
    .X(_0077_));
 sky130_fd_sc_hd__a22oi_1 _1644_ (.A1(\mem[12][8] ),
    .A2(_0850_),
    .B1(_0140_),
    .B2(\mem[13][8] ),
    .Y(_0643_));
 sky130_fd_sc_hd__a22oi_1 _1645_ (.A1(\mem[4][8] ),
    .A2(_0245_),
    .B1(_0163_),
    .B2(\mem[6][8] ),
    .Y(_0644_));
 sky130_fd_sc_hd__a21oi_1 _1646_ (.A1(_0247_),
    .A2(\mem[7][8] ),
    .B1(_0199_),
    .Y(_0645_));
 sky130_fd_sc_hd__a221oi_1 _1647_ (.A1(_0331_),
    .A2(_0643_),
    .B1(_0644_),
    .B2(_0645_),
    .C1(_0848_),
    .Y(_0646_));
 sky130_fd_sc_hd__mux2i_1 _1648_ (.A0(\mem[2][8] ),
    .A1(\mem[10][8] ),
    .S(_0199_),
    .Y(_0647_));
 sky130_fd_sc_hd__a22oi_1 _1649_ (.A1(_0149_),
    .A2(\mem[15][8] ),
    .B1(\mem[14][8] ),
    .B2(_0182_),
    .Y(_0648_));
 sky130_fd_sc_hd__o22ai_1 _1650_ (.A1(_0165_),
    .A2(_0647_),
    .B1(_0648_),
    .B2(_0857_),
    .Y(_0649_));
 sky130_fd_sc_hd__mux2i_1 _1651_ (.A0(\mem[3][8] ),
    .A1(\mem[11][8] ),
    .S(_0166_),
    .Y(_0650_));
 sky130_fd_sc_hd__nand3_1 _1652_ (.A(\mem[8][8] ),
    .B(_0838_),
    .C(_0174_),
    .Y(_0651_));
 sky130_fd_sc_hd__o21ai_0 _1653_ (.A1(_0282_),
    .A2(_0650_),
    .B1(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__nor3_1 _1654_ (.A(_0646_),
    .B(_0649_),
    .C(_0652_),
    .Y(_0653_));
 sky130_fd_sc_hd__mux2i_1 _1655_ (.A0(\mem[1][8] ),
    .A1(\mem[5][8] ),
    .S(_0867_),
    .Y(_0654_));
 sky130_fd_sc_hd__nand2_1 _1656_ (.A(\mem[9][8] ),
    .B(_0174_),
    .Y(_0655_));
 sky130_fd_sc_hd__o21ai_0 _1657_ (.A1(_0123_),
    .A2(_0654_),
    .B1(_0655_),
    .Y(_0656_));
 sky130_fd_sc_hd__a21oi_1 _1658_ (.A1(_0863_),
    .A2(_0656_),
    .B1(_0132_),
    .Y(_0657_));
 sky130_fd_sc_hd__nor2_1 _1659_ (.A(\mem[0][8] ),
    .B(_0129_),
    .Y(_0658_));
 sky130_fd_sc_hd__a21oi_4 _1660_ (.A1(_0653_),
    .A2(_0657_),
    .B1(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__a22o_1 _1661_ (.A1(net106),
    .A2(_0789_),
    .B1(_0793_),
    .B2(_0659_),
    .X(_0078_));
 sky130_fd_sc_hd__a32oi_1 _1662_ (.A1(_0832_),
    .A2(\mem[8][9] ),
    .A3(_0842_),
    .B1(_0243_),
    .B2(\mem[3][9] ),
    .Y(_0660_));
 sky130_fd_sc_hd__nand2_1 _1663_ (.A(_0884_),
    .B(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__a22oi_1 _1664_ (.A1(_0841_),
    .A2(\mem[7][9] ),
    .B1(\mem[4][9] ),
    .B2(_0842_),
    .Y(_0662_));
 sky130_fd_sc_hd__a21oi_1 _1665_ (.A1(\mem[5][9] ),
    .A2(_0226_),
    .B1(_0154_),
    .Y(_0663_));
 sky130_fd_sc_hd__a21oi_1 _1666_ (.A1(_0149_),
    .A2(\mem[15][9] ),
    .B1(_0857_),
    .Y(_0664_));
 sky130_fd_sc_hd__a21oi_1 _1667_ (.A1(_0662_),
    .A2(_0663_),
    .B1(_0664_),
    .Y(_0665_));
 sky130_fd_sc_hd__nand2_1 _1668_ (.A(\mem[12][9] ),
    .B(_0842_),
    .Y(_0666_));
 sky130_fd_sc_hd__a221oi_1 _1669_ (.A1(_0224_),
    .A2(\mem[11][9] ),
    .B1(\mem[10][9] ),
    .B2(_0859_),
    .C1(_0867_),
    .Y(_0667_));
 sky130_fd_sc_hd__a211oi_1 _1670_ (.A1(_0840_),
    .A2(_0666_),
    .B1(_0667_),
    .C1(_0869_),
    .Y(_0668_));
 sky130_fd_sc_hd__a21oi_1 _1671_ (.A1(_0661_),
    .A2(_0665_),
    .B1(_0668_),
    .Y(_0669_));
 sky130_fd_sc_hd__mux2i_1 _1672_ (.A0(\mem[9][9] ),
    .A1(\mem[13][9] ),
    .S(_0207_),
    .Y(_0670_));
 sky130_fd_sc_hd__nand2_1 _1673_ (.A(_0162_),
    .B(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__a21o_1 _1674_ (.A1(_0276_),
    .A2(\mem[1][9] ),
    .B1(_0832_),
    .X(_0672_));
 sky130_fd_sc_hd__mux2i_1 _1675_ (.A0(\mem[2][9] ),
    .A1(\mem[6][9] ),
    .S(_0867_),
    .Y(_0673_));
 sky130_fd_sc_hd__nand2_1 _1676_ (.A(\mem[14][9] ),
    .B(_0178_),
    .Y(_0674_));
 sky130_fd_sc_hd__o21ai_2 _1677_ (.A1(_0133_),
    .A2(_0673_),
    .B1(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__a32oi_4 _1678_ (.A1(_0193_),
    .A2(_0671_),
    .A3(_0672_),
    .B1(_0675_),
    .B2(_0860_),
    .Y(_0676_));
 sky130_fd_sc_hd__nor2_1 _1679_ (.A(\mem[0][9] ),
    .B(_0309_),
    .Y(_0677_));
 sky130_fd_sc_hd__a31oi_4 _1680_ (.A1(_0157_),
    .A2(_0669_),
    .A3(_0676_),
    .B1(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__a22o_1 _1681_ (.A1(net107),
    .A2(_0789_),
    .B1(_0793_),
    .B2(_0678_),
    .X(_0079_));
 sky130_fd_sc_hd__nand2b_1 _1682_ (.A_N(net72),
    .B(_0752_),
    .Y(_0679_));
 sky130_fd_sc_hd__clkbuf_2 _1683_ (.A(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__nand2_1 _1684_ (.A(net38),
    .B(_0759_),
    .Y(_0681_));
 sky130_fd_sc_hd__nor2_1 _1685_ (.A(_0680_),
    .B(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__mux2i_1 _1686_ (.A0(_0777_),
    .A1(_0878_),
    .S(_0753_),
    .Y(_0683_));
 sky130_fd_sc_hd__nand2_1 _1687_ (.A(_0754_),
    .B(_0786_),
    .Y(_0684_));
 sky130_fd_sc_hd__a31oi_4 _1688_ (.A1(_0744_),
    .A2(_0775_),
    .A3(_0776_),
    .B1(_0684_),
    .Y(_0685_));
 sky130_fd_sc_hd__and2_0 _1689_ (.A(_0825_),
    .B(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__a221o_1 _1690_ (.A1(net108),
    .A2(_0680_),
    .B1(_0682_),
    .B2(_0683_),
    .C1(_0686_),
    .X(_0080_));
 sky130_fd_sc_hd__nand3_4 _1691_ (.A(_0754_),
    .B(_0777_),
    .C(_0786_),
    .Y(_0687_));
 sky130_fd_sc_hd__clkbuf_4 _1692_ (.A(_0680_),
    .X(_0688_));
 sky130_fd_sc_hd__nand2_1 _1693_ (.A(net109),
    .B(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__o21ai_0 _1694_ (.A1(_0131_),
    .A2(_0687_),
    .B1(_0689_),
    .Y(_0081_));
 sky130_fd_sc_hd__clkbuf_4 _1695_ (.A(_0685_),
    .X(_0690_));
 sky130_fd_sc_hd__a22o_1 _1696_ (.A1(net110),
    .A2(_0688_),
    .B1(_0159_),
    .B2(_0690_),
    .X(_0082_));
 sky130_fd_sc_hd__a22o_1 _1697_ (.A1(net111),
    .A2(_0688_),
    .B1(_0189_),
    .B2(_0690_),
    .X(_0083_));
 sky130_fd_sc_hd__a22o_1 _1698_ (.A1(net112),
    .A2(_0688_),
    .B1(_0212_),
    .B2(_0690_),
    .X(_0084_));
 sky130_fd_sc_hd__a22o_1 _1699_ (.A1(net113),
    .A2(_0688_),
    .B1(_0230_),
    .B2(_0690_),
    .X(_0085_));
 sky130_fd_sc_hd__o21ai_0 _1700_ (.A1(\mem[0][15] ),
    .A2(_0831_),
    .B1(_0254_),
    .Y(_0691_));
 sky130_fd_sc_hd__nand2_1 _1701_ (.A(net114),
    .B(_0688_),
    .Y(_0692_));
 sky130_fd_sc_hd__o21ai_0 _1702_ (.A1(_0691_),
    .A2(_0687_),
    .B1(_0692_),
    .Y(_0086_));
 sky130_fd_sc_hd__buf_4 _1703_ (.A(_0680_),
    .X(_0693_));
 sky130_fd_sc_hd__a22o_1 _1704_ (.A1(net115),
    .A2(_0693_),
    .B1(_0270_),
    .B2(_0690_),
    .X(_0087_));
 sky130_fd_sc_hd__a22o_1 _1705_ (.A1(net116),
    .A2(_0693_),
    .B1(_0291_),
    .B2(_0690_),
    .X(_0088_));
 sky130_fd_sc_hd__a22o_1 _1706_ (.A1(net117),
    .A2(_0693_),
    .B1(_0311_),
    .B2(_0690_),
    .X(_0089_));
 sky130_fd_sc_hd__a22o_1 _1707_ (.A1(net118),
    .A2(_0693_),
    .B1(_0329_),
    .B2(_0690_),
    .X(_0090_));
 sky130_fd_sc_hd__nor3_1 _1708_ (.A(_0753_),
    .B(_0680_),
    .C(_0681_),
    .Y(_0694_));
 sky130_fd_sc_hd__nand3_1 _1709_ (.A(_0753_),
    .B(_0875_),
    .C(_0786_),
    .Y(_0695_));
 sky130_fd_sc_hd__nand2_1 _1710_ (.A(net119),
    .B(_0680_),
    .Y(_0696_));
 sky130_fd_sc_hd__o21ai_0 _1711_ (.A1(_0681_),
    .A2(_0695_),
    .B1(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__a221o_1 _1712_ (.A1(_0349_),
    .A2(_0685_),
    .B1(_0694_),
    .B2(net75),
    .C1(_0697_),
    .X(_0091_));
 sky130_fd_sc_hd__a22o_1 _1713_ (.A1(net120),
    .A2(_0693_),
    .B1(_0364_),
    .B2(_0690_),
    .X(_0092_));
 sky130_fd_sc_hd__a22o_1 _1714_ (.A1(net121),
    .A2(_0693_),
    .B1(_0379_),
    .B2(_0690_),
    .X(_0093_));
 sky130_fd_sc_hd__clkbuf_4 _1715_ (.A(_0685_),
    .X(_0698_));
 sky130_fd_sc_hd__a22o_1 _1716_ (.A1(net122),
    .A2(_0693_),
    .B1(_0395_),
    .B2(_0698_),
    .X(_0094_));
 sky130_fd_sc_hd__a22o_1 _1717_ (.A1(net123),
    .A2(_0693_),
    .B1(_0409_),
    .B2(_0698_),
    .X(_0095_));
 sky130_fd_sc_hd__a22o_1 _1718_ (.A1(net124),
    .A2(_0693_),
    .B1(_0423_),
    .B2(_0698_),
    .X(_0096_));
 sky130_fd_sc_hd__a22o_1 _1719_ (.A1(net125),
    .A2(_0693_),
    .B1(_0440_),
    .B2(_0698_),
    .X(_0097_));
 sky130_fd_sc_hd__clkbuf_4 _1720_ (.A(_0680_),
    .X(_0699_));
 sky130_fd_sc_hd__a22o_1 _1721_ (.A1(net126),
    .A2(_0699_),
    .B1(_0457_),
    .B2(_0698_),
    .X(_0098_));
 sky130_fd_sc_hd__o21ai_0 _1722_ (.A1(\mem[0][27] ),
    .A2(_0831_),
    .B1(_0471_),
    .Y(_0700_));
 sky130_fd_sc_hd__nand2_1 _1723_ (.A(net127),
    .B(_0688_),
    .Y(_0701_));
 sky130_fd_sc_hd__o21ai_0 _1724_ (.A1(_0700_),
    .A2(_0687_),
    .B1(_0701_),
    .Y(_0099_));
 sky130_fd_sc_hd__a22o_1 _1725_ (.A1(net128),
    .A2(_0699_),
    .B1(_0488_),
    .B2(_0698_),
    .X(_0100_));
 sky130_fd_sc_hd__a22o_1 _1726_ (.A1(net129),
    .A2(_0699_),
    .B1(_0508_),
    .B2(_0698_),
    .X(_0101_));
 sky130_fd_sc_hd__nand2_1 _1727_ (.A(net130),
    .B(_0680_),
    .Y(_0702_));
 sky130_fd_sc_hd__nor2_1 _1728_ (.A(_0758_),
    .B(_0699_),
    .Y(_0703_));
 sky130_fd_sc_hd__nand2_1 _1729_ (.A(_0759_),
    .B(_0703_),
    .Y(_0704_));
 sky130_fd_sc_hd__xor2_1 _1730_ (.A(_0878_),
    .B(_0875_),
    .X(_0705_));
 sky130_fd_sc_hd__nor4_1 _1731_ (.A(_0753_),
    .B(_0774_),
    .C(_0681_),
    .D(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hd__nand3_1 _1732_ (.A(net38),
    .B(_0753_),
    .C(_0759_),
    .Y(_0707_));
 sky130_fd_sc_hd__o21ai_0 _1733_ (.A1(_0745_),
    .A2(_0707_),
    .B1(_0702_),
    .Y(_0708_));
 sky130_fd_sc_hd__a31oi_1 _1734_ (.A1(_0744_),
    .A2(_0776_),
    .A3(_0706_),
    .B1(_0708_),
    .Y(_0709_));
 sky130_fd_sc_hd__nand3_1 _1735_ (.A(_0754_),
    .B(_0777_),
    .C(_0526_),
    .Y(_0710_));
 sky130_fd_sc_hd__a22oi_1 _1736_ (.A1(_0702_),
    .A2(_0704_),
    .B1(_0709_),
    .B2(_0710_),
    .Y(_0102_));
 sky130_fd_sc_hd__nand2_1 _1737_ (.A(net131),
    .B(_0688_),
    .Y(_0711_));
 sky130_fd_sc_hd__o21ai_0 _1738_ (.A1(_0540_),
    .A2(_0687_),
    .B1(_0711_),
    .Y(_0103_));
 sky130_fd_sc_hd__a22o_1 _1739_ (.A1(net132),
    .A2(_0699_),
    .B1(_0558_),
    .B2(_0698_),
    .X(_0104_));
 sky130_fd_sc_hd__a21oi_1 _1740_ (.A1(_0875_),
    .A2(_0774_),
    .B1(_0753_),
    .Y(_0712_));
 sky130_fd_sc_hd__o22ai_1 _1741_ (.A1(_0753_),
    .A2(_0744_),
    .B1(_0776_),
    .B2(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__a222oi_1 _1742_ (.A1(net133),
    .A2(_0699_),
    .B1(_0572_),
    .B2(_0685_),
    .C1(_0682_),
    .C2(_0713_),
    .Y(_0714_));
 sky130_fd_sc_hd__inv_1 _1743_ (.A(_0714_),
    .Y(_0105_));
 sky130_fd_sc_hd__nand2_1 _1744_ (.A(_0587_),
    .B(_0685_),
    .Y(_0715_));
 sky130_fd_sc_hd__nand2_1 _1745_ (.A(net134),
    .B(_0688_),
    .Y(_0716_));
 sky130_fd_sc_hd__o311ai_0 _1746_ (.A1(_0744_),
    .A2(_0680_),
    .A3(_0707_),
    .B1(_0715_),
    .C1(_0716_),
    .Y(_0106_));
 sky130_fd_sc_hd__a22o_1 _1747_ (.A1(net135),
    .A2(_0699_),
    .B1(_0606_),
    .B2(_0698_),
    .X(_0107_));
 sky130_fd_sc_hd__o21ai_0 _1748_ (.A1(\mem[0][6] ),
    .A2(_0831_),
    .B1(_0626_),
    .Y(_0717_));
 sky130_fd_sc_hd__nand2_1 _1749_ (.A(net136),
    .B(_0688_),
    .Y(_0718_));
 sky130_fd_sc_hd__o21ai_0 _1750_ (.A1(_0717_),
    .A2(_0687_),
    .B1(_0718_),
    .Y(_0108_));
 sky130_fd_sc_hd__a22o_1 _1751_ (.A1(net137),
    .A2(_0699_),
    .B1(_0642_),
    .B2(_0698_),
    .X(_0109_));
 sky130_fd_sc_hd__a22o_1 _1752_ (.A1(net138),
    .A2(_0699_),
    .B1(_0659_),
    .B2(_0685_),
    .X(_0110_));
 sky130_fd_sc_hd__a22o_1 _1753_ (.A1(net139),
    .A2(_0699_),
    .B1(_0678_),
    .B2(_0685_),
    .X(_0111_));
 sky130_fd_sc_hd__xnor2_1 _1754_ (.A(\rd_ptr[0] ),
    .B(_0827_),
    .Y(_0719_));
 sky130_fd_sc_hd__nor2_1 _1755_ (.A(_0764_),
    .B(_0719_),
    .Y(_0112_));
 sky130_fd_sc_hd__nand3_1 _1756_ (.A(_0889_),
    .B(_0826_),
    .C(_0231_),
    .Y(_0720_));
 sky130_fd_sc_hd__o31ai_1 _1757_ (.A1(_0872_),
    .A2(_0764_),
    .A3(_0231_),
    .B1(_0720_),
    .Y(_0113_));
 sky130_fd_sc_hd__a21o_1 _1758_ (.A1(_0218_),
    .A2(_0827_),
    .B1(_0884_),
    .X(_0721_));
 sky130_fd_sc_hd__nand3_1 _1759_ (.A(_0884_),
    .B(_0218_),
    .C(_0827_),
    .Y(_0722_));
 sky130_fd_sc_hd__a21oi_1 _1760_ (.A1(_0721_),
    .A2(_0722_),
    .B1(_0764_),
    .Y(_0114_));
 sky130_fd_sc_hd__nor2_1 _1761_ (.A(_0833_),
    .B(_0763_),
    .Y(_0723_));
 sky130_fd_sc_hd__nor2_1 _1762_ (.A(_0881_),
    .B(_0763_),
    .Y(_0724_));
 sky130_fd_sc_hd__nand4_1 _1763_ (.A(_0198_),
    .B(\rd_ptr[0] ),
    .C(\rd_ptr[1] ),
    .D(_0827_),
    .Y(_0725_));
 sky130_fd_sc_hd__mux2_1 _1764_ (.A0(_0723_),
    .A1(_0724_),
    .S(_0725_),
    .X(_0115_));
 sky130_fd_sc_hd__nor2_1 _1765_ (.A(\rd_ptr[4] ),
    .B(_0763_),
    .Y(_0726_));
 sky130_fd_sc_hd__nand2_1 _1766_ (.A(\rd_ptr[4] ),
    .B(_0791_),
    .Y(_0727_));
 sky130_fd_sc_hd__a21oi_1 _1767_ (.A1(_0827_),
    .A2(_0303_),
    .B1(_0727_),
    .Y(_0728_));
 sky130_fd_sc_hd__a31o_1 _1768_ (.A1(_0827_),
    .A2(_0303_),
    .A3(_0726_),
    .B1(_0728_),
    .X(_0116_));
 sky130_fd_sc_hd__xnor2_1 _1769_ (.A(_0876_),
    .B(_0756_),
    .Y(_0729_));
 sky130_fd_sc_hd__nor2_1 _1770_ (.A(_0764_),
    .B(_0729_),
    .Y(_0117_));
 sky130_fd_sc_hd__nand2_1 _1771_ (.A(_0898_),
    .B(_0791_),
    .Y(_0730_));
 sky130_fd_sc_hd__nand3_1 _1772_ (.A(\wr_ptr[1] ),
    .B(_0757_),
    .C(_0826_),
    .Y(_0731_));
 sky130_fd_sc_hd__o21ai_0 _1773_ (.A1(_0757_),
    .A2(_0730_),
    .B1(_0731_),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_1 _1774_ (.A(_0903_),
    .Y(_0732_));
 sky130_fd_sc_hd__o21ai_0 _1775_ (.A1(_0732_),
    .A2(_0756_),
    .B1(\wr_ptr[2] ),
    .Y(_0733_));
 sky130_fd_sc_hd__or3_1 _1776_ (.A(\wr_ptr[2] ),
    .B(_0732_),
    .C(_0756_),
    .X(_0734_));
 sky130_fd_sc_hd__a21oi_1 _1777_ (.A1(_0733_),
    .A2(_0734_),
    .B1(_0764_),
    .Y(_0119_));
 sky130_fd_sc_hd__nand3_1 _1778_ (.A(\wr_ptr[2] ),
    .B(\wr_ptr[0] ),
    .C(\wr_ptr[1] ),
    .Y(_0735_));
 sky130_fd_sc_hd__o21ai_0 _1779_ (.A1(_0756_),
    .A2(_0735_),
    .B1(_0766_),
    .Y(_0736_));
 sky130_fd_sc_hd__or3_1 _1780_ (.A(_0766_),
    .B(_0756_),
    .C(_0735_),
    .X(_0737_));
 sky130_fd_sc_hd__a21oi_1 _1781_ (.A1(_0736_),
    .A2(_0737_),
    .B1(_0764_),
    .Y(_0120_));
 sky130_fd_sc_hd__nand3_1 _1782_ (.A(\wr_ptr[2] ),
    .B(_0766_),
    .C(_0903_),
    .Y(_0738_));
 sky130_fd_sc_hd__o21ai_0 _1783_ (.A1(_0756_),
    .A2(_0738_),
    .B1(\wr_ptr[4] ),
    .Y(_0739_));
 sky130_fd_sc_hd__or3_1 _1784_ (.A(\wr_ptr[4] ),
    .B(_0756_),
    .C(_0738_),
    .X(_0740_));
 sky130_fd_sc_hd__a21oi_1 _1785_ (.A1(_0739_),
    .A2(_0740_),
    .B1(_0764_),
    .Y(_0121_));
 sky130_fd_sc_hd__fa_4 _1786_ (.A(_0872_),
    .B(\wr_ptr[1] ),
    .CIN(_0873_),
    .COUT(_0874_),
    .SUM(_0875_));
 sky130_fd_sc_hd__ha_1 _1787_ (.A(\rd_ptr[0] ),
    .B(_0876_),
    .COUT(_0877_),
    .SUM(_0878_));
 sky130_fd_sc_hd__ha_1 _1788_ (.A(_0872_),
    .B(\wr_ptr[1] ),
    .COUT(_0879_),
    .SUM(_0880_));
 sky130_fd_sc_hd__ha_2 _1789_ (.A(_0881_),
    .B(\wr_ptr[3] ),
    .COUT(_0882_),
    .SUM(_0883_));
 sky130_fd_sc_hd__ha_1 _1790_ (.A(_0884_),
    .B(\wr_ptr[2] ),
    .COUT(_0885_),
    .SUM(_0886_));
 sky130_fd_sc_hd__ha_2 _1791_ (.A(_0887_),
    .B(_0872_),
    .COUT(_0888_),
    .SUM(_0889_));
 sky130_fd_sc_hd__ha_1 _1792_ (.A(_0887_),
    .B(\rd_ptr[1] ),
    .COUT(_0890_),
    .SUM(_0891_));
 sky130_fd_sc_hd__ha_1 _1793_ (.A(\rd_ptr[0] ),
    .B(_0872_),
    .COUT(_0892_),
    .SUM(_0893_));
 sky130_fd_sc_hd__ha_2 _1794_ (.A(\rd_ptr[0] ),
    .B(\rd_ptr[1] ),
    .COUT(_0894_),
    .SUM(_0895_));
 sky130_fd_sc_hd__ha_1 _1795_ (.A(_0876_),
    .B(_0896_),
    .COUT(_0897_),
    .SUM(_0898_));
 sky130_fd_sc_hd__ha_1 _1796_ (.A(_0876_),
    .B(\wr_ptr[1] ),
    .COUT(_0899_),
    .SUM(_0900_));
 sky130_fd_sc_hd__ha_1 _1797_ (.A(\wr_ptr[0] ),
    .B(_0896_),
    .COUT(_0901_),
    .SUM(_0902_));
 sky130_fd_sc_hd__ha_1 _1798_ (.A(\wr_ptr[0] ),
    .B(\wr_ptr[1] ),
    .COUT(_0903_),
    .SUM(_0904_));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[0]$_DFFE_PN0P_  (.D(_0048_),
    .Q(net76),
    .RESET_B(net1),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[10]$_DFFE_PN0P_  (.D(_0049_),
    .Q(net77),
    .RESET_B(net1),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[11]$_DFFE_PN0P_  (.D(_0050_),
    .Q(net78),
    .RESET_B(net1),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[12]$_DFFE_PN0P_  (.D(_0051_),
    .Q(net79),
    .RESET_B(net1),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[13]$_DFFE_PN0P_  (.D(_0052_),
    .Q(net80),
    .RESET_B(net1),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[14]$_DFFE_PN0P_  (.D(_0053_),
    .Q(net81),
    .RESET_B(net1),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[15]$_DFFE_PN0P_  (.D(_0054_),
    .Q(net82),
    .RESET_B(net1),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[16]$_DFFE_PN0P_  (.D(_0055_),
    .Q(net83),
    .RESET_B(net1),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[17]$_DFFE_PN0P_  (.D(_0056_),
    .Q(net84),
    .RESET_B(net1),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[18]$_DFFE_PN0P_  (.D(_0057_),
    .Q(net85),
    .RESET_B(net1),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[19]$_DFFE_PN0P_  (.D(_0058_),
    .Q(net86),
    .RESET_B(net1),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[1]$_DFFE_PN0P_  (.D(_0059_),
    .Q(net87),
    .RESET_B(net1),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[20]$_DFFE_PN0P_  (.D(_0060_),
    .Q(net88),
    .RESET_B(net1),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[21]$_DFFE_PN0P_  (.D(_0061_),
    .Q(net89),
    .RESET_B(net1),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[22]$_DFFE_PN0P_  (.D(_0062_),
    .Q(net90),
    .RESET_B(net1),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[23]$_DFFE_PN0P_  (.D(_0063_),
    .Q(net91),
    .RESET_B(net1),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[24]$_DFFE_PN0P_  (.D(_0064_),
    .Q(net92),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[25]$_DFFE_PN0P_  (.D(_0065_),
    .Q(net93),
    .RESET_B(net1),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[26]$_DFFE_PN0P_  (.D(_0066_),
    .Q(net94),
    .RESET_B(net1),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[27]$_DFFE_PN0P_  (.D(_0067_),
    .Q(net95),
    .RESET_B(net1),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[28]$_DFFE_PN0P_  (.D(_0068_),
    .Q(net96),
    .RESET_B(net1),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[29]$_DFFE_PN0P_  (.D(_0069_),
    .Q(net97),
    .RESET_B(net1),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[2]$_DFFE_PN0P_  (.D(_0070_),
    .Q(net98),
    .RESET_B(net1),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[30]$_DFFE_PN0P_  (.D(_0071_),
    .Q(net99),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[31]$_DFFE_PN0P_  (.D(_0072_),
    .Q(net100),
    .RESET_B(net1),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[3]$_DFFE_PN0P_  (.D(_0073_),
    .Q(net101),
    .RESET_B(net1),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[4]$_DFFE_PN0P_  (.D(_0074_),
    .Q(net102),
    .RESET_B(net1),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[5]$_DFFE_PN0P_  (.D(_0075_),
    .Q(net103),
    .RESET_B(net1),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[6]$_DFFE_PN0P_  (.D(_0076_),
    .Q(net104),
    .RESET_B(net1),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[7]$_DFFE_PN0P_  (.D(_0077_),
    .Q(net105),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[8]$_DFFE_PN0P_  (.D(_0078_),
    .Q(net106),
    .RESET_B(net1),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \ext_data_reg[9]$_DFFE_PN0P_  (.D(_0079_),
    .Q(net107),
    .RESET_B(net1),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][0]$_DFFE_PP_  (.D(_0016_),
    .DE(_0015_),
    .Q(\mem[0][0] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][10]$_DFFE_PP_  (.D(_0017_),
    .DE(_0015_),
    .Q(\mem[0][10] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][11]$_DFFE_PP_  (.D(_0018_),
    .DE(_0015_),
    .Q(\mem[0][11] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][12]$_DFFE_PP_  (.D(_0019_),
    .DE(_0015_),
    .Q(\mem[0][12] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][13]$_DFFE_PP_  (.D(_0020_),
    .DE(_0015_),
    .Q(\mem[0][13] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][14]$_DFFE_PP_  (.D(_0021_),
    .DE(_0015_),
    .Q(\mem[0][14] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][15]$_DFFE_PP_  (.D(_0022_),
    .DE(_0015_),
    .Q(\mem[0][15] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][16]$_DFFE_PP_  (.D(_0023_),
    .DE(_0015_),
    .Q(\mem[0][16] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][17]$_DFFE_PP_  (.D(_0024_),
    .DE(_0015_),
    .Q(\mem[0][17] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][18]$_DFFE_PP_  (.D(_0025_),
    .DE(_0015_),
    .Q(\mem[0][18] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][19]$_DFFE_PP_  (.D(_0026_),
    .DE(_0015_),
    .Q(\mem[0][19] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][1]$_DFFE_PP_  (.D(_0027_),
    .DE(_0015_),
    .Q(\mem[0][1] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][20]$_DFFE_PP_  (.D(_0028_),
    .DE(_0015_),
    .Q(\mem[0][20] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][21]$_DFFE_PP_  (.D(_0029_),
    .DE(_0015_),
    .Q(\mem[0][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][22]$_DFFE_PP_  (.D(_0030_),
    .DE(_0015_),
    .Q(\mem[0][22] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][23]$_DFFE_PP_  (.D(_0031_),
    .DE(_0015_),
    .Q(\mem[0][23] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][24]$_DFFE_PP_  (.D(_0032_),
    .DE(_0015_),
    .Q(\mem[0][24] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][25]$_DFFE_PP_  (.D(_0033_),
    .DE(_0015_),
    .Q(\mem[0][25] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][26]$_DFFE_PP_  (.D(_0034_),
    .DE(_0015_),
    .Q(\mem[0][26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][27]$_DFFE_PP_  (.D(_0035_),
    .DE(_0015_),
    .Q(\mem[0][27] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][28]$_DFFE_PP_  (.D(_0036_),
    .DE(_0015_),
    .Q(\mem[0][28] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][29]$_DFFE_PP_  (.D(_0037_),
    .DE(_0015_),
    .Q(\mem[0][29] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][2]$_DFFE_PP_  (.D(_0038_),
    .DE(_0015_),
    .Q(\mem[0][2] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][30]$_DFFE_PP_  (.D(_0039_),
    .DE(_0015_),
    .Q(\mem[0][30] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][31]$_DFFE_PP_  (.D(_0040_),
    .DE(_0015_),
    .Q(\mem[0][31] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][3]$_DFFE_PP_  (.D(_0041_),
    .DE(_0015_),
    .Q(\mem[0][3] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][4]$_DFFE_PP_  (.D(_0042_),
    .DE(_0015_),
    .Q(\mem[0][4] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][5]$_DFFE_PP_  (.D(_0043_),
    .DE(_0015_),
    .Q(\mem[0][5] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][6]$_DFFE_PP_  (.D(_0044_),
    .DE(_0015_),
    .Q(\mem[0][6] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][7]$_DFFE_PP_  (.D(_0045_),
    .DE(_0015_),
    .Q(\mem[0][7] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][8]$_DFFE_PP_  (.D(_0046_),
    .DE(_0015_),
    .Q(\mem[0][8] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][9]$_DFFE_PP_  (.D(_0047_),
    .DE(_0015_),
    .Q(\mem[0][9] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][0]$_DFFE_PP_  (.D(_0016_),
    .DE(net155),
    .Q(\mem[10][0] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][10]$_DFFE_PP_  (.D(_0017_),
    .DE(net155),
    .Q(\mem[10][10] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][11]$_DFFE_PP_  (.D(_0018_),
    .DE(net154),
    .Q(\mem[10][11] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][12]$_DFFE_PP_  (.D(_0019_),
    .DE(net155),
    .Q(\mem[10][12] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][13]$_DFFE_PP_  (.D(_0020_),
    .DE(net153),
    .Q(\mem[10][13] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][14]$_DFFE_PP_  (.D(_0021_),
    .DE(net154),
    .Q(\mem[10][14] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][15]$_DFFE_PP_  (.D(_0022_),
    .DE(net154),
    .Q(\mem[10][15] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][16]$_DFFE_PP_  (.D(_0023_),
    .DE(net153),
    .Q(\mem[10][16] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][17]$_DFFE_PP_  (.D(_0024_),
    .DE(net153),
    .Q(\mem[10][17] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][18]$_DFFE_PP_  (.D(_0025_),
    .DE(net153),
    .Q(\mem[10][18] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][19]$_DFFE_PP_  (.D(_0026_),
    .DE(net155),
    .Q(\mem[10][19] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][1]$_DFFE_PP_  (.D(_0027_),
    .DE(_0005_),
    .Q(\mem[10][1] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][20]$_DFFE_PP_  (.D(_0028_),
    .DE(net154),
    .Q(\mem[10][20] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][21]$_DFFE_PP_  (.D(_0029_),
    .DE(_0005_),
    .Q(\mem[10][21] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][22]$_DFFE_PP_  (.D(_0030_),
    .DE(net154),
    .Q(\mem[10][22] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][23]$_DFFE_PP_  (.D(_0031_),
    .DE(_0005_),
    .Q(\mem[10][23] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][24]$_DFFE_PP_  (.D(_0032_),
    .DE(_0005_),
    .Q(\mem[10][24] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][25]$_DFFE_PP_  (.D(_0033_),
    .DE(net153),
    .Q(\mem[10][25] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][26]$_DFFE_PP_  (.D(_0034_),
    .DE(net153),
    .Q(\mem[10][26] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][27]$_DFFE_PP_  (.D(_0035_),
    .DE(net155),
    .Q(\mem[10][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][28]$_DFFE_PP_  (.D(_0036_),
    .DE(net153),
    .Q(\mem[10][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][29]$_DFFE_PP_  (.D(_0037_),
    .DE(net154),
    .Q(\mem[10][29] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][2]$_DFFE_PP_  (.D(_0038_),
    .DE(net155),
    .Q(\mem[10][2] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][30]$_DFFE_PP_  (.D(_0039_),
    .DE(net153),
    .Q(\mem[10][30] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][31]$_DFFE_PP_  (.D(_0040_),
    .DE(net154),
    .Q(\mem[10][31] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][3]$_DFFE_PP_  (.D(_0041_),
    .DE(_0005_),
    .Q(\mem[10][3] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][4]$_DFFE_PP_  (.D(_0042_),
    .DE(_0005_),
    .Q(\mem[10][4] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][5]$_DFFE_PP_  (.D(_0043_),
    .DE(net154),
    .Q(\mem[10][5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][6]$_DFFE_PP_  (.D(_0044_),
    .DE(net155),
    .Q(\mem[10][6] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][7]$_DFFE_PP_  (.D(_0045_),
    .DE(_0005_),
    .Q(\mem[10][7] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][8]$_DFFE_PP_  (.D(_0046_),
    .DE(net153),
    .Q(\mem[10][8] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][9]$_DFFE_PP_  (.D(_0047_),
    .DE(net154),
    .Q(\mem[10][9] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][0]$_DFFE_PP_  (.D(_0016_),
    .DE(_0004_),
    .Q(\mem[11][0] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][10]$_DFFE_PP_  (.D(_0017_),
    .DE(net156),
    .Q(\mem[11][10] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][11]$_DFFE_PP_  (.D(_0018_),
    .DE(net158),
    .Q(\mem[11][11] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][12]$_DFFE_PP_  (.D(_0019_),
    .DE(net158),
    .Q(\mem[11][12] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][13]$_DFFE_PP_  (.D(_0020_),
    .DE(net157),
    .Q(\mem[11][13] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][14]$_DFFE_PP_  (.D(_0021_),
    .DE(net156),
    .Q(\mem[11][14] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][15]$_DFFE_PP_  (.D(_0022_),
    .DE(net158),
    .Q(\mem[11][15] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][16]$_DFFE_PP_  (.D(_0023_),
    .DE(net157),
    .Q(\mem[11][16] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][17]$_DFFE_PP_  (.D(_0024_),
    .DE(net157),
    .Q(\mem[11][17] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][18]$_DFFE_PP_  (.D(_0025_),
    .DE(net156),
    .Q(\mem[11][18] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][19]$_DFFE_PP_  (.D(_0026_),
    .DE(net158),
    .Q(\mem[11][19] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][1]$_DFFE_PP_  (.D(_0027_),
    .DE(_0004_),
    .Q(\mem[11][1] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][20]$_DFFE_PP_  (.D(_0028_),
    .DE(_0004_),
    .Q(\mem[11][20] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][21]$_DFFE_PP_  (.D(_0029_),
    .DE(net157),
    .Q(\mem[11][21] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][22]$_DFFE_PP_  (.D(_0030_),
    .DE(net156),
    .Q(\mem[11][22] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][23]$_DFFE_PP_  (.D(_0031_),
    .DE(net156),
    .Q(\mem[11][23] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][24]$_DFFE_PP_  (.D(_0032_),
    .DE(net157),
    .Q(\mem[11][24] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][25]$_DFFE_PP_  (.D(_0033_),
    .DE(net157),
    .Q(\mem[11][25] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][26]$_DFFE_PP_  (.D(_0034_),
    .DE(net157),
    .Q(\mem[11][26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][27]$_DFFE_PP_  (.D(_0035_),
    .DE(net156),
    .Q(\mem[11][27] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][28]$_DFFE_PP_  (.D(_0036_),
    .DE(net157),
    .Q(\mem[11][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][29]$_DFFE_PP_  (.D(_0037_),
    .DE(net158),
    .Q(\mem[11][29] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][2]$_DFFE_PP_  (.D(_0038_),
    .DE(net158),
    .Q(\mem[11][2] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][30]$_DFFE_PP_  (.D(_0039_),
    .DE(net157),
    .Q(\mem[11][30] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][31]$_DFFE_PP_  (.D(_0040_),
    .DE(net158),
    .Q(\mem[11][31] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][3]$_DFFE_PP_  (.D(_0041_),
    .DE(_0004_),
    .Q(\mem[11][3] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][4]$_DFFE_PP_  (.D(_0042_),
    .DE(net157),
    .Q(\mem[11][4] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][5]$_DFFE_PP_  (.D(_0043_),
    .DE(net156),
    .Q(\mem[11][5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][6]$_DFFE_PP_  (.D(_0044_),
    .DE(net158),
    .Q(\mem[11][6] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][7]$_DFFE_PP_  (.D(_0045_),
    .DE(_0004_),
    .Q(\mem[11][7] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][8]$_DFFE_PP_  (.D(_0046_),
    .DE(net157),
    .Q(\mem[11][8] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][9]$_DFFE_PP_  (.D(_0047_),
    .DE(net156),
    .Q(\mem[11][9] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][0]$_DFFE_PP_  (.D(_0016_),
    .DE(net161),
    .Q(\mem[12][0] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][10]$_DFFE_PP_  (.D(_0017_),
    .DE(net159),
    .Q(\mem[12][10] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][11]$_DFFE_PP_  (.D(_0018_),
    .DE(net159),
    .Q(\mem[12][11] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][12]$_DFFE_PP_  (.D(_0019_),
    .DE(net159),
    .Q(\mem[12][12] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][13]$_DFFE_PP_  (.D(_0020_),
    .DE(net160),
    .Q(\mem[12][13] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][14]$_DFFE_PP_  (.D(_0021_),
    .DE(net159),
    .Q(\mem[12][14] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][15]$_DFFE_PP_  (.D(_0022_),
    .DE(net159),
    .Q(\mem[12][15] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][16]$_DFFE_PP_  (.D(_0023_),
    .DE(net160),
    .Q(\mem[12][16] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][17]$_DFFE_PP_  (.D(_0024_),
    .DE(net159),
    .Q(\mem[12][17] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][18]$_DFFE_PP_  (.D(_0025_),
    .DE(net160),
    .Q(\mem[12][18] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][19]$_DFFE_PP_  (.D(_0026_),
    .DE(net159),
    .Q(\mem[12][19] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][1]$_DFFE_PP_  (.D(_0027_),
    .DE(net161),
    .Q(\mem[12][1] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][20]$_DFFE_PP_  (.D(_0028_),
    .DE(_0003_),
    .Q(\mem[12][20] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][21]$_DFFE_PP_  (.D(_0029_),
    .DE(net161),
    .Q(\mem[12][21] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][22]$_DFFE_PP_  (.D(_0030_),
    .DE(net160),
    .Q(\mem[12][22] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][23]$_DFFE_PP_  (.D(_0031_),
    .DE(net161),
    .Q(\mem[12][23] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][24]$_DFFE_PP_  (.D(_0032_),
    .DE(net161),
    .Q(\mem[12][24] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][25]$_DFFE_PP_  (.D(_0033_),
    .DE(net160),
    .Q(\mem[12][25] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][26]$_DFFE_PP_  (.D(_0034_),
    .DE(net160),
    .Q(\mem[12][26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][27]$_DFFE_PP_  (.D(_0035_),
    .DE(net159),
    .Q(\mem[12][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][28]$_DFFE_PP_  (.D(_0036_),
    .DE(net160),
    .Q(\mem[12][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][29]$_DFFE_PP_  (.D(_0037_),
    .DE(net160),
    .Q(\mem[12][29] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][2]$_DFFE_PP_  (.D(_0038_),
    .DE(net159),
    .Q(\mem[12][2] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][30]$_DFFE_PP_  (.D(_0039_),
    .DE(net161),
    .Q(\mem[12][30] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][31]$_DFFE_PP_  (.D(_0040_),
    .DE(net161),
    .Q(\mem[12][31] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][3]$_DFFE_PP_  (.D(_0041_),
    .DE(net161),
    .Q(\mem[12][3] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][4]$_DFFE_PP_  (.D(_0042_),
    .DE(net161),
    .Q(\mem[12][4] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][5]$_DFFE_PP_  (.D(_0043_),
    .DE(_0003_),
    .Q(\mem[12][5] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][6]$_DFFE_PP_  (.D(_0044_),
    .DE(net159),
    .Q(\mem[12][6] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][7]$_DFFE_PP_  (.D(_0045_),
    .DE(net161),
    .Q(\mem[12][7] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][8]$_DFFE_PP_  (.D(_0046_),
    .DE(net159),
    .Q(\mem[12][8] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][9]$_DFFE_PP_  (.D(_0047_),
    .DE(net160),
    .Q(\mem[12][9] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][0]$_DFFE_PP_  (.D(_0016_),
    .DE(net149),
    .Q(\mem[13][0] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][10]$_DFFE_PP_  (.D(_0017_),
    .DE(net148),
    .Q(\mem[13][10] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][11]$_DFFE_PP_  (.D(_0018_),
    .DE(net148),
    .Q(\mem[13][11] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][12]$_DFFE_PP_  (.D(_0019_),
    .DE(net148),
    .Q(\mem[13][12] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][13]$_DFFE_PP_  (.D(_0020_),
    .DE(net147),
    .Q(\mem[13][13] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][14]$_DFFE_PP_  (.D(_0021_),
    .DE(_0002_),
    .Q(\mem[13][14] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][15]$_DFFE_PP_  (.D(_0022_),
    .DE(net148),
    .Q(\mem[13][15] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][16]$_DFFE_PP_  (.D(_0023_),
    .DE(net147),
    .Q(\mem[13][16] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][17]$_DFFE_PP_  (.D(_0024_),
    .DE(net148),
    .Q(\mem[13][17] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][18]$_DFFE_PP_  (.D(_0025_),
    .DE(net147),
    .Q(\mem[13][18] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][19]$_DFFE_PP_  (.D(_0026_),
    .DE(net148),
    .Q(\mem[13][19] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][1]$_DFFE_PP_  (.D(_0027_),
    .DE(_0002_),
    .Q(\mem[13][1] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][20]$_DFFE_PP_  (.D(_0028_),
    .DE(_0002_),
    .Q(\mem[13][20] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][21]$_DFFE_PP_  (.D(_0029_),
    .DE(net147),
    .Q(\mem[13][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][22]$_DFFE_PP_  (.D(_0030_),
    .DE(net147),
    .Q(\mem[13][22] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][23]$_DFFE_PP_  (.D(_0031_),
    .DE(net149),
    .Q(\mem[13][23] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][24]$_DFFE_PP_  (.D(_0032_),
    .DE(net149),
    .Q(\mem[13][24] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][25]$_DFFE_PP_  (.D(_0033_),
    .DE(net147),
    .Q(\mem[13][25] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][26]$_DFFE_PP_  (.D(_0034_),
    .DE(net147),
    .Q(\mem[13][26] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][27]$_DFFE_PP_  (.D(_0035_),
    .DE(net148),
    .Q(\mem[13][27] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][28]$_DFFE_PP_  (.D(_0036_),
    .DE(net147),
    .Q(\mem[13][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][29]$_DFFE_PP_  (.D(_0037_),
    .DE(_0002_),
    .Q(\mem[13][29] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][2]$_DFFE_PP_  (.D(_0038_),
    .DE(net148),
    .Q(\mem[13][2] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][30]$_DFFE_PP_  (.D(_0039_),
    .DE(net149),
    .Q(\mem[13][30] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][31]$_DFFE_PP_  (.D(_0040_),
    .DE(net149),
    .Q(\mem[13][31] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][3]$_DFFE_PP_  (.D(_0041_),
    .DE(net149),
    .Q(\mem[13][3] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][4]$_DFFE_PP_  (.D(_0042_),
    .DE(net149),
    .Q(\mem[13][4] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][5]$_DFFE_PP_  (.D(_0043_),
    .DE(_0002_),
    .Q(\mem[13][5] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][6]$_DFFE_PP_  (.D(_0044_),
    .DE(net148),
    .Q(\mem[13][6] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][7]$_DFFE_PP_  (.D(_0045_),
    .DE(net147),
    .Q(\mem[13][7] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][8]$_DFFE_PP_  (.D(_0046_),
    .DE(net147),
    .Q(\mem[13][8] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][9]$_DFFE_PP_  (.D(_0047_),
    .DE(net148),
    .Q(\mem[13][9] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][0]$_DFFE_PP_  (.D(_0016_),
    .DE(_0001_),
    .Q(\mem[14][0] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][10]$_DFFE_PP_  (.D(_0017_),
    .DE(net141),
    .Q(\mem[14][10] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][11]$_DFFE_PP_  (.D(_0018_),
    .DE(net142),
    .Q(\mem[14][11] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][12]$_DFFE_PP_  (.D(_0019_),
    .DE(net142),
    .Q(\mem[14][12] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][13]$_DFFE_PP_  (.D(_0020_),
    .DE(net141),
    .Q(\mem[14][13] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][14]$_DFFE_PP_  (.D(_0021_),
    .DE(net142),
    .Q(\mem[14][14] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][15]$_DFFE_PP_  (.D(_0022_),
    .DE(net142),
    .Q(\mem[14][15] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][16]$_DFFE_PP_  (.D(_0023_),
    .DE(net141),
    .Q(\mem[14][16] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][17]$_DFFE_PP_  (.D(_0024_),
    .DE(net141),
    .Q(\mem[14][17] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][18]$_DFFE_PP_  (.D(_0025_),
    .DE(net141),
    .Q(\mem[14][18] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][19]$_DFFE_PP_  (.D(_0026_),
    .DE(net142),
    .Q(\mem[14][19] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][1]$_DFFE_PP_  (.D(_0027_),
    .DE(net143),
    .Q(\mem[14][1] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][20]$_DFFE_PP_  (.D(_0028_),
    .DE(net143),
    .Q(\mem[14][20] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][21]$_DFFE_PP_  (.D(_0029_),
    .DE(net141),
    .Q(\mem[14][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][22]$_DFFE_PP_  (.D(_0030_),
    .DE(net143),
    .Q(\mem[14][22] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][23]$_DFFE_PP_  (.D(_0031_),
    .DE(net143),
    .Q(\mem[14][23] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][24]$_DFFE_PP_  (.D(_0032_),
    .DE(net143),
    .Q(\mem[14][24] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][25]$_DFFE_PP_  (.D(_0033_),
    .DE(net141),
    .Q(\mem[14][25] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][26]$_DFFE_PP_  (.D(_0034_),
    .DE(net141),
    .Q(\mem[14][26] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][27]$_DFFE_PP_  (.D(_0035_),
    .DE(net141),
    .Q(\mem[14][27] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][28]$_DFFE_PP_  (.D(_0036_),
    .DE(net141),
    .Q(\mem[14][28] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][29]$_DFFE_PP_  (.D(_0037_),
    .DE(net142),
    .Q(\mem[14][29] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][2]$_DFFE_PP_  (.D(_0038_),
    .DE(net142),
    .Q(\mem[14][2] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][30]$_DFFE_PP_  (.D(_0039_),
    .DE(net143),
    .Q(\mem[14][30] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][31]$_DFFE_PP_  (.D(_0040_),
    .DE(net143),
    .Q(\mem[14][31] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][3]$_DFFE_PP_  (.D(_0041_),
    .DE(net143),
    .Q(\mem[14][3] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][4]$_DFFE_PP_  (.D(_0042_),
    .DE(net143),
    .Q(\mem[14][4] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][5]$_DFFE_PP_  (.D(_0043_),
    .DE(net142),
    .Q(\mem[14][5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][6]$_DFFE_PP_  (.D(_0044_),
    .DE(net142),
    .Q(\mem[14][6] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][7]$_DFFE_PP_  (.D(_0045_),
    .DE(net143),
    .Q(\mem[14][7] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][8]$_DFFE_PP_  (.D(_0046_),
    .DE(net141),
    .Q(\mem[14][8] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][9]$_DFFE_PP_  (.D(_0047_),
    .DE(net141),
    .Q(\mem[14][9] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][0]$_DFFE_PP_  (.D(_0016_),
    .DE(_0000_),
    .Q(\mem[15][0] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][10]$_DFFE_PP_  (.D(_0017_),
    .DE(net144),
    .Q(\mem[15][10] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][11]$_DFFE_PP_  (.D(_0018_),
    .DE(net146),
    .Q(\mem[15][11] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][12]$_DFFE_PP_  (.D(_0019_),
    .DE(net146),
    .Q(\mem[15][12] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][13]$_DFFE_PP_  (.D(_0020_),
    .DE(net144),
    .Q(\mem[15][13] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][14]$_DFFE_PP_  (.D(_0021_),
    .DE(net146),
    .Q(\mem[15][14] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][15]$_DFFE_PP_  (.D(_0022_),
    .DE(net144),
    .Q(\mem[15][15] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][16]$_DFFE_PP_  (.D(_0023_),
    .DE(net145),
    .Q(\mem[15][16] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][17]$_DFFE_PP_  (.D(_0024_),
    .DE(net144),
    .Q(\mem[15][17] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][18]$_DFFE_PP_  (.D(_0025_),
    .DE(net145),
    .Q(\mem[15][18] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][19]$_DFFE_PP_  (.D(_0026_),
    .DE(net146),
    .Q(\mem[15][19] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][1]$_DFFE_PP_  (.D(_0027_),
    .DE(net146),
    .Q(\mem[15][1] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][20]$_DFFE_PP_  (.D(_0028_),
    .DE(net146),
    .Q(\mem[15][20] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][21]$_DFFE_PP_  (.D(_0029_),
    .DE(net145),
    .Q(\mem[15][21] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][22]$_DFFE_PP_  (.D(_0030_),
    .DE(_0000_),
    .Q(\mem[15][22] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][23]$_DFFE_PP_  (.D(_0031_),
    .DE(_0000_),
    .Q(\mem[15][23] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][24]$_DFFE_PP_  (.D(_0032_),
    .DE(_0000_),
    .Q(\mem[15][24] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][25]$_DFFE_PP_  (.D(_0033_),
    .DE(net145),
    .Q(\mem[15][25] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][26]$_DFFE_PP_  (.D(_0034_),
    .DE(net144),
    .Q(\mem[15][26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][27]$_DFFE_PP_  (.D(_0035_),
    .DE(net146),
    .Q(\mem[15][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][28]$_DFFE_PP_  (.D(_0036_),
    .DE(net145),
    .Q(\mem[15][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][29]$_DFFE_PP_  (.D(_0037_),
    .DE(net146),
    .Q(\mem[15][29] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][2]$_DFFE_PP_  (.D(_0038_),
    .DE(net146),
    .Q(\mem[15][2] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][30]$_DFFE_PP_  (.D(_0039_),
    .DE(_0000_),
    .Q(\mem[15][30] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][31]$_DFFE_PP_  (.D(_0040_),
    .DE(net145),
    .Q(\mem[15][31] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][3]$_DFFE_PP_  (.D(_0041_),
    .DE(_0000_),
    .Q(\mem[15][3] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][4]$_DFFE_PP_  (.D(_0042_),
    .DE(_0000_),
    .Q(\mem[15][4] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][5]$_DFFE_PP_  (.D(_0043_),
    .DE(net144),
    .Q(\mem[15][5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][6]$_DFFE_PP_  (.D(_0044_),
    .DE(net146),
    .Q(\mem[15][6] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][7]$_DFFE_PP_  (.D(_0045_),
    .DE(net145),
    .Q(\mem[15][7] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][8]$_DFFE_PP_  (.D(_0046_),
    .DE(net144),
    .Q(\mem[15][8] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][9]$_DFFE_PP_  (.D(_0047_),
    .DE(net144),
    .Q(\mem[15][9] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][0]$_DFFE_PP_  (.D(_0016_),
    .DE(_0014_),
    .Q(\mem[1][0] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][10]$_DFFE_PP_  (.D(_0017_),
    .DE(_0014_),
    .Q(\mem[1][10] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][11]$_DFFE_PP_  (.D(_0018_),
    .DE(_0014_),
    .Q(\mem[1][11] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][12]$_DFFE_PP_  (.D(_0019_),
    .DE(_0014_),
    .Q(\mem[1][12] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][13]$_DFFE_PP_  (.D(_0020_),
    .DE(_0014_),
    .Q(\mem[1][13] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][14]$_DFFE_PP_  (.D(_0021_),
    .DE(_0014_),
    .Q(\mem[1][14] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][15]$_DFFE_PP_  (.D(_0022_),
    .DE(_0014_),
    .Q(\mem[1][15] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][16]$_DFFE_PP_  (.D(_0023_),
    .DE(_0014_),
    .Q(\mem[1][16] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][17]$_DFFE_PP_  (.D(_0024_),
    .DE(_0014_),
    .Q(\mem[1][17] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][18]$_DFFE_PP_  (.D(_0025_),
    .DE(_0014_),
    .Q(\mem[1][18] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][19]$_DFFE_PP_  (.D(_0026_),
    .DE(_0014_),
    .Q(\mem[1][19] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][1]$_DFFE_PP_  (.D(_0027_),
    .DE(_0014_),
    .Q(\mem[1][1] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][20]$_DFFE_PP_  (.D(_0028_),
    .DE(_0014_),
    .Q(\mem[1][20] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][21]$_DFFE_PP_  (.D(_0029_),
    .DE(_0014_),
    .Q(\mem[1][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][22]$_DFFE_PP_  (.D(_0030_),
    .DE(_0014_),
    .Q(\mem[1][22] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][23]$_DFFE_PP_  (.D(_0031_),
    .DE(_0014_),
    .Q(\mem[1][23] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][24]$_DFFE_PP_  (.D(_0032_),
    .DE(_0014_),
    .Q(\mem[1][24] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][25]$_DFFE_PP_  (.D(_0033_),
    .DE(_0014_),
    .Q(\mem[1][25] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][26]$_DFFE_PP_  (.D(_0034_),
    .DE(_0014_),
    .Q(\mem[1][26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][27]$_DFFE_PP_  (.D(_0035_),
    .DE(_0014_),
    .Q(\mem[1][27] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][28]$_DFFE_PP_  (.D(_0036_),
    .DE(_0014_),
    .Q(\mem[1][28] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][29]$_DFFE_PP_  (.D(_0037_),
    .DE(_0014_),
    .Q(\mem[1][29] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][2]$_DFFE_PP_  (.D(_0038_),
    .DE(_0014_),
    .Q(\mem[1][2] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][30]$_DFFE_PP_  (.D(_0039_),
    .DE(_0014_),
    .Q(\mem[1][30] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][31]$_DFFE_PP_  (.D(_0040_),
    .DE(_0014_),
    .Q(\mem[1][31] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][3]$_DFFE_PP_  (.D(_0041_),
    .DE(_0014_),
    .Q(\mem[1][3] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][4]$_DFFE_PP_  (.D(_0042_),
    .DE(_0014_),
    .Q(\mem[1][4] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][5]$_DFFE_PP_  (.D(_0043_),
    .DE(_0014_),
    .Q(\mem[1][5] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][6]$_DFFE_PP_  (.D(_0044_),
    .DE(_0014_),
    .Q(\mem[1][6] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][7]$_DFFE_PP_  (.D(_0045_),
    .DE(_0014_),
    .Q(\mem[1][7] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][8]$_DFFE_PP_  (.D(_0046_),
    .DE(_0014_),
    .Q(\mem[1][8] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][9]$_DFFE_PP_  (.D(_0047_),
    .DE(_0014_),
    .Q(\mem[1][9] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][0]$_DFFE_PP_  (.D(_0016_),
    .DE(_0013_),
    .Q(\mem[2][0] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][10]$_DFFE_PP_  (.D(_0017_),
    .DE(_0013_),
    .Q(\mem[2][10] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][11]$_DFFE_PP_  (.D(_0018_),
    .DE(_0013_),
    .Q(\mem[2][11] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][12]$_DFFE_PP_  (.D(_0019_),
    .DE(_0013_),
    .Q(\mem[2][12] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][13]$_DFFE_PP_  (.D(_0020_),
    .DE(_0013_),
    .Q(\mem[2][13] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][14]$_DFFE_PP_  (.D(_0021_),
    .DE(_0013_),
    .Q(\mem[2][14] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][15]$_DFFE_PP_  (.D(_0022_),
    .DE(_0013_),
    .Q(\mem[2][15] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][16]$_DFFE_PP_  (.D(_0023_),
    .DE(_0013_),
    .Q(\mem[2][16] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][17]$_DFFE_PP_  (.D(_0024_),
    .DE(_0013_),
    .Q(\mem[2][17] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][18]$_DFFE_PP_  (.D(_0025_),
    .DE(_0013_),
    .Q(\mem[2][18] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][19]$_DFFE_PP_  (.D(_0026_),
    .DE(_0013_),
    .Q(\mem[2][19] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][1]$_DFFE_PP_  (.D(_0027_),
    .DE(_0013_),
    .Q(\mem[2][1] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][20]$_DFFE_PP_  (.D(_0028_),
    .DE(_0013_),
    .Q(\mem[2][20] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][21]$_DFFE_PP_  (.D(_0029_),
    .DE(_0013_),
    .Q(\mem[2][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][22]$_DFFE_PP_  (.D(_0030_),
    .DE(_0013_),
    .Q(\mem[2][22] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][23]$_DFFE_PP_  (.D(_0031_),
    .DE(_0013_),
    .Q(\mem[2][23] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][24]$_DFFE_PP_  (.D(_0032_),
    .DE(_0013_),
    .Q(\mem[2][24] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][25]$_DFFE_PP_  (.D(_0033_),
    .DE(_0013_),
    .Q(\mem[2][25] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][26]$_DFFE_PP_  (.D(_0034_),
    .DE(_0013_),
    .Q(\mem[2][26] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][27]$_DFFE_PP_  (.D(_0035_),
    .DE(_0013_),
    .Q(\mem[2][27] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][28]$_DFFE_PP_  (.D(_0036_),
    .DE(_0013_),
    .Q(\mem[2][28] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][29]$_DFFE_PP_  (.D(_0037_),
    .DE(_0013_),
    .Q(\mem[2][29] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][2]$_DFFE_PP_  (.D(_0038_),
    .DE(_0013_),
    .Q(\mem[2][2] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][30]$_DFFE_PP_  (.D(_0039_),
    .DE(_0013_),
    .Q(\mem[2][30] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][31]$_DFFE_PP_  (.D(_0040_),
    .DE(_0013_),
    .Q(\mem[2][31] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][3]$_DFFE_PP_  (.D(_0041_),
    .DE(_0013_),
    .Q(\mem[2][3] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][4]$_DFFE_PP_  (.D(_0042_),
    .DE(_0013_),
    .Q(\mem[2][4] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][5]$_DFFE_PP_  (.D(_0043_),
    .DE(_0013_),
    .Q(\mem[2][5] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][6]$_DFFE_PP_  (.D(_0044_),
    .DE(_0013_),
    .Q(\mem[2][6] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][7]$_DFFE_PP_  (.D(_0045_),
    .DE(_0013_),
    .Q(\mem[2][7] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][8]$_DFFE_PP_  (.D(_0046_),
    .DE(_0013_),
    .Q(\mem[2][8] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][9]$_DFFE_PP_  (.D(_0047_),
    .DE(_0013_),
    .Q(\mem[2][9] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][0]$_DFFE_PP_  (.D(_0016_),
    .DE(_0012_),
    .Q(\mem[3][0] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][10]$_DFFE_PP_  (.D(_0017_),
    .DE(_0012_),
    .Q(\mem[3][10] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][11]$_DFFE_PP_  (.D(_0018_),
    .DE(_0012_),
    .Q(\mem[3][11] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][12]$_DFFE_PP_  (.D(_0019_),
    .DE(_0012_),
    .Q(\mem[3][12] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][13]$_DFFE_PP_  (.D(_0020_),
    .DE(_0012_),
    .Q(\mem[3][13] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][14]$_DFFE_PP_  (.D(_0021_),
    .DE(_0012_),
    .Q(\mem[3][14] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][15]$_DFFE_PP_  (.D(_0022_),
    .DE(_0012_),
    .Q(\mem[3][15] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][16]$_DFFE_PP_  (.D(_0023_),
    .DE(_0012_),
    .Q(\mem[3][16] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][17]$_DFFE_PP_  (.D(_0024_),
    .DE(_0012_),
    .Q(\mem[3][17] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][18]$_DFFE_PP_  (.D(_0025_),
    .DE(_0012_),
    .Q(\mem[3][18] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][19]$_DFFE_PP_  (.D(_0026_),
    .DE(_0012_),
    .Q(\mem[3][19] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][1]$_DFFE_PP_  (.D(_0027_),
    .DE(_0012_),
    .Q(\mem[3][1] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][20]$_DFFE_PP_  (.D(_0028_),
    .DE(_0012_),
    .Q(\mem[3][20] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][21]$_DFFE_PP_  (.D(_0029_),
    .DE(_0012_),
    .Q(\mem[3][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][22]$_DFFE_PP_  (.D(_0030_),
    .DE(_0012_),
    .Q(\mem[3][22] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][23]$_DFFE_PP_  (.D(_0031_),
    .DE(_0012_),
    .Q(\mem[3][23] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][24]$_DFFE_PP_  (.D(_0032_),
    .DE(_0012_),
    .Q(\mem[3][24] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][25]$_DFFE_PP_  (.D(_0033_),
    .DE(_0012_),
    .Q(\mem[3][25] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][26]$_DFFE_PP_  (.D(_0034_),
    .DE(_0012_),
    .Q(\mem[3][26] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][27]$_DFFE_PP_  (.D(_0035_),
    .DE(_0012_),
    .Q(\mem[3][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][28]$_DFFE_PP_  (.D(_0036_),
    .DE(_0012_),
    .Q(\mem[3][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][29]$_DFFE_PP_  (.D(_0037_),
    .DE(_0012_),
    .Q(\mem[3][29] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][2]$_DFFE_PP_  (.D(_0038_),
    .DE(_0012_),
    .Q(\mem[3][2] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][30]$_DFFE_PP_  (.D(_0039_),
    .DE(_0012_),
    .Q(\mem[3][30] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][31]$_DFFE_PP_  (.D(_0040_),
    .DE(_0012_),
    .Q(\mem[3][31] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][3]$_DFFE_PP_  (.D(_0041_),
    .DE(_0012_),
    .Q(\mem[3][3] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][4]$_DFFE_PP_  (.D(_0042_),
    .DE(_0012_),
    .Q(\mem[3][4] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][5]$_DFFE_PP_  (.D(_0043_),
    .DE(_0012_),
    .Q(\mem[3][5] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][6]$_DFFE_PP_  (.D(_0044_),
    .DE(_0012_),
    .Q(\mem[3][6] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][7]$_DFFE_PP_  (.D(_0045_),
    .DE(_0012_),
    .Q(\mem[3][7] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][8]$_DFFE_PP_  (.D(_0046_),
    .DE(_0012_),
    .Q(\mem[3][8] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][9]$_DFFE_PP_  (.D(_0047_),
    .DE(_0012_),
    .Q(\mem[3][9] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][0]$_DFFE_PP_  (.D(_0016_),
    .DE(_0011_),
    .Q(\mem[4][0] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][10]$_DFFE_PP_  (.D(_0017_),
    .DE(_0011_),
    .Q(\mem[4][10] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][11]$_DFFE_PP_  (.D(_0018_),
    .DE(_0011_),
    .Q(\mem[4][11] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][12]$_DFFE_PP_  (.D(_0019_),
    .DE(_0011_),
    .Q(\mem[4][12] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][13]$_DFFE_PP_  (.D(_0020_),
    .DE(_0011_),
    .Q(\mem[4][13] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][14]$_DFFE_PP_  (.D(_0021_),
    .DE(_0011_),
    .Q(\mem[4][14] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][15]$_DFFE_PP_  (.D(_0022_),
    .DE(_0011_),
    .Q(\mem[4][15] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][16]$_DFFE_PP_  (.D(_0023_),
    .DE(_0011_),
    .Q(\mem[4][16] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][17]$_DFFE_PP_  (.D(_0024_),
    .DE(_0011_),
    .Q(\mem[4][17] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][18]$_DFFE_PP_  (.D(_0025_),
    .DE(_0011_),
    .Q(\mem[4][18] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][19]$_DFFE_PP_  (.D(_0026_),
    .DE(_0011_),
    .Q(\mem[4][19] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][1]$_DFFE_PP_  (.D(_0027_),
    .DE(_0011_),
    .Q(\mem[4][1] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][20]$_DFFE_PP_  (.D(_0028_),
    .DE(_0011_),
    .Q(\mem[4][20] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][21]$_DFFE_PP_  (.D(_0029_),
    .DE(_0011_),
    .Q(\mem[4][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][22]$_DFFE_PP_  (.D(_0030_),
    .DE(_0011_),
    .Q(\mem[4][22] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][23]$_DFFE_PP_  (.D(_0031_),
    .DE(_0011_),
    .Q(\mem[4][23] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][24]$_DFFE_PP_  (.D(_0032_),
    .DE(_0011_),
    .Q(\mem[4][24] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][25]$_DFFE_PP_  (.D(_0033_),
    .DE(_0011_),
    .Q(\mem[4][25] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][26]$_DFFE_PP_  (.D(_0034_),
    .DE(_0011_),
    .Q(\mem[4][26] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][27]$_DFFE_PP_  (.D(_0035_),
    .DE(_0011_),
    .Q(\mem[4][27] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][28]$_DFFE_PP_  (.D(_0036_),
    .DE(_0011_),
    .Q(\mem[4][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][29]$_DFFE_PP_  (.D(_0037_),
    .DE(_0011_),
    .Q(\mem[4][29] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][2]$_DFFE_PP_  (.D(_0038_),
    .DE(_0011_),
    .Q(\mem[4][2] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][30]$_DFFE_PP_  (.D(_0039_),
    .DE(_0011_),
    .Q(\mem[4][30] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][31]$_DFFE_PP_  (.D(_0040_),
    .DE(_0011_),
    .Q(\mem[4][31] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][3]$_DFFE_PP_  (.D(_0041_),
    .DE(_0011_),
    .Q(\mem[4][3] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][4]$_DFFE_PP_  (.D(_0042_),
    .DE(_0011_),
    .Q(\mem[4][4] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][5]$_DFFE_PP_  (.D(_0043_),
    .DE(_0011_),
    .Q(\mem[4][5] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][6]$_DFFE_PP_  (.D(_0044_),
    .DE(_0011_),
    .Q(\mem[4][6] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][7]$_DFFE_PP_  (.D(_0045_),
    .DE(_0011_),
    .Q(\mem[4][7] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][8]$_DFFE_PP_  (.D(_0046_),
    .DE(_0011_),
    .Q(\mem[4][8] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][9]$_DFFE_PP_  (.D(_0047_),
    .DE(_0011_),
    .Q(\mem[4][9] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][0]$_DFFE_PP_  (.D(_0016_),
    .DE(_0010_),
    .Q(\mem[5][0] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][10]$_DFFE_PP_  (.D(_0017_),
    .DE(_0010_),
    .Q(\mem[5][10] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][11]$_DFFE_PP_  (.D(_0018_),
    .DE(_0010_),
    .Q(\mem[5][11] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][12]$_DFFE_PP_  (.D(_0019_),
    .DE(_0010_),
    .Q(\mem[5][12] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][13]$_DFFE_PP_  (.D(_0020_),
    .DE(_0010_),
    .Q(\mem[5][13] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][14]$_DFFE_PP_  (.D(_0021_),
    .DE(_0010_),
    .Q(\mem[5][14] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][15]$_DFFE_PP_  (.D(_0022_),
    .DE(_0010_),
    .Q(\mem[5][15] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][16]$_DFFE_PP_  (.D(_0023_),
    .DE(_0010_),
    .Q(\mem[5][16] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][17]$_DFFE_PP_  (.D(_0024_),
    .DE(_0010_),
    .Q(\mem[5][17] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][18]$_DFFE_PP_  (.D(_0025_),
    .DE(_0010_),
    .Q(\mem[5][18] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][19]$_DFFE_PP_  (.D(_0026_),
    .DE(_0010_),
    .Q(\mem[5][19] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][1]$_DFFE_PP_  (.D(_0027_),
    .DE(_0010_),
    .Q(\mem[5][1] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][20]$_DFFE_PP_  (.D(_0028_),
    .DE(_0010_),
    .Q(\mem[5][20] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][21]$_DFFE_PP_  (.D(_0029_),
    .DE(_0010_),
    .Q(\mem[5][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][22]$_DFFE_PP_  (.D(_0030_),
    .DE(_0010_),
    .Q(\mem[5][22] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][23]$_DFFE_PP_  (.D(_0031_),
    .DE(_0010_),
    .Q(\mem[5][23] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][24]$_DFFE_PP_  (.D(_0032_),
    .DE(_0010_),
    .Q(\mem[5][24] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][25]$_DFFE_PP_  (.D(_0033_),
    .DE(_0010_),
    .Q(\mem[5][25] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][26]$_DFFE_PP_  (.D(_0034_),
    .DE(_0010_),
    .Q(\mem[5][26] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][27]$_DFFE_PP_  (.D(_0035_),
    .DE(_0010_),
    .Q(\mem[5][27] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][28]$_DFFE_PP_  (.D(_0036_),
    .DE(_0010_),
    .Q(\mem[5][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][29]$_DFFE_PP_  (.D(_0037_),
    .DE(_0010_),
    .Q(\mem[5][29] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][2]$_DFFE_PP_  (.D(_0038_),
    .DE(_0010_),
    .Q(\mem[5][2] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][30]$_DFFE_PP_  (.D(_0039_),
    .DE(_0010_),
    .Q(\mem[5][30] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][31]$_DFFE_PP_  (.D(_0040_),
    .DE(_0010_),
    .Q(\mem[5][31] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][3]$_DFFE_PP_  (.D(_0041_),
    .DE(_0010_),
    .Q(\mem[5][3] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][4]$_DFFE_PP_  (.D(_0042_),
    .DE(_0010_),
    .Q(\mem[5][4] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][5]$_DFFE_PP_  (.D(_0043_),
    .DE(_0010_),
    .Q(\mem[5][5] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][6]$_DFFE_PP_  (.D(_0044_),
    .DE(_0010_),
    .Q(\mem[5][6] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][7]$_DFFE_PP_  (.D(_0045_),
    .DE(_0010_),
    .Q(\mem[5][7] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][8]$_DFFE_PP_  (.D(_0046_),
    .DE(_0010_),
    .Q(\mem[5][8] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][9]$_DFFE_PP_  (.D(_0047_),
    .DE(_0010_),
    .Q(\mem[5][9] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][0]$_DFFE_PP_  (.D(_0016_),
    .DE(_0009_),
    .Q(\mem[6][0] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][10]$_DFFE_PP_  (.D(_0017_),
    .DE(_0009_),
    .Q(\mem[6][10] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][11]$_DFFE_PP_  (.D(_0018_),
    .DE(_0009_),
    .Q(\mem[6][11] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][12]$_DFFE_PP_  (.D(_0019_),
    .DE(_0009_),
    .Q(\mem[6][12] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][13]$_DFFE_PP_  (.D(_0020_),
    .DE(_0009_),
    .Q(\mem[6][13] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][14]$_DFFE_PP_  (.D(_0021_),
    .DE(_0009_),
    .Q(\mem[6][14] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][15]$_DFFE_PP_  (.D(_0022_),
    .DE(_0009_),
    .Q(\mem[6][15] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][16]$_DFFE_PP_  (.D(_0023_),
    .DE(_0009_),
    .Q(\mem[6][16] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][17]$_DFFE_PP_  (.D(_0024_),
    .DE(_0009_),
    .Q(\mem[6][17] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][18]$_DFFE_PP_  (.D(_0025_),
    .DE(_0009_),
    .Q(\mem[6][18] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][19]$_DFFE_PP_  (.D(_0026_),
    .DE(_0009_),
    .Q(\mem[6][19] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][1]$_DFFE_PP_  (.D(_0027_),
    .DE(_0009_),
    .Q(\mem[6][1] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][20]$_DFFE_PP_  (.D(_0028_),
    .DE(_0009_),
    .Q(\mem[6][20] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][21]$_DFFE_PP_  (.D(_0029_),
    .DE(_0009_),
    .Q(\mem[6][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][22]$_DFFE_PP_  (.D(_0030_),
    .DE(_0009_),
    .Q(\mem[6][22] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][23]$_DFFE_PP_  (.D(_0031_),
    .DE(_0009_),
    .Q(\mem[6][23] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][24]$_DFFE_PP_  (.D(_0032_),
    .DE(_0009_),
    .Q(\mem[6][24] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][25]$_DFFE_PP_  (.D(_0033_),
    .DE(_0009_),
    .Q(\mem[6][25] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][26]$_DFFE_PP_  (.D(_0034_),
    .DE(_0009_),
    .Q(\mem[6][26] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][27]$_DFFE_PP_  (.D(_0035_),
    .DE(_0009_),
    .Q(\mem[6][27] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][28]$_DFFE_PP_  (.D(_0036_),
    .DE(_0009_),
    .Q(\mem[6][28] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][29]$_DFFE_PP_  (.D(_0037_),
    .DE(_0009_),
    .Q(\mem[6][29] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][2]$_DFFE_PP_  (.D(_0038_),
    .DE(_0009_),
    .Q(\mem[6][2] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][30]$_DFFE_PP_  (.D(_0039_),
    .DE(_0009_),
    .Q(\mem[6][30] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][31]$_DFFE_PP_  (.D(_0040_),
    .DE(_0009_),
    .Q(\mem[6][31] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][3]$_DFFE_PP_  (.D(_0041_),
    .DE(_0009_),
    .Q(\mem[6][3] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][4]$_DFFE_PP_  (.D(_0042_),
    .DE(_0009_),
    .Q(\mem[6][4] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][5]$_DFFE_PP_  (.D(_0043_),
    .DE(_0009_),
    .Q(\mem[6][5] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][6]$_DFFE_PP_  (.D(_0044_),
    .DE(_0009_),
    .Q(\mem[6][6] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][7]$_DFFE_PP_  (.D(_0045_),
    .DE(_0009_),
    .Q(\mem[6][7] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][8]$_DFFE_PP_  (.D(_0046_),
    .DE(_0009_),
    .Q(\mem[6][8] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][9]$_DFFE_PP_  (.D(_0047_),
    .DE(_0009_),
    .Q(\mem[6][9] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][0]$_DFFE_PP_  (.D(_0016_),
    .DE(_0008_),
    .Q(\mem[7][0] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][10]$_DFFE_PP_  (.D(_0017_),
    .DE(_0008_),
    .Q(\mem[7][10] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][11]$_DFFE_PP_  (.D(_0018_),
    .DE(_0008_),
    .Q(\mem[7][11] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][12]$_DFFE_PP_  (.D(_0019_),
    .DE(_0008_),
    .Q(\mem[7][12] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][13]$_DFFE_PP_  (.D(_0020_),
    .DE(_0008_),
    .Q(\mem[7][13] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][14]$_DFFE_PP_  (.D(_0021_),
    .DE(_0008_),
    .Q(\mem[7][14] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][15]$_DFFE_PP_  (.D(_0022_),
    .DE(_0008_),
    .Q(\mem[7][15] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][16]$_DFFE_PP_  (.D(_0023_),
    .DE(_0008_),
    .Q(\mem[7][16] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][17]$_DFFE_PP_  (.D(_0024_),
    .DE(_0008_),
    .Q(\mem[7][17] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][18]$_DFFE_PP_  (.D(_0025_),
    .DE(_0008_),
    .Q(\mem[7][18] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][19]$_DFFE_PP_  (.D(_0026_),
    .DE(_0008_),
    .Q(\mem[7][19] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][1]$_DFFE_PP_  (.D(_0027_),
    .DE(_0008_),
    .Q(\mem[7][1] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][20]$_DFFE_PP_  (.D(_0028_),
    .DE(_0008_),
    .Q(\mem[7][20] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][21]$_DFFE_PP_  (.D(_0029_),
    .DE(_0008_),
    .Q(\mem[7][21] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][22]$_DFFE_PP_  (.D(_0030_),
    .DE(_0008_),
    .Q(\mem[7][22] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][23]$_DFFE_PP_  (.D(_0031_),
    .DE(_0008_),
    .Q(\mem[7][23] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][24]$_DFFE_PP_  (.D(_0032_),
    .DE(_0008_),
    .Q(\mem[7][24] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][25]$_DFFE_PP_  (.D(_0033_),
    .DE(_0008_),
    .Q(\mem[7][25] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][26]$_DFFE_PP_  (.D(_0034_),
    .DE(_0008_),
    .Q(\mem[7][26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][27]$_DFFE_PP_  (.D(_0035_),
    .DE(_0008_),
    .Q(\mem[7][27] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][28]$_DFFE_PP_  (.D(_0036_),
    .DE(_0008_),
    .Q(\mem[7][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][29]$_DFFE_PP_  (.D(_0037_),
    .DE(_0008_),
    .Q(\mem[7][29] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][2]$_DFFE_PP_  (.D(_0038_),
    .DE(_0008_),
    .Q(\mem[7][2] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][30]$_DFFE_PP_  (.D(_0039_),
    .DE(_0008_),
    .Q(\mem[7][30] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][31]$_DFFE_PP_  (.D(_0040_),
    .DE(_0008_),
    .Q(\mem[7][31] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][3]$_DFFE_PP_  (.D(_0041_),
    .DE(_0008_),
    .Q(\mem[7][3] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][4]$_DFFE_PP_  (.D(_0042_),
    .DE(_0008_),
    .Q(\mem[7][4] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][5]$_DFFE_PP_  (.D(_0043_),
    .DE(_0008_),
    .Q(\mem[7][5] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][6]$_DFFE_PP_  (.D(_0044_),
    .DE(_0008_),
    .Q(\mem[7][6] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][7]$_DFFE_PP_  (.D(_0045_),
    .DE(_0008_),
    .Q(\mem[7][7] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][8]$_DFFE_PP_  (.D(_0046_),
    .DE(_0008_),
    .Q(\mem[7][8] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][9]$_DFFE_PP_  (.D(_0047_),
    .DE(_0008_),
    .Q(\mem[7][9] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][0]$_DFFE_PP_  (.D(_0016_),
    .DE(_0007_),
    .Q(\mem[8][0] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][10]$_DFFE_PP_  (.D(_0017_),
    .DE(net163),
    .Q(\mem[8][10] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][11]$_DFFE_PP_  (.D(_0018_),
    .DE(net162),
    .Q(\mem[8][11] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][12]$_DFFE_PP_  (.D(_0019_),
    .DE(net163),
    .Q(\mem[8][12] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][13]$_DFFE_PP_  (.D(_0020_),
    .DE(net162),
    .Q(\mem[8][13] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][14]$_DFFE_PP_  (.D(_0021_),
    .DE(net162),
    .Q(\mem[8][14] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][15]$_DFFE_PP_  (.D(_0022_),
    .DE(net163),
    .Q(\mem[8][15] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][16]$_DFFE_PP_  (.D(_0023_),
    .DE(net164),
    .Q(\mem[8][16] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][17]$_DFFE_PP_  (.D(_0024_),
    .DE(net162),
    .Q(\mem[8][17] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][18]$_DFFE_PP_  (.D(_0025_),
    .DE(net164),
    .Q(\mem[8][18] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][19]$_DFFE_PP_  (.D(_0026_),
    .DE(net163),
    .Q(\mem[8][19] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][1]$_DFFE_PP_  (.D(_0027_),
    .DE(net164),
    .Q(\mem[8][1] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][20]$_DFFE_PP_  (.D(_0028_),
    .DE(net164),
    .Q(\mem[8][20] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][21]$_DFFE_PP_  (.D(_0029_),
    .DE(_0007_),
    .Q(\mem[8][21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][22]$_DFFE_PP_  (.D(_0030_),
    .DE(net164),
    .Q(\mem[8][22] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][23]$_DFFE_PP_  (.D(_0031_),
    .DE(net164),
    .Q(\mem[8][23] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][24]$_DFFE_PP_  (.D(_0032_),
    .DE(net164),
    .Q(\mem[8][24] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][25]$_DFFE_PP_  (.D(_0033_),
    .DE(net162),
    .Q(\mem[8][25] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][26]$_DFFE_PP_  (.D(_0034_),
    .DE(net162),
    .Q(\mem[8][26] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][27]$_DFFE_PP_  (.D(_0035_),
    .DE(net163),
    .Q(\mem[8][27] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][28]$_DFFE_PP_  (.D(_0036_),
    .DE(net162),
    .Q(\mem[8][28] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][29]$_DFFE_PP_  (.D(_0037_),
    .DE(net163),
    .Q(\mem[8][29] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][2]$_DFFE_PP_  (.D(_0038_),
    .DE(net162),
    .Q(\mem[8][2] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][30]$_DFFE_PP_  (.D(_0039_),
    .DE(net164),
    .Q(\mem[8][30] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][31]$_DFFE_PP_  (.D(_0040_),
    .DE(net164),
    .Q(\mem[8][31] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][3]$_DFFE_PP_  (.D(_0041_),
    .DE(net164),
    .Q(\mem[8][3] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][4]$_DFFE_PP_  (.D(_0042_),
    .DE(net164),
    .Q(\mem[8][4] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][5]$_DFFE_PP_  (.D(_0043_),
    .DE(net163),
    .Q(\mem[8][5] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][6]$_DFFE_PP_  (.D(_0044_),
    .DE(net163),
    .Q(\mem[8][6] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][7]$_DFFE_PP_  (.D(_0045_),
    .DE(_0007_),
    .Q(\mem[8][7] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][8]$_DFFE_PP_  (.D(_0046_),
    .DE(net163),
    .Q(\mem[8][8] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][9]$_DFFE_PP_  (.D(_0047_),
    .DE(net162),
    .Q(\mem[8][9] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][0]$_DFFE_PP_  (.D(_0016_),
    .DE(_0006_),
    .Q(\mem[9][0] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][10]$_DFFE_PP_  (.D(_0017_),
    .DE(net151),
    .Q(\mem[9][10] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][11]$_DFFE_PP_  (.D(_0018_),
    .DE(net151),
    .Q(\mem[9][11] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][12]$_DFFE_PP_  (.D(_0019_),
    .DE(net151),
    .Q(\mem[9][12] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][13]$_DFFE_PP_  (.D(_0020_),
    .DE(net150),
    .Q(\mem[9][13] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][14]$_DFFE_PP_  (.D(_0021_),
    .DE(_0006_),
    .Q(\mem[9][14] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][15]$_DFFE_PP_  (.D(_0022_),
    .DE(net151),
    .Q(\mem[9][15] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][16]$_DFFE_PP_  (.D(_0023_),
    .DE(net150),
    .Q(\mem[9][16] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][17]$_DFFE_PP_  (.D(_0024_),
    .DE(net151),
    .Q(\mem[9][17] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][18]$_DFFE_PP_  (.D(_0025_),
    .DE(net152),
    .Q(\mem[9][18] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][19]$_DFFE_PP_  (.D(_0026_),
    .DE(net151),
    .Q(\mem[9][19] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][1]$_DFFE_PP_  (.D(_0027_),
    .DE(net150),
    .Q(\mem[9][1] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][20]$_DFFE_PP_  (.D(_0028_),
    .DE(_0006_),
    .Q(\mem[9][20] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][21]$_DFFE_PP_  (.D(_0029_),
    .DE(net150),
    .Q(\mem[9][21] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][22]$_DFFE_PP_  (.D(_0030_),
    .DE(net150),
    .Q(\mem[9][22] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][23]$_DFFE_PP_  (.D(_0031_),
    .DE(net150),
    .Q(\mem[9][23] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][24]$_DFFE_PP_  (.D(_0032_),
    .DE(net150),
    .Q(\mem[9][24] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][25]$_DFFE_PP_  (.D(_0033_),
    .DE(net152),
    .Q(\mem[9][25] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][26]$_DFFE_PP_  (.D(_0034_),
    .DE(net152),
    .Q(\mem[9][26] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][27]$_DFFE_PP_  (.D(_0035_),
    .DE(net151),
    .Q(\mem[9][27] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][28]$_DFFE_PP_  (.D(_0036_),
    .DE(net152),
    .Q(\mem[9][28] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][29]$_DFFE_PP_  (.D(_0037_),
    .DE(_0006_),
    .Q(\mem[9][29] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][2]$_DFFE_PP_  (.D(_0038_),
    .DE(_0006_),
    .Q(\mem[9][2] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][30]$_DFFE_PP_  (.D(_0039_),
    .DE(net150),
    .Q(\mem[9][30] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][31]$_DFFE_PP_  (.D(_0040_),
    .DE(_0006_),
    .Q(\mem[9][31] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][3]$_DFFE_PP_  (.D(_0041_),
    .DE(net150),
    .Q(\mem[9][3] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][4]$_DFFE_PP_  (.D(_0042_),
    .DE(net150),
    .Q(\mem[9][4] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][5]$_DFFE_PP_  (.D(_0043_),
    .DE(net152),
    .Q(\mem[9][5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][6]$_DFFE_PP_  (.D(_0044_),
    .DE(net151),
    .Q(\mem[9][6] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][7]$_DFFE_PP_  (.D(_0045_),
    .DE(net150),
    .Q(\mem[9][7] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][8]$_DFFE_PP_  (.D(_0046_),
    .DE(net151),
    .Q(\mem[9][8] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][9]$_DFFE_PP_  (.D(_0047_),
    .DE(net151),
    .Q(\mem[9][9] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[0]$_DFFE_PN0P_  (.D(_0080_),
    .Q(net108),
    .RESET_B(net1),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[10]$_DFFE_PN0P_  (.D(_0081_),
    .Q(net109),
    .RESET_B(net1),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[11]$_DFFE_PN0P_  (.D(_0082_),
    .Q(net110),
    .RESET_B(net1),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[12]$_DFFE_PN0P_  (.D(_0083_),
    .Q(net111),
    .RESET_B(net1),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[13]$_DFFE_PN0P_  (.D(_0084_),
    .Q(net112),
    .RESET_B(net1),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[14]$_DFFE_PN0P_  (.D(_0085_),
    .Q(net113),
    .RESET_B(net1),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[15]$_DFFE_PN0P_  (.D(_0086_),
    .Q(net114),
    .RESET_B(net1),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[16]$_DFFE_PN0P_  (.D(_0087_),
    .Q(net115),
    .RESET_B(net1),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[17]$_DFFE_PN0P_  (.D(_0088_),
    .Q(net116),
    .RESET_B(net1),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[18]$_DFFE_PN0P_  (.D(_0089_),
    .Q(net117),
    .RESET_B(net1),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[19]$_DFFE_PN0P_  (.D(_0090_),
    .Q(net118),
    .RESET_B(net1),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[1]$_DFFE_PN0P_  (.D(_0091_),
    .Q(net119),
    .RESET_B(net1),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[20]$_DFFE_PN0P_  (.D(_0092_),
    .Q(net120),
    .RESET_B(net1),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[21]$_DFFE_PN0P_  (.D(_0093_),
    .Q(net121),
    .RESET_B(net1),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[22]$_DFFE_PN0P_  (.D(_0094_),
    .Q(net122),
    .RESET_B(net1),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[23]$_DFFE_PN0P_  (.D(_0095_),
    .Q(net123),
    .RESET_B(net1),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[24]$_DFFE_PN0P_  (.D(_0096_),
    .Q(net124),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[25]$_DFFE_PN0P_  (.D(_0097_),
    .Q(net125),
    .RESET_B(net1),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[26]$_DFFE_PN0P_  (.D(_0098_),
    .Q(net126),
    .RESET_B(net1),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[27]$_DFFE_PN0P_  (.D(_0099_),
    .Q(net127),
    .RESET_B(net1),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[28]$_DFFE_PN0P_  (.D(_0100_),
    .Q(net128),
    .RESET_B(net1),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[29]$_DFFE_PN0P_  (.D(_0101_),
    .Q(net129),
    .RESET_B(net1),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[2]$_DFFE_PN0P_  (.D(_0102_),
    .Q(net130),
    .RESET_B(net1),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[30]$_DFFE_PN0P_  (.D(_0103_),
    .Q(net131),
    .RESET_B(net1),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[31]$_DFFE_PN0P_  (.D(_0104_),
    .Q(net132),
    .RESET_B(net1),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[3]$_DFFE_PN0P_  (.D(_0105_),
    .Q(net133),
    .RESET_B(net1),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[4]$_DFFE_PN0P_  (.D(_0106_),
    .Q(net134),
    .RESET_B(net1),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[5]$_DFFE_PN0P_  (.D(_0107_),
    .Q(net135),
    .RESET_B(net1),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[6]$_DFFE_PN0P_  (.D(_0108_),
    .Q(net136),
    .RESET_B(net1),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[7]$_DFFE_PN0P_  (.D(_0109_),
    .Q(net137),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[8]$_DFFE_PN0P_  (.D(_0110_),
    .Q(net138),
    .RESET_B(net1),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_rdata[9]$_DFFE_PN0P_  (.D(_0111_),
    .Q(net139),
    .RESET_B(net1),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfrtp_1 \mem_ready$_DFF_PN0_  (.D(net39),
    .Q(net140),
    .RESET_B(net1),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_2 \rd_ptr[0]$_DFFE_PN0P_  (.D(_0112_),
    .Q(\rd_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_2 \rd_ptr[1]$_DFFE_PN0P_  (.D(_0113_),
    .Q(\rd_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_2 \rd_ptr[2]$_DFFE_PN0P_  (.D(_0114_),
    .Q(\rd_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[3]$_DFFE_PN0P_  (.D(_0115_),
    .Q(\rd_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr[4]$_DFFE_PN0P_  (.D(_0116_),
    .Q(\rd_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[0]$_DFFE_PN0P_  (.D(_0117_),
    .Q(\wr_ptr[0] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_4 \wr_ptr[1]$_DFFE_PN0P_  (.D(_0118_),
    .Q(\wr_ptr[1] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfrtp_4 \wr_ptr[2]$_DFFE_PN0P_  (.D(_0119_),
    .Q(\wr_ptr[2] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[3]$_DFFE_PN0P_  (.D(_0120_),
    .Q(\wr_ptr[3] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr[4]$_DFFE_PN0P_  (.D(_0121_),
    .Q(\wr_ptr[4] ),
    .RESET_B(net1),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__buf_16 hold1 (.A(net73),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_538 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(ext_rd_en),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(ext_wr_data[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ext_wr_data[10]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(ext_wr_data[11]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ext_wr_data[12]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(ext_wr_data[13]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(ext_wr_data[14]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(ext_wr_data[15]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(ext_wr_data[16]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(ext_wr_data[17]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(ext_wr_data[18]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(ext_wr_data[19]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(ext_wr_data[1]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(ext_wr_data[20]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(ext_wr_data[21]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(ext_wr_data[22]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(ext_wr_data[23]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(ext_wr_data[24]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(ext_wr_data[25]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(ext_wr_data[26]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(ext_wr_data[27]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(ext_wr_data[28]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(ext_wr_data[29]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(ext_wr_data[2]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(ext_wr_data[30]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(ext_wr_data[31]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(ext_wr_data[3]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(ext_wr_data[4]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(ext_wr_data[5]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(ext_wr_data[6]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(ext_wr_data[7]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(ext_wr_data[8]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(ext_wr_data[9]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(ext_wr_en),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(mem_addr[0]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(mem_addr[1]),
    .X(net37));
 sky130_fd_sc_hd__dlymetal6s2s_1 input37 (.A(mem_addr[2]),
    .X(net38));
 sky130_fd_sc_hd__dlymetal6s2s_1 input38 (.A(net166),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(mem_wdata[0]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(mem_wdata[10]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(mem_wdata[11]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(mem_wdata[12]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(mem_wdata[13]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(mem_wdata[14]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(mem_wdata[15]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(mem_wdata[16]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(mem_wdata[17]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(mem_wdata[18]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(mem_wdata[19]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(mem_wdata[1]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(mem_wdata[20]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(mem_wdata[21]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(mem_wdata[22]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(mem_wdata[23]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(mem_wdata[24]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(mem_wdata[25]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(mem_wdata[26]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(mem_wdata[27]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(mem_wdata[28]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(mem_wdata[29]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(mem_wdata[2]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(mem_wdata[30]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(mem_wdata[31]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(mem_wdata[3]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(mem_wdata[4]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(mem_wdata[5]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(mem_wdata[6]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(mem_wdata[7]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(mem_wdata[8]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(mem_wdata[9]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 input71 (.A(mem_write),
    .X(net72));
 sky130_fd_sc_hd__buf_2 input72 (.A(net165),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net74),
    .X(ext_empty));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net75),
    .X(ext_full));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net76),
    .X(ext_rd_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net77),
    .X(ext_rd_data[10]));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net78),
    .X(ext_rd_data[11]));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net79),
    .X(ext_rd_data[12]));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net80),
    .X(ext_rd_data[13]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net81),
    .X(ext_rd_data[14]));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net82),
    .X(ext_rd_data[15]));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net83),
    .X(ext_rd_data[16]));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net84),
    .X(ext_rd_data[17]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net85),
    .X(ext_rd_data[18]));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(net86),
    .X(ext_rd_data[19]));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(net87),
    .X(ext_rd_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(net88),
    .X(ext_rd_data[20]));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(net89),
    .X(ext_rd_data[21]));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net90),
    .X(ext_rd_data[22]));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(net91),
    .X(ext_rd_data[23]));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(net92),
    .X(ext_rd_data[24]));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(net93),
    .X(ext_rd_data[25]));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(net94),
    .X(ext_rd_data[26]));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net95),
    .X(ext_rd_data[27]));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(net96),
    .X(ext_rd_data[28]));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(net97),
    .X(ext_rd_data[29]));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(net98),
    .X(ext_rd_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(net99),
    .X(ext_rd_data[30]));
 sky130_fd_sc_hd__clkbuf_1 output99 (.A(net100),
    .X(ext_rd_data[31]));
 sky130_fd_sc_hd__clkbuf_1 output100 (.A(net101),
    .X(ext_rd_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(net102),
    .X(ext_rd_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net103),
    .X(ext_rd_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(net104),
    .X(ext_rd_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output104 (.A(net105),
    .X(ext_rd_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output105 (.A(net106),
    .X(ext_rd_data[8]));
 sky130_fd_sc_hd__clkbuf_1 output106 (.A(net107),
    .X(ext_rd_data[9]));
 sky130_fd_sc_hd__clkbuf_1 output107 (.A(net108),
    .X(mem_rdata[0]));
 sky130_fd_sc_hd__clkbuf_1 output108 (.A(net109),
    .X(mem_rdata[10]));
 sky130_fd_sc_hd__clkbuf_1 output109 (.A(net110),
    .X(mem_rdata[11]));
 sky130_fd_sc_hd__clkbuf_1 output110 (.A(net111),
    .X(mem_rdata[12]));
 sky130_fd_sc_hd__clkbuf_1 output111 (.A(net112),
    .X(mem_rdata[13]));
 sky130_fd_sc_hd__clkbuf_1 output112 (.A(net113),
    .X(mem_rdata[14]));
 sky130_fd_sc_hd__clkbuf_1 output113 (.A(net114),
    .X(mem_rdata[15]));
 sky130_fd_sc_hd__clkbuf_1 output114 (.A(net115),
    .X(mem_rdata[16]));
 sky130_fd_sc_hd__clkbuf_1 output115 (.A(net116),
    .X(mem_rdata[17]));
 sky130_fd_sc_hd__clkbuf_1 output116 (.A(net117),
    .X(mem_rdata[18]));
 sky130_fd_sc_hd__clkbuf_1 output117 (.A(net118),
    .X(mem_rdata[19]));
 sky130_fd_sc_hd__clkbuf_1 output118 (.A(net119),
    .X(mem_rdata[1]));
 sky130_fd_sc_hd__clkbuf_1 output119 (.A(net120),
    .X(mem_rdata[20]));
 sky130_fd_sc_hd__clkbuf_1 output120 (.A(net121),
    .X(mem_rdata[21]));
 sky130_fd_sc_hd__clkbuf_1 output121 (.A(net122),
    .X(mem_rdata[22]));
 sky130_fd_sc_hd__clkbuf_1 output122 (.A(net123),
    .X(mem_rdata[23]));
 sky130_fd_sc_hd__clkbuf_1 output123 (.A(net124),
    .X(mem_rdata[24]));
 sky130_fd_sc_hd__clkbuf_1 output124 (.A(net125),
    .X(mem_rdata[25]));
 sky130_fd_sc_hd__clkbuf_1 output125 (.A(net126),
    .X(mem_rdata[26]));
 sky130_fd_sc_hd__clkbuf_1 output126 (.A(net127),
    .X(mem_rdata[27]));
 sky130_fd_sc_hd__clkbuf_1 output127 (.A(net128),
    .X(mem_rdata[28]));
 sky130_fd_sc_hd__clkbuf_1 output128 (.A(net129),
    .X(mem_rdata[29]));
 sky130_fd_sc_hd__clkbuf_1 output129 (.A(net130),
    .X(mem_rdata[2]));
 sky130_fd_sc_hd__clkbuf_1 output130 (.A(net131),
    .X(mem_rdata[30]));
 sky130_fd_sc_hd__clkbuf_1 output131 (.A(net132),
    .X(mem_rdata[31]));
 sky130_fd_sc_hd__clkbuf_1 output132 (.A(net133),
    .X(mem_rdata[3]));
 sky130_fd_sc_hd__clkbuf_1 output133 (.A(net134),
    .X(mem_rdata[4]));
 sky130_fd_sc_hd__clkbuf_1 output134 (.A(net135),
    .X(mem_rdata[5]));
 sky130_fd_sc_hd__clkbuf_1 output135 (.A(net136),
    .X(mem_rdata[6]));
 sky130_fd_sc_hd__clkbuf_1 output136 (.A(net137),
    .X(mem_rdata[7]));
 sky130_fd_sc_hd__clkbuf_1 output137 (.A(net138),
    .X(mem_rdata[8]));
 sky130_fd_sc_hd__clkbuf_1 output138 (.A(net139),
    .X(mem_rdata[9]));
 sky130_fd_sc_hd__clkbuf_1 output139 (.A(net140),
    .X(mem_ready));
 sky130_fd_sc_hd__buf_6 load_slew140 (.A(net142),
    .X(net141));
 sky130_fd_sc_hd__buf_6 load_slew141 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__buf_6 wire142 (.A(_0001_),
    .X(net143));
 sky130_fd_sc_hd__buf_6 load_slew143 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__buf_8 load_slew144 (.A(_0000_),
    .X(net145));
 sky130_fd_sc_hd__buf_16 max_cap145 (.A(_0000_),
    .X(net146));
 sky130_fd_sc_hd__buf_6 wire146 (.A(_0002_),
    .X(net147));
 sky130_fd_sc_hd__buf_6 load_slew147 (.A(_0002_),
    .X(net148));
 sky130_fd_sc_hd__buf_8 load_slew148 (.A(_0002_),
    .X(net149));
 sky130_fd_sc_hd__buf_6 wire149 (.A(_0006_),
    .X(net150));
 sky130_fd_sc_hd__buf_6 load_slew150 (.A(_0006_),
    .X(net151));
 sky130_fd_sc_hd__buf_6 load_slew151 (.A(_0006_),
    .X(net152));
 sky130_fd_sc_hd__buf_6 load_slew152 (.A(_0005_),
    .X(net153));
 sky130_fd_sc_hd__buf_8 max_cap153 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__buf_8 max_cap154 (.A(_0005_),
    .X(net155));
 sky130_fd_sc_hd__buf_8 max_cap155 (.A(net158),
    .X(net156));
 sky130_fd_sc_hd__buf_6 wire156 (.A(_0004_),
    .X(net157));
 sky130_fd_sc_hd__buf_8 load_slew157 (.A(_0004_),
    .X(net158));
 sky130_fd_sc_hd__buf_16 max_cap158 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__buf_6 wire159 (.A(_0003_),
    .X(net160));
 sky130_fd_sc_hd__buf_8 load_slew160 (.A(_0003_),
    .X(net161));
 sky130_fd_sc_hd__buf_8 max_cap161 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__buf_6 wire162 (.A(_0007_),
    .X(net163));
 sky130_fd_sc_hd__buf_6 wire163 (.A(_0007_),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_2_1__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_2_3__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_2_2__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_2_0__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload0 (.A(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload1 (.A(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkinv_1 clkload2 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload3 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload4 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkinv_1 clkload5 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload6 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkinv_1 clkload7 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkinv_2 clkload8 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkinv_1 clkload9 (.A(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkinv_2 clkload10 (.A(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkinv_1 clkload11 (.A(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkinv_1 clkload12 (.A(clknet_leaf_51_clk));
 sky130_fd_sc_hd__inv_6 clkload13 (.A(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload14 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload15 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkinv_1 clkload16 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkinv_1 clkload17 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkinv_2 clkload18 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload19 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload20 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload21 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkinv_1 clkload22 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkinv_2 clkload23 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload24 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload25 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload26 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload27 (.A(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload28 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkinv_1 clkload29 (.A(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkinv_1 clkload30 (.A(clknet_leaf_38_clk));
 sky130_fd_sc_hd__bufinv_16 clkload31 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload32 (.A(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload33 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload34 (.A(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload35 (.A(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload36 (.A(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload37 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload38 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload39 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload40 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload41 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload42 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload43 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload44 (.A(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload45 (.A(clknet_leaf_28_clk));
 sky130_fd_sc_hd__bufinv_16 clkload46 (.A(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload47 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload48 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(mem_valid),
    .X(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0133_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0181_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0320_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_0143_));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_242 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_374 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_420 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_21 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_387 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_417 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_354 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_444 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_314 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_5 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_64 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_87 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_372 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_22 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_372 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_362 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_30 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_390 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_353 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_445 ();
endmodule
