module parameterized_crc_generator (clk,
    crc_init,
    data_valid,
    rst_n,
    crc_out,
    data_in);
 input clk;
 input crc_init;
 input data_valid;
 input rst_n;
 output [7:0] crc_out;
 input [7:0] data_in;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire _34_;
 wire _35_;
 wire _36_;
 wire _37_;
 wire _38_;
 wire _39_;
 wire _40_;
 wire _41_;
 wire \crc_reflected[0] ;
 wire \crc_reflected[1] ;
 wire \crc_reflected[2] ;
 wire \crc_reflected[3] ;
 wire \crc_reflected[4] ;
 wire \crc_reflected[5] ;
 wire \crc_reflected[6] ;
 wire \crc_reflected[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net20;

 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _42_ (.A1(net9),
    .A2(\crc_reflected[6] ),
    .ZN(_08_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _43_ (.A1(\crc_reflected[0] ),
    .A2(net3),
    .ZN(_09_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _44_ (.A1(_08_),
    .A2(_09_),
    .Z(_10_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _45_ (.A1(net10),
    .A2(\crc_reflected[7] ),
    .A3(_10_),
    .ZN(_11_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _46_ (.A1(net11),
    .A2(\crc_reflected[0] ),
    .ZN(_12_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _47_ (.A1(net11),
    .A2(_11_),
    .B(_12_),
    .C(net2),
    .ZN(_00_));
 gf180mcu_fd_sc_mcu9t5v0__inv_2 _48_ (.I(net2),
    .ZN(_13_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _49_ (.A1(_13_),
    .A2(\crc_reflected[1] ),
    .Z(_14_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _50_ (.A1(net2),
    .A2(\crc_reflected[1] ),
    .ZN(_15_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _51_ (.A1(net4),
    .A2(_08_),
    .A3(_09_),
    .Z(_16_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _52_ (.A1(net11),
    .A2(_16_),
    .Z(_17_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _53_ (.I0(_14_),
    .I1(_15_),
    .S(_17_),
    .Z(_01_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _54_ (.A1(net5),
    .A2(\crc_reflected[2] ),
    .Z(_18_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _55_ (.A1(\crc_reflected[1] ),
    .A2(net4),
    .ZN(_19_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _56_ (.A1(_10_),
    .A2(_18_),
    .A3(_19_),
    .Z(_20_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _57_ (.A1(net11),
    .A2(\crc_reflected[2] ),
    .ZN(_21_));
 gf180mcu_fd_sc_mcu9t5v0__aoi211_2 _58_ (.A1(net11),
    .A2(_20_),
    .B(_21_),
    .C(net2),
    .ZN(_02_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _59_ (.A1(_13_),
    .A2(\crc_reflected[3] ),
    .Z(_22_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _60_ (.A1(net2),
    .A2(\crc_reflected[3] ),
    .ZN(_23_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _61_ (.A1(net10),
    .A2(\crc_reflected[7] ),
    .A3(net6),
    .Z(_24_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _62_ (.A1(_18_),
    .A2(_19_),
    .A3(_24_),
    .ZN(_25_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _63_ (.A1(net11),
    .A2(_25_),
    .Z(_26_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _64_ (.I0(_22_),
    .I1(_23_),
    .S(_26_),
    .Z(_03_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _65_ (.A1(net7),
    .A2(\crc_reflected[4] ),
    .Z(_27_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _66_ (.A1(net6),
    .A2(\crc_reflected[3] ),
    .ZN(_28_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _67_ (.A1(_18_),
    .A2(_27_),
    .A3(_28_),
    .ZN(_29_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _68_ (.I0(\crc_reflected[4] ),
    .I1(_29_),
    .S(net11),
    .Z(_30_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _69_ (.A1(_13_),
    .A2(_30_),
    .Z(_04_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _70_ (.A1(_13_),
    .A2(\crc_reflected[5] ),
    .Z(_31_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _71_ (.A1(net2),
    .A2(\crc_reflected[5] ),
    .ZN(_32_));
 gf180mcu_fd_sc_mcu9t5v0__xnor3_2 _72_ (.A1(net8),
    .A2(_27_),
    .A3(_28_),
    .ZN(_33_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _73_ (.A1(net11),
    .A2(_33_),
    .Z(_34_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _74_ (.I0(_31_),
    .I1(_32_),
    .S(_34_),
    .Z(_05_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _75_ (.A1(net8),
    .A2(\crc_reflected[5] ),
    .ZN(_35_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _76_ (.A1(_08_),
    .A2(_27_),
    .A3(_35_),
    .Z(_36_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _77_ (.I0(\crc_reflected[6] ),
    .I1(_36_),
    .S(net11),
    .Z(_37_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _78_ (.A1(_13_),
    .A2(_37_),
    .Z(_06_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _79_ (.A1(_13_),
    .A2(\crc_reflected[7] ),
    .Z(_38_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _80_ (.A1(net2),
    .A2(\crc_reflected[7] ),
    .ZN(_39_));
 gf180mcu_fd_sc_mcu9t5v0__xor3_2 _81_ (.A1(net10),
    .A2(_08_),
    .A3(_35_),
    .Z(_40_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _82_ (.A1(net11),
    .A2(_40_),
    .Z(_41_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _83_ (.I0(_38_),
    .I1(_39_),
    .S(_41_),
    .Z(_07_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \crc_out[0]$_DFF_PN0_  (.D(\crc_reflected[0] ),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net12));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \crc_out[1]$_DFF_PN0_  (.D(\crc_reflected[1] ),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net13));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \crc_out[2]$_DFF_PN0_  (.D(\crc_reflected[2] ),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(net14));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \crc_out[3]$_DFF_PN0_  (.D(\crc_reflected[3] ),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net15));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \crc_out[4]$_DFF_PN0_  (.D(\crc_reflected[4] ),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net16));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \crc_out[5]$_DFF_PN0_  (.D(\crc_reflected[5] ),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net17));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \crc_out[6]$_DFF_PN0_  (.D(\crc_reflected[6] ),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \crc_out[7]$_DFF_PN0_  (.D(\crc_reflected[7] ),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \crc_reg[0]$_DFFE_PN0P_  (.D(_00_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\crc_reflected[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \crc_reg[1]$_DFFE_PN0P_  (.D(_01_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\crc_reflected[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \crc_reg[2]$_DFFE_PN0P_  (.D(_02_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\crc_reflected[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \crc_reg[3]$_DFFE_PN0P_  (.D(_03_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\crc_reflected[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \crc_reg[4]$_DFFE_PN0P_  (.D(_04_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\crc_reflected[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \crc_reg[5]$_DFFE_PN0P_  (.D(_05_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\crc_reflected[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \crc_reg[6]$_DFFE_PN0P_  (.D(_06_),
    .RN(net1),
    .CLK(clknet_1_1__leaf_clk),
    .Q(\crc_reflected[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \crc_reg[7]$_DFFE_PN0P_  (.D(_07_),
    .RN(net1),
    .CLK(clknet_1_0__leaf_clk),
    .Q(\crc_reflected[7] ));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 hold1 (.I(net20),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_57 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_58 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_59 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_60 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_61 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_62 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_63 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_64 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_65 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_67 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_68 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_69 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_70 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_71 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_72 ();
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 input1 (.I(crc_init),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(data_in[0]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(data_in[1]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(data_in[2]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(data_in[3]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(data_in[4]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(data_in[5]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(data_in[6]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(data_in[7]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input10 (.I(data_valid),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output11 (.I(net12),
    .Z(crc_out[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output12 (.I(net13),
    .Z(crc_out[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output13 (.I(net14),
    .Z(crc_out[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output14 (.I(net15),
    .Z(crc_out[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output15 (.I(net16),
    .Z(crc_out[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output16 (.I(net17),
    .Z(crc_out[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output17 (.I(net18),
    .Z(crc_out[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output18 (.I(net19),
    .Z(crc_out[7]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_1_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload0 (.I(clknet_1_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_253 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_128 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_256 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_220 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_259 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_35 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_255 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_263 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_260 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_264 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_266 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_27_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_265 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_259 ();
endmodule
