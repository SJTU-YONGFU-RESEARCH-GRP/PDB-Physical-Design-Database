module wishbone_master (clk,
    read_done,
    read_err,
    read_req,
    rst_n,
    wb_ack_i,
    wb_cyc_o,
    wb_err_i,
    wb_rty_i,
    wb_stb_o,
    wb_tgd_i,
    wb_tgd_o,
    wb_we_o,
    write_done,
    write_err,
    write_req,
    read_addr,
    read_data,
    read_sel,
    wb_adr_o,
    wb_dat_i,
    wb_dat_o,
    wb_sel_o,
    write_addr,
    write_data,
    write_sel);
 input clk;
 output read_done;
 output read_err;
 input read_req;
 input rst_n;
 input wb_ack_i;
 output wb_cyc_o;
 input wb_err_i;
 input wb_rty_i;
 output wb_stb_o;
 input wb_tgd_i;
 output wb_tgd_o;
 output wb_we_o;
 output write_done;
 output write_err;
 input write_req;
 input [31:0] read_addr;
 output [31:0] read_data;
 input [3:0] read_sel;
 output [31:0] wb_adr_o;
 input [31:0] wb_dat_i;
 output [31:0] wb_dat_o;
 output [3:0] wb_sel_o;
 input [31:0] write_addr;
 input [31:0] write_data;
 input [3:0] write_sel;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire clknet_0_clk;
 wire _270_;
 wire \retry_count[0] ;
 wire \retry_count[1] ;
 wire \retry_count[2] ;
 wire \retry_count[3] ;
 wire \state[0] ;
 wire \state[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net250;

 sky130_fd_sc_hd__buf_4 _271_ (.A(_253_),
    .X(_111_));
 sky130_fd_sc_hd__nor4b_1 _272_ (.A(net39),
    .B(net72),
    .C(net73),
    .D_N(_254_),
    .Y(_112_));
 sky130_fd_sc_hd__nor2b_1 _273_ (.A(\retry_count[3] ),
    .B_N(_261_),
    .Y(_113_));
 sky130_fd_sc_hd__buf_4 _274_ (.A(write_req),
    .X(_114_));
 sky130_fd_sc_hd__nand2b_1 _275_ (.A_N(_114_),
    .B(_111_),
    .Y(_115_));
 sky130_fd_sc_hd__o32a_1 _276_ (.A1(_111_),
    .A2(_112_),
    .A3(_113_),
    .B1(net34),
    .B2(_115_),
    .X(_270_));
 sky130_fd_sc_hd__inv_1 _277_ (.A(\state[0] ),
    .Y(_251_));
 sky130_fd_sc_hd__inv_1 _278_ (.A(\retry_count[0] ),
    .Y(_263_));
 sky130_fd_sc_hd__inv_1 _279_ (.A(\state[1] ),
    .Y(_252_));
 sky130_fd_sc_hd__inv_1 _280_ (.A(\retry_count[1] ),
    .Y(_264_));
 sky130_fd_sc_hd__nand2_4 _281_ (.A(net39),
    .B(_255_),
    .Y(_116_));
 sky130_fd_sc_hd__buf_6 _282_ (.A(_116_),
    .X(_117_));
 sky130_fd_sc_hd__mux2_1 _283_ (.A0(net40),
    .A1(net142),
    .S(_117_),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _284_ (.A0(net41),
    .A1(net143),
    .S(_117_),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _285_ (.A0(net42),
    .A1(net144),
    .S(_117_),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _286_ (.A0(net43),
    .A1(net145),
    .S(_117_),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _287_ (.A0(net44),
    .A1(net146),
    .S(_117_),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _288_ (.A0(net45),
    .A1(net147),
    .S(_117_),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _289_ (.A0(net46),
    .A1(net148),
    .S(_117_),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _290_ (.A0(net47),
    .A1(net149),
    .S(_117_),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _291_ (.A0(net48),
    .A1(net150),
    .S(_117_),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _292_ (.A0(net49),
    .A1(net151),
    .S(_117_),
    .X(_009_));
 sky130_fd_sc_hd__buf_6 _293_ (.A(_116_),
    .X(_118_));
 sky130_fd_sc_hd__mux2_1 _294_ (.A0(net50),
    .A1(net152),
    .S(_118_),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _295_ (.A0(net51),
    .A1(net153),
    .S(_118_),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _296_ (.A0(net52),
    .A1(net154),
    .S(_118_),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _297_ (.A0(net53),
    .A1(net155),
    .S(_118_),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _298_ (.A0(net54),
    .A1(net156),
    .S(_118_),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _299_ (.A0(net55),
    .A1(net157),
    .S(_118_),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _300_ (.A0(net56),
    .A1(net158),
    .S(_118_),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _301_ (.A0(net57),
    .A1(net159),
    .S(_118_),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _302_ (.A0(net58),
    .A1(net160),
    .S(_118_),
    .X(_018_));
 sky130_fd_sc_hd__mux2_1 _303_ (.A0(net59),
    .A1(net161),
    .S(_118_),
    .X(_019_));
 sky130_fd_sc_hd__buf_6 _304_ (.A(_116_),
    .X(_119_));
 sky130_fd_sc_hd__mux2_1 _305_ (.A0(net60),
    .A1(net162),
    .S(_119_),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _306_ (.A0(net61),
    .A1(net163),
    .S(_119_),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _307_ (.A0(net62),
    .A1(net164),
    .S(_119_),
    .X(_022_));
 sky130_fd_sc_hd__mux2_1 _308_ (.A0(net63),
    .A1(net165),
    .S(_119_),
    .X(_023_));
 sky130_fd_sc_hd__mux2_1 _309_ (.A0(net64),
    .A1(net166),
    .S(_119_),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _310_ (.A0(net65),
    .A1(net167),
    .S(_119_),
    .X(_025_));
 sky130_fd_sc_hd__mux2_1 _311_ (.A0(net66),
    .A1(net168),
    .S(_119_),
    .X(_026_));
 sky130_fd_sc_hd__mux2_1 _312_ (.A0(net67),
    .A1(net169),
    .S(_119_),
    .X(_027_));
 sky130_fd_sc_hd__mux2_1 _313_ (.A0(net68),
    .A1(net170),
    .S(_119_),
    .X(_028_));
 sky130_fd_sc_hd__mux2_1 _314_ (.A0(net69),
    .A1(net171),
    .S(_119_),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _315_ (.A0(net70),
    .A1(net172),
    .S(_116_),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _316_ (.A0(net71),
    .A1(net173),
    .S(_116_),
    .X(_031_));
 sky130_fd_sc_hd__nand2b_1 _317_ (.A_N(_114_),
    .B(net34),
    .Y(_120_));
 sky130_fd_sc_hd__mux2i_1 _318_ (.A0(_255_),
    .A1(net174),
    .S(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__a21oi_1 _319_ (.A1(net39),
    .A2(_255_),
    .B1(net174),
    .Y(_122_));
 sky130_fd_sc_hd__a21oi_1 _320_ (.A1(_111_),
    .A2(_121_),
    .B1(_122_),
    .Y(_032_));
 sky130_fd_sc_hd__buf_2 _321_ (.A(_254_),
    .X(_123_));
 sky130_fd_sc_hd__inv_1 _322_ (.A(net175),
    .Y(_124_));
 sky130_fd_sc_hd__buf_2 _323_ (.A(_261_),
    .X(_125_));
 sky130_fd_sc_hd__a211oi_1 _324_ (.A1(_111_),
    .A2(_120_),
    .B1(_123_),
    .C1(_125_),
    .Y(_126_));
 sky130_fd_sc_hd__a21oi_1 _325_ (.A1(_123_),
    .A2(_124_),
    .B1(_126_),
    .Y(_127_));
 sky130_fd_sc_hd__inv_1 _326_ (.A(net246),
    .Y(_128_));
 sky130_fd_sc_hd__nand2_1 _327_ (.A(\retry_count[3] ),
    .B(_128_),
    .Y(_129_));
 sky130_fd_sc_hd__nand2b_1 _328_ (.A_N(net39),
    .B(net72),
    .Y(_130_));
 sky130_fd_sc_hd__a222oi_1 _329_ (.A1(_111_),
    .A2(_120_),
    .B1(_129_),
    .B2(_125_),
    .C1(_130_),
    .C2(_255_),
    .Y(_131_));
 sky130_fd_sc_hd__o22a_1 _330_ (.A1(_255_),
    .A2(_127_),
    .B1(_131_),
    .B2(net175),
    .X(_033_));
 sky130_fd_sc_hd__nor2_1 _331_ (.A(net39),
    .B(net72),
    .Y(_132_));
 sky130_fd_sc_hd__nand2_1 _332_ (.A(net73),
    .B(_132_),
    .Y(_133_));
 sky130_fd_sc_hd__a21oi_1 _333_ (.A1(_123_),
    .A2(_133_),
    .B1(_125_),
    .Y(_134_));
 sky130_fd_sc_hd__nor3b_1 _334_ (.A(net39),
    .B(net72),
    .C_N(net73),
    .Y(_135_));
 sky130_fd_sc_hd__nand3b_1 _335_ (.A_N(_125_),
    .B(_123_),
    .C(_135_),
    .Y(_136_));
 sky130_fd_sc_hd__mux2i_1 _336_ (.A0(_134_),
    .A1(_136_),
    .S(_263_),
    .Y(_034_));
 sky130_fd_sc_hd__inv_1 _337_ (.A(_266_),
    .Y(_137_));
 sky130_fd_sc_hd__o22ai_1 _338_ (.A1(_264_),
    .A2(_134_),
    .B1(_136_),
    .B2(_137_),
    .Y(_035_));
 sky130_fd_sc_hd__nand2_1 _339_ (.A(_267_),
    .B(_135_),
    .Y(_138_));
 sky130_fd_sc_hd__nor2_1 _340_ (.A(\retry_count[2] ),
    .B(_125_),
    .Y(_139_));
 sky130_fd_sc_hd__nand2_1 _341_ (.A(_123_),
    .B(_139_),
    .Y(_140_));
 sky130_fd_sc_hd__a21oi_1 _342_ (.A1(_123_),
    .A2(_138_),
    .B1(_125_),
    .Y(_141_));
 sky130_fd_sc_hd__inv_1 _343_ (.A(\retry_count[2] ),
    .Y(_142_));
 sky130_fd_sc_hd__o22ai_1 _344_ (.A1(_138_),
    .A2(_140_),
    .B1(_141_),
    .B2(_142_),
    .Y(_036_));
 sky130_fd_sc_hd__nand4_1 _345_ (.A(\retry_count[2] ),
    .B(\retry_count[0] ),
    .C(\retry_count[1] ),
    .D(_135_),
    .Y(_143_));
 sky130_fd_sc_hd__nor2_1 _346_ (.A(\retry_count[3] ),
    .B(_125_),
    .Y(_144_));
 sky130_fd_sc_hd__nand2_1 _347_ (.A(_123_),
    .B(_144_),
    .Y(_145_));
 sky130_fd_sc_hd__a21oi_1 _348_ (.A1(_123_),
    .A2(_143_),
    .B1(_125_),
    .Y(_146_));
 sky130_fd_sc_hd__inv_1 _349_ (.A(\retry_count[3] ),
    .Y(_147_));
 sky130_fd_sc_hd__o22ai_1 _350_ (.A1(_143_),
    .A2(_145_),
    .B1(_146_),
    .B2(_147_),
    .Y(_037_));
 sky130_fd_sc_hd__buf_6 _351_ (.A(_114_),
    .X(_148_));
 sky130_fd_sc_hd__nor2b_1 _352_ (.A(_148_),
    .B_N(_111_),
    .Y(_149_));
 sky130_fd_sc_hd__a221oi_1 _353_ (.A1(_123_),
    .A2(_132_),
    .B1(_113_),
    .B2(net246),
    .C1(_111_),
    .Y(_150_));
 sky130_fd_sc_hd__o21bai_1 _354_ (.A1(net34),
    .A2(_115_),
    .B1_N(_112_),
    .Y(_151_));
 sky130_fd_sc_hd__nand2_1 _355_ (.A(\state[0] ),
    .B(_151_),
    .Y(_152_));
 sky130_fd_sc_hd__o31ai_1 _356_ (.A1(_149_),
    .A2(_112_),
    .A3(_150_),
    .B1(_152_),
    .Y(_038_));
 sky130_fd_sc_hd__a221oi_1 _357_ (.A1(_123_),
    .A2(_132_),
    .B1(_113_),
    .B2(_128_),
    .C1(_111_),
    .Y(_153_));
 sky130_fd_sc_hd__nand2_4 _358_ (.A(_111_),
    .B(_114_),
    .Y(_154_));
 sky130_fd_sc_hd__nand2b_1 _359_ (.A_N(_151_),
    .B(_154_),
    .Y(_155_));
 sky130_fd_sc_hd__nand2_1 _360_ (.A(\state[1] ),
    .B(_151_),
    .Y(_156_));
 sky130_fd_sc_hd__o21ai_0 _361_ (.A1(_153_),
    .A2(_155_),
    .B1(_156_),
    .Y(_039_));
 sky130_fd_sc_hd__o21ai_4 _362_ (.A1(_114_),
    .A2(net34),
    .B1(_253_),
    .Y(_157_));
 sky130_fd_sc_hd__clkbuf_4 _363_ (.A(_157_),
    .X(_158_));
 sky130_fd_sc_hd__buf_6 _364_ (.A(_148_),
    .X(_159_));
 sky130_fd_sc_hd__mux2i_1 _365_ (.A0(net2),
    .A1(net74),
    .S(_159_),
    .Y(_160_));
 sky130_fd_sc_hd__buf_2 _366_ (.A(_157_),
    .X(_161_));
 sky130_fd_sc_hd__nand2_1 _367_ (.A(net176),
    .B(_161_),
    .Y(_162_));
 sky130_fd_sc_hd__o21ai_0 _368_ (.A1(_158_),
    .A2(_160_),
    .B1(_162_),
    .Y(_040_));
 sky130_fd_sc_hd__mux2i_2 _369_ (.A0(net3),
    .A1(net75),
    .S(_159_),
    .Y(_163_));
 sky130_fd_sc_hd__nand2_1 _370_ (.A(net177),
    .B(_161_),
    .Y(_164_));
 sky130_fd_sc_hd__o21ai_0 _371_ (.A1(_158_),
    .A2(_163_),
    .B1(_164_),
    .Y(_041_));
 sky130_fd_sc_hd__mux2i_1 _372_ (.A0(net4),
    .A1(net76),
    .S(_159_),
    .Y(_165_));
 sky130_fd_sc_hd__nand2_1 _373_ (.A(net178),
    .B(_161_),
    .Y(_166_));
 sky130_fd_sc_hd__o21ai_0 _374_ (.A1(_158_),
    .A2(_165_),
    .B1(_166_),
    .Y(_042_));
 sky130_fd_sc_hd__mux2i_1 _375_ (.A0(net5),
    .A1(net77),
    .S(_159_),
    .Y(_167_));
 sky130_fd_sc_hd__nand2_1 _376_ (.A(net179),
    .B(_161_),
    .Y(_168_));
 sky130_fd_sc_hd__o21ai_0 _377_ (.A1(_158_),
    .A2(_167_),
    .B1(_168_),
    .Y(_043_));
 sky130_fd_sc_hd__buf_2 _378_ (.A(_157_),
    .X(_169_));
 sky130_fd_sc_hd__mux2i_1 _379_ (.A0(net6),
    .A1(net78),
    .S(_159_),
    .Y(_170_));
 sky130_fd_sc_hd__nand2_1 _380_ (.A(net180),
    .B(_161_),
    .Y(_171_));
 sky130_fd_sc_hd__o21ai_0 _381_ (.A1(_169_),
    .A2(_170_),
    .B1(_171_),
    .Y(_044_));
 sky130_fd_sc_hd__mux2i_1 _382_ (.A0(net7),
    .A1(net79),
    .S(_159_),
    .Y(_172_));
 sky130_fd_sc_hd__nand2_1 _383_ (.A(net181),
    .B(_161_),
    .Y(_173_));
 sky130_fd_sc_hd__o21ai_0 _384_ (.A1(_169_),
    .A2(_172_),
    .B1(_173_),
    .Y(_045_));
 sky130_fd_sc_hd__mux2i_1 _385_ (.A0(net8),
    .A1(net80),
    .S(_159_),
    .Y(_174_));
 sky130_fd_sc_hd__nand2_1 _386_ (.A(net182),
    .B(_161_),
    .Y(_175_));
 sky130_fd_sc_hd__o21ai_0 _387_ (.A1(_169_),
    .A2(_174_),
    .B1(_175_),
    .Y(_046_));
 sky130_fd_sc_hd__mux2i_1 _388_ (.A0(net9),
    .A1(net81),
    .S(_159_),
    .Y(_176_));
 sky130_fd_sc_hd__nand2_1 _389_ (.A(net183),
    .B(_161_),
    .Y(_177_));
 sky130_fd_sc_hd__o21ai_0 _390_ (.A1(_169_),
    .A2(_176_),
    .B1(_177_),
    .Y(_047_));
 sky130_fd_sc_hd__mux2i_1 _391_ (.A0(net10),
    .A1(net82),
    .S(_159_),
    .Y(_178_));
 sky130_fd_sc_hd__nand2_1 _392_ (.A(net184),
    .B(_161_),
    .Y(_179_));
 sky130_fd_sc_hd__o21ai_0 _393_ (.A1(_169_),
    .A2(_178_),
    .B1(_179_),
    .Y(_048_));
 sky130_fd_sc_hd__mux2i_1 _394_ (.A0(net11),
    .A1(net83),
    .S(_159_),
    .Y(_180_));
 sky130_fd_sc_hd__nand2_1 _395_ (.A(net185),
    .B(_161_),
    .Y(_181_));
 sky130_fd_sc_hd__o21ai_0 _396_ (.A1(_169_),
    .A2(_180_),
    .B1(_181_),
    .Y(_049_));
 sky130_fd_sc_hd__buf_6 _397_ (.A(_148_),
    .X(_182_));
 sky130_fd_sc_hd__mux2i_1 _398_ (.A0(net12),
    .A1(net84),
    .S(_182_),
    .Y(_183_));
 sky130_fd_sc_hd__buf_2 _399_ (.A(_157_),
    .X(_184_));
 sky130_fd_sc_hd__nand2_1 _400_ (.A(net186),
    .B(_184_),
    .Y(_185_));
 sky130_fd_sc_hd__o21ai_0 _401_ (.A1(_169_),
    .A2(_183_),
    .B1(_185_),
    .Y(_050_));
 sky130_fd_sc_hd__mux2i_1 _402_ (.A0(net13),
    .A1(net85),
    .S(_182_),
    .Y(_186_));
 sky130_fd_sc_hd__nand2_1 _403_ (.A(net187),
    .B(_184_),
    .Y(_187_));
 sky130_fd_sc_hd__o21ai_0 _404_ (.A1(_169_),
    .A2(_186_),
    .B1(_187_),
    .Y(_051_));
 sky130_fd_sc_hd__mux2i_1 _405_ (.A0(net14),
    .A1(net86),
    .S(_182_),
    .Y(_188_));
 sky130_fd_sc_hd__nand2_1 _406_ (.A(net188),
    .B(_184_),
    .Y(_189_));
 sky130_fd_sc_hd__o21ai_0 _407_ (.A1(_169_),
    .A2(_188_),
    .B1(_189_),
    .Y(_052_));
 sky130_fd_sc_hd__mux2i_1 _408_ (.A0(net15),
    .A1(net87),
    .S(_182_),
    .Y(_190_));
 sky130_fd_sc_hd__nand2_1 _409_ (.A(net189),
    .B(_184_),
    .Y(_191_));
 sky130_fd_sc_hd__o21ai_0 _410_ (.A1(_169_),
    .A2(_190_),
    .B1(_191_),
    .Y(_053_));
 sky130_fd_sc_hd__clkbuf_2 _411_ (.A(_157_),
    .X(_192_));
 sky130_fd_sc_hd__mux2i_1 _412_ (.A0(net16),
    .A1(net88),
    .S(_182_),
    .Y(_193_));
 sky130_fd_sc_hd__nand2_1 _413_ (.A(net190),
    .B(_184_),
    .Y(_194_));
 sky130_fd_sc_hd__o21ai_0 _414_ (.A1(_192_),
    .A2(_193_),
    .B1(_194_),
    .Y(_054_));
 sky130_fd_sc_hd__mux2i_1 _415_ (.A0(net17),
    .A1(net89),
    .S(_182_),
    .Y(_195_));
 sky130_fd_sc_hd__nand2_1 _416_ (.A(net191),
    .B(_184_),
    .Y(_196_));
 sky130_fd_sc_hd__o21ai_0 _417_ (.A1(_192_),
    .A2(_195_),
    .B1(_196_),
    .Y(_055_));
 sky130_fd_sc_hd__mux2i_1 _418_ (.A0(net18),
    .A1(net90),
    .S(_182_),
    .Y(_197_));
 sky130_fd_sc_hd__nand2_1 _419_ (.A(net192),
    .B(_184_),
    .Y(_198_));
 sky130_fd_sc_hd__o21ai_0 _420_ (.A1(_192_),
    .A2(_197_),
    .B1(_198_),
    .Y(_056_));
 sky130_fd_sc_hd__mux2i_1 _421_ (.A0(net19),
    .A1(net91),
    .S(_182_),
    .Y(_199_));
 sky130_fd_sc_hd__nand2_1 _422_ (.A(net193),
    .B(_184_),
    .Y(_200_));
 sky130_fd_sc_hd__o21ai_0 _423_ (.A1(_192_),
    .A2(_199_),
    .B1(_200_),
    .Y(_057_));
 sky130_fd_sc_hd__mux2i_1 _424_ (.A0(net20),
    .A1(net92),
    .S(_182_),
    .Y(_201_));
 sky130_fd_sc_hd__nand2_1 _425_ (.A(net194),
    .B(_184_),
    .Y(_202_));
 sky130_fd_sc_hd__o21ai_0 _426_ (.A1(_192_),
    .A2(_201_),
    .B1(_202_),
    .Y(_058_));
 sky130_fd_sc_hd__mux2i_1 _427_ (.A0(net21),
    .A1(net93),
    .S(_182_),
    .Y(_203_));
 sky130_fd_sc_hd__nand2_1 _428_ (.A(net195),
    .B(_184_),
    .Y(_204_));
 sky130_fd_sc_hd__o21ai_0 _429_ (.A1(_192_),
    .A2(_203_),
    .B1(_204_),
    .Y(_059_));
 sky130_fd_sc_hd__buf_6 _430_ (.A(_148_),
    .X(_205_));
 sky130_fd_sc_hd__mux2i_1 _431_ (.A0(net22),
    .A1(net94),
    .S(_205_),
    .Y(_206_));
 sky130_fd_sc_hd__buf_2 _432_ (.A(_157_),
    .X(_207_));
 sky130_fd_sc_hd__nand2_1 _433_ (.A(net196),
    .B(_207_),
    .Y(_208_));
 sky130_fd_sc_hd__o21ai_0 _434_ (.A1(_192_),
    .A2(_206_),
    .B1(_208_),
    .Y(_060_));
 sky130_fd_sc_hd__mux2i_1 _435_ (.A0(net23),
    .A1(net95),
    .S(_205_),
    .Y(_209_));
 sky130_fd_sc_hd__nand2_1 _436_ (.A(net197),
    .B(_207_),
    .Y(_210_));
 sky130_fd_sc_hd__o21ai_0 _437_ (.A1(_192_),
    .A2(_209_),
    .B1(_210_),
    .Y(_061_));
 sky130_fd_sc_hd__mux2i_1 _438_ (.A0(net24),
    .A1(net96),
    .S(_205_),
    .Y(_211_));
 sky130_fd_sc_hd__nand2_1 _439_ (.A(net198),
    .B(_207_),
    .Y(_212_));
 sky130_fd_sc_hd__o21ai_0 _440_ (.A1(_192_),
    .A2(_211_),
    .B1(_212_),
    .Y(_062_));
 sky130_fd_sc_hd__mux2i_1 _441_ (.A0(net25),
    .A1(net97),
    .S(_205_),
    .Y(_213_));
 sky130_fd_sc_hd__nand2_1 _442_ (.A(net199),
    .B(_207_),
    .Y(_214_));
 sky130_fd_sc_hd__o21ai_0 _443_ (.A1(_192_),
    .A2(_213_),
    .B1(_214_),
    .Y(_063_));
 sky130_fd_sc_hd__buf_2 _444_ (.A(_157_),
    .X(_215_));
 sky130_fd_sc_hd__mux2i_1 _445_ (.A0(net26),
    .A1(net98),
    .S(_205_),
    .Y(_216_));
 sky130_fd_sc_hd__nand2_1 _446_ (.A(net200),
    .B(_207_),
    .Y(_217_));
 sky130_fd_sc_hd__o21ai_0 _447_ (.A1(_215_),
    .A2(_216_),
    .B1(_217_),
    .Y(_064_));
 sky130_fd_sc_hd__mux2i_1 _448_ (.A0(net27),
    .A1(net99),
    .S(_205_),
    .Y(_218_));
 sky130_fd_sc_hd__nand2_1 _449_ (.A(net201),
    .B(_207_),
    .Y(_219_));
 sky130_fd_sc_hd__o21ai_0 _450_ (.A1(_215_),
    .A2(_218_),
    .B1(_219_),
    .Y(_065_));
 sky130_fd_sc_hd__mux2i_1 _451_ (.A0(net28),
    .A1(net100),
    .S(_205_),
    .Y(_220_));
 sky130_fd_sc_hd__nand2_1 _452_ (.A(net202),
    .B(_207_),
    .Y(_221_));
 sky130_fd_sc_hd__o21ai_0 _453_ (.A1(_215_),
    .A2(_220_),
    .B1(_221_),
    .Y(_066_));
 sky130_fd_sc_hd__mux2i_1 _454_ (.A0(net29),
    .A1(net101),
    .S(_205_),
    .Y(_222_));
 sky130_fd_sc_hd__nand2_1 _455_ (.A(net203),
    .B(_207_),
    .Y(_223_));
 sky130_fd_sc_hd__o21ai_0 _456_ (.A1(_215_),
    .A2(_222_),
    .B1(_223_),
    .Y(_067_));
 sky130_fd_sc_hd__mux2i_1 _457_ (.A0(net30),
    .A1(net102),
    .S(_205_),
    .Y(_224_));
 sky130_fd_sc_hd__nand2_1 _458_ (.A(net204),
    .B(_207_),
    .Y(_225_));
 sky130_fd_sc_hd__o21ai_0 _459_ (.A1(_215_),
    .A2(_224_),
    .B1(_225_),
    .Y(_068_));
 sky130_fd_sc_hd__mux2i_1 _460_ (.A0(net31),
    .A1(net103),
    .S(_205_),
    .Y(_226_));
 sky130_fd_sc_hd__nand2_1 _461_ (.A(net205),
    .B(_207_),
    .Y(_227_));
 sky130_fd_sc_hd__o21ai_0 _462_ (.A1(_215_),
    .A2(_226_),
    .B1(_227_),
    .Y(_069_));
 sky130_fd_sc_hd__mux2i_1 _463_ (.A0(net32),
    .A1(net104),
    .S(_148_),
    .Y(_228_));
 sky130_fd_sc_hd__nand2_1 _464_ (.A(net206),
    .B(_158_),
    .Y(_229_));
 sky130_fd_sc_hd__o21ai_0 _465_ (.A1(_215_),
    .A2(_228_),
    .B1(_229_),
    .Y(_070_));
 sky130_fd_sc_hd__mux2i_1 _466_ (.A0(net33),
    .A1(net105),
    .S(_148_),
    .Y(_230_));
 sky130_fd_sc_hd__nand2_1 _467_ (.A(net207),
    .B(_158_),
    .Y(_231_));
 sky130_fd_sc_hd__o21ai_0 _468_ (.A1(_215_),
    .A2(_230_),
    .B1(_231_),
    .Y(_071_));
 sky130_fd_sc_hd__buf_6 _469_ (.A(_154_),
    .X(_232_));
 sky130_fd_sc_hd__mux2_1 _470_ (.A0(net106),
    .A1(net209),
    .S(_232_),
    .X(_072_));
 sky130_fd_sc_hd__mux2_1 _471_ (.A0(net107),
    .A1(net210),
    .S(_232_),
    .X(_073_));
 sky130_fd_sc_hd__mux2_1 _472_ (.A0(net108),
    .A1(net211),
    .S(_232_),
    .X(_074_));
 sky130_fd_sc_hd__mux2_1 _473_ (.A0(net109),
    .A1(net212),
    .S(_232_),
    .X(_075_));
 sky130_fd_sc_hd__mux2_1 _474_ (.A0(net110),
    .A1(net213),
    .S(_232_),
    .X(_076_));
 sky130_fd_sc_hd__mux2_1 _475_ (.A0(net111),
    .A1(net214),
    .S(_232_),
    .X(_077_));
 sky130_fd_sc_hd__mux2_1 _476_ (.A0(net112),
    .A1(net215),
    .S(_232_),
    .X(_078_));
 sky130_fd_sc_hd__mux2_1 _477_ (.A0(net113),
    .A1(net216),
    .S(_232_),
    .X(_079_));
 sky130_fd_sc_hd__buf_6 _478_ (.A(_154_),
    .X(_233_));
 sky130_fd_sc_hd__mux2_1 _479_ (.A0(net114),
    .A1(net217),
    .S(_233_),
    .X(_080_));
 sky130_fd_sc_hd__mux2_1 _480_ (.A0(net115),
    .A1(net218),
    .S(_233_),
    .X(_081_));
 sky130_fd_sc_hd__mux2_1 _481_ (.A0(net116),
    .A1(net219),
    .S(_233_),
    .X(_082_));
 sky130_fd_sc_hd__mux2_1 _482_ (.A0(net117),
    .A1(net220),
    .S(_233_),
    .X(_083_));
 sky130_fd_sc_hd__mux2_1 _483_ (.A0(net118),
    .A1(net221),
    .S(_233_),
    .X(_084_));
 sky130_fd_sc_hd__mux2_1 _484_ (.A0(net119),
    .A1(net222),
    .S(_233_),
    .X(_085_));
 sky130_fd_sc_hd__mux2_1 _485_ (.A0(net120),
    .A1(net223),
    .S(_233_),
    .X(_086_));
 sky130_fd_sc_hd__mux2_1 _486_ (.A0(net121),
    .A1(net224),
    .S(_233_),
    .X(_087_));
 sky130_fd_sc_hd__mux2_1 _487_ (.A0(net122),
    .A1(net225),
    .S(_233_),
    .X(_088_));
 sky130_fd_sc_hd__mux2_1 _488_ (.A0(net123),
    .A1(net226),
    .S(_233_),
    .X(_089_));
 sky130_fd_sc_hd__buf_6 _489_ (.A(_154_),
    .X(_234_));
 sky130_fd_sc_hd__mux2_1 _490_ (.A0(net124),
    .A1(net227),
    .S(_234_),
    .X(_090_));
 sky130_fd_sc_hd__mux2_1 _491_ (.A0(net125),
    .A1(net228),
    .S(_234_),
    .X(_091_));
 sky130_fd_sc_hd__mux2_1 _492_ (.A0(net126),
    .A1(net229),
    .S(_234_),
    .X(_092_));
 sky130_fd_sc_hd__mux2_1 _493_ (.A0(net127),
    .A1(net230),
    .S(_234_),
    .X(_093_));
 sky130_fd_sc_hd__mux2_1 _494_ (.A0(net128),
    .A1(net231),
    .S(_234_),
    .X(_094_));
 sky130_fd_sc_hd__mux2_1 _495_ (.A0(net129),
    .A1(net232),
    .S(_234_),
    .X(_095_));
 sky130_fd_sc_hd__mux2_1 _496_ (.A0(net130),
    .A1(net233),
    .S(_234_),
    .X(_096_));
 sky130_fd_sc_hd__mux2_1 _497_ (.A0(net131),
    .A1(net234),
    .S(_234_),
    .X(_097_));
 sky130_fd_sc_hd__mux2_1 _498_ (.A0(net132),
    .A1(net235),
    .S(_234_),
    .X(_098_));
 sky130_fd_sc_hd__mux2_1 _499_ (.A0(net133),
    .A1(net236),
    .S(_234_),
    .X(_099_));
 sky130_fd_sc_hd__mux2_1 _500_ (.A0(net134),
    .A1(net237),
    .S(_154_),
    .X(_100_));
 sky130_fd_sc_hd__mux2_1 _501_ (.A0(net135),
    .A1(net238),
    .S(_154_),
    .X(_101_));
 sky130_fd_sc_hd__mux2_1 _502_ (.A0(net136),
    .A1(net239),
    .S(_154_),
    .X(_102_));
 sky130_fd_sc_hd__mux2_1 _503_ (.A0(net137),
    .A1(net240),
    .S(_154_),
    .X(_103_));
 sky130_fd_sc_hd__mux2i_1 _504_ (.A0(net35),
    .A1(net138),
    .S(_148_),
    .Y(_235_));
 sky130_fd_sc_hd__nand2_1 _505_ (.A(net241),
    .B(_158_),
    .Y(_236_));
 sky130_fd_sc_hd__o21ai_0 _506_ (.A1(_215_),
    .A2(_235_),
    .B1(_236_),
    .Y(_104_));
 sky130_fd_sc_hd__mux2i_1 _507_ (.A0(net36),
    .A1(net139),
    .S(_148_),
    .Y(_237_));
 sky130_fd_sc_hd__nand2_1 _508_ (.A(net242),
    .B(_158_),
    .Y(_238_));
 sky130_fd_sc_hd__o21ai_0 _509_ (.A1(_215_),
    .A2(_237_),
    .B1(_238_),
    .Y(_105_));
 sky130_fd_sc_hd__mux2i_1 _510_ (.A0(net37),
    .A1(net140),
    .S(_148_),
    .Y(_239_));
 sky130_fd_sc_hd__nand2_1 _511_ (.A(net243),
    .B(_158_),
    .Y(_240_));
 sky130_fd_sc_hd__o21ai_0 _512_ (.A1(_157_),
    .A2(_239_),
    .B1(_240_),
    .Y(_106_));
 sky130_fd_sc_hd__mux2i_2 _513_ (.A0(net38),
    .A1(net141),
    .S(_148_),
    .Y(_241_));
 sky130_fd_sc_hd__nand2_1 _514_ (.A(net244),
    .B(_158_),
    .Y(_242_));
 sky130_fd_sc_hd__o21ai_0 _515_ (.A1(_157_),
    .A2(_241_),
    .B1(_242_),
    .Y(_107_));
 sky130_fd_sc_hd__and2_0 _516_ (.A(_111_),
    .B(net34),
    .X(_243_));
 sky130_fd_sc_hd__o21ai_0 _517_ (.A1(_128_),
    .A2(_243_),
    .B1(_232_),
    .Y(_108_));
 sky130_fd_sc_hd__a21oi_1 _518_ (.A1(net39),
    .A2(_115_),
    .B1(net247),
    .Y(_244_));
 sky130_fd_sc_hd__a21oi_1 _519_ (.A1(net247),
    .A2(_232_),
    .B1(_259_),
    .Y(_245_));
 sky130_fd_sc_hd__nor2_1 _520_ (.A(_244_),
    .B(_245_),
    .Y(_109_));
 sky130_fd_sc_hd__nor2_1 _521_ (.A(_257_),
    .B(_149_),
    .Y(_246_));
 sky130_fd_sc_hd__nor2_1 _522_ (.A(_259_),
    .B(_125_),
    .Y(_247_));
 sky130_fd_sc_hd__o21ai_0 _523_ (.A1(_147_),
    .A2(_128_),
    .B1(_125_),
    .Y(_248_));
 sky130_fd_sc_hd__nand2_1 _524_ (.A(_259_),
    .B(_130_),
    .Y(_249_));
 sky130_fd_sc_hd__a31oi_1 _525_ (.A1(_248_),
    .A2(_249_),
    .A3(_246_),
    .B1(net248),
    .Y(_250_));
 sky130_fd_sc_hd__a21oi_1 _526_ (.A1(_246_),
    .A2(_247_),
    .B1(_250_),
    .Y(_110_));
 sky130_fd_sc_hd__ha_1 _527_ (.A(_251_),
    .B(_252_),
    .COUT(_253_),
    .SUM(_254_));
 sky130_fd_sc_hd__ha_2 _528_ (.A(_251_),
    .B(\state[1] ),
    .COUT(_255_),
    .SUM(_256_));
 sky130_fd_sc_hd__ha_1 _529_ (.A(_251_),
    .B(\state[1] ),
    .COUT(_257_),
    .SUM(_258_));
 sky130_fd_sc_hd__ha_1 _530_ (.A(\state[0] ),
    .B(_252_),
    .COUT(_259_),
    .SUM(_260_));
 sky130_fd_sc_hd__ha_1 _531_ (.A(\state[0] ),
    .B(\state[1] ),
    .COUT(_261_),
    .SUM(_262_));
 sky130_fd_sc_hd__ha_1 _532_ (.A(_263_),
    .B(_264_),
    .COUT(_265_),
    .SUM(_266_));
 sky130_fd_sc_hd__ha_1 _533_ (.A(\retry_count[0] ),
    .B(\retry_count[1] ),
    .COUT(_267_),
    .SUM(_268_));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_1 _535_ (.A(net208),
    .X(net245));
 sky130_fd_sc_hd__buf_4 _536_ (.A(net249),
    .X(wb_tgd_o));
 sky130_fd_sc_hd__dfrtp_1 \read_data[0]$_DFFE_PN0P_  (.D(_000_),
    .Q(net142),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[10]$_DFFE_PN0P_  (.D(_001_),
    .Q(net143),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[11]$_DFFE_PN0P_  (.D(_002_),
    .Q(net144),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[12]$_DFFE_PN0P_  (.D(_003_),
    .Q(net145),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[13]$_DFFE_PN0P_  (.D(_004_),
    .Q(net146),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[14]$_DFFE_PN0P_  (.D(_005_),
    .Q(net147),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[15]$_DFFE_PN0P_  (.D(_006_),
    .Q(net148),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[16]$_DFFE_PN0P_  (.D(_007_),
    .Q(net149),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[17]$_DFFE_PN0P_  (.D(_008_),
    .Q(net150),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[18]$_DFFE_PN0P_  (.D(_009_),
    .Q(net151),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[19]$_DFFE_PN0P_  (.D(_010_),
    .Q(net152),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[1]$_DFFE_PN0P_  (.D(_011_),
    .Q(net153),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[20]$_DFFE_PN0P_  (.D(_012_),
    .Q(net154),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[21]$_DFFE_PN0P_  (.D(_013_),
    .Q(net155),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[22]$_DFFE_PN0P_  (.D(_014_),
    .Q(net156),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[23]$_DFFE_PN0P_  (.D(_015_),
    .Q(net157),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[24]$_DFFE_PN0P_  (.D(_016_),
    .Q(net158),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[25]$_DFFE_PN0P_  (.D(_017_),
    .Q(net159),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[26]$_DFFE_PN0P_  (.D(_018_),
    .Q(net160),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[27]$_DFFE_PN0P_  (.D(_019_),
    .Q(net161),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[28]$_DFFE_PN0P_  (.D(_020_),
    .Q(net162),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[29]$_DFFE_PN0P_  (.D(_021_),
    .Q(net163),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[2]$_DFFE_PN0P_  (.D(_022_),
    .Q(net164),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[30]$_DFFE_PN0P_  (.D(_023_),
    .Q(net165),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[31]$_DFFE_PN0P_  (.D(_024_),
    .Q(net166),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[3]$_DFFE_PN0P_  (.D(_025_),
    .Q(net167),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[4]$_DFFE_PN0P_  (.D(_026_),
    .Q(net168),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[5]$_DFFE_PN0P_  (.D(_027_),
    .Q(net169),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[6]$_DFFE_PN0P_  (.D(_028_),
    .Q(net170),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[7]$_DFFE_PN0P_  (.D(_029_),
    .Q(net171),
    .RESET_B(net1),
    .CLK(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[8]$_DFFE_PN0P_  (.D(_030_),
    .Q(net172),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_data[9]$_DFFE_PN0P_  (.D(_031_),
    .Q(net173),
    .RESET_B(net1),
    .CLK(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_done$_DFFE_PN0P_  (.D(_032_),
    .Q(net174),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \read_err$_DFFE_PN0P_  (.D(_033_),
    .Q(net175),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \retry_count[0]$_DFFE_PN0P_  (.D(_034_),
    .Q(\retry_count[0] ),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \retry_count[1]$_DFFE_PN0P_  (.D(_035_),
    .Q(\retry_count[1] ),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \retry_count[2]$_DFFE_PN0P_  (.D(_036_),
    .Q(\retry_count[2] ),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \retry_count[3]$_DFFE_PN0P_  (.D(_037_),
    .Q(\retry_count[3] ),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \state[0]$_DFFE_PN0P_  (.D(_038_),
    .Q(\state[0] ),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \state[1]$_DFFE_PN0P_  (.D(_039_),
    .Q(\state[1] ),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[0]$_DFFE_PN0P_  (.D(_040_),
    .Q(net176),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[10]$_DFFE_PN0P_  (.D(_041_),
    .Q(net177),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[11]$_DFFE_PN0P_  (.D(_042_),
    .Q(net178),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[12]$_DFFE_PN0P_  (.D(_043_),
    .Q(net179),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[13]$_DFFE_PN0P_  (.D(_044_),
    .Q(net180),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[14]$_DFFE_PN0P_  (.D(_045_),
    .Q(net181),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[15]$_DFFE_PN0P_  (.D(_046_),
    .Q(net182),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[16]$_DFFE_PN0P_  (.D(_047_),
    .Q(net183),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[17]$_DFFE_PN0P_  (.D(_048_),
    .Q(net184),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[18]$_DFFE_PN0P_  (.D(_049_),
    .Q(net185),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[19]$_DFFE_PN0P_  (.D(_050_),
    .Q(net186),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[1]$_DFFE_PN0P_  (.D(_051_),
    .Q(net187),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[20]$_DFFE_PN0P_  (.D(_052_),
    .Q(net188),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[21]$_DFFE_PN0P_  (.D(_053_),
    .Q(net189),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[22]$_DFFE_PN0P_  (.D(_054_),
    .Q(net190),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[23]$_DFFE_PN0P_  (.D(_055_),
    .Q(net191),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[24]$_DFFE_PN0P_  (.D(_056_),
    .Q(net192),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[25]$_DFFE_PN0P_  (.D(_057_),
    .Q(net193),
    .RESET_B(net1),
    .CLK(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[26]$_DFFE_PN0P_  (.D(_058_),
    .Q(net194),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[27]$_DFFE_PN0P_  (.D(_059_),
    .Q(net195),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[28]$_DFFE_PN0P_  (.D(_060_),
    .Q(net196),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[29]$_DFFE_PN0P_  (.D(_061_),
    .Q(net197),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[2]$_DFFE_PN0P_  (.D(_062_),
    .Q(net198),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[30]$_DFFE_PN0P_  (.D(_063_),
    .Q(net199),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[31]$_DFFE_PN0P_  (.D(_064_),
    .Q(net200),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[3]$_DFFE_PN0P_  (.D(_065_),
    .Q(net201),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[4]$_DFFE_PN0P_  (.D(_066_),
    .Q(net202),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[5]$_DFFE_PN0P_  (.D(_067_),
    .Q(net203),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[6]$_DFFE_PN0P_  (.D(_068_),
    .Q(net204),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[7]$_DFFE_PN0P_  (.D(_069_),
    .Q(net205),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[8]$_DFFE_PN0P_  (.D(_070_),
    .Q(net206),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_adr_o[9]$_DFFE_PN0P_  (.D(_071_),
    .Q(net207),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_cyc_o$_DFF_PN0_  (.D(_270_),
    .Q(net208),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[0]$_DFFE_PN0P_  (.D(_072_),
    .Q(net209),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[10]$_DFFE_PN0P_  (.D(_073_),
    .Q(net210),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[11]$_DFFE_PN0P_  (.D(_074_),
    .Q(net211),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[12]$_DFFE_PN0P_  (.D(_075_),
    .Q(net212),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[13]$_DFFE_PN0P_  (.D(_076_),
    .Q(net213),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[14]$_DFFE_PN0P_  (.D(_077_),
    .Q(net214),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[15]$_DFFE_PN0P_  (.D(_078_),
    .Q(net215),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[16]$_DFFE_PN0P_  (.D(_079_),
    .Q(net216),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[17]$_DFFE_PN0P_  (.D(_080_),
    .Q(net217),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[18]$_DFFE_PN0P_  (.D(_081_),
    .Q(net218),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[19]$_DFFE_PN0P_  (.D(_082_),
    .Q(net219),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[1]$_DFFE_PN0P_  (.D(_083_),
    .Q(net220),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[20]$_DFFE_PN0P_  (.D(_084_),
    .Q(net221),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[21]$_DFFE_PN0P_  (.D(_085_),
    .Q(net222),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[22]$_DFFE_PN0P_  (.D(_086_),
    .Q(net223),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[23]$_DFFE_PN0P_  (.D(_087_),
    .Q(net224),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[24]$_DFFE_PN0P_  (.D(_088_),
    .Q(net225),
    .RESET_B(net1),
    .CLK(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[25]$_DFFE_PN0P_  (.D(_089_),
    .Q(net226),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[26]$_DFFE_PN0P_  (.D(_090_),
    .Q(net227),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[27]$_DFFE_PN0P_  (.D(_091_),
    .Q(net228),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[28]$_DFFE_PN0P_  (.D(_092_),
    .Q(net229),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[29]$_DFFE_PN0P_  (.D(_093_),
    .Q(net230),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[2]$_DFFE_PN0P_  (.D(_094_),
    .Q(net231),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[30]$_DFFE_PN0P_  (.D(_095_),
    .Q(net232),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[31]$_DFFE_PN0P_  (.D(_096_),
    .Q(net233),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[3]$_DFFE_PN0P_  (.D(_097_),
    .Q(net234),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[4]$_DFFE_PN0P_  (.D(_098_),
    .Q(net235),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[5]$_DFFE_PN0P_  (.D(_099_),
    .Q(net236),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[6]$_DFFE_PN0P_  (.D(_100_),
    .Q(net237),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[7]$_DFFE_PN0P_  (.D(_101_),
    .Q(net238),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[8]$_DFFE_PN0P_  (.D(_102_),
    .Q(net239),
    .RESET_B(net1),
    .CLK(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_dat_o[9]$_DFFE_PN0P_  (.D(_103_),
    .Q(net240),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_sel_o[0]$_DFFE_PN0P_  (.D(_104_),
    .Q(net241),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_sel_o[1]$_DFFE_PN0P_  (.D(_105_),
    .Q(net242),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_sel_o[2]$_DFFE_PN0P_  (.D(_106_),
    .Q(net243),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_sel_o[3]$_DFFE_PN0P_  (.D(_107_),
    .Q(net244),
    .RESET_B(net1),
    .CLK(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \wb_we_o$_DFFE_PN0P_  (.D(_108_),
    .Q(net246),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \write_done$_DFFE_PN0P_  (.D(_109_),
    .Q(net247),
    .RESET_B(net1),
    .CLK(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \write_err$_DFFE_PN0P_  (.D(_110_),
    .Q(net248),
    .RESET_B(net1),
    .CLK(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__buf_16 hold1 (.A(net250),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_107 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(read_addr[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(read_addr[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(read_addr[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(read_addr[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(read_addr[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(read_addr[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(read_addr[15]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(read_addr[16]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(read_addr[17]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(read_addr[18]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(read_addr[19]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(read_addr[1]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(read_addr[20]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(read_addr[21]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(read_addr[22]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(read_addr[23]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(read_addr[24]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(read_addr[25]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(read_addr[26]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(read_addr[27]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(read_addr[28]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(read_addr[29]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(read_addr[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(read_addr[30]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(read_addr[31]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(read_addr[3]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(read_addr[4]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(read_addr[5]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(read_addr[6]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(read_addr[7]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(read_addr[8]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(read_addr[9]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(read_req),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(read_sel[0]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(read_sel[1]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(read_sel[2]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(read_sel[3]),
    .X(net38));
 sky130_fd_sc_hd__buf_2 input38 (.A(wb_ack_i),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(wb_dat_i[0]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(wb_dat_i[10]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(wb_dat_i[11]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(wb_dat_i[12]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(wb_dat_i[13]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(wb_dat_i[14]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(wb_dat_i[15]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(wb_dat_i[16]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(wb_dat_i[17]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(wb_dat_i[18]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(wb_dat_i[19]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(wb_dat_i[1]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(wb_dat_i[20]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(wb_dat_i[21]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(wb_dat_i[22]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(wb_dat_i[23]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(wb_dat_i[24]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(wb_dat_i[25]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(wb_dat_i[26]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(wb_dat_i[27]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(wb_dat_i[28]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(wb_dat_i[29]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(wb_dat_i[2]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(wb_dat_i[30]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(wb_dat_i[31]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(wb_dat_i[3]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(wb_dat_i[4]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(wb_dat_i[5]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(wb_dat_i[6]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(wb_dat_i[7]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(wb_dat_i[8]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(wb_dat_i[9]),
    .X(net71));
 sky130_fd_sc_hd__dlymetal6s2s_1 input71 (.A(wb_err_i),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(wb_rty_i),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(write_addr[0]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(write_addr[10]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(write_addr[11]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(write_addr[12]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(write_addr[13]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(write_addr[14]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(write_addr[15]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(write_addr[16]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(write_addr[17]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(write_addr[18]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(write_addr[19]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(write_addr[1]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(write_addr[20]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(write_addr[21]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(write_addr[22]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(write_addr[23]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(write_addr[24]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(write_addr[25]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(write_addr[26]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(write_addr[27]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(write_addr[28]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(write_addr[29]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(write_addr[2]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(write_addr[30]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(write_addr[31]),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 input98 (.A(write_addr[3]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 input99 (.A(write_addr[4]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(write_addr[5]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input101 (.A(write_addr[6]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(write_addr[7]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 input103 (.A(write_addr[8]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input104 (.A(write_addr[9]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(write_data[0]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(write_data[10]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_1 input107 (.A(write_data[11]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 input108 (.A(write_data[12]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 input109 (.A(write_data[13]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_1 input110 (.A(write_data[14]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 input111 (.A(write_data[15]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_1 input112 (.A(write_data[16]),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_1 input113 (.A(write_data[17]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_1 input114 (.A(write_data[18]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_1 input115 (.A(write_data[19]),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_1 input116 (.A(write_data[1]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_1 input117 (.A(write_data[20]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 input118 (.A(write_data[21]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_1 input119 (.A(write_data[22]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_1 input120 (.A(write_data[23]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input121 (.A(write_data[24]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(write_data[25]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(write_data[26]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(write_data[27]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input125 (.A(write_data[28]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(write_data[29]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(write_data[2]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 input128 (.A(write_data[30]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 input129 (.A(write_data[31]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 input130 (.A(write_data[3]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input131 (.A(write_data[4]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(write_data[5]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 input133 (.A(write_data[6]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 input134 (.A(write_data[7]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 input135 (.A(write_data[8]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 input136 (.A(write_data[9]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 input137 (.A(write_sel[0]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 input138 (.A(write_sel[1]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 input139 (.A(write_sel[2]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 input140 (.A(write_sel[3]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 output141 (.A(net142),
    .X(read_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output142 (.A(net143),
    .X(read_data[10]));
 sky130_fd_sc_hd__clkbuf_1 output143 (.A(net144),
    .X(read_data[11]));
 sky130_fd_sc_hd__clkbuf_1 output144 (.A(net145),
    .X(read_data[12]));
 sky130_fd_sc_hd__clkbuf_1 output145 (.A(net146),
    .X(read_data[13]));
 sky130_fd_sc_hd__clkbuf_1 output146 (.A(net147),
    .X(read_data[14]));
 sky130_fd_sc_hd__clkbuf_1 output147 (.A(net148),
    .X(read_data[15]));
 sky130_fd_sc_hd__clkbuf_1 output148 (.A(net149),
    .X(read_data[16]));
 sky130_fd_sc_hd__clkbuf_1 output149 (.A(net150),
    .X(read_data[17]));
 sky130_fd_sc_hd__clkbuf_1 output150 (.A(net151),
    .X(read_data[18]));
 sky130_fd_sc_hd__clkbuf_1 output151 (.A(net152),
    .X(read_data[19]));
 sky130_fd_sc_hd__clkbuf_1 output152 (.A(net153),
    .X(read_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output153 (.A(net154),
    .X(read_data[20]));
 sky130_fd_sc_hd__clkbuf_1 output154 (.A(net155),
    .X(read_data[21]));
 sky130_fd_sc_hd__clkbuf_1 output155 (.A(net156),
    .X(read_data[22]));
 sky130_fd_sc_hd__clkbuf_1 output156 (.A(net157),
    .X(read_data[23]));
 sky130_fd_sc_hd__clkbuf_1 output157 (.A(net158),
    .X(read_data[24]));
 sky130_fd_sc_hd__clkbuf_1 output158 (.A(net159),
    .X(read_data[25]));
 sky130_fd_sc_hd__clkbuf_1 output159 (.A(net160),
    .X(read_data[26]));
 sky130_fd_sc_hd__clkbuf_1 output160 (.A(net161),
    .X(read_data[27]));
 sky130_fd_sc_hd__clkbuf_1 output161 (.A(net162),
    .X(read_data[28]));
 sky130_fd_sc_hd__clkbuf_1 output162 (.A(net163),
    .X(read_data[29]));
 sky130_fd_sc_hd__clkbuf_1 output163 (.A(net164),
    .X(read_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output164 (.A(net165),
    .X(read_data[30]));
 sky130_fd_sc_hd__clkbuf_1 output165 (.A(net166),
    .X(read_data[31]));
 sky130_fd_sc_hd__clkbuf_1 output166 (.A(net167),
    .X(read_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output167 (.A(net168),
    .X(read_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output168 (.A(net169),
    .X(read_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output169 (.A(net170),
    .X(read_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output170 (.A(net171),
    .X(read_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output171 (.A(net172),
    .X(read_data[8]));
 sky130_fd_sc_hd__clkbuf_1 output172 (.A(net173),
    .X(read_data[9]));
 sky130_fd_sc_hd__clkbuf_1 output173 (.A(net174),
    .X(read_done));
 sky130_fd_sc_hd__clkbuf_1 output174 (.A(net175),
    .X(read_err));
 sky130_fd_sc_hd__clkbuf_1 output175 (.A(net176),
    .X(wb_adr_o[0]));
 sky130_fd_sc_hd__clkbuf_1 output176 (.A(net177),
    .X(wb_adr_o[10]));
 sky130_fd_sc_hd__clkbuf_1 output177 (.A(net178),
    .X(wb_adr_o[11]));
 sky130_fd_sc_hd__clkbuf_1 output178 (.A(net179),
    .X(wb_adr_o[12]));
 sky130_fd_sc_hd__clkbuf_1 output179 (.A(net180),
    .X(wb_adr_o[13]));
 sky130_fd_sc_hd__clkbuf_1 output180 (.A(net181),
    .X(wb_adr_o[14]));
 sky130_fd_sc_hd__clkbuf_1 output181 (.A(net182),
    .X(wb_adr_o[15]));
 sky130_fd_sc_hd__clkbuf_1 output182 (.A(net183),
    .X(wb_adr_o[16]));
 sky130_fd_sc_hd__clkbuf_1 output183 (.A(net184),
    .X(wb_adr_o[17]));
 sky130_fd_sc_hd__clkbuf_1 output184 (.A(net185),
    .X(wb_adr_o[18]));
 sky130_fd_sc_hd__clkbuf_1 output185 (.A(net186),
    .X(wb_adr_o[19]));
 sky130_fd_sc_hd__clkbuf_1 output186 (.A(net187),
    .X(wb_adr_o[1]));
 sky130_fd_sc_hd__clkbuf_1 output187 (.A(net188),
    .X(wb_adr_o[20]));
 sky130_fd_sc_hd__clkbuf_1 output188 (.A(net189),
    .X(wb_adr_o[21]));
 sky130_fd_sc_hd__clkbuf_1 output189 (.A(net190),
    .X(wb_adr_o[22]));
 sky130_fd_sc_hd__clkbuf_1 output190 (.A(net191),
    .X(wb_adr_o[23]));
 sky130_fd_sc_hd__clkbuf_1 output191 (.A(net192),
    .X(wb_adr_o[24]));
 sky130_fd_sc_hd__clkbuf_1 output192 (.A(net193),
    .X(wb_adr_o[25]));
 sky130_fd_sc_hd__clkbuf_1 output193 (.A(net194),
    .X(wb_adr_o[26]));
 sky130_fd_sc_hd__clkbuf_1 output194 (.A(net195),
    .X(wb_adr_o[27]));
 sky130_fd_sc_hd__clkbuf_1 output195 (.A(net196),
    .X(wb_adr_o[28]));
 sky130_fd_sc_hd__clkbuf_1 output196 (.A(net197),
    .X(wb_adr_o[29]));
 sky130_fd_sc_hd__clkbuf_1 output197 (.A(net198),
    .X(wb_adr_o[2]));
 sky130_fd_sc_hd__clkbuf_1 output198 (.A(net199),
    .X(wb_adr_o[30]));
 sky130_fd_sc_hd__clkbuf_1 output199 (.A(net200),
    .X(wb_adr_o[31]));
 sky130_fd_sc_hd__clkbuf_1 output200 (.A(net201),
    .X(wb_adr_o[3]));
 sky130_fd_sc_hd__clkbuf_1 output201 (.A(net202),
    .X(wb_adr_o[4]));
 sky130_fd_sc_hd__clkbuf_1 output202 (.A(net203),
    .X(wb_adr_o[5]));
 sky130_fd_sc_hd__clkbuf_1 output203 (.A(net204),
    .X(wb_adr_o[6]));
 sky130_fd_sc_hd__clkbuf_1 output204 (.A(net205),
    .X(wb_adr_o[7]));
 sky130_fd_sc_hd__clkbuf_1 output205 (.A(net206),
    .X(wb_adr_o[8]));
 sky130_fd_sc_hd__clkbuf_1 output206 (.A(net207),
    .X(wb_adr_o[9]));
 sky130_fd_sc_hd__clkbuf_1 output207 (.A(net208),
    .X(wb_cyc_o));
 sky130_fd_sc_hd__clkbuf_1 output208 (.A(net209),
    .X(wb_dat_o[0]));
 sky130_fd_sc_hd__clkbuf_1 output209 (.A(net210),
    .X(wb_dat_o[10]));
 sky130_fd_sc_hd__clkbuf_1 output210 (.A(net211),
    .X(wb_dat_o[11]));
 sky130_fd_sc_hd__clkbuf_1 output211 (.A(net212),
    .X(wb_dat_o[12]));
 sky130_fd_sc_hd__clkbuf_1 output212 (.A(net213),
    .X(wb_dat_o[13]));
 sky130_fd_sc_hd__clkbuf_1 output213 (.A(net214),
    .X(wb_dat_o[14]));
 sky130_fd_sc_hd__clkbuf_1 output214 (.A(net215),
    .X(wb_dat_o[15]));
 sky130_fd_sc_hd__clkbuf_1 output215 (.A(net216),
    .X(wb_dat_o[16]));
 sky130_fd_sc_hd__clkbuf_1 output216 (.A(net217),
    .X(wb_dat_o[17]));
 sky130_fd_sc_hd__clkbuf_1 output217 (.A(net218),
    .X(wb_dat_o[18]));
 sky130_fd_sc_hd__clkbuf_1 output218 (.A(net219),
    .X(wb_dat_o[19]));
 sky130_fd_sc_hd__clkbuf_1 output219 (.A(net220),
    .X(wb_dat_o[1]));
 sky130_fd_sc_hd__clkbuf_1 output220 (.A(net221),
    .X(wb_dat_o[20]));
 sky130_fd_sc_hd__clkbuf_1 output221 (.A(net222),
    .X(wb_dat_o[21]));
 sky130_fd_sc_hd__clkbuf_1 output222 (.A(net223),
    .X(wb_dat_o[22]));
 sky130_fd_sc_hd__clkbuf_1 output223 (.A(net224),
    .X(wb_dat_o[23]));
 sky130_fd_sc_hd__clkbuf_1 output224 (.A(net225),
    .X(wb_dat_o[24]));
 sky130_fd_sc_hd__clkbuf_1 output225 (.A(net226),
    .X(wb_dat_o[25]));
 sky130_fd_sc_hd__clkbuf_1 output226 (.A(net227),
    .X(wb_dat_o[26]));
 sky130_fd_sc_hd__clkbuf_1 output227 (.A(net228),
    .X(wb_dat_o[27]));
 sky130_fd_sc_hd__clkbuf_1 output228 (.A(net229),
    .X(wb_dat_o[28]));
 sky130_fd_sc_hd__clkbuf_1 output229 (.A(net230),
    .X(wb_dat_o[29]));
 sky130_fd_sc_hd__clkbuf_1 output230 (.A(net231),
    .X(wb_dat_o[2]));
 sky130_fd_sc_hd__clkbuf_1 output231 (.A(net232),
    .X(wb_dat_o[30]));
 sky130_fd_sc_hd__clkbuf_1 output232 (.A(net233),
    .X(wb_dat_o[31]));
 sky130_fd_sc_hd__clkbuf_1 output233 (.A(net234),
    .X(wb_dat_o[3]));
 sky130_fd_sc_hd__clkbuf_1 output234 (.A(net235),
    .X(wb_dat_o[4]));
 sky130_fd_sc_hd__clkbuf_1 output235 (.A(net236),
    .X(wb_dat_o[5]));
 sky130_fd_sc_hd__clkbuf_1 output236 (.A(net237),
    .X(wb_dat_o[6]));
 sky130_fd_sc_hd__clkbuf_1 output237 (.A(net238),
    .X(wb_dat_o[7]));
 sky130_fd_sc_hd__clkbuf_1 output238 (.A(net239),
    .X(wb_dat_o[8]));
 sky130_fd_sc_hd__clkbuf_1 output239 (.A(net240),
    .X(wb_dat_o[9]));
 sky130_fd_sc_hd__clkbuf_1 output240 (.A(net241),
    .X(wb_sel_o[0]));
 sky130_fd_sc_hd__clkbuf_1 output241 (.A(net242),
    .X(wb_sel_o[1]));
 sky130_fd_sc_hd__clkbuf_1 output242 (.A(net243),
    .X(wb_sel_o[2]));
 sky130_fd_sc_hd__clkbuf_1 output243 (.A(net244),
    .X(wb_sel_o[3]));
 sky130_fd_sc_hd__clkbuf_1 output244 (.A(net245),
    .X(wb_stb_o));
 sky130_fd_sc_hd__clkbuf_1 output245 (.A(net246),
    .X(wb_we_o));
 sky130_fd_sc_hd__clkbuf_1 output246 (.A(net247),
    .X(write_done));
 sky130_fd_sc_hd__clkbuf_1 output247 (.A(net248),
    .X(write_err));
 sky130_fd_sc_hd__conb_1 _536__248 (.LO(net249));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__bufinv_16 clkload0 (.A(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload1 (.A(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload2 (.A(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload3 (.A(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload4 (.A(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload5 (.A(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload6 (.A(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net250));
 sky130_fd_sc_hd__fill_1 FILLER_0_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_102 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_94 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_126 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_14 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_188 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_128 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_173 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_203 ();
endmodule
