module bidirectional_fifo (a_almost_empty,
    a_almost_full,
    a_empty,
    a_full,
    a_rd_en,
    a_wr_en,
    b_almost_empty,
    b_almost_full,
    b_empty,
    b_full,
    b_rd_en,
    b_wr_en,
    clk,
    rst_n,
    a_rd_data,
    a_to_b_count,
    a_wr_data,
    b_rd_data,
    b_to_a_count,
    b_wr_data);
 output a_almost_empty;
 output a_almost_full;
 output a_empty;
 output a_full;
 input a_rd_en;
 input a_wr_en;
 output b_almost_empty;
 output b_almost_full;
 output b_empty;
 output b_full;
 input b_rd_en;
 input b_wr_en;
 input clk;
 input rst_n;
 output [7:0] a_rd_data;
 output [4:0] a_to_b_count;
 input [7:0] a_wr_data;
 output [7:0] b_rd_data;
 output [4:0] b_to_a_count;
 input [7:0] b_wr_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire net42;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire net40;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire \a_rd_ptr[0] ;
 wire \a_rd_ptr[1] ;
 wire \a_rd_ptr[2] ;
 wire \a_rd_ptr[3] ;
 wire \a_rd_ptr[4] ;
 wire \a_to_b_mem[0][0] ;
 wire \a_to_b_mem[0][1] ;
 wire \a_to_b_mem[0][2] ;
 wire \a_to_b_mem[0][3] ;
 wire \a_to_b_mem[0][4] ;
 wire \a_to_b_mem[0][5] ;
 wire \a_to_b_mem[0][6] ;
 wire \a_to_b_mem[0][7] ;
 wire \a_to_b_mem[10][0] ;
 wire \a_to_b_mem[10][1] ;
 wire \a_to_b_mem[10][2] ;
 wire \a_to_b_mem[10][3] ;
 wire \a_to_b_mem[10][4] ;
 wire \a_to_b_mem[10][5] ;
 wire \a_to_b_mem[10][6] ;
 wire \a_to_b_mem[10][7] ;
 wire \a_to_b_mem[11][0] ;
 wire \a_to_b_mem[11][1] ;
 wire \a_to_b_mem[11][2] ;
 wire \a_to_b_mem[11][3] ;
 wire \a_to_b_mem[11][4] ;
 wire \a_to_b_mem[11][5] ;
 wire \a_to_b_mem[11][6] ;
 wire \a_to_b_mem[11][7] ;
 wire \a_to_b_mem[12][0] ;
 wire \a_to_b_mem[12][1] ;
 wire \a_to_b_mem[12][2] ;
 wire \a_to_b_mem[12][3] ;
 wire \a_to_b_mem[12][4] ;
 wire \a_to_b_mem[12][5] ;
 wire \a_to_b_mem[12][6] ;
 wire \a_to_b_mem[12][7] ;
 wire \a_to_b_mem[13][0] ;
 wire \a_to_b_mem[13][1] ;
 wire \a_to_b_mem[13][2] ;
 wire \a_to_b_mem[13][3] ;
 wire \a_to_b_mem[13][4] ;
 wire \a_to_b_mem[13][5] ;
 wire \a_to_b_mem[13][6] ;
 wire \a_to_b_mem[13][7] ;
 wire \a_to_b_mem[14][0] ;
 wire \a_to_b_mem[14][1] ;
 wire \a_to_b_mem[14][2] ;
 wire \a_to_b_mem[14][3] ;
 wire \a_to_b_mem[14][4] ;
 wire \a_to_b_mem[14][5] ;
 wire \a_to_b_mem[14][6] ;
 wire \a_to_b_mem[14][7] ;
 wire \a_to_b_mem[15][0] ;
 wire \a_to_b_mem[15][1] ;
 wire \a_to_b_mem[15][2] ;
 wire \a_to_b_mem[15][3] ;
 wire \a_to_b_mem[15][4] ;
 wire \a_to_b_mem[15][5] ;
 wire \a_to_b_mem[15][6] ;
 wire \a_to_b_mem[15][7] ;
 wire \a_to_b_mem[1][0] ;
 wire \a_to_b_mem[1][1] ;
 wire \a_to_b_mem[1][2] ;
 wire \a_to_b_mem[1][3] ;
 wire \a_to_b_mem[1][4] ;
 wire \a_to_b_mem[1][5] ;
 wire \a_to_b_mem[1][6] ;
 wire \a_to_b_mem[1][7] ;
 wire \a_to_b_mem[2][0] ;
 wire \a_to_b_mem[2][1] ;
 wire \a_to_b_mem[2][2] ;
 wire \a_to_b_mem[2][3] ;
 wire \a_to_b_mem[2][4] ;
 wire \a_to_b_mem[2][5] ;
 wire \a_to_b_mem[2][6] ;
 wire \a_to_b_mem[2][7] ;
 wire \a_to_b_mem[3][0] ;
 wire \a_to_b_mem[3][1] ;
 wire \a_to_b_mem[3][2] ;
 wire \a_to_b_mem[3][3] ;
 wire \a_to_b_mem[3][4] ;
 wire \a_to_b_mem[3][5] ;
 wire \a_to_b_mem[3][6] ;
 wire \a_to_b_mem[3][7] ;
 wire \a_to_b_mem[4][0] ;
 wire \a_to_b_mem[4][1] ;
 wire \a_to_b_mem[4][2] ;
 wire \a_to_b_mem[4][3] ;
 wire \a_to_b_mem[4][4] ;
 wire \a_to_b_mem[4][5] ;
 wire \a_to_b_mem[4][6] ;
 wire \a_to_b_mem[4][7] ;
 wire \a_to_b_mem[5][0] ;
 wire \a_to_b_mem[5][1] ;
 wire \a_to_b_mem[5][2] ;
 wire \a_to_b_mem[5][3] ;
 wire \a_to_b_mem[5][4] ;
 wire \a_to_b_mem[5][5] ;
 wire \a_to_b_mem[5][6] ;
 wire \a_to_b_mem[5][7] ;
 wire \a_to_b_mem[6][0] ;
 wire \a_to_b_mem[6][1] ;
 wire \a_to_b_mem[6][2] ;
 wire \a_to_b_mem[6][3] ;
 wire \a_to_b_mem[6][4] ;
 wire \a_to_b_mem[6][5] ;
 wire \a_to_b_mem[6][6] ;
 wire \a_to_b_mem[6][7] ;
 wire \a_to_b_mem[7][0] ;
 wire \a_to_b_mem[7][1] ;
 wire \a_to_b_mem[7][2] ;
 wire \a_to_b_mem[7][3] ;
 wire \a_to_b_mem[7][4] ;
 wire \a_to_b_mem[7][5] ;
 wire \a_to_b_mem[7][6] ;
 wire \a_to_b_mem[7][7] ;
 wire \a_to_b_mem[8][0] ;
 wire \a_to_b_mem[8][1] ;
 wire \a_to_b_mem[8][2] ;
 wire \a_to_b_mem[8][3] ;
 wire \a_to_b_mem[8][4] ;
 wire \a_to_b_mem[8][5] ;
 wire \a_to_b_mem[8][6] ;
 wire \a_to_b_mem[8][7] ;
 wire \a_to_b_mem[9][0] ;
 wire \a_to_b_mem[9][1] ;
 wire \a_to_b_mem[9][2] ;
 wire \a_to_b_mem[9][3] ;
 wire \a_to_b_mem[9][4] ;
 wire \a_to_b_mem[9][5] ;
 wire \a_to_b_mem[9][6] ;
 wire \a_to_b_mem[9][7] ;
 wire \a_wr_ptr[0] ;
 wire \a_wr_ptr[1] ;
 wire \a_wr_ptr[2] ;
 wire \a_wr_ptr[3] ;
 wire \a_wr_ptr[4] ;
 wire \b_rd_ptr[0] ;
 wire \b_rd_ptr[1] ;
 wire \b_rd_ptr[2] ;
 wire \b_rd_ptr[3] ;
 wire \b_rd_ptr[4] ;
 wire \b_to_a_mem[0][0] ;
 wire \b_to_a_mem[0][1] ;
 wire \b_to_a_mem[0][2] ;
 wire \b_to_a_mem[0][3] ;
 wire \b_to_a_mem[0][4] ;
 wire \b_to_a_mem[0][5] ;
 wire \b_to_a_mem[0][6] ;
 wire \b_to_a_mem[0][7] ;
 wire \b_to_a_mem[10][0] ;
 wire \b_to_a_mem[10][1] ;
 wire \b_to_a_mem[10][2] ;
 wire \b_to_a_mem[10][3] ;
 wire \b_to_a_mem[10][4] ;
 wire \b_to_a_mem[10][5] ;
 wire \b_to_a_mem[10][6] ;
 wire \b_to_a_mem[10][7] ;
 wire \b_to_a_mem[11][0] ;
 wire \b_to_a_mem[11][1] ;
 wire \b_to_a_mem[11][2] ;
 wire \b_to_a_mem[11][3] ;
 wire \b_to_a_mem[11][4] ;
 wire \b_to_a_mem[11][5] ;
 wire \b_to_a_mem[11][6] ;
 wire \b_to_a_mem[11][7] ;
 wire \b_to_a_mem[12][0] ;
 wire \b_to_a_mem[12][1] ;
 wire \b_to_a_mem[12][2] ;
 wire \b_to_a_mem[12][3] ;
 wire \b_to_a_mem[12][4] ;
 wire \b_to_a_mem[12][5] ;
 wire \b_to_a_mem[12][6] ;
 wire \b_to_a_mem[12][7] ;
 wire \b_to_a_mem[13][0] ;
 wire \b_to_a_mem[13][1] ;
 wire \b_to_a_mem[13][2] ;
 wire \b_to_a_mem[13][3] ;
 wire \b_to_a_mem[13][4] ;
 wire \b_to_a_mem[13][5] ;
 wire \b_to_a_mem[13][6] ;
 wire \b_to_a_mem[13][7] ;
 wire \b_to_a_mem[14][0] ;
 wire \b_to_a_mem[14][1] ;
 wire \b_to_a_mem[14][2] ;
 wire \b_to_a_mem[14][3] ;
 wire \b_to_a_mem[14][4] ;
 wire \b_to_a_mem[14][5] ;
 wire \b_to_a_mem[14][6] ;
 wire \b_to_a_mem[14][7] ;
 wire \b_to_a_mem[15][0] ;
 wire \b_to_a_mem[15][1] ;
 wire \b_to_a_mem[15][2] ;
 wire \b_to_a_mem[15][3] ;
 wire \b_to_a_mem[15][4] ;
 wire \b_to_a_mem[15][5] ;
 wire \b_to_a_mem[15][6] ;
 wire \b_to_a_mem[15][7] ;
 wire \b_to_a_mem[1][0] ;
 wire \b_to_a_mem[1][1] ;
 wire \b_to_a_mem[1][2] ;
 wire \b_to_a_mem[1][3] ;
 wire \b_to_a_mem[1][4] ;
 wire \b_to_a_mem[1][5] ;
 wire \b_to_a_mem[1][6] ;
 wire \b_to_a_mem[1][7] ;
 wire \b_to_a_mem[2][0] ;
 wire \b_to_a_mem[2][1] ;
 wire \b_to_a_mem[2][2] ;
 wire \b_to_a_mem[2][3] ;
 wire \b_to_a_mem[2][4] ;
 wire \b_to_a_mem[2][5] ;
 wire \b_to_a_mem[2][6] ;
 wire \b_to_a_mem[2][7] ;
 wire \b_to_a_mem[3][0] ;
 wire \b_to_a_mem[3][1] ;
 wire \b_to_a_mem[3][2] ;
 wire \b_to_a_mem[3][3] ;
 wire \b_to_a_mem[3][4] ;
 wire \b_to_a_mem[3][5] ;
 wire \b_to_a_mem[3][6] ;
 wire \b_to_a_mem[3][7] ;
 wire \b_to_a_mem[4][0] ;
 wire \b_to_a_mem[4][1] ;
 wire \b_to_a_mem[4][2] ;
 wire \b_to_a_mem[4][3] ;
 wire \b_to_a_mem[4][4] ;
 wire \b_to_a_mem[4][5] ;
 wire \b_to_a_mem[4][6] ;
 wire \b_to_a_mem[4][7] ;
 wire \b_to_a_mem[5][0] ;
 wire \b_to_a_mem[5][1] ;
 wire \b_to_a_mem[5][2] ;
 wire \b_to_a_mem[5][3] ;
 wire \b_to_a_mem[5][4] ;
 wire \b_to_a_mem[5][5] ;
 wire \b_to_a_mem[5][6] ;
 wire \b_to_a_mem[5][7] ;
 wire \b_to_a_mem[6][0] ;
 wire \b_to_a_mem[6][1] ;
 wire \b_to_a_mem[6][2] ;
 wire \b_to_a_mem[6][3] ;
 wire \b_to_a_mem[6][4] ;
 wire \b_to_a_mem[6][5] ;
 wire \b_to_a_mem[6][6] ;
 wire \b_to_a_mem[6][7] ;
 wire \b_to_a_mem[7][0] ;
 wire \b_to_a_mem[7][1] ;
 wire \b_to_a_mem[7][2] ;
 wire \b_to_a_mem[7][3] ;
 wire \b_to_a_mem[7][4] ;
 wire \b_to_a_mem[7][5] ;
 wire \b_to_a_mem[7][6] ;
 wire \b_to_a_mem[7][7] ;
 wire \b_to_a_mem[8][0] ;
 wire \b_to_a_mem[8][1] ;
 wire \b_to_a_mem[8][2] ;
 wire \b_to_a_mem[8][3] ;
 wire \b_to_a_mem[8][4] ;
 wire \b_to_a_mem[8][5] ;
 wire \b_to_a_mem[8][6] ;
 wire \b_to_a_mem[8][7] ;
 wire \b_to_a_mem[9][0] ;
 wire \b_to_a_mem[9][1] ;
 wire \b_to_a_mem[9][2] ;
 wire \b_to_a_mem[9][3] ;
 wire \b_to_a_mem[9][4] ;
 wire \b_to_a_mem[9][5] ;
 wire \b_to_a_mem[9][6] ;
 wire \b_to_a_mem[9][7] ;
 wire \b_wr_ptr[0] ;
 wire \b_wr_ptr[1] ;
 wire \b_wr_ptr[2] ;
 wire \b_wr_ptr[3] ;
 wire \b_wr_ptr[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net41;
 wire net43;

 BUF_X2 _1257_ (.A(_1226_),
    .Z(_0787_));
 AND2_X1 _1258_ (.A1(_1231_),
    .A2(_1228_),
    .ZN(_0788_));
 INV_X1 _1259_ (.A(_1253_),
    .ZN(_1214_));
 AOI221_X2 _1260_ (.A(_1230_),
    .B1(_0788_),
    .B2(_1214_),
    .C1(_1227_),
    .C2(_1231_),
    .ZN(_0789_));
 XOR2_X2 _1261_ (.A(_0787_),
    .B(_0789_),
    .Z(_0790_));
 INV_X4 _1262_ (.A(_0790_),
    .ZN(net16));
 AND2_X1 _1263_ (.A1(_0787_),
    .A2(_1231_),
    .ZN(_0791_));
 AOI221_X2 _1264_ (.A(_1225_),
    .B1(_1230_),
    .B2(_0787_),
    .C1(_1215_),
    .C2(_0791_),
    .ZN(_0792_));
 XNOR2_X2 _1265_ (.A(\a_wr_ptr[4] ),
    .B(\b_rd_ptr[4] ),
    .ZN(_0793_));
 XOR2_X2 _1266_ (.A(_0792_),
    .B(_0793_),
    .Z(_0794_));
 INV_X8 _1267_ (.A(_0794_),
    .ZN(_0795_));
 INV_X4 clone1 (.A(net43),
    .ZN(net42));
 FILLCELL_X32 FILLER_0_1 ();
 INV_X4 _1270_ (.A(_1254_),
    .ZN(net13));
 XNOR2_X2 _1271_ (.A(_1215_),
    .B(_1231_),
    .ZN(_0797_));
 INV_X4 _1272_ (.A(_0797_),
    .ZN(net15));
 INV_X4 _1273_ (.A(_1256_),
    .ZN(net30));
 XNOR2_X2 _1274_ (.A(_1218_),
    .B(_1234_),
    .ZN(_0798_));
 INV_X4 _1275_ (.A(_0798_),
    .ZN(net32));
 BUF_X2 _1276_ (.A(_1221_),
    .Z(_0799_));
 AND2_X1 _1277_ (.A1(_1234_),
    .A2(_1223_),
    .ZN(_0800_));
 INV_X1 _1278_ (.A(_1255_),
    .ZN(_1217_));
 AOI221_X2 _1279_ (.A(_1233_),
    .B1(_0800_),
    .B2(_1217_),
    .C1(_1222_),
    .C2(_1234_),
    .ZN(_0801_));
 XOR2_X2 _1280_ (.A(_0799_),
    .B(_0801_),
    .Z(_0802_));
 INV_X4 _1281_ (.A(_0802_),
    .ZN(net33));
 AND2_X1 _1282_ (.A1(_0799_),
    .A2(_1234_),
    .ZN(_0803_));
 AOI221_X2 _1283_ (.A(_1220_),
    .B1(_1233_),
    .B2(_0799_),
    .C1(net38),
    .C2(_0803_),
    .ZN(_0804_));
 XNOR2_X1 _1284_ (.A(\b_wr_ptr[4] ),
    .B(\a_rd_ptr[4] ),
    .ZN(_0805_));
 XOR2_X2 _1285_ (.A(_0805_),
    .B(_0804_),
    .Z(_0806_));
 INV_X4 _1286_ (.A(_0806_),
    .ZN(_0807_));
 BUF_X8 _1287_ (.A(_0807_),
    .Z(_0808_));
 BUF_X8 _1288_ (.A(_0808_),
    .Z(net34));
 BUF_X8 _1289_ (.A(net37),
    .Z(_0809_));
 BUF_X8 _1290_ (.A(_0809_),
    .Z(_0810_));
 CLKBUF_X2 _1291_ (.A(net14),
    .Z(_0811_));
 INV_X1 _1292_ (.A(_0811_),
    .ZN(_0812_));
 NAND4_X1 _1293_ (.A1(_0787_),
    .A2(_1254_),
    .A3(_0812_),
    .A4(_0797_),
    .ZN(_0813_));
 OR4_X1 _1294_ (.A1(_0787_),
    .A2(net13),
    .A3(_0811_),
    .A4(net15),
    .ZN(_0814_));
 MUX2_X1 _1295_ (.A(_0813_),
    .B(_0814_),
    .S(_0789_),
    .Z(_0815_));
 BUF_X8 _1296_ (.A(_0815_),
    .Z(_0816_));
 BUF_X8 _1297_ (.A(_0816_),
    .Z(_0817_));
 NOR2_X1 _1298_ (.A1(_0810_),
    .A2(_0817_),
    .ZN(net21));
 BUF_X8 _1299_ (.A(_0806_),
    .Z(_0818_));
 BUF_X4 _1300_ (.A(_0818_),
    .Z(_0819_));
 CLKBUF_X2 _1301_ (.A(net31),
    .Z(_0820_));
 INV_X1 _1302_ (.A(_0820_),
    .ZN(_0821_));
 NAND4_X1 _1303_ (.A1(_0799_),
    .A2(_1256_),
    .A3(_0821_),
    .A4(_0798_),
    .ZN(_0822_));
 OR4_X1 _1304_ (.A1(_0799_),
    .A2(net30),
    .A3(_0820_),
    .A4(net32),
    .ZN(_0823_));
 MUX2_X1 _1305_ (.A(_0822_),
    .B(_0823_),
    .S(_0801_),
    .Z(_0824_));
 BUF_X8 _1306_ (.A(_0824_),
    .Z(_0825_));
 BUF_X1 rebuffer6 (.A(net14),
    .Z(net40));
 NOR2_X4 _1308_ (.A1(_0819_),
    .A2(_0825_),
    .ZN(net4));
 NOR2_X4 _1309_ (.A1(_0825_),
    .A2(net34),
    .ZN(net3));
 NOR2_X1 _1310_ (.A1(_0795_),
    .A2(_0817_),
    .ZN(net20));
 BUF_X1 _1311_ (.A(a_wr_data[0]),
    .Z(_0827_));
 BUF_X2 _1312_ (.A(_0827_),
    .Z(_0828_));
 INV_X4 _1313_ (.A(\a_wr_ptr[2] ),
    .ZN(_0829_));
 BUF_X2 _1314_ (.A(a_wr_en),
    .Z(_0830_));
 INV_X4 _1315_ (.A(_0830_),
    .ZN(_0831_));
 BUF_X4 _1316_ (.A(\a_wr_ptr[3] ),
    .Z(_0832_));
 NOR2_X4 _1317_ (.A1(_0831_),
    .A2(_0832_),
    .ZN(_0833_));
 NAND3_X2 _1318_ (.A1(_0829_),
    .A2(_1246_),
    .A3(_0833_),
    .ZN(_0834_));
 AND4_X1 _1319_ (.A1(_0787_),
    .A2(_1254_),
    .A3(_0812_),
    .A4(_0797_),
    .ZN(_0835_));
 NOR4_X1 _1320_ (.A1(_0787_),
    .A2(net13),
    .A3(_0811_),
    .A4(net15),
    .ZN(_0836_));
 MUX2_X2 _1321_ (.A(_0835_),
    .B(_0836_),
    .S(_0789_),
    .Z(_0837_));
 BUF_X8 _1322_ (.A(_0837_),
    .Z(_0838_));
 AOI21_X4 _1323_ (.A(_0834_),
    .B1(_0838_),
    .B2(_0795_),
    .ZN(_0839_));
 MUX2_X1 _1324_ (.A(\a_to_b_mem[0][0] ),
    .B(_0828_),
    .S(_0839_),
    .Z(_0021_));
 CLKBUF_X2 _1325_ (.A(a_wr_data[1]),
    .Z(_0840_));
 BUF_X2 _1326_ (.A(_0840_),
    .Z(_0841_));
 MUX2_X1 _1327_ (.A(\a_to_b_mem[0][1] ),
    .B(_0841_),
    .S(_0839_),
    .Z(_0022_));
 CLKBUF_X2 _1328_ (.A(a_wr_data[2]),
    .Z(_0842_));
 BUF_X2 _1329_ (.A(_0842_),
    .Z(_0843_));
 MUX2_X1 _1330_ (.A(\a_to_b_mem[0][2] ),
    .B(_0843_),
    .S(_0839_),
    .Z(_0023_));
 CLKBUF_X2 _1331_ (.A(a_wr_data[3]),
    .Z(_0844_));
 BUF_X2 _1332_ (.A(_0844_),
    .Z(_0845_));
 MUX2_X1 _1333_ (.A(\a_to_b_mem[0][3] ),
    .B(_0845_),
    .S(_0839_),
    .Z(_0024_));
 CLKBUF_X2 _1334_ (.A(a_wr_data[4]),
    .Z(_0846_));
 BUF_X2 _1335_ (.A(_0846_),
    .Z(_0847_));
 MUX2_X1 _1336_ (.A(\a_to_b_mem[0][4] ),
    .B(_0847_),
    .S(_0839_),
    .Z(_0025_));
 CLKBUF_X2 _1337_ (.A(a_wr_data[5]),
    .Z(_0848_));
 BUF_X2 _1338_ (.A(_0848_),
    .Z(_0849_));
 MUX2_X1 _1339_ (.A(\a_to_b_mem[0][5] ),
    .B(_0849_),
    .S(_0839_),
    .Z(_0026_));
 CLKBUF_X2 _1340_ (.A(a_wr_data[6]),
    .Z(_0850_));
 BUF_X2 _1341_ (.A(_0850_),
    .Z(_0851_));
 MUX2_X1 _1342_ (.A(\a_to_b_mem[0][6] ),
    .B(_0851_),
    .S(_0839_),
    .Z(_0027_));
 CLKBUF_X2 _1343_ (.A(a_wr_data[7]),
    .Z(_0852_));
 BUF_X2 _1344_ (.A(_0852_),
    .Z(_0853_));
 MUX2_X1 _1345_ (.A(\a_to_b_mem[0][7] ),
    .B(_0853_),
    .S(_0839_),
    .Z(_0028_));
 BUF_X4 _1346_ (.A(\a_wr_ptr[2] ),
    .Z(_0854_));
 INV_X1 _1347_ (.A(_1247_),
    .ZN(_0855_));
 NAND2_X1 _1348_ (.A1(_0830_),
    .A2(_0832_),
    .ZN(_0856_));
 NOR3_X2 _1349_ (.A1(_0854_),
    .A2(_0855_),
    .A3(_0856_),
    .ZN(_0857_));
 OAI21_X4 _1350_ (.A(_0857_),
    .B1(_0816_),
    .B2(_0809_),
    .ZN(_0858_));
 MUX2_X1 _1351_ (.A(_0828_),
    .B(\a_to_b_mem[10][0] ),
    .S(_0858_),
    .Z(_0029_));
 MUX2_X1 _1352_ (.A(_0841_),
    .B(\a_to_b_mem[10][1] ),
    .S(_0858_),
    .Z(_0030_));
 MUX2_X1 _1353_ (.A(_0843_),
    .B(\a_to_b_mem[10][2] ),
    .S(_0858_),
    .Z(_0031_));
 MUX2_X1 _1354_ (.A(_0845_),
    .B(\a_to_b_mem[10][3] ),
    .S(_0858_),
    .Z(_0032_));
 MUX2_X1 _1355_ (.A(_0847_),
    .B(\a_to_b_mem[10][4] ),
    .S(_0858_),
    .Z(_0033_));
 MUX2_X1 _1356_ (.A(_0849_),
    .B(\a_to_b_mem[10][5] ),
    .S(_0858_),
    .Z(_0034_));
 MUX2_X1 _1357_ (.A(_0851_),
    .B(\a_to_b_mem[10][6] ),
    .S(_0858_),
    .Z(_0035_));
 MUX2_X1 _1358_ (.A(_0853_),
    .B(\a_to_b_mem[10][7] ),
    .S(_0858_),
    .Z(_0036_));
 INV_X1 _1359_ (.A(_1251_),
    .ZN(_0859_));
 NOR3_X2 _1360_ (.A1(_0854_),
    .A2(_0859_),
    .A3(_0856_),
    .ZN(_0860_));
 OAI21_X4 _1361_ (.A(_0860_),
    .B1(_0816_),
    .B2(_0809_),
    .ZN(_0861_));
 MUX2_X1 _1362_ (.A(_0828_),
    .B(\a_to_b_mem[11][0] ),
    .S(_0861_),
    .Z(_0037_));
 MUX2_X1 _1363_ (.A(_0841_),
    .B(\a_to_b_mem[11][1] ),
    .S(_0861_),
    .Z(_0038_));
 MUX2_X1 _1364_ (.A(_0843_),
    .B(\a_to_b_mem[11][2] ),
    .S(_0861_),
    .Z(_0039_));
 MUX2_X1 _1365_ (.A(_0845_),
    .B(\a_to_b_mem[11][3] ),
    .S(_0861_),
    .Z(_0040_));
 MUX2_X1 _1366_ (.A(_0847_),
    .B(\a_to_b_mem[11][4] ),
    .S(_0861_),
    .Z(_0041_));
 MUX2_X1 _1367_ (.A(_0849_),
    .B(\a_to_b_mem[11][5] ),
    .S(_0861_),
    .Z(_0042_));
 MUX2_X1 _1368_ (.A(_0851_),
    .B(\a_to_b_mem[11][6] ),
    .S(_0861_),
    .Z(_0043_));
 MUX2_X1 _1369_ (.A(_0853_),
    .B(\a_to_b_mem[11][7] ),
    .S(_0861_),
    .Z(_0044_));
 AND2_X2 _1370_ (.A1(_0830_),
    .A2(_0832_),
    .ZN(_0862_));
 NAND3_X2 _1371_ (.A1(_0854_),
    .A2(_1246_),
    .A3(_0862_),
    .ZN(_0863_));
 AOI21_X4 _1372_ (.A(_0863_),
    .B1(_0838_),
    .B2(_0795_),
    .ZN(_0864_));
 MUX2_X1 _1373_ (.A(\a_to_b_mem[12][0] ),
    .B(_0828_),
    .S(_0864_),
    .Z(_0045_));
 MUX2_X1 _1374_ (.A(\a_to_b_mem[12][1] ),
    .B(_0841_),
    .S(_0864_),
    .Z(_0046_));
 MUX2_X1 _1375_ (.A(\a_to_b_mem[12][2] ),
    .B(_0843_),
    .S(_0864_),
    .Z(_0047_));
 MUX2_X1 _1376_ (.A(\a_to_b_mem[12][3] ),
    .B(_0845_),
    .S(_0864_),
    .Z(_0048_));
 MUX2_X1 _1377_ (.A(\a_to_b_mem[12][4] ),
    .B(_0847_),
    .S(_0864_),
    .Z(_0049_));
 MUX2_X1 _1378_ (.A(\a_to_b_mem[12][5] ),
    .B(_0849_),
    .S(_0864_),
    .Z(_0050_));
 MUX2_X1 _1379_ (.A(\a_to_b_mem[12][6] ),
    .B(_0851_),
    .S(_0864_),
    .Z(_0051_));
 MUX2_X1 _1380_ (.A(\a_to_b_mem[12][7] ),
    .B(_0853_),
    .S(_0864_),
    .Z(_0052_));
 NAND3_X2 _1381_ (.A1(_0854_),
    .A2(_1249_),
    .A3(_0862_),
    .ZN(_0865_));
 AOI21_X4 _1382_ (.A(_0865_),
    .B1(_0838_),
    .B2(_0795_),
    .ZN(_0866_));
 MUX2_X1 _1383_ (.A(\a_to_b_mem[13][0] ),
    .B(_0828_),
    .S(_0866_),
    .Z(_0053_));
 MUX2_X1 _1384_ (.A(\a_to_b_mem[13][1] ),
    .B(_0841_),
    .S(_0866_),
    .Z(_0054_));
 MUX2_X1 _1385_ (.A(\a_to_b_mem[13][2] ),
    .B(_0843_),
    .S(_0866_),
    .Z(_0055_));
 MUX2_X1 _1386_ (.A(\a_to_b_mem[13][3] ),
    .B(_0845_),
    .S(_0866_),
    .Z(_0056_));
 MUX2_X1 _1387_ (.A(\a_to_b_mem[13][4] ),
    .B(_0847_),
    .S(_0866_),
    .Z(_0057_));
 MUX2_X1 _1388_ (.A(\a_to_b_mem[13][5] ),
    .B(_0849_),
    .S(_0866_),
    .Z(_0058_));
 MUX2_X1 _1389_ (.A(\a_to_b_mem[13][6] ),
    .B(_0851_),
    .S(_0866_),
    .Z(_0059_));
 MUX2_X1 _1390_ (.A(\a_to_b_mem[13][7] ),
    .B(_0853_),
    .S(_0866_),
    .Z(_0060_));
 NAND3_X2 _1391_ (.A1(_0854_),
    .A2(_1247_),
    .A3(_0862_),
    .ZN(_0867_));
 AOI21_X4 _1392_ (.A(_0867_),
    .B1(_0838_),
    .B2(_0795_),
    .ZN(_0868_));
 MUX2_X1 _1393_ (.A(\a_to_b_mem[14][0] ),
    .B(_0828_),
    .S(_0868_),
    .Z(_0061_));
 MUX2_X1 _1394_ (.A(\a_to_b_mem[14][1] ),
    .B(_0841_),
    .S(_0868_),
    .Z(_0062_));
 MUX2_X1 _1395_ (.A(\a_to_b_mem[14][2] ),
    .B(_0843_),
    .S(_0868_),
    .Z(_0063_));
 MUX2_X1 _1396_ (.A(\a_to_b_mem[14][3] ),
    .B(_0845_),
    .S(_0868_),
    .Z(_0064_));
 MUX2_X1 _1397_ (.A(\a_to_b_mem[14][4] ),
    .B(_0847_),
    .S(_0868_),
    .Z(_0065_));
 MUX2_X1 _1398_ (.A(\a_to_b_mem[14][5] ),
    .B(_0849_),
    .S(_0868_),
    .Z(_0066_));
 MUX2_X1 _1399_ (.A(\a_to_b_mem[14][6] ),
    .B(_0851_),
    .S(_0868_),
    .Z(_0067_));
 MUX2_X1 _1400_ (.A(\a_to_b_mem[14][7] ),
    .B(_0853_),
    .S(_0868_),
    .Z(_0068_));
 NAND3_X1 _1401_ (.A1(_0854_),
    .A2(_1251_),
    .A3(_0862_),
    .ZN(_0869_));
 AOI21_X4 _1402_ (.A(_0869_),
    .B1(_0837_),
    .B2(_0795_),
    .ZN(_0870_));
 MUX2_X1 _1403_ (.A(\a_to_b_mem[15][0] ),
    .B(_0828_),
    .S(_0870_),
    .Z(_0069_));
 MUX2_X1 _1404_ (.A(\a_to_b_mem[15][1] ),
    .B(_0841_),
    .S(_0870_),
    .Z(_0070_));
 MUX2_X1 _1405_ (.A(\a_to_b_mem[15][2] ),
    .B(_0843_),
    .S(_0870_),
    .Z(_0071_));
 MUX2_X1 _1406_ (.A(\a_to_b_mem[15][3] ),
    .B(_0845_),
    .S(_0870_),
    .Z(_0072_));
 MUX2_X1 _1407_ (.A(\a_to_b_mem[15][4] ),
    .B(_0847_),
    .S(_0870_),
    .Z(_0073_));
 MUX2_X1 _1408_ (.A(\a_to_b_mem[15][5] ),
    .B(_0849_),
    .S(_0870_),
    .Z(_0074_));
 MUX2_X1 _1409_ (.A(\a_to_b_mem[15][6] ),
    .B(_0851_),
    .S(_0870_),
    .Z(_0075_));
 MUX2_X1 _1410_ (.A(\a_to_b_mem[15][7] ),
    .B(_0853_),
    .S(_0870_),
    .Z(_0076_));
 NAND3_X1 _1411_ (.A1(_0829_),
    .A2(_1249_),
    .A3(_0833_),
    .ZN(_0871_));
 AOI21_X4 _1412_ (.A(_0871_),
    .B1(_0838_),
    .B2(_0795_),
    .ZN(_0872_));
 MUX2_X1 _1413_ (.A(\a_to_b_mem[1][0] ),
    .B(_0828_),
    .S(_0872_),
    .Z(_0077_));
 MUX2_X1 _1414_ (.A(\a_to_b_mem[1][1] ),
    .B(_0841_),
    .S(_0872_),
    .Z(_0078_));
 MUX2_X1 _1415_ (.A(\a_to_b_mem[1][2] ),
    .B(_0843_),
    .S(_0872_),
    .Z(_0079_));
 MUX2_X1 _1416_ (.A(\a_to_b_mem[1][3] ),
    .B(_0845_),
    .S(_0872_),
    .Z(_0080_));
 MUX2_X1 _1417_ (.A(\a_to_b_mem[1][4] ),
    .B(_0847_),
    .S(_0872_),
    .Z(_0081_));
 MUX2_X1 _1418_ (.A(\a_to_b_mem[1][5] ),
    .B(_0849_),
    .S(_0872_),
    .Z(_0082_));
 MUX2_X1 _1419_ (.A(\a_to_b_mem[1][6] ),
    .B(_0851_),
    .S(_0872_),
    .Z(_0083_));
 MUX2_X1 _1420_ (.A(\a_to_b_mem[1][7] ),
    .B(_0853_),
    .S(_0872_),
    .Z(_0084_));
 NAND3_X2 _1421_ (.A1(_0829_),
    .A2(_1247_),
    .A3(_0833_),
    .ZN(_0873_));
 AOI21_X4 _1422_ (.A(_0873_),
    .B1(_0838_),
    .B2(net42),
    .ZN(_0874_));
 MUX2_X1 _1423_ (.A(\a_to_b_mem[2][0] ),
    .B(_0828_),
    .S(_0874_),
    .Z(_0085_));
 MUX2_X1 _1424_ (.A(\a_to_b_mem[2][1] ),
    .B(_0841_),
    .S(_0874_),
    .Z(_0086_));
 MUX2_X1 _1425_ (.A(\a_to_b_mem[2][2] ),
    .B(_0843_),
    .S(_0874_),
    .Z(_0087_));
 MUX2_X1 _1426_ (.A(\a_to_b_mem[2][3] ),
    .B(_0845_),
    .S(_0874_),
    .Z(_0088_));
 MUX2_X1 _1427_ (.A(\a_to_b_mem[2][4] ),
    .B(_0847_),
    .S(_0874_),
    .Z(_0089_));
 MUX2_X1 _1428_ (.A(\a_to_b_mem[2][5] ),
    .B(_0849_),
    .S(_0874_),
    .Z(_0090_));
 MUX2_X1 _1429_ (.A(\a_to_b_mem[2][6] ),
    .B(_0851_),
    .S(_0874_),
    .Z(_0091_));
 MUX2_X1 _1430_ (.A(\a_to_b_mem[2][7] ),
    .B(_0853_),
    .S(_0874_),
    .Z(_0092_));
 NAND3_X1 _1431_ (.A1(_0829_),
    .A2(_1251_),
    .A3(_0833_),
    .ZN(_0875_));
 AOI21_X4 _1432_ (.A(_0875_),
    .B1(_0837_),
    .B2(net42),
    .ZN(_0876_));
 MUX2_X1 _1433_ (.A(\a_to_b_mem[3][0] ),
    .B(_0828_),
    .S(_0876_),
    .Z(_0093_));
 MUX2_X1 _1434_ (.A(\a_to_b_mem[3][1] ),
    .B(_0841_),
    .S(_0876_),
    .Z(_0094_));
 MUX2_X1 _1435_ (.A(\a_to_b_mem[3][2] ),
    .B(_0843_),
    .S(_0876_),
    .Z(_0095_));
 MUX2_X1 _1436_ (.A(\a_to_b_mem[3][3] ),
    .B(_0845_),
    .S(_0876_),
    .Z(_0096_));
 MUX2_X1 _1437_ (.A(\a_to_b_mem[3][4] ),
    .B(_0847_),
    .S(_0876_),
    .Z(_0097_));
 MUX2_X1 _1438_ (.A(\a_to_b_mem[3][5] ),
    .B(_0849_),
    .S(_0876_),
    .Z(_0098_));
 MUX2_X1 _1439_ (.A(\a_to_b_mem[3][6] ),
    .B(_0851_),
    .S(_0876_),
    .Z(_0099_));
 MUX2_X1 _1440_ (.A(\a_to_b_mem[3][7] ),
    .B(_0853_),
    .S(_0876_),
    .Z(_0100_));
 AND3_X1 _1441_ (.A1(_0854_),
    .A2(_1246_),
    .A3(_0833_),
    .ZN(_0877_));
 OAI21_X4 _1442_ (.A(_0877_),
    .B1(_0816_),
    .B2(_0809_),
    .ZN(_0878_));
 MUX2_X1 _1443_ (.A(_0827_),
    .B(\a_to_b_mem[4][0] ),
    .S(_0878_),
    .Z(_0101_));
 MUX2_X1 _1444_ (.A(_0840_),
    .B(\a_to_b_mem[4][1] ),
    .S(_0878_),
    .Z(_0102_));
 MUX2_X1 _1445_ (.A(_0842_),
    .B(\a_to_b_mem[4][2] ),
    .S(_0878_),
    .Z(_0103_));
 MUX2_X1 _1446_ (.A(_0844_),
    .B(\a_to_b_mem[4][3] ),
    .S(_0878_),
    .Z(_0104_));
 MUX2_X1 _1447_ (.A(_0846_),
    .B(\a_to_b_mem[4][4] ),
    .S(_0878_),
    .Z(_0105_));
 MUX2_X1 _1448_ (.A(_0848_),
    .B(\a_to_b_mem[4][5] ),
    .S(_0878_),
    .Z(_0106_));
 MUX2_X1 _1449_ (.A(_0850_),
    .B(\a_to_b_mem[4][6] ),
    .S(_0878_),
    .Z(_0107_));
 MUX2_X1 _1450_ (.A(_0852_),
    .B(\a_to_b_mem[4][7] ),
    .S(_0878_),
    .Z(_0108_));
 AND3_X1 _1451_ (.A1(_0854_),
    .A2(_1249_),
    .A3(_0833_),
    .ZN(_0879_));
 OAI21_X4 _1452_ (.A(_0879_),
    .B1(_0816_),
    .B2(_0809_),
    .ZN(_0880_));
 MUX2_X1 _1453_ (.A(_0827_),
    .B(\a_to_b_mem[5][0] ),
    .S(_0880_),
    .Z(_0109_));
 MUX2_X1 _1454_ (.A(_0840_),
    .B(\a_to_b_mem[5][1] ),
    .S(_0880_),
    .Z(_0110_));
 MUX2_X1 _1455_ (.A(_0842_),
    .B(\a_to_b_mem[5][2] ),
    .S(_0880_),
    .Z(_0111_));
 MUX2_X1 _1456_ (.A(_0844_),
    .B(\a_to_b_mem[5][3] ),
    .S(_0880_),
    .Z(_0112_));
 MUX2_X1 _1457_ (.A(_0846_),
    .B(\a_to_b_mem[5][4] ),
    .S(_0880_),
    .Z(_0113_));
 MUX2_X1 _1458_ (.A(_0848_),
    .B(\a_to_b_mem[5][5] ),
    .S(_0880_),
    .Z(_0114_));
 MUX2_X1 _1459_ (.A(_0850_),
    .B(\a_to_b_mem[5][6] ),
    .S(_0880_),
    .Z(_0115_));
 MUX2_X1 _1460_ (.A(_0852_),
    .B(\a_to_b_mem[5][7] ),
    .S(_0880_),
    .Z(_0116_));
 NOR4_X4 _1461_ (.A1(_0831_),
    .A2(_0832_),
    .A3(_0829_),
    .A4(_0855_),
    .ZN(_0881_));
 OAI21_X4 _1462_ (.A(_0881_),
    .B1(_0816_),
    .B2(_0809_),
    .ZN(_0882_));
 MUX2_X1 _1463_ (.A(_0827_),
    .B(\a_to_b_mem[6][0] ),
    .S(_0882_),
    .Z(_0117_));
 MUX2_X1 _1464_ (.A(_0840_),
    .B(\a_to_b_mem[6][1] ),
    .S(_0882_),
    .Z(_0118_));
 MUX2_X1 _1465_ (.A(_0842_),
    .B(\a_to_b_mem[6][2] ),
    .S(_0882_),
    .Z(_0119_));
 MUX2_X1 _1466_ (.A(_0844_),
    .B(\a_to_b_mem[6][3] ),
    .S(_0882_),
    .Z(_0120_));
 MUX2_X1 _1467_ (.A(_0846_),
    .B(\a_to_b_mem[6][4] ),
    .S(_0882_),
    .Z(_0121_));
 MUX2_X1 _1468_ (.A(_0848_),
    .B(\a_to_b_mem[6][5] ),
    .S(_0882_),
    .Z(_0122_));
 MUX2_X1 _1469_ (.A(_0850_),
    .B(\a_to_b_mem[6][6] ),
    .S(_0882_),
    .Z(_0123_));
 MUX2_X1 _1470_ (.A(_0852_),
    .B(\a_to_b_mem[6][7] ),
    .S(_0882_),
    .Z(_0124_));
 NOR4_X4 _1471_ (.A1(_0831_),
    .A2(_0832_),
    .A3(_0829_),
    .A4(_0859_),
    .ZN(_0883_));
 OAI21_X4 _1472_ (.A(_0883_),
    .B1(_0816_),
    .B2(_0809_),
    .ZN(_0884_));
 MUX2_X1 _1473_ (.A(_0827_),
    .B(\a_to_b_mem[7][0] ),
    .S(_0884_),
    .Z(_0125_));
 MUX2_X1 _1474_ (.A(_0840_),
    .B(\a_to_b_mem[7][1] ),
    .S(_0884_),
    .Z(_0126_));
 MUX2_X1 _1475_ (.A(_0842_),
    .B(\a_to_b_mem[7][2] ),
    .S(_0884_),
    .Z(_0127_));
 MUX2_X1 _1476_ (.A(_0844_),
    .B(\a_to_b_mem[7][3] ),
    .S(_0884_),
    .Z(_0128_));
 MUX2_X1 _1477_ (.A(_0846_),
    .B(\a_to_b_mem[7][4] ),
    .S(_0884_),
    .Z(_0129_));
 MUX2_X1 _1478_ (.A(_0848_),
    .B(\a_to_b_mem[7][5] ),
    .S(_0884_),
    .Z(_0130_));
 MUX2_X1 _1479_ (.A(_0850_),
    .B(\a_to_b_mem[7][6] ),
    .S(_0884_),
    .Z(_0131_));
 MUX2_X1 _1480_ (.A(_0852_),
    .B(\a_to_b_mem[7][7] ),
    .S(_0884_),
    .Z(_0132_));
 AND3_X1 _1481_ (.A1(_0829_),
    .A2(_1246_),
    .A3(_0862_),
    .ZN(_0885_));
 OAI21_X4 _1482_ (.A(_0885_),
    .B1(_0816_),
    .B2(net37),
    .ZN(_0886_));
 MUX2_X1 _1483_ (.A(_0827_),
    .B(\a_to_b_mem[8][0] ),
    .S(_0886_),
    .Z(_0133_));
 MUX2_X1 _1484_ (.A(_0840_),
    .B(\a_to_b_mem[8][1] ),
    .S(_0886_),
    .Z(_0134_));
 MUX2_X1 _1485_ (.A(_0842_),
    .B(\a_to_b_mem[8][2] ),
    .S(_0886_),
    .Z(_0135_));
 MUX2_X1 _1486_ (.A(_0844_),
    .B(\a_to_b_mem[8][3] ),
    .S(_0886_),
    .Z(_0136_));
 MUX2_X1 _1487_ (.A(_0846_),
    .B(\a_to_b_mem[8][4] ),
    .S(_0886_),
    .Z(_0137_));
 MUX2_X1 _1488_ (.A(_0848_),
    .B(\a_to_b_mem[8][5] ),
    .S(_0886_),
    .Z(_0138_));
 MUX2_X1 _1489_ (.A(_0850_),
    .B(\a_to_b_mem[8][6] ),
    .S(_0886_),
    .Z(_0139_));
 MUX2_X1 _1490_ (.A(_0852_),
    .B(\a_to_b_mem[8][7] ),
    .S(_0886_),
    .Z(_0140_));
 AND3_X1 _1491_ (.A1(_0829_),
    .A2(_1249_),
    .A3(_0862_),
    .ZN(_0887_));
 OAI21_X4 _1492_ (.A(_0887_),
    .B1(_0816_),
    .B2(net37),
    .ZN(_0888_));
 MUX2_X1 _1493_ (.A(_0827_),
    .B(\a_to_b_mem[9][0] ),
    .S(_0888_),
    .Z(_0141_));
 MUX2_X1 _1494_ (.A(_0840_),
    .B(\a_to_b_mem[9][1] ),
    .S(_0888_),
    .Z(_0142_));
 MUX2_X1 _1495_ (.A(_0842_),
    .B(\a_to_b_mem[9][2] ),
    .S(_0888_),
    .Z(_0143_));
 MUX2_X1 _1496_ (.A(_0844_),
    .B(\a_to_b_mem[9][3] ),
    .S(_0888_),
    .Z(_0144_));
 MUX2_X1 _1497_ (.A(_0846_),
    .B(\a_to_b_mem[9][4] ),
    .S(_0888_),
    .Z(_0145_));
 MUX2_X1 _1498_ (.A(_0848_),
    .B(\a_to_b_mem[9][5] ),
    .S(_0888_),
    .Z(_0146_));
 MUX2_X1 _1499_ (.A(_0850_),
    .B(\a_to_b_mem[9][6] ),
    .S(_0888_),
    .Z(_0147_));
 MUX2_X1 _1500_ (.A(_0852_),
    .B(\a_to_b_mem[9][7] ),
    .S(_0888_),
    .Z(_0148_));
 CLKBUF_X2 _1501_ (.A(b_wr_data[0]),
    .Z(_0889_));
 BUF_X2 _1502_ (.A(_0889_),
    .Z(_0890_));
 INV_X4 _1503_ (.A(\b_wr_ptr[2] ),
    .ZN(_0891_));
 BUF_X2 _1504_ (.A(b_wr_en),
    .Z(_0892_));
 INV_X4 _1505_ (.A(_0892_),
    .ZN(_0893_));
 BUF_X4 _1506_ (.A(\b_wr_ptr[3] ),
    .Z(_0894_));
 NOR2_X4 _1507_ (.A1(_0893_),
    .A2(_0894_),
    .ZN(_0895_));
 NAND3_X2 _1508_ (.A1(_0891_),
    .A2(_1237_),
    .A3(_0895_),
    .ZN(_0896_));
 AND4_X1 _1509_ (.A1(_0799_),
    .A2(_1256_),
    .A3(_0821_),
    .A4(_0798_),
    .ZN(_0897_));
 NOR4_X1 _1510_ (.A1(_0799_),
    .A2(net30),
    .A3(_0820_),
    .A4(net32),
    .ZN(_0898_));
 MUX2_X2 _1511_ (.A(_0897_),
    .B(_0898_),
    .S(_0801_),
    .Z(_0899_));
 BUF_X8 _1512_ (.A(_0899_),
    .Z(_0900_));
 AOI21_X4 _1513_ (.A(_0896_),
    .B1(_0900_),
    .B2(_0808_),
    .ZN(_0901_));
 MUX2_X1 _1514_ (.A(\b_to_a_mem[0][0] ),
    .B(_0890_),
    .S(_0901_),
    .Z(_0167_));
 CLKBUF_X2 _1515_ (.A(b_wr_data[1]),
    .Z(_0902_));
 BUF_X2 _1516_ (.A(_0902_),
    .Z(_0903_));
 MUX2_X1 _1517_ (.A(\b_to_a_mem[0][1] ),
    .B(_0903_),
    .S(_0901_),
    .Z(_0168_));
 CLKBUF_X2 _1518_ (.A(b_wr_data[2]),
    .Z(_0904_));
 BUF_X2 _1519_ (.A(_0904_),
    .Z(_0905_));
 MUX2_X1 _1520_ (.A(\b_to_a_mem[0][2] ),
    .B(_0905_),
    .S(_0901_),
    .Z(_0169_));
 CLKBUF_X2 _1521_ (.A(b_wr_data[3]),
    .Z(_0906_));
 BUF_X2 _1522_ (.A(_0906_),
    .Z(_0907_));
 MUX2_X1 _1523_ (.A(\b_to_a_mem[0][3] ),
    .B(_0907_),
    .S(_0901_),
    .Z(_0170_));
 BUF_X2 _1524_ (.A(b_wr_data[4]),
    .Z(_0908_));
 BUF_X2 _1525_ (.A(_0908_),
    .Z(_0909_));
 MUX2_X1 _1526_ (.A(\b_to_a_mem[0][4] ),
    .B(_0909_),
    .S(_0901_),
    .Z(_0171_));
 BUF_X2 _1527_ (.A(b_wr_data[5]),
    .Z(_0910_));
 BUF_X2 _1528_ (.A(_0910_),
    .Z(_0911_));
 MUX2_X1 _1529_ (.A(\b_to_a_mem[0][5] ),
    .B(_0911_),
    .S(_0901_),
    .Z(_0172_));
 BUF_X2 _1530_ (.A(b_wr_data[6]),
    .Z(_0912_));
 BUF_X2 _1531_ (.A(_0912_),
    .Z(_0913_));
 MUX2_X1 _1532_ (.A(\b_to_a_mem[0][6] ),
    .B(_0913_),
    .S(_0901_),
    .Z(_0173_));
 CLKBUF_X2 _1533_ (.A(b_wr_data[7]),
    .Z(_0914_));
 BUF_X2 _1534_ (.A(_0914_),
    .Z(_0915_));
 MUX2_X1 _1535_ (.A(\b_to_a_mem[0][7] ),
    .B(_0915_),
    .S(_0901_),
    .Z(_0174_));
 BUF_X4 _1536_ (.A(\b_wr_ptr[2] ),
    .Z(_0916_));
 INV_X1 _1537_ (.A(_1238_),
    .ZN(_0917_));
 NAND2_X1 _1538_ (.A1(_0892_),
    .A2(_0894_),
    .ZN(_0918_));
 NOR3_X2 _1539_ (.A1(_0916_),
    .A2(_0917_),
    .A3(_0918_),
    .ZN(_0919_));
 OAI21_X4 _1540_ (.A(_0919_),
    .B1(_0825_),
    .B2(_0818_),
    .ZN(_0920_));
 MUX2_X1 _1541_ (.A(_0890_),
    .B(\b_to_a_mem[10][0] ),
    .S(_0920_),
    .Z(_0175_));
 MUX2_X1 _1542_ (.A(_0903_),
    .B(\b_to_a_mem[10][1] ),
    .S(_0920_),
    .Z(_0176_));
 MUX2_X1 _1543_ (.A(_0905_),
    .B(\b_to_a_mem[10][2] ),
    .S(_0920_),
    .Z(_0177_));
 MUX2_X1 _1544_ (.A(_0907_),
    .B(\b_to_a_mem[10][3] ),
    .S(_0920_),
    .Z(_0178_));
 MUX2_X1 _1545_ (.A(_0909_),
    .B(\b_to_a_mem[10][4] ),
    .S(_0920_),
    .Z(_0179_));
 MUX2_X1 _1546_ (.A(_0911_),
    .B(\b_to_a_mem[10][5] ),
    .S(_0920_),
    .Z(_0180_));
 MUX2_X1 _1547_ (.A(_0913_),
    .B(\b_to_a_mem[10][6] ),
    .S(_0920_),
    .Z(_0181_));
 MUX2_X1 _1548_ (.A(_0915_),
    .B(\b_to_a_mem[10][7] ),
    .S(_0920_),
    .Z(_0182_));
 INV_X1 _1549_ (.A(_1242_),
    .ZN(_0921_));
 NOR3_X2 _1550_ (.A1(_0916_),
    .A2(_0921_),
    .A3(_0918_),
    .ZN(_0922_));
 OAI21_X4 _1551_ (.A(_0922_),
    .B1(_0825_),
    .B2(_0818_),
    .ZN(_0923_));
 MUX2_X1 _1552_ (.A(_0890_),
    .B(\b_to_a_mem[11][0] ),
    .S(_0923_),
    .Z(_0183_));
 MUX2_X1 _1553_ (.A(_0903_),
    .B(\b_to_a_mem[11][1] ),
    .S(_0923_),
    .Z(_0184_));
 MUX2_X1 _1554_ (.A(_0905_),
    .B(\b_to_a_mem[11][2] ),
    .S(_0923_),
    .Z(_0185_));
 MUX2_X1 _1555_ (.A(_0907_),
    .B(\b_to_a_mem[11][3] ),
    .S(_0923_),
    .Z(_0186_));
 MUX2_X1 _1556_ (.A(_0909_),
    .B(\b_to_a_mem[11][4] ),
    .S(_0923_),
    .Z(_0187_));
 MUX2_X1 _1557_ (.A(_0911_),
    .B(\b_to_a_mem[11][5] ),
    .S(_0923_),
    .Z(_0188_));
 MUX2_X1 _1558_ (.A(_0913_),
    .B(\b_to_a_mem[11][6] ),
    .S(_0923_),
    .Z(_0189_));
 MUX2_X1 _1559_ (.A(_0915_),
    .B(\b_to_a_mem[11][7] ),
    .S(_0923_),
    .Z(_0190_));
 AND2_X2 _1560_ (.A1(_0892_),
    .A2(_0894_),
    .ZN(_0924_));
 NAND3_X2 _1561_ (.A1(_0916_),
    .A2(_1237_),
    .A3(_0924_),
    .ZN(_0925_));
 AOI21_X4 _1562_ (.A(_0925_),
    .B1(_0900_),
    .B2(_0808_),
    .ZN(_0926_));
 MUX2_X1 _1563_ (.A(\b_to_a_mem[12][0] ),
    .B(_0890_),
    .S(_0926_),
    .Z(_0191_));
 MUX2_X1 _1564_ (.A(\b_to_a_mem[12][1] ),
    .B(_0903_),
    .S(_0926_),
    .Z(_0192_));
 MUX2_X1 _1565_ (.A(\b_to_a_mem[12][2] ),
    .B(_0905_),
    .S(_0926_),
    .Z(_0193_));
 MUX2_X1 _1566_ (.A(\b_to_a_mem[12][3] ),
    .B(_0907_),
    .S(_0926_),
    .Z(_0194_));
 MUX2_X1 _1567_ (.A(\b_to_a_mem[12][4] ),
    .B(_0909_),
    .S(_0926_),
    .Z(_0195_));
 MUX2_X1 _1568_ (.A(\b_to_a_mem[12][5] ),
    .B(_0911_),
    .S(_0926_),
    .Z(_0196_));
 MUX2_X1 _1569_ (.A(\b_to_a_mem[12][6] ),
    .B(_0913_),
    .S(_0926_),
    .Z(_0197_));
 MUX2_X1 _1570_ (.A(\b_to_a_mem[12][7] ),
    .B(_0915_),
    .S(_0926_),
    .Z(_0198_));
 NAND3_X2 _1571_ (.A1(_0916_),
    .A2(_1240_),
    .A3(_0924_),
    .ZN(_0927_));
 AOI21_X4 _1572_ (.A(_0927_),
    .B1(_0900_),
    .B2(_0808_),
    .ZN(_0928_));
 MUX2_X1 _1573_ (.A(\b_to_a_mem[13][0] ),
    .B(_0890_),
    .S(_0928_),
    .Z(_0199_));
 MUX2_X1 _1574_ (.A(\b_to_a_mem[13][1] ),
    .B(_0903_),
    .S(_0928_),
    .Z(_0200_));
 MUX2_X1 _1575_ (.A(\b_to_a_mem[13][2] ),
    .B(_0905_),
    .S(_0928_),
    .Z(_0201_));
 MUX2_X1 _1576_ (.A(\b_to_a_mem[13][3] ),
    .B(_0907_),
    .S(_0928_),
    .Z(_0202_));
 MUX2_X1 _1577_ (.A(\b_to_a_mem[13][4] ),
    .B(_0909_),
    .S(_0928_),
    .Z(_0203_));
 MUX2_X1 _1578_ (.A(\b_to_a_mem[13][5] ),
    .B(_0911_),
    .S(_0928_),
    .Z(_0204_));
 MUX2_X1 _1579_ (.A(\b_to_a_mem[13][6] ),
    .B(_0913_),
    .S(_0928_),
    .Z(_0205_));
 MUX2_X1 _1580_ (.A(\b_to_a_mem[13][7] ),
    .B(_0915_),
    .S(_0928_),
    .Z(_0206_));
 NAND3_X2 _1581_ (.A1(_0916_),
    .A2(_1238_),
    .A3(_0924_),
    .ZN(_0929_));
 AOI21_X4 _1582_ (.A(_0929_),
    .B1(_0900_),
    .B2(_0808_),
    .ZN(_0930_));
 MUX2_X1 _1583_ (.A(\b_to_a_mem[14][0] ),
    .B(_0890_),
    .S(_0930_),
    .Z(_0207_));
 MUX2_X1 _1584_ (.A(\b_to_a_mem[14][1] ),
    .B(_0903_),
    .S(_0930_),
    .Z(_0208_));
 MUX2_X1 _1585_ (.A(\b_to_a_mem[14][2] ),
    .B(_0905_),
    .S(_0930_),
    .Z(_0209_));
 MUX2_X1 _1586_ (.A(\b_to_a_mem[14][3] ),
    .B(_0907_),
    .S(_0930_),
    .Z(_0210_));
 MUX2_X1 _1587_ (.A(\b_to_a_mem[14][4] ),
    .B(_0909_),
    .S(_0930_),
    .Z(_0211_));
 MUX2_X1 _1588_ (.A(\b_to_a_mem[14][5] ),
    .B(_0911_),
    .S(_0930_),
    .Z(_0212_));
 MUX2_X1 _1589_ (.A(\b_to_a_mem[14][6] ),
    .B(_0913_),
    .S(_0930_),
    .Z(_0213_));
 MUX2_X1 _1590_ (.A(\b_to_a_mem[14][7] ),
    .B(_0915_),
    .S(_0930_),
    .Z(_0214_));
 NAND3_X1 _1591_ (.A1(_0916_),
    .A2(_1242_),
    .A3(_0924_),
    .ZN(_0931_));
 AOI21_X4 _1592_ (.A(_0931_),
    .B1(_0899_),
    .B2(_0807_),
    .ZN(_0932_));
 MUX2_X1 _1593_ (.A(\b_to_a_mem[15][0] ),
    .B(_0890_),
    .S(_0932_),
    .Z(_0215_));
 MUX2_X1 _1594_ (.A(\b_to_a_mem[15][1] ),
    .B(_0903_),
    .S(_0932_),
    .Z(_0216_));
 MUX2_X1 _1595_ (.A(\b_to_a_mem[15][2] ),
    .B(_0905_),
    .S(_0932_),
    .Z(_0217_));
 MUX2_X1 _1596_ (.A(\b_to_a_mem[15][3] ),
    .B(_0907_),
    .S(_0932_),
    .Z(_0218_));
 MUX2_X1 _1597_ (.A(\b_to_a_mem[15][4] ),
    .B(_0909_),
    .S(_0932_),
    .Z(_0219_));
 MUX2_X1 _1598_ (.A(\b_to_a_mem[15][5] ),
    .B(_0911_),
    .S(_0932_),
    .Z(_0220_));
 MUX2_X1 _1599_ (.A(\b_to_a_mem[15][6] ),
    .B(_0913_),
    .S(_0932_),
    .Z(_0221_));
 MUX2_X1 _1600_ (.A(\b_to_a_mem[15][7] ),
    .B(_0915_),
    .S(_0932_),
    .Z(_0222_));
 NAND3_X2 _1601_ (.A1(_0891_),
    .A2(_1240_),
    .A3(_0895_),
    .ZN(_0300_));
 AOI21_X4 _1602_ (.A(_0300_),
    .B1(_0900_),
    .B2(_0807_),
    .ZN(_0301_));
 MUX2_X1 _1603_ (.A(\b_to_a_mem[1][0] ),
    .B(_0890_),
    .S(_0301_),
    .Z(_0223_));
 MUX2_X1 _1604_ (.A(\b_to_a_mem[1][1] ),
    .B(_0903_),
    .S(_0301_),
    .Z(_0224_));
 MUX2_X1 _1605_ (.A(\b_to_a_mem[1][2] ),
    .B(_0905_),
    .S(_0301_),
    .Z(_0225_));
 MUX2_X1 _1606_ (.A(\b_to_a_mem[1][3] ),
    .B(_0907_),
    .S(_0301_),
    .Z(_0226_));
 MUX2_X1 _1607_ (.A(\b_to_a_mem[1][4] ),
    .B(_0909_),
    .S(_0301_),
    .Z(_0227_));
 MUX2_X1 _1608_ (.A(\b_to_a_mem[1][5] ),
    .B(_0911_),
    .S(_0301_),
    .Z(_0228_));
 MUX2_X1 _1609_ (.A(\b_to_a_mem[1][6] ),
    .B(_0913_),
    .S(_0301_),
    .Z(_0229_));
 MUX2_X1 _1610_ (.A(\b_to_a_mem[1][7] ),
    .B(_0915_),
    .S(_0301_),
    .Z(_0230_));
 NAND3_X1 _1611_ (.A1(_0891_),
    .A2(_1238_),
    .A3(_0895_),
    .ZN(_0302_));
 AOI21_X4 _1612_ (.A(_0302_),
    .B1(_0900_),
    .B2(_0807_),
    .ZN(_0303_));
 MUX2_X1 _1613_ (.A(\b_to_a_mem[2][0] ),
    .B(_0890_),
    .S(_0303_),
    .Z(_0231_));
 MUX2_X1 _1614_ (.A(\b_to_a_mem[2][1] ),
    .B(_0903_),
    .S(_0303_),
    .Z(_0232_));
 MUX2_X1 _1615_ (.A(\b_to_a_mem[2][2] ),
    .B(_0905_),
    .S(_0303_),
    .Z(_0233_));
 MUX2_X1 _1616_ (.A(\b_to_a_mem[2][3] ),
    .B(_0907_),
    .S(_0303_),
    .Z(_0234_));
 MUX2_X1 _1617_ (.A(\b_to_a_mem[2][4] ),
    .B(_0909_),
    .S(_0303_),
    .Z(_0235_));
 MUX2_X1 _1618_ (.A(\b_to_a_mem[2][5] ),
    .B(_0911_),
    .S(_0303_),
    .Z(_0236_));
 MUX2_X1 _1619_ (.A(\b_to_a_mem[2][6] ),
    .B(_0913_),
    .S(_0303_),
    .Z(_0237_));
 MUX2_X1 _1620_ (.A(\b_to_a_mem[2][7] ),
    .B(_0915_),
    .S(_0303_),
    .Z(_0238_));
 NAND3_X2 _1621_ (.A1(_0891_),
    .A2(_1242_),
    .A3(_0895_),
    .ZN(_0304_));
 AOI21_X4 _1622_ (.A(_0304_),
    .B1(_0899_),
    .B2(_0807_),
    .ZN(_0305_));
 MUX2_X1 _1623_ (.A(\b_to_a_mem[3][0] ),
    .B(_0890_),
    .S(_0305_),
    .Z(_0239_));
 MUX2_X1 _1624_ (.A(\b_to_a_mem[3][1] ),
    .B(_0903_),
    .S(_0305_),
    .Z(_0240_));
 MUX2_X1 _1625_ (.A(\b_to_a_mem[3][2] ),
    .B(_0905_),
    .S(_0305_),
    .Z(_0241_));
 MUX2_X1 _1626_ (.A(\b_to_a_mem[3][3] ),
    .B(_0907_),
    .S(_0305_),
    .Z(_0242_));
 MUX2_X1 _1627_ (.A(\b_to_a_mem[3][4] ),
    .B(_0909_),
    .S(_0305_),
    .Z(_0243_));
 MUX2_X1 _1628_ (.A(\b_to_a_mem[3][5] ),
    .B(_0911_),
    .S(_0305_),
    .Z(_0244_));
 MUX2_X1 _1629_ (.A(\b_to_a_mem[3][6] ),
    .B(_0913_),
    .S(_0305_),
    .Z(_0245_));
 MUX2_X1 _1630_ (.A(\b_to_a_mem[3][7] ),
    .B(_0915_),
    .S(_0305_),
    .Z(_0246_));
 AND3_X1 _1631_ (.A1(_0916_),
    .A2(_1237_),
    .A3(_0895_),
    .ZN(_0306_));
 OAI21_X4 _1632_ (.A(_0306_),
    .B1(_0825_),
    .B2(_0818_),
    .ZN(_0307_));
 MUX2_X1 _1633_ (.A(_0889_),
    .B(\b_to_a_mem[4][0] ),
    .S(_0307_),
    .Z(_0247_));
 MUX2_X1 _1634_ (.A(_0902_),
    .B(\b_to_a_mem[4][1] ),
    .S(_0307_),
    .Z(_0248_));
 MUX2_X1 _1635_ (.A(_0904_),
    .B(\b_to_a_mem[4][2] ),
    .S(_0307_),
    .Z(_0249_));
 MUX2_X1 _1636_ (.A(_0906_),
    .B(\b_to_a_mem[4][3] ),
    .S(_0307_),
    .Z(_0250_));
 MUX2_X1 _1637_ (.A(_0908_),
    .B(\b_to_a_mem[4][4] ),
    .S(_0307_),
    .Z(_0251_));
 MUX2_X1 _1638_ (.A(_0910_),
    .B(\b_to_a_mem[4][5] ),
    .S(_0307_),
    .Z(_0252_));
 MUX2_X1 _1639_ (.A(_0912_),
    .B(\b_to_a_mem[4][6] ),
    .S(_0307_),
    .Z(_0253_));
 MUX2_X1 _1640_ (.A(_0914_),
    .B(\b_to_a_mem[4][7] ),
    .S(_0307_),
    .Z(_0254_));
 AND3_X1 _1641_ (.A1(_0916_),
    .A2(_1240_),
    .A3(_0895_),
    .ZN(_0308_));
 OAI21_X4 _1642_ (.A(_0308_),
    .B1(_0825_),
    .B2(_0818_),
    .ZN(_0309_));
 MUX2_X1 _1643_ (.A(_0889_),
    .B(\b_to_a_mem[5][0] ),
    .S(_0309_),
    .Z(_0255_));
 MUX2_X1 _1644_ (.A(_0902_),
    .B(\b_to_a_mem[5][1] ),
    .S(_0309_),
    .Z(_0256_));
 MUX2_X1 _1645_ (.A(_0904_),
    .B(\b_to_a_mem[5][2] ),
    .S(_0309_),
    .Z(_0257_));
 MUX2_X1 _1646_ (.A(_0906_),
    .B(\b_to_a_mem[5][3] ),
    .S(_0309_),
    .Z(_0258_));
 MUX2_X1 _1647_ (.A(_0908_),
    .B(\b_to_a_mem[5][4] ),
    .S(_0309_),
    .Z(_0259_));
 MUX2_X1 _1648_ (.A(_0910_),
    .B(\b_to_a_mem[5][5] ),
    .S(_0309_),
    .Z(_0260_));
 MUX2_X1 _1649_ (.A(_0912_),
    .B(\b_to_a_mem[5][6] ),
    .S(_0309_),
    .Z(_0261_));
 MUX2_X1 _1650_ (.A(_0914_),
    .B(\b_to_a_mem[5][7] ),
    .S(_0309_),
    .Z(_0262_));
 NOR4_X4 _1651_ (.A1(_0893_),
    .A2(_0894_),
    .A3(_0891_),
    .A4(_0917_),
    .ZN(_0310_));
 OAI21_X4 _1652_ (.A(_0310_),
    .B1(_0825_),
    .B2(_0818_),
    .ZN(_0311_));
 MUX2_X1 _1653_ (.A(_0889_),
    .B(\b_to_a_mem[6][0] ),
    .S(_0311_),
    .Z(_0263_));
 MUX2_X1 _1654_ (.A(_0902_),
    .B(\b_to_a_mem[6][1] ),
    .S(_0311_),
    .Z(_0264_));
 MUX2_X1 _1655_ (.A(_0904_),
    .B(\b_to_a_mem[6][2] ),
    .S(_0311_),
    .Z(_0265_));
 MUX2_X1 _1656_ (.A(_0906_),
    .B(\b_to_a_mem[6][3] ),
    .S(_0311_),
    .Z(_0266_));
 MUX2_X1 _1657_ (.A(_0908_),
    .B(\b_to_a_mem[6][4] ),
    .S(_0311_),
    .Z(_0267_));
 MUX2_X1 _1658_ (.A(_0910_),
    .B(\b_to_a_mem[6][5] ),
    .S(_0311_),
    .Z(_0268_));
 MUX2_X1 _1659_ (.A(_0912_),
    .B(\b_to_a_mem[6][6] ),
    .S(_0311_),
    .Z(_0269_));
 MUX2_X1 _1660_ (.A(_0914_),
    .B(\b_to_a_mem[6][7] ),
    .S(_0311_),
    .Z(_0270_));
 NOR4_X4 _1661_ (.A1(_0893_),
    .A2(_0894_),
    .A3(_0891_),
    .A4(_0921_),
    .ZN(_0312_));
 OAI21_X4 _1662_ (.A(_0312_),
    .B1(_0825_),
    .B2(_0818_),
    .ZN(_0313_));
 MUX2_X1 _1663_ (.A(_0889_),
    .B(\b_to_a_mem[7][0] ),
    .S(_0313_),
    .Z(_0271_));
 MUX2_X1 _1664_ (.A(_0902_),
    .B(\b_to_a_mem[7][1] ),
    .S(_0313_),
    .Z(_0272_));
 MUX2_X1 _1665_ (.A(_0904_),
    .B(\b_to_a_mem[7][2] ),
    .S(_0313_),
    .Z(_0273_));
 MUX2_X1 _1666_ (.A(_0906_),
    .B(\b_to_a_mem[7][3] ),
    .S(_0313_),
    .Z(_0274_));
 MUX2_X1 _1667_ (.A(_0908_),
    .B(\b_to_a_mem[7][4] ),
    .S(_0313_),
    .Z(_0275_));
 MUX2_X1 _1668_ (.A(_0910_),
    .B(\b_to_a_mem[7][5] ),
    .S(_0313_),
    .Z(_0276_));
 MUX2_X1 _1669_ (.A(_0912_),
    .B(\b_to_a_mem[7][6] ),
    .S(_0313_),
    .Z(_0277_));
 MUX2_X1 _1670_ (.A(_0914_),
    .B(\b_to_a_mem[7][7] ),
    .S(_0313_),
    .Z(_0278_));
 AND3_X1 _1671_ (.A1(_0891_),
    .A2(_1237_),
    .A3(_0924_),
    .ZN(_0314_));
 OAI21_X4 _1672_ (.A(_0314_),
    .B1(_0825_),
    .B2(net36),
    .ZN(_0315_));
 MUX2_X1 _1673_ (.A(_0889_),
    .B(\b_to_a_mem[8][0] ),
    .S(_0315_),
    .Z(_0279_));
 MUX2_X1 _1674_ (.A(_0902_),
    .B(\b_to_a_mem[8][1] ),
    .S(_0315_),
    .Z(_0280_));
 MUX2_X1 _1675_ (.A(_0904_),
    .B(\b_to_a_mem[8][2] ),
    .S(_0315_),
    .Z(_0281_));
 MUX2_X1 _1676_ (.A(_0906_),
    .B(\b_to_a_mem[8][3] ),
    .S(_0315_),
    .Z(_0282_));
 MUX2_X1 _1677_ (.A(_0908_),
    .B(\b_to_a_mem[8][4] ),
    .S(_0315_),
    .Z(_0283_));
 MUX2_X1 _1678_ (.A(_0910_),
    .B(\b_to_a_mem[8][5] ),
    .S(_0315_),
    .Z(_0284_));
 MUX2_X1 _1679_ (.A(_0912_),
    .B(\b_to_a_mem[8][6] ),
    .S(_0315_),
    .Z(_0285_));
 MUX2_X1 _1680_ (.A(_0914_),
    .B(\b_to_a_mem[8][7] ),
    .S(_0315_),
    .Z(_0286_));
 AND3_X1 _1681_ (.A1(_0891_),
    .A2(_1240_),
    .A3(_0924_),
    .ZN(_0316_));
 OAI21_X4 _1682_ (.A(_0316_),
    .B1(_0825_),
    .B2(net36),
    .ZN(_0317_));
 MUX2_X1 _1683_ (.A(_0889_),
    .B(\b_to_a_mem[9][0] ),
    .S(_0317_),
    .Z(_0287_));
 MUX2_X1 _1684_ (.A(_0902_),
    .B(\b_to_a_mem[9][1] ),
    .S(_0317_),
    .Z(_0288_));
 MUX2_X1 _1685_ (.A(_0904_),
    .B(\b_to_a_mem[9][2] ),
    .S(_0317_),
    .Z(_0289_));
 MUX2_X1 _1686_ (.A(_0906_),
    .B(\b_to_a_mem[9][3] ),
    .S(_0317_),
    .Z(_0290_));
 MUX2_X1 _1687_ (.A(_0908_),
    .B(\b_to_a_mem[9][4] ),
    .S(_0317_),
    .Z(_0291_));
 MUX2_X1 _1688_ (.A(_0910_),
    .B(\b_to_a_mem[9][5] ),
    .S(_0317_),
    .Z(_0292_));
 MUX2_X1 _1689_ (.A(_0912_),
    .B(\b_to_a_mem[9][6] ),
    .S(_0317_),
    .Z(_0293_));
 MUX2_X1 _1690_ (.A(_0914_),
    .B(\b_to_a_mem[9][7] ),
    .S(_0317_),
    .Z(_0294_));
 CLKBUF_X3 _1691_ (.A(a_rd_en),
    .Z(_0318_));
 INV_X2 _1692_ (.A(_0318_),
    .ZN(_0319_));
 BUF_X2 _1693_ (.A(rst_n),
    .Z(_0320_));
 INV_X2 _1694_ (.A(_0320_),
    .ZN(_0321_));
 NOR2_X4 _1695_ (.A1(_0319_),
    .A2(_0321_),
    .ZN(_0322_));
 BUF_X2 _1696_ (.A(\a_rd_ptr[0] ),
    .Z(_0323_));
 CLKBUF_X3 _1697_ (.A(_0323_),
    .Z(_0324_));
 BUF_X2 _1698_ (.A(\a_rd_ptr[1] ),
    .Z(_0325_));
 BUF_X4 _1699_ (.A(_0325_),
    .Z(_0326_));
 BUF_X4 _1700_ (.A(_0326_),
    .Z(_0327_));
 MUX2_X1 _1701_ (.A(\b_to_a_mem[4][0] ),
    .B(\b_to_a_mem[6][0] ),
    .S(_0327_),
    .Z(_0328_));
 NOR2_X1 _1702_ (.A1(_0324_),
    .A2(_0328_),
    .ZN(_0329_));
 INV_X2 _1703_ (.A(_0323_),
    .ZN(_0330_));
 CLKBUF_X3 _1704_ (.A(_0330_),
    .Z(_0331_));
 MUX2_X1 _1705_ (.A(\b_to_a_mem[5][0] ),
    .B(\b_to_a_mem[7][0] ),
    .S(_0327_),
    .Z(_0332_));
 NOR2_X1 _1706_ (.A1(_0331_),
    .A2(_0332_),
    .ZN(_0333_));
 CLKBUF_X3 _1707_ (.A(\a_rd_ptr[2] ),
    .Z(_0334_));
 CLKBUF_X3 _1708_ (.A(\a_rd_ptr[3] ),
    .Z(_0335_));
 INV_X2 _1709_ (.A(_0335_),
    .ZN(_0336_));
 NAND2_X4 _1710_ (.A1(_0334_),
    .A2(_0336_),
    .ZN(_0337_));
 NAND2_X4 _1711_ (.A1(_0334_),
    .A2(_0335_),
    .ZN(_0338_));
 BUF_X4 _1712_ (.A(_0325_),
    .Z(_0339_));
 MUX2_X1 _1713_ (.A(\b_to_a_mem[12][0] ),
    .B(\b_to_a_mem[14][0] ),
    .S(_0339_),
    .Z(_0340_));
 NOR2_X1 _1714_ (.A1(_0323_),
    .A2(_0340_),
    .ZN(_0341_));
 CLKBUF_X3 _1715_ (.A(_0330_),
    .Z(_0342_));
 BUF_X4 _1716_ (.A(_0325_),
    .Z(_0343_));
 MUX2_X1 _1717_ (.A(\b_to_a_mem[13][0] ),
    .B(\b_to_a_mem[15][0] ),
    .S(_0343_),
    .Z(_0344_));
 NOR2_X1 _1718_ (.A1(_0342_),
    .A2(_0344_),
    .ZN(_0345_));
 OAI33_X1 _1719_ (.A1(_0329_),
    .A2(_0333_),
    .A3(_0337_),
    .B1(_0338_),
    .B2(_0341_),
    .B3(_0345_),
    .ZN(_0346_));
 MUX2_X1 _1720_ (.A(\b_to_a_mem[0][0] ),
    .B(\b_to_a_mem[2][0] ),
    .S(_0327_),
    .Z(_0347_));
 NOR2_X1 _1721_ (.A1(_0324_),
    .A2(_0347_),
    .ZN(_0348_));
 BUF_X4 _1722_ (.A(_0326_),
    .Z(_0349_));
 MUX2_X1 _1723_ (.A(\b_to_a_mem[1][0] ),
    .B(\b_to_a_mem[3][0] ),
    .S(_0349_),
    .Z(_0350_));
 NOR2_X1 _1724_ (.A1(_0331_),
    .A2(_0350_),
    .ZN(_0351_));
 INV_X2 _1725_ (.A(_0334_),
    .ZN(_0352_));
 NAND2_X4 _1726_ (.A1(_0352_),
    .A2(_0336_),
    .ZN(_0353_));
 NAND2_X4 _1727_ (.A1(_0352_),
    .A2(_0335_),
    .ZN(_0354_));
 MUX2_X1 _1728_ (.A(\b_to_a_mem[8][0] ),
    .B(\b_to_a_mem[10][0] ),
    .S(_0343_),
    .Z(_0355_));
 NOR2_X1 _1729_ (.A1(_0323_),
    .A2(_0355_),
    .ZN(_0356_));
 MUX2_X1 _1730_ (.A(\b_to_a_mem[9][0] ),
    .B(\b_to_a_mem[11][0] ),
    .S(_0326_),
    .Z(_0357_));
 NOR2_X1 _1731_ (.A1(_0330_),
    .A2(_0357_),
    .ZN(_0358_));
 OAI33_X1 _1732_ (.A1(_0348_),
    .A2(_0351_),
    .A3(_0353_),
    .B1(_0354_),
    .B2(_0356_),
    .B3(_0358_),
    .ZN(_0359_));
 OAI221_X1 _1733_ (.A(_0322_),
    .B1(_0346_),
    .B2(_0359_),
    .C1(net34),
    .C2(_0825_),
    .ZN(_0360_));
 CLKBUF_X3 _1734_ (.A(_0320_),
    .Z(_0361_));
 CLKBUF_X3 _1735_ (.A(_0899_),
    .Z(_0362_));
 NAND4_X1 _1736_ (.A1(net5),
    .A2(_0361_),
    .A3(_0819_),
    .A4(_0362_),
    .ZN(_0363_));
 CLKBUF_X3 _1737_ (.A(_0320_),
    .Z(_0364_));
 CLKBUF_X3 _1738_ (.A(_0364_),
    .Z(_0365_));
 NAND3_X1 _1739_ (.A1(_0319_),
    .A2(net5),
    .A3(_0365_),
    .ZN(_0366_));
 NAND3_X1 _1740_ (.A1(_0360_),
    .A2(_0363_),
    .A3(_0366_),
    .ZN(_0008_));
 MUX2_X1 _1741_ (.A(\b_to_a_mem[8][1] ),
    .B(\b_to_a_mem[10][1] ),
    .S(_0327_),
    .Z(_0367_));
 NOR2_X1 _1742_ (.A1(_0324_),
    .A2(_0367_),
    .ZN(_0368_));
 MUX2_X1 _1743_ (.A(\b_to_a_mem[9][1] ),
    .B(\b_to_a_mem[11][1] ),
    .S(_0349_),
    .Z(_0369_));
 NOR2_X1 _1744_ (.A1(_0331_),
    .A2(_0369_),
    .ZN(_0370_));
 CLKBUF_X3 _1745_ (.A(_0323_),
    .Z(_0371_));
 BUF_X4 _1746_ (.A(_0326_),
    .Z(_0372_));
 MUX2_X1 _1747_ (.A(\b_to_a_mem[0][1] ),
    .B(\b_to_a_mem[2][1] ),
    .S(_0372_),
    .Z(_0373_));
 NOR2_X1 _1748_ (.A1(_0371_),
    .A2(_0373_),
    .ZN(_0374_));
 CLKBUF_X3 _1749_ (.A(_0330_),
    .Z(_0375_));
 MUX2_X1 _1750_ (.A(\b_to_a_mem[1][1] ),
    .B(\b_to_a_mem[3][1] ),
    .S(_0339_),
    .Z(_0376_));
 NOR2_X1 _1751_ (.A1(_0375_),
    .A2(_0376_),
    .ZN(_0377_));
 OAI33_X1 _1752_ (.A1(_0354_),
    .A2(_0368_),
    .A3(_0370_),
    .B1(_0374_),
    .B2(_0377_),
    .B3(_0353_),
    .ZN(_0378_));
 MUX2_X1 _1753_ (.A(\b_to_a_mem[12][1] ),
    .B(\b_to_a_mem[14][1] ),
    .S(_0372_),
    .Z(_0379_));
 NOR2_X1 _1754_ (.A1(_0371_),
    .A2(_0379_),
    .ZN(_0380_));
 BUF_X4 _1755_ (.A(_0326_),
    .Z(_0381_));
 MUX2_X1 _1756_ (.A(\b_to_a_mem[13][1] ),
    .B(\b_to_a_mem[15][1] ),
    .S(_0381_),
    .Z(_0382_));
 NOR2_X1 _1757_ (.A1(_0375_),
    .A2(_0382_),
    .ZN(_0383_));
 CLKBUF_X3 _1758_ (.A(_0323_),
    .Z(_0384_));
 MUX2_X1 _1759_ (.A(\b_to_a_mem[4][1] ),
    .B(\b_to_a_mem[6][1] ),
    .S(_0339_),
    .Z(_0385_));
 NOR2_X1 _1760_ (.A1(_0384_),
    .A2(_0385_),
    .ZN(_0386_));
 MUX2_X1 _1761_ (.A(\b_to_a_mem[5][1] ),
    .B(\b_to_a_mem[7][1] ),
    .S(_0343_),
    .Z(_0387_));
 NOR2_X1 _1762_ (.A1(_0342_),
    .A2(_0387_),
    .ZN(_0388_));
 OAI33_X1 _1763_ (.A1(_0338_),
    .A2(_0380_),
    .A3(_0383_),
    .B1(_0386_),
    .B2(_0388_),
    .B3(_0337_),
    .ZN(_0389_));
 OAI221_X2 _1764_ (.A(_0322_),
    .B1(_0378_),
    .B2(_0389_),
    .C1(_0825_),
    .C2(net34),
    .ZN(_0390_));
 NAND4_X1 _1765_ (.A1(net6),
    .A2(_0361_),
    .A3(_0819_),
    .A4(_0362_),
    .ZN(_0391_));
 NAND3_X1 _1766_ (.A1(_0319_),
    .A2(net6),
    .A3(_0365_),
    .ZN(_0392_));
 NAND3_X1 _1767_ (.A1(_0390_),
    .A2(_0391_),
    .A3(_0392_),
    .ZN(_0009_));
 MUX2_X1 _1768_ (.A(\b_to_a_mem[8][2] ),
    .B(\b_to_a_mem[10][2] ),
    .S(_0327_),
    .Z(_0393_));
 NOR2_X1 _1769_ (.A1(_0324_),
    .A2(_0393_),
    .ZN(_0394_));
 MUX2_X1 _1770_ (.A(\b_to_a_mem[9][2] ),
    .B(\b_to_a_mem[11][2] ),
    .S(_0349_),
    .Z(_0395_));
 NOR2_X1 _1771_ (.A1(_0331_),
    .A2(_0395_),
    .ZN(_0396_));
 MUX2_X1 _1772_ (.A(\b_to_a_mem[0][2] ),
    .B(\b_to_a_mem[2][2] ),
    .S(_0372_),
    .Z(_0397_));
 NOR2_X1 _1773_ (.A1(_0371_),
    .A2(_0397_),
    .ZN(_0398_));
 MUX2_X1 _1774_ (.A(\b_to_a_mem[1][2] ),
    .B(\b_to_a_mem[3][2] ),
    .S(_0343_),
    .Z(_0399_));
 NOR2_X1 _1775_ (.A1(_0375_),
    .A2(_0399_),
    .ZN(_0400_));
 OAI33_X1 _1776_ (.A1(_0354_),
    .A2(_0394_),
    .A3(_0396_),
    .B1(_0398_),
    .B2(_0400_),
    .B3(_0353_),
    .ZN(_0401_));
 MUX2_X1 _1777_ (.A(\b_to_a_mem[12][2] ),
    .B(\b_to_a_mem[14][2] ),
    .S(_0372_),
    .Z(_0402_));
 NOR2_X1 _1778_ (.A1(_0371_),
    .A2(_0402_),
    .ZN(_0403_));
 MUX2_X1 _1779_ (.A(\b_to_a_mem[13][2] ),
    .B(\b_to_a_mem[15][2] ),
    .S(_0381_),
    .Z(_0404_));
 NOR2_X1 _1780_ (.A1(_0375_),
    .A2(_0404_),
    .ZN(_0405_));
 MUX2_X1 _1781_ (.A(\b_to_a_mem[4][2] ),
    .B(\b_to_a_mem[6][2] ),
    .S(_0339_),
    .Z(_0406_));
 NOR2_X1 _1782_ (.A1(_0384_),
    .A2(_0406_),
    .ZN(_0407_));
 MUX2_X1 _1783_ (.A(\b_to_a_mem[5][2] ),
    .B(\b_to_a_mem[7][2] ),
    .S(_0343_),
    .Z(_0408_));
 NOR2_X1 _1784_ (.A1(_0342_),
    .A2(_0408_),
    .ZN(_0409_));
 OAI33_X1 _1785_ (.A1(_0338_),
    .A2(_0403_),
    .A3(_0405_),
    .B1(_0407_),
    .B2(_0409_),
    .B3(_0337_),
    .ZN(_0410_));
 OAI221_X2 _1786_ (.A(_0322_),
    .B1(_0401_),
    .B2(_0410_),
    .C1(_0825_),
    .C2(net34),
    .ZN(_0411_));
 NAND4_X1 _1787_ (.A1(net7),
    .A2(_0361_),
    .A3(_0819_),
    .A4(_0362_),
    .ZN(_0412_));
 NAND3_X1 _1788_ (.A1(_0319_),
    .A2(net7),
    .A3(_0365_),
    .ZN(_0413_));
 NAND3_X1 _1789_ (.A1(_0411_),
    .A2(_0412_),
    .A3(_0413_),
    .ZN(_0010_));
 MUX2_X1 _1790_ (.A(\b_to_a_mem[8][3] ),
    .B(\b_to_a_mem[10][3] ),
    .S(_0327_),
    .Z(_0414_));
 NOR2_X1 _1791_ (.A1(_0324_),
    .A2(_0414_),
    .ZN(_0415_));
 MUX2_X1 _1792_ (.A(\b_to_a_mem[9][3] ),
    .B(\b_to_a_mem[11][3] ),
    .S(_0349_),
    .Z(_0416_));
 NOR2_X1 _1793_ (.A1(_0331_),
    .A2(_0416_),
    .ZN(_0417_));
 MUX2_X1 _1794_ (.A(\b_to_a_mem[0][3] ),
    .B(\b_to_a_mem[2][3] ),
    .S(_0372_),
    .Z(_0418_));
 NOR2_X1 _1795_ (.A1(_0371_),
    .A2(_0418_),
    .ZN(_0419_));
 MUX2_X1 _1796_ (.A(\b_to_a_mem[1][3] ),
    .B(\b_to_a_mem[3][3] ),
    .S(_0343_),
    .Z(_0420_));
 NOR2_X1 _1797_ (.A1(_0375_),
    .A2(_0420_),
    .ZN(_0421_));
 OAI33_X1 _1798_ (.A1(_0354_),
    .A2(_0415_),
    .A3(_0417_),
    .B1(_0419_),
    .B2(_0421_),
    .B3(_0353_),
    .ZN(_0422_));
 MUX2_X1 _1799_ (.A(\b_to_a_mem[12][3] ),
    .B(\b_to_a_mem[14][3] ),
    .S(_0372_),
    .Z(_0423_));
 NOR2_X1 _1800_ (.A1(_0371_),
    .A2(_0423_),
    .ZN(_0424_));
 MUX2_X1 _1801_ (.A(\b_to_a_mem[13][3] ),
    .B(\b_to_a_mem[15][3] ),
    .S(_0381_),
    .Z(_0425_));
 NOR2_X1 _1802_ (.A1(_0375_),
    .A2(_0425_),
    .ZN(_0426_));
 MUX2_X1 _1803_ (.A(\b_to_a_mem[4][3] ),
    .B(\b_to_a_mem[6][3] ),
    .S(_0339_),
    .Z(_0427_));
 NOR2_X1 _1804_ (.A1(_0384_),
    .A2(_0427_),
    .ZN(_0428_));
 MUX2_X1 _1805_ (.A(\b_to_a_mem[5][3] ),
    .B(\b_to_a_mem[7][3] ),
    .S(_0326_),
    .Z(_0429_));
 NOR2_X1 _1806_ (.A1(_0342_),
    .A2(_0429_),
    .ZN(_0430_));
 OAI33_X1 _1807_ (.A1(_0338_),
    .A2(_0424_),
    .A3(_0426_),
    .B1(_0428_),
    .B2(_0430_),
    .B3(_0337_),
    .ZN(_0431_));
 OAI221_X2 _1808_ (.A(_0322_),
    .B1(_0422_),
    .B2(_0431_),
    .C1(_0825_),
    .C2(net34),
    .ZN(_0432_));
 NAND4_X1 _1809_ (.A1(net8),
    .A2(_0361_),
    .A3(_0819_),
    .A4(_0362_),
    .ZN(_0433_));
 NAND3_X1 _1810_ (.A1(_0319_),
    .A2(net8),
    .A3(_0365_),
    .ZN(_0434_));
 NAND3_X1 _1811_ (.A1(_0432_),
    .A2(_0433_),
    .A3(_0434_),
    .ZN(_0011_));
 MUX2_X1 _1812_ (.A(\b_to_a_mem[8][4] ),
    .B(\b_to_a_mem[10][4] ),
    .S(_0327_),
    .Z(_0435_));
 NOR2_X1 _1813_ (.A1(_0324_),
    .A2(_0435_),
    .ZN(_0436_));
 MUX2_X1 _1814_ (.A(\b_to_a_mem[9][4] ),
    .B(\b_to_a_mem[11][4] ),
    .S(_0349_),
    .Z(_0437_));
 NOR2_X1 _1815_ (.A1(_0331_),
    .A2(_0437_),
    .ZN(_0438_));
 MUX2_X1 _1816_ (.A(\b_to_a_mem[0][4] ),
    .B(\b_to_a_mem[2][4] ),
    .S(_0381_),
    .Z(_0439_));
 NOR2_X1 _1817_ (.A1(_0384_),
    .A2(_0439_),
    .ZN(_0440_));
 MUX2_X1 _1818_ (.A(\b_to_a_mem[1][4] ),
    .B(\b_to_a_mem[3][4] ),
    .S(_0343_),
    .Z(_0441_));
 NOR2_X1 _1819_ (.A1(_0342_),
    .A2(_0441_),
    .ZN(_0442_));
 OAI33_X1 _1820_ (.A1(_0354_),
    .A2(_0436_),
    .A3(_0438_),
    .B1(_0440_),
    .B2(_0442_),
    .B3(_0353_),
    .ZN(_0443_));
 MUX2_X1 _1821_ (.A(\b_to_a_mem[12][4] ),
    .B(\b_to_a_mem[14][4] ),
    .S(_0372_),
    .Z(_0444_));
 NOR2_X1 _1822_ (.A1(_0371_),
    .A2(_0444_),
    .ZN(_0445_));
 MUX2_X1 _1823_ (.A(\b_to_a_mem[13][4] ),
    .B(\b_to_a_mem[15][4] ),
    .S(_0381_),
    .Z(_0446_));
 NOR2_X1 _1824_ (.A1(_0375_),
    .A2(_0446_),
    .ZN(_0447_));
 MUX2_X1 _1825_ (.A(\b_to_a_mem[4][4] ),
    .B(\b_to_a_mem[6][4] ),
    .S(_0339_),
    .Z(_0448_));
 NOR2_X1 _1826_ (.A1(_0384_),
    .A2(_0448_),
    .ZN(_0449_));
 MUX2_X1 _1827_ (.A(\b_to_a_mem[5][4] ),
    .B(\b_to_a_mem[7][4] ),
    .S(_0326_),
    .Z(_0450_));
 NOR2_X1 _1828_ (.A1(_0342_),
    .A2(_0450_),
    .ZN(_0451_));
 OAI33_X1 _1829_ (.A1(_0338_),
    .A2(_0445_),
    .A3(_0447_),
    .B1(_0449_),
    .B2(_0451_),
    .B3(_0337_),
    .ZN(_0452_));
 OAI221_X2 _1830_ (.A(_0322_),
    .B1(_0443_),
    .B2(_0452_),
    .C1(_0825_),
    .C2(net34),
    .ZN(_0453_));
 CLKBUF_X3 _1831_ (.A(_0320_),
    .Z(_0454_));
 NAND4_X1 _1832_ (.A1(net9),
    .A2(_0454_),
    .A3(_0819_),
    .A4(_0362_),
    .ZN(_0455_));
 NAND3_X1 _1833_ (.A1(_0319_),
    .A2(net9),
    .A3(_0365_),
    .ZN(_0456_));
 NAND3_X1 _1834_ (.A1(_0453_),
    .A2(_0455_),
    .A3(_0456_),
    .ZN(_0012_));
 MUX2_X1 _1835_ (.A(\b_to_a_mem[8][5] ),
    .B(\b_to_a_mem[10][5] ),
    .S(_0327_),
    .Z(_0457_));
 NOR2_X1 _1836_ (.A1(_0324_),
    .A2(_0457_),
    .ZN(_0458_));
 MUX2_X1 _1837_ (.A(\b_to_a_mem[9][5] ),
    .B(\b_to_a_mem[11][5] ),
    .S(_0349_),
    .Z(_0459_));
 NOR2_X1 _1838_ (.A1(_0331_),
    .A2(_0459_),
    .ZN(_0460_));
 MUX2_X1 _1839_ (.A(\b_to_a_mem[0][5] ),
    .B(\b_to_a_mem[2][5] ),
    .S(_0381_),
    .Z(_0461_));
 NOR2_X1 _1840_ (.A1(_0384_),
    .A2(_0461_),
    .ZN(_0462_));
 MUX2_X1 _1841_ (.A(\b_to_a_mem[1][5] ),
    .B(\b_to_a_mem[3][5] ),
    .S(_0343_),
    .Z(_0463_));
 NOR2_X1 _1842_ (.A1(_0342_),
    .A2(_0463_),
    .ZN(_0464_));
 OAI33_X1 _1843_ (.A1(_0354_),
    .A2(_0458_),
    .A3(_0460_),
    .B1(_0462_),
    .B2(_0464_),
    .B3(_0353_),
    .ZN(_0465_));
 MUX2_X1 _1844_ (.A(\b_to_a_mem[12][5] ),
    .B(\b_to_a_mem[14][5] ),
    .S(_0372_),
    .Z(_0466_));
 NOR2_X1 _1845_ (.A1(_0371_),
    .A2(_0466_),
    .ZN(_0467_));
 MUX2_X1 _1846_ (.A(\b_to_a_mem[13][5] ),
    .B(\b_to_a_mem[15][5] ),
    .S(_0381_),
    .Z(_0468_));
 NOR2_X1 _1847_ (.A1(_0375_),
    .A2(_0468_),
    .ZN(_0469_));
 MUX2_X1 _1848_ (.A(\b_to_a_mem[4][5] ),
    .B(\b_to_a_mem[6][5] ),
    .S(_0339_),
    .Z(_0470_));
 NOR2_X1 _1849_ (.A1(_0384_),
    .A2(_0470_),
    .ZN(_0471_));
 MUX2_X1 _1850_ (.A(\b_to_a_mem[5][5] ),
    .B(\b_to_a_mem[7][5] ),
    .S(_0326_),
    .Z(_0472_));
 NOR2_X1 _1851_ (.A1(_0342_),
    .A2(_0472_),
    .ZN(_0473_));
 OAI33_X1 _1852_ (.A1(_0338_),
    .A2(_0467_),
    .A3(_0469_),
    .B1(_0471_),
    .B2(_0473_),
    .B3(_0337_),
    .ZN(_0474_));
 OAI221_X2 _1853_ (.A(_0322_),
    .B1(_0465_),
    .B2(_0474_),
    .C1(_0825_),
    .C2(net34),
    .ZN(_0475_));
 NAND4_X1 _1854_ (.A1(net10),
    .A2(_0454_),
    .A3(_0819_),
    .A4(_0362_),
    .ZN(_0476_));
 NAND3_X1 _1855_ (.A1(_0319_),
    .A2(net10),
    .A3(_0365_),
    .ZN(_0477_));
 NAND3_X1 _1856_ (.A1(_0475_),
    .A2(_0476_),
    .A3(_0477_),
    .ZN(_0013_));
 MUX2_X1 _1857_ (.A(\b_to_a_mem[8][6] ),
    .B(\b_to_a_mem[10][6] ),
    .S(_0349_),
    .Z(_0478_));
 NOR2_X1 _1858_ (.A1(_0324_),
    .A2(_0478_),
    .ZN(_0479_));
 MUX2_X1 _1859_ (.A(\b_to_a_mem[9][6] ),
    .B(\b_to_a_mem[11][6] ),
    .S(_0349_),
    .Z(_0480_));
 NOR2_X1 _1860_ (.A1(_0331_),
    .A2(_0480_),
    .ZN(_0481_));
 MUX2_X1 _1861_ (.A(\b_to_a_mem[0][6] ),
    .B(\b_to_a_mem[2][6] ),
    .S(_0381_),
    .Z(_0482_));
 NOR2_X1 _1862_ (.A1(_0384_),
    .A2(_0482_),
    .ZN(_0483_));
 MUX2_X1 _1863_ (.A(\b_to_a_mem[1][6] ),
    .B(\b_to_a_mem[3][6] ),
    .S(_0343_),
    .Z(_0484_));
 NOR2_X1 _1864_ (.A1(_0342_),
    .A2(_0484_),
    .ZN(_0485_));
 OAI33_X1 _1865_ (.A1(_0354_),
    .A2(_0479_),
    .A3(_0481_),
    .B1(_0483_),
    .B2(_0485_),
    .B3(_0353_),
    .ZN(_0486_));
 MUX2_X1 _1866_ (.A(\b_to_a_mem[12][6] ),
    .B(\b_to_a_mem[14][6] ),
    .S(_0372_),
    .Z(_0487_));
 NOR2_X1 _1867_ (.A1(_0371_),
    .A2(_0487_),
    .ZN(_0488_));
 MUX2_X1 _1868_ (.A(\b_to_a_mem[13][6] ),
    .B(\b_to_a_mem[15][6] ),
    .S(_0381_),
    .Z(_0489_));
 NOR2_X1 _1869_ (.A1(_0375_),
    .A2(_0489_),
    .ZN(_0490_));
 MUX2_X1 _1870_ (.A(\b_to_a_mem[4][6] ),
    .B(\b_to_a_mem[6][6] ),
    .S(_0339_),
    .Z(_0491_));
 NOR2_X1 _1871_ (.A1(_0384_),
    .A2(_0491_),
    .ZN(_0492_));
 MUX2_X1 _1872_ (.A(\b_to_a_mem[5][6] ),
    .B(\b_to_a_mem[7][6] ),
    .S(_0326_),
    .Z(_0493_));
 NOR2_X1 _1873_ (.A1(_0330_),
    .A2(_0493_),
    .ZN(_0494_));
 OAI33_X1 _1874_ (.A1(_0338_),
    .A2(_0488_),
    .A3(_0490_),
    .B1(_0492_),
    .B2(_0494_),
    .B3(_0337_),
    .ZN(_0495_));
 OAI221_X2 _1875_ (.A(_0322_),
    .B1(_0486_),
    .B2(_0495_),
    .C1(_0825_),
    .C2(net34),
    .ZN(_0496_));
 NAND4_X1 _1876_ (.A1(net11),
    .A2(_0454_),
    .A3(_0819_),
    .A4(_0362_),
    .ZN(_0497_));
 NAND3_X1 _1877_ (.A1(_0319_),
    .A2(net11),
    .A3(_0365_),
    .ZN(_0498_));
 NAND3_X1 _1878_ (.A1(_0496_),
    .A2(_0497_),
    .A3(_0498_),
    .ZN(_0014_));
 MUX2_X1 _1879_ (.A(\b_to_a_mem[8][7] ),
    .B(\b_to_a_mem[10][7] ),
    .S(_0349_),
    .Z(_0499_));
 NOR2_X1 _1880_ (.A1(_0324_),
    .A2(_0499_),
    .ZN(_0500_));
 MUX2_X1 _1881_ (.A(\b_to_a_mem[9][7] ),
    .B(\b_to_a_mem[11][7] ),
    .S(_0349_),
    .Z(_0501_));
 NOR2_X1 _1882_ (.A1(_0331_),
    .A2(_0501_),
    .ZN(_0502_));
 MUX2_X1 _1883_ (.A(\b_to_a_mem[0][7] ),
    .B(\b_to_a_mem[2][7] ),
    .S(_0381_),
    .Z(_0503_));
 NOR2_X1 _1884_ (.A1(_0384_),
    .A2(_0503_),
    .ZN(_0504_));
 MUX2_X1 _1885_ (.A(\b_to_a_mem[1][7] ),
    .B(\b_to_a_mem[3][7] ),
    .S(_0343_),
    .Z(_0505_));
 NOR2_X1 _1886_ (.A1(_0342_),
    .A2(_0505_),
    .ZN(_0506_));
 OAI33_X1 _1887_ (.A1(_0354_),
    .A2(_0500_),
    .A3(_0502_),
    .B1(_0504_),
    .B2(_0506_),
    .B3(_0353_),
    .ZN(_0507_));
 MUX2_X1 _1888_ (.A(\b_to_a_mem[12][7] ),
    .B(\b_to_a_mem[14][7] ),
    .S(_0372_),
    .Z(_0508_));
 NOR2_X1 _1889_ (.A1(_0371_),
    .A2(_0508_),
    .ZN(_0509_));
 MUX2_X1 _1890_ (.A(\b_to_a_mem[13][7] ),
    .B(\b_to_a_mem[15][7] ),
    .S(_0339_),
    .Z(_0510_));
 NOR2_X1 _1891_ (.A1(_0375_),
    .A2(_0510_),
    .ZN(_0511_));
 MUX2_X1 _1892_ (.A(\b_to_a_mem[4][7] ),
    .B(\b_to_a_mem[6][7] ),
    .S(_0339_),
    .Z(_0512_));
 NOR2_X1 _1893_ (.A1(_0323_),
    .A2(_0512_),
    .ZN(_0513_));
 MUX2_X1 _1894_ (.A(\b_to_a_mem[5][7] ),
    .B(\b_to_a_mem[7][7] ),
    .S(_0326_),
    .Z(_0514_));
 NOR2_X1 _1895_ (.A1(_0330_),
    .A2(_0514_),
    .ZN(_0515_));
 OAI33_X1 _1896_ (.A1(_0338_),
    .A2(_0509_),
    .A3(_0511_),
    .B1(_0513_),
    .B2(_0515_),
    .B3(_0337_),
    .ZN(_0516_));
 OAI221_X2 _1897_ (.A(_0322_),
    .B1(_0507_),
    .B2(_0516_),
    .C1(_0825_),
    .C2(net34),
    .ZN(_0517_));
 NAND4_X1 _1898_ (.A1(net12),
    .A2(_0454_),
    .A3(_0819_),
    .A4(_0362_),
    .ZN(_0518_));
 NAND3_X1 _1899_ (.A1(_0319_),
    .A2(net12),
    .A3(_0365_),
    .ZN(_0519_));
 NAND3_X1 _1900_ (.A1(_0517_),
    .A2(_0518_),
    .A3(_0519_),
    .ZN(_0015_));
 AND2_X1 _1901_ (.A1(_0006_),
    .A2(_0364_),
    .ZN(_0520_));
 CLKBUF_X3 _1902_ (.A(_0321_),
    .Z(_0521_));
 NOR2_X1 _1903_ (.A1(_0331_),
    .A2(_0521_),
    .ZN(_0522_));
 OAI21_X1 _1904_ (.A(_0318_),
    .B1(_0808_),
    .B2(_0825_),
    .ZN(_0523_));
 MUX2_X1 _1905_ (.A(_0520_),
    .B(_0522_),
    .S(_0523_),
    .Z(_0016_));
 BUF_X2 _1906_ (.A(_0320_),
    .Z(_0524_));
 AND2_X1 _1907_ (.A1(_0007_),
    .A2(_0524_),
    .ZN(_0525_));
 AND2_X1 _1908_ (.A1(_0327_),
    .A2(_0364_),
    .ZN(_0526_));
 MUX2_X1 _1909_ (.A(_0525_),
    .B(_0526_),
    .S(_0523_),
    .Z(_0017_));
 CLKBUF_X3 _1910_ (.A(_0321_),
    .Z(_0527_));
 NOR2_X1 _1911_ (.A1(_0352_),
    .A2(_0527_),
    .ZN(_0528_));
 NOR2_X1 _1912_ (.A1(_0334_),
    .A2(_0521_),
    .ZN(_0529_));
 NAND2_X1 _1913_ (.A1(_0318_),
    .A2(_1244_),
    .ZN(_0530_));
 AOI21_X1 _1914_ (.A(_0530_),
    .B1(_0362_),
    .B2(_0818_),
    .ZN(_0531_));
 MUX2_X1 _1915_ (.A(_0528_),
    .B(_0529_),
    .S(_0531_),
    .Z(_0018_));
 NOR2_X1 _1916_ (.A1(_0336_),
    .A2(_0527_),
    .ZN(_0532_));
 NOR2_X1 _1917_ (.A1(_0335_),
    .A2(_0521_),
    .ZN(_0533_));
 NAND4_X1 _1918_ (.A1(_0318_),
    .A2(_0324_),
    .A3(_0327_),
    .A4(_0334_),
    .ZN(_0534_));
 AOI21_X1 _1919_ (.A(_0534_),
    .B1(_0362_),
    .B2(_0818_),
    .ZN(_0535_));
 MUX2_X1 _1920_ (.A(_0532_),
    .B(_0533_),
    .S(_0535_),
    .Z(_0019_));
 AND2_X1 _1921_ (.A1(\a_rd_ptr[4] ),
    .A2(_0524_),
    .ZN(_0536_));
 NOR2_X1 _1922_ (.A1(\a_rd_ptr[4] ),
    .A2(_0521_),
    .ZN(_0537_));
 NAND4_X1 _1923_ (.A1(_0318_),
    .A2(_0334_),
    .A3(_0335_),
    .A4(_1244_),
    .ZN(_0538_));
 AOI21_X1 _1924_ (.A(_0538_),
    .B1(_0900_),
    .B2(_0818_),
    .ZN(_0539_));
 MUX2_X1 _1925_ (.A(_0536_),
    .B(_0537_),
    .S(_0539_),
    .Z(_0020_));
 AND2_X1 _1926_ (.A1(\a_wr_ptr[0] ),
    .A2(_0524_),
    .ZN(_0540_));
 AND2_X1 _1927_ (.A1(_0000_),
    .A2(_0364_),
    .ZN(_0541_));
 AOI21_X2 _1928_ (.A(_0831_),
    .B1(net42),
    .B2(_0838_),
    .ZN(_0542_));
 MUX2_X1 _1929_ (.A(_0540_),
    .B(_0541_),
    .S(_0542_),
    .Z(_0149_));
 AND2_X1 _1930_ (.A1(\a_wr_ptr[1] ),
    .A2(_0524_),
    .ZN(_0543_));
 AND2_X1 _1931_ (.A1(_0001_),
    .A2(_0364_),
    .ZN(_0544_));
 MUX2_X1 _1932_ (.A(_0543_),
    .B(_0544_),
    .S(_0542_),
    .Z(_0150_));
 NOR2_X1 _1933_ (.A1(_0829_),
    .A2(_0527_),
    .ZN(_0545_));
 NOR2_X1 _1934_ (.A1(_0854_),
    .A2(_0521_),
    .ZN(_0546_));
 NAND2_X1 _1935_ (.A1(_0830_),
    .A2(_1251_),
    .ZN(_0547_));
 CLKBUF_X3 _1936_ (.A(_0837_),
    .Z(_0548_));
 AOI21_X1 _1937_ (.A(_0547_),
    .B1(_0548_),
    .B2(net42),
    .ZN(_0549_));
 MUX2_X1 _1938_ (.A(_0545_),
    .B(_0546_),
    .S(_0549_),
    .Z(_0151_));
 AND2_X1 _1939_ (.A1(_0832_),
    .A2(_0524_),
    .ZN(_0550_));
 NOR2_X1 _1940_ (.A1(_0832_),
    .A2(_0521_),
    .ZN(_0551_));
 NAND4_X1 _1941_ (.A1(_0830_),
    .A2(_0854_),
    .A3(\a_wr_ptr[1] ),
    .A4(\a_wr_ptr[0] ),
    .ZN(_0552_));
 AOI21_X1 _1942_ (.A(_0552_),
    .B1(_0548_),
    .B2(net42),
    .ZN(_0553_));
 MUX2_X1 _1943_ (.A(_0550_),
    .B(_0551_),
    .S(_0553_),
    .Z(_0152_));
 AND2_X1 _1944_ (.A1(\a_wr_ptr[4] ),
    .A2(_0524_),
    .ZN(_0554_));
 NOR2_X1 _1945_ (.A1(\a_wr_ptr[4] ),
    .A2(_0521_),
    .ZN(_0555_));
 MUX2_X1 _1946_ (.A(_0554_),
    .B(_0555_),
    .S(_0870_),
    .Z(_0153_));
 BUF_X2 _1947_ (.A(b_rd_en),
    .Z(_0556_));
 INV_X4 _1948_ (.A(_0556_),
    .ZN(_0557_));
 NOR2_X4 _1949_ (.A1(_0557_),
    .A2(_0321_),
    .ZN(_0558_));
 CLKBUF_X3 _1950_ (.A(\b_rd_ptr[0] ),
    .Z(_0559_));
 CLKBUF_X3 _1951_ (.A(_0559_),
    .Z(_0560_));
 CLKBUF_X2 _1952_ (.A(\b_rd_ptr[1] ),
    .Z(_0561_));
 BUF_X4 _1953_ (.A(_0561_),
    .Z(_0562_));
 BUF_X4 _1954_ (.A(_0562_),
    .Z(_0563_));
 MUX2_X1 _1955_ (.A(\a_to_b_mem[4][0] ),
    .B(\a_to_b_mem[6][0] ),
    .S(_0563_),
    .Z(_0564_));
 NOR2_X1 _1956_ (.A1(_0560_),
    .A2(_0564_),
    .ZN(_0565_));
 INV_X2 _1957_ (.A(_0559_),
    .ZN(_0566_));
 CLKBUF_X3 _1958_ (.A(_0566_),
    .Z(_0567_));
 MUX2_X1 _1959_ (.A(\a_to_b_mem[5][0] ),
    .B(\a_to_b_mem[7][0] ),
    .S(_0563_),
    .Z(_0568_));
 NOR2_X1 _1960_ (.A1(_0567_),
    .A2(_0568_),
    .ZN(_0569_));
 CLKBUF_X3 _1961_ (.A(\b_rd_ptr[2] ),
    .Z(_0570_));
 CLKBUF_X3 _1962_ (.A(\b_rd_ptr[3] ),
    .Z(_0571_));
 INV_X2 _1963_ (.A(_0571_),
    .ZN(_0572_));
 NAND2_X4 _1964_ (.A1(_0570_),
    .A2(_0572_),
    .ZN(_0573_));
 NAND2_X4 _1965_ (.A1(_0570_),
    .A2(_0571_),
    .ZN(_0574_));
 BUF_X4 _1966_ (.A(_0561_),
    .Z(_0575_));
 MUX2_X1 _1967_ (.A(\a_to_b_mem[12][0] ),
    .B(\a_to_b_mem[14][0] ),
    .S(_0575_),
    .Z(_0576_));
 NOR2_X1 _1968_ (.A1(_0559_),
    .A2(_0576_),
    .ZN(_0577_));
 CLKBUF_X3 _1969_ (.A(_0566_),
    .Z(_0578_));
 BUF_X4 _1970_ (.A(_0561_),
    .Z(_0579_));
 MUX2_X1 _1971_ (.A(\a_to_b_mem[13][0] ),
    .B(\a_to_b_mem[15][0] ),
    .S(_0579_),
    .Z(_0580_));
 NOR2_X1 _1972_ (.A1(_0578_),
    .A2(_0580_),
    .ZN(_0581_));
 OAI33_X1 _1973_ (.A1(_0565_),
    .A2(_0569_),
    .A3(_0573_),
    .B1(_0574_),
    .B2(_0577_),
    .B3(_0581_),
    .ZN(_0582_));
 MUX2_X1 _1974_ (.A(\a_to_b_mem[0][0] ),
    .B(\a_to_b_mem[2][0] ),
    .S(_0563_),
    .Z(_0583_));
 NOR2_X1 _1975_ (.A1(_0560_),
    .A2(_0583_),
    .ZN(_0584_));
 BUF_X4 _1976_ (.A(_0562_),
    .Z(_0585_));
 MUX2_X1 _1977_ (.A(\a_to_b_mem[1][0] ),
    .B(\a_to_b_mem[3][0] ),
    .S(_0585_),
    .Z(_0586_));
 NOR2_X1 _1978_ (.A1(_0567_),
    .A2(_0586_),
    .ZN(_0587_));
 INV_X1 _1979_ (.A(_0570_),
    .ZN(_0588_));
 NAND2_X2 _1980_ (.A1(_0588_),
    .A2(_0572_),
    .ZN(_0589_));
 NAND2_X2 _1981_ (.A1(_0588_),
    .A2(_0571_),
    .ZN(_0590_));
 MUX2_X1 _1982_ (.A(\a_to_b_mem[8][0] ),
    .B(\a_to_b_mem[10][0] ),
    .S(_0579_),
    .Z(_0591_));
 NOR2_X1 _1983_ (.A1(_0559_),
    .A2(_0591_),
    .ZN(_0592_));
 MUX2_X1 _1984_ (.A(\a_to_b_mem[9][0] ),
    .B(\a_to_b_mem[11][0] ),
    .S(_0562_),
    .Z(_0593_));
 NOR2_X1 _1985_ (.A1(_0566_),
    .A2(_0593_),
    .ZN(_0594_));
 OAI33_X1 _1986_ (.A1(_0584_),
    .A2(_0587_),
    .A3(_0589_),
    .B1(_0590_),
    .B2(_0592_),
    .B3(_0594_),
    .ZN(_0595_));
 OAI221_X2 _1987_ (.A(_0558_),
    .B1(_0582_),
    .B2(_0595_),
    .C1(_0795_),
    .C2(_0817_),
    .ZN(_0596_));
 NAND4_X1 _1988_ (.A1(net22),
    .A2(_0454_),
    .A3(_0810_),
    .A4(_0548_),
    .ZN(_0597_));
 NAND3_X1 _1989_ (.A1(_0557_),
    .A2(net22),
    .A3(_0365_),
    .ZN(_0598_));
 NAND3_X1 _1990_ (.A1(_0596_),
    .A2(_0597_),
    .A3(_0598_),
    .ZN(_0154_));
 MUX2_X1 _1991_ (.A(\a_to_b_mem[8][1] ),
    .B(\a_to_b_mem[10][1] ),
    .S(_0563_),
    .Z(_0599_));
 NOR2_X1 _1992_ (.A1(_0560_),
    .A2(_0599_),
    .ZN(_0600_));
 MUX2_X1 _1993_ (.A(\a_to_b_mem[9][1] ),
    .B(\a_to_b_mem[11][1] ),
    .S(_0585_),
    .Z(_0601_));
 NOR2_X1 _1994_ (.A1(_0567_),
    .A2(_0601_),
    .ZN(_0602_));
 CLKBUF_X3 _1995_ (.A(_0559_),
    .Z(_0603_));
 BUF_X4 _1996_ (.A(_0562_),
    .Z(_0604_));
 MUX2_X1 _1997_ (.A(\a_to_b_mem[0][1] ),
    .B(\a_to_b_mem[2][1] ),
    .S(_0604_),
    .Z(_0605_));
 NOR2_X1 _1998_ (.A1(_0603_),
    .A2(_0605_),
    .ZN(_0606_));
 CLKBUF_X3 _1999_ (.A(_0566_),
    .Z(_0607_));
 MUX2_X1 _2000_ (.A(\a_to_b_mem[1][1] ),
    .B(\a_to_b_mem[3][1] ),
    .S(_0575_),
    .Z(_0608_));
 NOR2_X1 _2001_ (.A1(_0607_),
    .A2(_0608_),
    .ZN(_0609_));
 OAI33_X1 _2002_ (.A1(_0590_),
    .A2(_0600_),
    .A3(_0602_),
    .B1(_0606_),
    .B2(_0609_),
    .B3(_0589_),
    .ZN(_0610_));
 MUX2_X1 _2003_ (.A(\a_to_b_mem[12][1] ),
    .B(\a_to_b_mem[14][1] ),
    .S(_0604_),
    .Z(_0611_));
 NOR2_X1 _2004_ (.A1(_0603_),
    .A2(_0611_),
    .ZN(_0612_));
 BUF_X4 _2005_ (.A(_0562_),
    .Z(_0613_));
 MUX2_X1 _2006_ (.A(\a_to_b_mem[13][1] ),
    .B(\a_to_b_mem[15][1] ),
    .S(_0613_),
    .Z(_0614_));
 NOR2_X1 _2007_ (.A1(_0607_),
    .A2(_0614_),
    .ZN(_0615_));
 CLKBUF_X3 _2008_ (.A(_0559_),
    .Z(_0616_));
 MUX2_X1 _2009_ (.A(\a_to_b_mem[4][1] ),
    .B(\a_to_b_mem[6][1] ),
    .S(_0575_),
    .Z(_0617_));
 NOR2_X1 _2010_ (.A1(_0616_),
    .A2(_0617_),
    .ZN(_0618_));
 MUX2_X1 _2011_ (.A(\a_to_b_mem[5][1] ),
    .B(\a_to_b_mem[7][1] ),
    .S(_0579_),
    .Z(_0619_));
 NOR2_X1 _2012_ (.A1(_0578_),
    .A2(_0619_),
    .ZN(_0620_));
 OAI33_X1 _2013_ (.A1(_0574_),
    .A2(_0612_),
    .A3(_0615_),
    .B1(_0618_),
    .B2(_0620_),
    .B3(_0573_),
    .ZN(_0621_));
 OAI221_X2 _2014_ (.A(_0558_),
    .B1(_0610_),
    .B2(_0621_),
    .C1(_0817_),
    .C2(_0795_),
    .ZN(_0622_));
 NAND4_X1 _2015_ (.A1(net23),
    .A2(_0454_),
    .A3(_0810_),
    .A4(_0548_),
    .ZN(_0623_));
 NAND3_X1 _2016_ (.A1(_0557_),
    .A2(net23),
    .A3(_0365_),
    .ZN(_0624_));
 NAND3_X1 _2017_ (.A1(_0622_),
    .A2(_0623_),
    .A3(_0624_),
    .ZN(_0155_));
 MUX2_X1 _2018_ (.A(\a_to_b_mem[8][2] ),
    .B(\a_to_b_mem[10][2] ),
    .S(_0563_),
    .Z(_0625_));
 NOR2_X1 _2019_ (.A1(_0560_),
    .A2(_0625_),
    .ZN(_0626_));
 MUX2_X1 _2020_ (.A(\a_to_b_mem[9][2] ),
    .B(\a_to_b_mem[11][2] ),
    .S(_0585_),
    .Z(_0627_));
 NOR2_X1 _2021_ (.A1(_0567_),
    .A2(_0627_),
    .ZN(_0628_));
 MUX2_X1 _2022_ (.A(\a_to_b_mem[0][2] ),
    .B(\a_to_b_mem[2][2] ),
    .S(_0604_),
    .Z(_0629_));
 NOR2_X1 _2023_ (.A1(_0603_),
    .A2(_0629_),
    .ZN(_0630_));
 MUX2_X1 _2024_ (.A(\a_to_b_mem[1][2] ),
    .B(\a_to_b_mem[3][2] ),
    .S(_0579_),
    .Z(_0631_));
 NOR2_X1 _2025_ (.A1(_0607_),
    .A2(_0631_),
    .ZN(_0632_));
 OAI33_X1 _2026_ (.A1(_0590_),
    .A2(_0626_),
    .A3(_0628_),
    .B1(_0630_),
    .B2(_0632_),
    .B3(_0589_),
    .ZN(_0633_));
 MUX2_X1 _2027_ (.A(\a_to_b_mem[12][2] ),
    .B(\a_to_b_mem[14][2] ),
    .S(_0604_),
    .Z(_0634_));
 NOR2_X1 _2028_ (.A1(_0603_),
    .A2(_0634_),
    .ZN(_0635_));
 MUX2_X1 _2029_ (.A(\a_to_b_mem[13][2] ),
    .B(\a_to_b_mem[15][2] ),
    .S(_0613_),
    .Z(_0636_));
 NOR2_X1 _2030_ (.A1(_0607_),
    .A2(_0636_),
    .ZN(_0637_));
 MUX2_X1 _2031_ (.A(\a_to_b_mem[4][2] ),
    .B(\a_to_b_mem[6][2] ),
    .S(_0575_),
    .Z(_0638_));
 NOR2_X1 _2032_ (.A1(_0616_),
    .A2(_0638_),
    .ZN(_0639_));
 MUX2_X1 _2033_ (.A(\a_to_b_mem[5][2] ),
    .B(\a_to_b_mem[7][2] ),
    .S(_0579_),
    .Z(_0640_));
 NOR2_X1 _2034_ (.A1(_0578_),
    .A2(_0640_),
    .ZN(_0641_));
 OAI33_X1 _2035_ (.A1(_0574_),
    .A2(_0635_),
    .A3(_0637_),
    .B1(_0639_),
    .B2(_0641_),
    .B3(_0573_),
    .ZN(_0642_));
 OAI221_X2 _2036_ (.A(_0558_),
    .B1(_0633_),
    .B2(_0642_),
    .C1(_0817_),
    .C2(_0795_),
    .ZN(_0643_));
 NAND4_X1 _2037_ (.A1(net24),
    .A2(_0454_),
    .A3(_0810_),
    .A4(_0548_),
    .ZN(_0644_));
 NAND3_X1 _2038_ (.A1(_0557_),
    .A2(net24),
    .A3(_0361_),
    .ZN(_0645_));
 NAND3_X1 _2039_ (.A1(_0643_),
    .A2(_0644_),
    .A3(_0645_),
    .ZN(_0156_));
 MUX2_X1 _2040_ (.A(\a_to_b_mem[8][3] ),
    .B(\a_to_b_mem[10][3] ),
    .S(_0563_),
    .Z(_0646_));
 NOR2_X1 _2041_ (.A1(_0560_),
    .A2(_0646_),
    .ZN(_0647_));
 MUX2_X1 _2042_ (.A(\a_to_b_mem[9][3] ),
    .B(\a_to_b_mem[11][3] ),
    .S(_0585_),
    .Z(_0648_));
 NOR2_X1 _2043_ (.A1(_0567_),
    .A2(_0648_),
    .ZN(_0649_));
 MUX2_X1 _2044_ (.A(\a_to_b_mem[0][3] ),
    .B(\a_to_b_mem[2][3] ),
    .S(_0604_),
    .Z(_0650_));
 NOR2_X1 _2045_ (.A1(_0603_),
    .A2(_0650_),
    .ZN(_0651_));
 MUX2_X1 _2046_ (.A(\a_to_b_mem[1][3] ),
    .B(\a_to_b_mem[3][3] ),
    .S(_0579_),
    .Z(_0652_));
 NOR2_X1 _2047_ (.A1(_0607_),
    .A2(_0652_),
    .ZN(_0653_));
 OAI33_X1 _2048_ (.A1(_0590_),
    .A2(_0647_),
    .A3(_0649_),
    .B1(_0651_),
    .B2(_0653_),
    .B3(_0589_),
    .ZN(_0654_));
 MUX2_X1 _2049_ (.A(\a_to_b_mem[12][3] ),
    .B(\a_to_b_mem[14][3] ),
    .S(_0604_),
    .Z(_0655_));
 NOR2_X1 _2050_ (.A1(_0603_),
    .A2(_0655_),
    .ZN(_0656_));
 MUX2_X1 _2051_ (.A(\a_to_b_mem[13][3] ),
    .B(\a_to_b_mem[15][3] ),
    .S(_0613_),
    .Z(_0657_));
 NOR2_X1 _2052_ (.A1(_0607_),
    .A2(_0657_),
    .ZN(_0658_));
 MUX2_X1 _2053_ (.A(\a_to_b_mem[4][3] ),
    .B(\a_to_b_mem[6][3] ),
    .S(_0575_),
    .Z(_0659_));
 NOR2_X1 _2054_ (.A1(_0616_),
    .A2(_0659_),
    .ZN(_0660_));
 MUX2_X1 _2055_ (.A(\a_to_b_mem[5][3] ),
    .B(\a_to_b_mem[7][3] ),
    .S(_0562_),
    .Z(_0661_));
 NOR2_X1 _2056_ (.A1(_0578_),
    .A2(_0661_),
    .ZN(_0662_));
 OAI33_X1 _2057_ (.A1(_0574_),
    .A2(_0656_),
    .A3(_0658_),
    .B1(_0660_),
    .B2(_0662_),
    .B3(_0573_),
    .ZN(_0663_));
 OAI221_X2 _2058_ (.A(_0558_),
    .B1(_0654_),
    .B2(_0663_),
    .C1(_0817_),
    .C2(_0795_),
    .ZN(_0664_));
 NAND4_X1 _2059_ (.A1(net25),
    .A2(_0454_),
    .A3(_0810_),
    .A4(_0548_),
    .ZN(_0665_));
 NAND3_X1 _2060_ (.A1(_0557_),
    .A2(net25),
    .A3(_0361_),
    .ZN(_0666_));
 NAND3_X1 _2061_ (.A1(_0664_),
    .A2(_0665_),
    .A3(_0666_),
    .ZN(_0157_));
 MUX2_X1 _2062_ (.A(\a_to_b_mem[8][4] ),
    .B(\a_to_b_mem[10][4] ),
    .S(_0563_),
    .Z(_0667_));
 NOR2_X1 _2063_ (.A1(_0560_),
    .A2(_0667_),
    .ZN(_0668_));
 MUX2_X1 _2064_ (.A(\a_to_b_mem[9][4] ),
    .B(\a_to_b_mem[11][4] ),
    .S(_0585_),
    .Z(_0669_));
 NOR2_X1 _2065_ (.A1(_0567_),
    .A2(_0669_),
    .ZN(_0670_));
 MUX2_X1 _2066_ (.A(\a_to_b_mem[0][4] ),
    .B(\a_to_b_mem[2][4] ),
    .S(_0613_),
    .Z(_0671_));
 NOR2_X1 _2067_ (.A1(_0616_),
    .A2(_0671_),
    .ZN(_0672_));
 MUX2_X1 _2068_ (.A(\a_to_b_mem[1][4] ),
    .B(\a_to_b_mem[3][4] ),
    .S(_0579_),
    .Z(_0673_));
 NOR2_X1 _2069_ (.A1(_0578_),
    .A2(_0673_),
    .ZN(_0674_));
 OAI33_X1 _2070_ (.A1(_0590_),
    .A2(_0668_),
    .A3(_0670_),
    .B1(_0672_),
    .B2(_0674_),
    .B3(_0589_),
    .ZN(_0675_));
 MUX2_X1 _2071_ (.A(\a_to_b_mem[12][4] ),
    .B(\a_to_b_mem[14][4] ),
    .S(_0604_),
    .Z(_0676_));
 NOR2_X1 _2072_ (.A1(_0603_),
    .A2(_0676_),
    .ZN(_0677_));
 MUX2_X1 _2073_ (.A(\a_to_b_mem[13][4] ),
    .B(\a_to_b_mem[15][4] ),
    .S(_0613_),
    .Z(_0678_));
 NOR2_X1 _2074_ (.A1(_0607_),
    .A2(_0678_),
    .ZN(_0679_));
 MUX2_X1 _2075_ (.A(\a_to_b_mem[4][4] ),
    .B(\a_to_b_mem[6][4] ),
    .S(_0575_),
    .Z(_0680_));
 NOR2_X1 _2076_ (.A1(_0616_),
    .A2(_0680_),
    .ZN(_0681_));
 MUX2_X1 _2077_ (.A(\a_to_b_mem[5][4] ),
    .B(\a_to_b_mem[7][4] ),
    .S(_0562_),
    .Z(_0682_));
 NOR2_X1 _2078_ (.A1(_0578_),
    .A2(_0682_),
    .ZN(_0683_));
 OAI33_X1 _2079_ (.A1(_0574_),
    .A2(_0677_),
    .A3(_0679_),
    .B1(_0681_),
    .B2(_0683_),
    .B3(_0573_),
    .ZN(_0684_));
 OAI221_X2 _2080_ (.A(_0558_),
    .B1(_0675_),
    .B2(_0684_),
    .C1(_0817_),
    .C2(_0795_),
    .ZN(_0685_));
 NAND4_X1 _2081_ (.A1(net26),
    .A2(_0454_),
    .A3(_0810_),
    .A4(_0548_),
    .ZN(_0686_));
 NAND3_X1 _2082_ (.A1(_0557_),
    .A2(net26),
    .A3(_0361_),
    .ZN(_0687_));
 NAND3_X1 _2083_ (.A1(_0685_),
    .A2(_0686_),
    .A3(_0687_),
    .ZN(_0158_));
 MUX2_X1 _2084_ (.A(\a_to_b_mem[8][5] ),
    .B(\a_to_b_mem[10][5] ),
    .S(_0563_),
    .Z(_0688_));
 NOR2_X1 _2085_ (.A1(_0560_),
    .A2(_0688_),
    .ZN(_0689_));
 MUX2_X1 _2086_ (.A(\a_to_b_mem[9][5] ),
    .B(\a_to_b_mem[11][5] ),
    .S(_0585_),
    .Z(_0690_));
 NOR2_X1 _2087_ (.A1(_0567_),
    .A2(_0690_),
    .ZN(_0691_));
 MUX2_X1 _2088_ (.A(\a_to_b_mem[0][5] ),
    .B(\a_to_b_mem[2][5] ),
    .S(_0613_),
    .Z(_0692_));
 NOR2_X1 _2089_ (.A1(_0616_),
    .A2(_0692_),
    .ZN(_0693_));
 MUX2_X1 _2090_ (.A(\a_to_b_mem[1][5] ),
    .B(\a_to_b_mem[3][5] ),
    .S(_0579_),
    .Z(_0694_));
 NOR2_X1 _2091_ (.A1(_0578_),
    .A2(_0694_),
    .ZN(_0695_));
 OAI33_X1 _2092_ (.A1(_0590_),
    .A2(_0689_),
    .A3(_0691_),
    .B1(_0693_),
    .B2(_0695_),
    .B3(_0589_),
    .ZN(_0696_));
 MUX2_X1 _2093_ (.A(\a_to_b_mem[12][5] ),
    .B(\a_to_b_mem[14][5] ),
    .S(_0604_),
    .Z(_0697_));
 NOR2_X1 _2094_ (.A1(_0603_),
    .A2(_0697_),
    .ZN(_0698_));
 MUX2_X1 _2095_ (.A(\a_to_b_mem[13][5] ),
    .B(\a_to_b_mem[15][5] ),
    .S(_0613_),
    .Z(_0699_));
 NOR2_X1 _2096_ (.A1(_0607_),
    .A2(_0699_),
    .ZN(_0700_));
 MUX2_X1 _2097_ (.A(\a_to_b_mem[4][5] ),
    .B(\a_to_b_mem[6][5] ),
    .S(_0575_),
    .Z(_0701_));
 NOR2_X1 _2098_ (.A1(_0616_),
    .A2(_0701_),
    .ZN(_0702_));
 MUX2_X1 _2099_ (.A(\a_to_b_mem[5][5] ),
    .B(\a_to_b_mem[7][5] ),
    .S(_0562_),
    .Z(_0703_));
 NOR2_X1 _2100_ (.A1(_0578_),
    .A2(_0703_),
    .ZN(_0704_));
 OAI33_X1 _2101_ (.A1(_0574_),
    .A2(_0698_),
    .A3(_0700_),
    .B1(_0702_),
    .B2(_0704_),
    .B3(_0573_),
    .ZN(_0705_));
 OAI221_X2 _2102_ (.A(_0558_),
    .B1(_0696_),
    .B2(_0705_),
    .C1(_0817_),
    .C2(_0795_),
    .ZN(_0706_));
 NAND4_X1 _2103_ (.A1(net27),
    .A2(_0454_),
    .A3(_0810_),
    .A4(_0548_),
    .ZN(_0707_));
 NAND3_X1 _2104_ (.A1(_0557_),
    .A2(net27),
    .A3(_0361_),
    .ZN(_0708_));
 NAND3_X1 _2105_ (.A1(_0706_),
    .A2(_0707_),
    .A3(_0708_),
    .ZN(_0159_));
 MUX2_X1 _2106_ (.A(\a_to_b_mem[8][6] ),
    .B(\a_to_b_mem[10][6] ),
    .S(_0585_),
    .Z(_0709_));
 NOR2_X1 _2107_ (.A1(_0560_),
    .A2(_0709_),
    .ZN(_0710_));
 MUX2_X1 _2108_ (.A(\a_to_b_mem[9][6] ),
    .B(\a_to_b_mem[11][6] ),
    .S(_0585_),
    .Z(_0711_));
 NOR2_X1 _2109_ (.A1(_0567_),
    .A2(_0711_),
    .ZN(_0712_));
 MUX2_X1 _2110_ (.A(\a_to_b_mem[0][6] ),
    .B(\a_to_b_mem[2][6] ),
    .S(_0613_),
    .Z(_0713_));
 NOR2_X1 _2111_ (.A1(_0616_),
    .A2(_0713_),
    .ZN(_0714_));
 MUX2_X1 _2112_ (.A(\a_to_b_mem[1][6] ),
    .B(\a_to_b_mem[3][6] ),
    .S(_0579_),
    .Z(_0715_));
 NOR2_X1 _2113_ (.A1(_0578_),
    .A2(_0715_),
    .ZN(_0716_));
 OAI33_X1 _2114_ (.A1(_0590_),
    .A2(_0710_),
    .A3(_0712_),
    .B1(_0714_),
    .B2(_0716_),
    .B3(_0589_),
    .ZN(_0717_));
 MUX2_X1 _2115_ (.A(\a_to_b_mem[12][6] ),
    .B(\a_to_b_mem[14][6] ),
    .S(_0604_),
    .Z(_0718_));
 NOR2_X1 _2116_ (.A1(_0603_),
    .A2(_0718_),
    .ZN(_0719_));
 MUX2_X1 _2117_ (.A(\a_to_b_mem[13][6] ),
    .B(\a_to_b_mem[15][6] ),
    .S(_0613_),
    .Z(_0720_));
 NOR2_X1 _2118_ (.A1(_0607_),
    .A2(_0720_),
    .ZN(_0721_));
 MUX2_X1 _2119_ (.A(\a_to_b_mem[4][6] ),
    .B(\a_to_b_mem[6][6] ),
    .S(_0575_),
    .Z(_0722_));
 NOR2_X1 _2120_ (.A1(_0616_),
    .A2(_0722_),
    .ZN(_0723_));
 MUX2_X1 _2121_ (.A(\a_to_b_mem[5][6] ),
    .B(\a_to_b_mem[7][6] ),
    .S(_0562_),
    .Z(_0724_));
 NOR2_X1 _2122_ (.A1(_0566_),
    .A2(_0724_),
    .ZN(_0725_));
 OAI33_X1 _2123_ (.A1(_0574_),
    .A2(_0719_),
    .A3(_0721_),
    .B1(_0723_),
    .B2(_0725_),
    .B3(_0573_),
    .ZN(_0726_));
 OAI221_X2 _2124_ (.A(_0558_),
    .B1(_0717_),
    .B2(_0726_),
    .C1(_0817_),
    .C2(_0795_),
    .ZN(_0727_));
 NAND4_X1 _2125_ (.A1(net28),
    .A2(_0364_),
    .A3(_0810_),
    .A4(_0548_),
    .ZN(_0728_));
 NAND3_X1 _2126_ (.A1(_0557_),
    .A2(net28),
    .A3(_0361_),
    .ZN(_0729_));
 NAND3_X1 _2127_ (.A1(_0727_),
    .A2(_0728_),
    .A3(_0729_),
    .ZN(_0160_));
 MUX2_X1 _2128_ (.A(\a_to_b_mem[8][7] ),
    .B(\a_to_b_mem[10][7] ),
    .S(_0585_),
    .Z(_0730_));
 NOR2_X1 _2129_ (.A1(_0560_),
    .A2(_0730_),
    .ZN(_0731_));
 MUX2_X1 _2130_ (.A(\a_to_b_mem[9][7] ),
    .B(\a_to_b_mem[11][7] ),
    .S(_0585_),
    .Z(_0732_));
 NOR2_X1 _2131_ (.A1(_0567_),
    .A2(_0732_),
    .ZN(_0733_));
 MUX2_X1 _2132_ (.A(\a_to_b_mem[0][7] ),
    .B(\a_to_b_mem[2][7] ),
    .S(_0613_),
    .Z(_0734_));
 NOR2_X1 _2133_ (.A1(_0616_),
    .A2(_0734_),
    .ZN(_0735_));
 MUX2_X1 _2134_ (.A(\a_to_b_mem[1][7] ),
    .B(\a_to_b_mem[3][7] ),
    .S(_0579_),
    .Z(_0736_));
 NOR2_X1 _2135_ (.A1(_0578_),
    .A2(_0736_),
    .ZN(_0737_));
 OAI33_X1 _2136_ (.A1(_0590_),
    .A2(_0731_),
    .A3(_0733_),
    .B1(_0735_),
    .B2(_0737_),
    .B3(_0589_),
    .ZN(_0738_));
 MUX2_X1 _2137_ (.A(\a_to_b_mem[12][7] ),
    .B(\a_to_b_mem[14][7] ),
    .S(_0604_),
    .Z(_0739_));
 NOR2_X1 _2138_ (.A1(_0603_),
    .A2(_0739_),
    .ZN(_0740_));
 MUX2_X1 _2139_ (.A(\a_to_b_mem[13][7] ),
    .B(\a_to_b_mem[15][7] ),
    .S(_0575_),
    .Z(_0741_));
 NOR2_X1 _2140_ (.A1(_0607_),
    .A2(_0741_),
    .ZN(_0742_));
 MUX2_X1 _2141_ (.A(\a_to_b_mem[4][7] ),
    .B(\a_to_b_mem[6][7] ),
    .S(_0575_),
    .Z(_0743_));
 NOR2_X1 _2142_ (.A1(_0559_),
    .A2(_0743_),
    .ZN(_0744_));
 MUX2_X1 _2143_ (.A(\a_to_b_mem[5][7] ),
    .B(\a_to_b_mem[7][7] ),
    .S(_0562_),
    .Z(_0745_));
 NOR2_X1 _2144_ (.A1(_0566_),
    .A2(_0745_),
    .ZN(_0746_));
 OAI33_X1 _2145_ (.A1(_0574_),
    .A2(_0740_),
    .A3(_0742_),
    .B1(_0744_),
    .B2(_0746_),
    .B3(_0573_),
    .ZN(_0747_));
 OAI221_X2 _2146_ (.A(_0558_),
    .B1(_0738_),
    .B2(_0747_),
    .C1(_0817_),
    .C2(net42),
    .ZN(_0748_));
 NAND4_X1 _2147_ (.A1(net29),
    .A2(_0364_),
    .A3(_0810_),
    .A4(_0548_),
    .ZN(_0749_));
 NAND3_X1 _2148_ (.A1(_0557_),
    .A2(net29),
    .A3(_0361_),
    .ZN(_0750_));
 NAND3_X1 _2149_ (.A1(_0748_),
    .A2(_0749_),
    .A3(_0750_),
    .ZN(_0161_));
 AND2_X1 _2150_ (.A1(_0002_),
    .A2(_0524_),
    .ZN(_0751_));
 NOR2_X1 _2151_ (.A1(_0567_),
    .A2(_0521_),
    .ZN(_0752_));
 OAI21_X1 _2152_ (.A(_0556_),
    .B1(net42),
    .B2(_0816_),
    .ZN(_0753_));
 MUX2_X1 _2153_ (.A(_0751_),
    .B(_0752_),
    .S(_0753_),
    .Z(_0162_));
 AND2_X1 _2154_ (.A1(_0003_),
    .A2(_0524_),
    .ZN(_0754_));
 AND2_X1 _2155_ (.A1(_0563_),
    .A2(_0364_),
    .ZN(_0755_));
 MUX2_X1 _2156_ (.A(_0754_),
    .B(_0755_),
    .S(_0753_),
    .Z(_0163_));
 NOR2_X1 _2157_ (.A1(_0588_),
    .A2(_0527_),
    .ZN(_0756_));
 NOR2_X1 _2158_ (.A1(_0570_),
    .A2(_0521_),
    .ZN(_0757_));
 NAND2_X1 _2159_ (.A1(_0556_),
    .A2(_1235_),
    .ZN(_0758_));
 AOI21_X1 _2160_ (.A(_0758_),
    .B1(_0838_),
    .B2(_0809_),
    .ZN(_0759_));
 MUX2_X1 _2161_ (.A(_0756_),
    .B(_0757_),
    .S(_0759_),
    .Z(_0164_));
 NOR2_X1 _2162_ (.A1(_0572_),
    .A2(_0527_),
    .ZN(_0760_));
 NOR2_X1 _2163_ (.A1(_0571_),
    .A2(_0521_),
    .ZN(_0761_));
 NAND4_X1 _2164_ (.A1(_0556_),
    .A2(_0560_),
    .A3(_0563_),
    .A4(_0570_),
    .ZN(_0762_));
 AOI21_X1 _2165_ (.A(_0762_),
    .B1(_0838_),
    .B2(_0809_),
    .ZN(_0763_));
 MUX2_X1 _2166_ (.A(_0760_),
    .B(_0761_),
    .S(_0763_),
    .Z(_0165_));
 AND2_X1 _2167_ (.A1(\b_rd_ptr[4] ),
    .A2(_0524_),
    .ZN(_0764_));
 NOR2_X1 _2168_ (.A1(\b_rd_ptr[4] ),
    .A2(_0527_),
    .ZN(_0765_));
 NAND4_X1 _2169_ (.A1(_0556_),
    .A2(_0570_),
    .A3(_0571_),
    .A4(_1235_),
    .ZN(_0766_));
 AOI21_X1 _2170_ (.A(_0766_),
    .B1(_0838_),
    .B2(_0809_),
    .ZN(_0767_));
 MUX2_X1 _2171_ (.A(_0764_),
    .B(_0765_),
    .S(_0767_),
    .Z(_0166_));
 AND2_X1 _2172_ (.A1(\b_wr_ptr[0] ),
    .A2(_0524_),
    .ZN(_0768_));
 AND2_X1 _2173_ (.A1(_0004_),
    .A2(_0364_),
    .ZN(_0769_));
 AOI21_X2 _2174_ (.A(_0893_),
    .B1(_0808_),
    .B2(_0900_),
    .ZN(_0770_));
 MUX2_X1 _2175_ (.A(_0768_),
    .B(_0769_),
    .S(_0770_),
    .Z(_0295_));
 AND2_X1 _2176_ (.A1(\b_wr_ptr[1] ),
    .A2(_0320_),
    .ZN(_0771_));
 AND2_X1 _2177_ (.A1(_0005_),
    .A2(_0364_),
    .ZN(_0772_));
 MUX2_X1 _2178_ (.A(_0771_),
    .B(_0772_),
    .S(_0770_),
    .Z(_0296_));
 NOR2_X1 _2179_ (.A1(_0891_),
    .A2(_0527_),
    .ZN(_0773_));
 NOR2_X1 _2180_ (.A1(_0916_),
    .A2(_0527_),
    .ZN(_0774_));
 NAND2_X1 _2181_ (.A1(_0892_),
    .A2(_1242_),
    .ZN(_0775_));
 AOI21_X1 _2182_ (.A(_0775_),
    .B1(_0900_),
    .B2(_0808_),
    .ZN(_0776_));
 MUX2_X1 _2183_ (.A(_0773_),
    .B(_0774_),
    .S(_0776_),
    .Z(_0297_));
 AND2_X1 _2184_ (.A1(_0894_),
    .A2(_0320_),
    .ZN(_0777_));
 NOR2_X1 _2185_ (.A1(_0894_),
    .A2(_0527_),
    .ZN(_0778_));
 NAND4_X1 _2186_ (.A1(_0892_),
    .A2(_0916_),
    .A3(\b_wr_ptr[1] ),
    .A4(\b_wr_ptr[0] ),
    .ZN(_0779_));
 AOI21_X1 _2187_ (.A(_0779_),
    .B1(_0900_),
    .B2(_0808_),
    .ZN(_0780_));
 MUX2_X1 _2188_ (.A(_0777_),
    .B(_0778_),
    .S(_0780_),
    .Z(_0298_));
 AND2_X1 _2189_ (.A1(\b_wr_ptr[4] ),
    .A2(_0320_),
    .ZN(_0781_));
 NOR2_X1 _2190_ (.A1(\b_wr_ptr[4] ),
    .A2(_0527_),
    .ZN(_0782_));
 MUX2_X1 _2191_ (.A(_0781_),
    .B(_0782_),
    .S(_0932_),
    .Z(_0299_));
 XOR2_X2 _2192_ (.A(_1256_),
    .B(_0820_),
    .Z(_0783_));
 NOR4_X4 _2193_ (.A1(_0808_),
    .A2(net33),
    .A3(net32),
    .A4(_0783_),
    .ZN(net1));
 NAND2_X1 _2194_ (.A1(_0820_),
    .A2(net32),
    .ZN(_0784_));
 OAI21_X4 _2195_ (.A(_0819_),
    .B1(_0784_),
    .B2(_0802_),
    .ZN(net2));
 XOR2_X2 _2196_ (.A(_1254_),
    .B(_0811_),
    .Z(_0785_));
 NOR4_X4 _2197_ (.A1(net15),
    .A2(net16),
    .A3(_0795_),
    .A4(_0785_),
    .ZN(net18));
 NAND2_X1 _2198_ (.A1(_0811_),
    .A2(net15),
    .ZN(_0786_));
 OAI21_X4 _2199_ (.A(_0810_),
    .B1(_0786_),
    .B2(_0790_),
    .ZN(net19));
 FA_X1 _2200_ (.A(_1214_),
    .B(\a_wr_ptr[1] ),
    .CI(_1213_),
    .CO(_1215_),
    .S(net14));
 FA_X1 _2201_ (.A(_1216_),
    .B(_1217_),
    .CI(\b_wr_ptr[1] ),
    .CO(_1218_),
    .S(net31));
 HA_X1 _2202_ (.A(_1219_),
    .B(\b_wr_ptr[3] ),
    .CO(_1220_),
    .S(_1221_));
 HA_X1 _2203_ (.A(_1216_),
    .B(\b_wr_ptr[1] ),
    .CO(_1222_),
    .S(_1223_));
 HA_X1 _2204_ (.A(\a_wr_ptr[3] ),
    .B(_1224_),
    .CO(_1225_),
    .S(_1226_));
 HA_X1 _2205_ (.A(\a_wr_ptr[1] ),
    .B(_1213_),
    .CO(_1227_),
    .S(_1228_));
 HA_X1 _2206_ (.A(\a_wr_ptr[2] ),
    .B(_1229_),
    .CO(_1230_),
    .S(_1231_));
 HA_X1 _2207_ (.A(_1232_),
    .B(\b_wr_ptr[2] ),
    .CO(_1233_),
    .S(_1234_));
 HA_X1 _2208_ (.A(\b_rd_ptr[0] ),
    .B(\b_rd_ptr[1] ),
    .CO(_1235_),
    .S(_0003_));
 HA_X1 _2209_ (.A(_0004_),
    .B(_1236_),
    .CO(_1237_),
    .S(_0005_));
 HA_X1 _2210_ (.A(_0004_),
    .B(\b_wr_ptr[1] ),
    .CO(_1238_),
    .S(_1239_));
 HA_X1 _2211_ (.A(\b_wr_ptr[0] ),
    .B(_1236_),
    .CO(_1240_),
    .S(_1241_));
 HA_X1 _2212_ (.A(\b_wr_ptr[0] ),
    .B(\b_wr_ptr[1] ),
    .CO(_1242_),
    .S(_1243_));
 HA_X1 _2213_ (.A(\a_rd_ptr[0] ),
    .B(\a_rd_ptr[1] ),
    .CO(_1244_),
    .S(_0007_));
 HA_X1 _2214_ (.A(_0000_),
    .B(_1245_),
    .CO(_1246_),
    .S(_0001_));
 HA_X1 _2215_ (.A(_0000_),
    .B(\a_wr_ptr[1] ),
    .CO(_1247_),
    .S(_1248_));
 HA_X1 _2216_ (.A(\a_wr_ptr[0] ),
    .B(_1245_),
    .CO(_1249_),
    .S(_1250_));
 HA_X1 _2217_ (.A(\a_wr_ptr[0] ),
    .B(\a_wr_ptr[1] ),
    .CO(_1251_),
    .S(_1252_));
 HA_X1 _2218_ (.A(_0000_),
    .B(\b_rd_ptr[0] ),
    .CO(_1253_),
    .S(_1254_));
 HA_X1 _2219_ (.A(\a_rd_ptr[0] ),
    .B(_0004_),
    .CO(_1255_),
    .S(_1256_));
 DFF_X2 \a_rd_data_reg[0]$_SDFFE_PN0P_  (.D(_0008_),
    .CK(clknet_leaf_26_clk),
    .Q(net5),
    .QN(_1212_));
 DFF_X2 \a_rd_data_reg[1]$_SDFFE_PN0P_  (.D(_0009_),
    .CK(clknet_leaf_38_clk),
    .Q(net6),
    .QN(_1211_));
 DFF_X2 \a_rd_data_reg[2]$_SDFFE_PN0P_  (.D(_0010_),
    .CK(clknet_leaf_39_clk),
    .Q(net7),
    .QN(_1210_));
 DFF_X2 \a_rd_data_reg[3]$_SDFFE_PN0P_  (.D(_0011_),
    .CK(clknet_leaf_27_clk),
    .Q(net8),
    .QN(_1209_));
 DFF_X2 \a_rd_data_reg[4]$_SDFFE_PN0P_  (.D(_0012_),
    .CK(clknet_leaf_39_clk),
    .Q(net9),
    .QN(_1208_));
 DFF_X2 \a_rd_data_reg[5]$_SDFFE_PN0P_  (.D(_0013_),
    .CK(clknet_leaf_39_clk),
    .Q(net10),
    .QN(_1207_));
 DFF_X2 \a_rd_data_reg[6]$_SDFFE_PN0P_  (.D(_0014_),
    .CK(clknet_leaf_39_clk),
    .Q(net11),
    .QN(_1206_));
 DFF_X2 \a_rd_data_reg[7]$_SDFFE_PN0P_  (.D(_0015_),
    .CK(clknet_leaf_39_clk),
    .Q(net12),
    .QN(_1205_));
 DFF_X2 \a_rd_ptr[0]$_SDFFE_PN0P_  (.D(_0016_),
    .CK(clknet_leaf_39_clk),
    .Q(\a_rd_ptr[0] ),
    .QN(_0006_));
 DFF_X1 \a_rd_ptr[1]$_SDFFE_PN0P_  (.D(_0017_),
    .CK(clknet_leaf_37_clk),
    .Q(\a_rd_ptr[1] ),
    .QN(_1216_));
 DFF_X1 \a_rd_ptr[2]$_SDFFE_PN0P_  (.D(_0018_),
    .CK(clknet_leaf_37_clk),
    .Q(\a_rd_ptr[2] ),
    .QN(_1232_));
 DFF_X1 \a_rd_ptr[3]$_SDFFE_PN0P_  (.D(_0019_),
    .CK(clknet_leaf_39_clk),
    .Q(\a_rd_ptr[3] ),
    .QN(_1219_));
 DFF_X1 \a_rd_ptr[4]$_SDFFE_PN0P_  (.D(_0020_),
    .CK(clknet_leaf_41_clk),
    .Q(\a_rd_ptr[4] ),
    .QN(_1204_));
 DFF_X1 \a_to_b_mem[0][0]$_DFFE_PP_  (.D(_0021_),
    .CK(clknet_leaf_6_clk),
    .Q(\a_to_b_mem[0][0] ),
    .QN(_1203_));
 DFF_X1 \a_to_b_mem[0][1]$_DFFE_PP_  (.D(_0022_),
    .CK(clknet_leaf_2_clk),
    .Q(\a_to_b_mem[0][1] ),
    .QN(_1202_));
 DFF_X1 \a_to_b_mem[0][2]$_DFFE_PP_  (.D(_0023_),
    .CK(clknet_leaf_2_clk),
    .Q(\a_to_b_mem[0][2] ),
    .QN(_1201_));
 DFF_X1 \a_to_b_mem[0][3]$_DFFE_PP_  (.D(_0024_),
    .CK(clknet_leaf_3_clk),
    .Q(\a_to_b_mem[0][3] ),
    .QN(_1200_));
 DFF_X1 \a_to_b_mem[0][4]$_DFFE_PP_  (.D(_0025_),
    .CK(clknet_leaf_4_clk),
    .Q(\a_to_b_mem[0][4] ),
    .QN(_1199_));
 DFF_X1 \a_to_b_mem[0][5]$_DFFE_PP_  (.D(_0026_),
    .CK(clknet_leaf_7_clk),
    .Q(\a_to_b_mem[0][5] ),
    .QN(_1198_));
 DFF_X1 \a_to_b_mem[0][6]$_DFFE_PP_  (.D(_0027_),
    .CK(clknet_leaf_0_clk),
    .Q(\a_to_b_mem[0][6] ),
    .QN(_1197_));
 DFF_X1 \a_to_b_mem[0][7]$_DFFE_PP_  (.D(_0028_),
    .CK(clknet_leaf_2_clk),
    .Q(\a_to_b_mem[0][7] ),
    .QN(_1196_));
 DFF_X1 \a_to_b_mem[10][0]$_DFFE_PP_  (.D(_0029_),
    .CK(clknet_leaf_18_clk),
    .Q(\a_to_b_mem[10][0] ),
    .QN(_1195_));
 DFF_X1 \a_to_b_mem[10][1]$_DFFE_PP_  (.D(_0030_),
    .CK(clknet_leaf_11_clk),
    .Q(\a_to_b_mem[10][1] ),
    .QN(_1194_));
 DFF_X1 \a_to_b_mem[10][2]$_DFFE_PP_  (.D(_0031_),
    .CK(clknet_leaf_11_clk),
    .Q(\a_to_b_mem[10][2] ),
    .QN(_1193_));
 DFF_X1 \a_to_b_mem[10][3]$_DFFE_PP_  (.D(_0032_),
    .CK(clknet_leaf_15_clk),
    .Q(\a_to_b_mem[10][3] ),
    .QN(_1192_));
 DFF_X1 \a_to_b_mem[10][4]$_DFFE_PP_  (.D(_0033_),
    .CK(clknet_leaf_16_clk),
    .Q(\a_to_b_mem[10][4] ),
    .QN(_1191_));
 DFF_X1 \a_to_b_mem[10][5]$_DFFE_PP_  (.D(_0034_),
    .CK(clknet_leaf_16_clk),
    .Q(\a_to_b_mem[10][5] ),
    .QN(_1190_));
 DFF_X1 \a_to_b_mem[10][6]$_DFFE_PP_  (.D(_0035_),
    .CK(clknet_leaf_15_clk),
    .Q(\a_to_b_mem[10][6] ),
    .QN(_1189_));
 DFF_X1 \a_to_b_mem[10][7]$_DFFE_PP_  (.D(_0036_),
    .CK(clknet_leaf_11_clk),
    .Q(\a_to_b_mem[10][7] ),
    .QN(_1188_));
 DFF_X1 \a_to_b_mem[11][0]$_DFFE_PP_  (.D(_0037_),
    .CK(clknet_leaf_18_clk),
    .Q(\a_to_b_mem[11][0] ),
    .QN(_1187_));
 DFF_X1 \a_to_b_mem[11][1]$_DFFE_PP_  (.D(_0038_),
    .CK(clknet_leaf_10_clk),
    .Q(\a_to_b_mem[11][1] ),
    .QN(_1186_));
 DFF_X1 \a_to_b_mem[11][2]$_DFFE_PP_  (.D(_0039_),
    .CK(clknet_leaf_10_clk),
    .Q(\a_to_b_mem[11][2] ),
    .QN(_1185_));
 DFF_X1 \a_to_b_mem[11][3]$_DFFE_PP_  (.D(_0040_),
    .CK(clknet_leaf_12_clk),
    .Q(\a_to_b_mem[11][3] ),
    .QN(_1184_));
 DFF_X1 \a_to_b_mem[11][4]$_DFFE_PP_  (.D(_0041_),
    .CK(clknet_leaf_18_clk),
    .Q(\a_to_b_mem[11][4] ),
    .QN(_1183_));
 DFF_X1 \a_to_b_mem[11][5]$_DFFE_PP_  (.D(_0042_),
    .CK(clknet_leaf_15_clk),
    .Q(\a_to_b_mem[11][5] ),
    .QN(_1182_));
 DFF_X1 \a_to_b_mem[11][6]$_DFFE_PP_  (.D(_0043_),
    .CK(clknet_leaf_12_clk),
    .Q(\a_to_b_mem[11][6] ),
    .QN(_1181_));
 DFF_X1 \a_to_b_mem[11][7]$_DFFE_PP_  (.D(_0044_),
    .CK(clknet_leaf_12_clk),
    .Q(\a_to_b_mem[11][7] ),
    .QN(_1180_));
 DFF_X1 \a_to_b_mem[12][0]$_DFFE_PP_  (.D(_0045_),
    .CK(clknet_leaf_5_clk),
    .Q(\a_to_b_mem[12][0] ),
    .QN(_1179_));
 DFF_X1 \a_to_b_mem[12][1]$_DFFE_PP_  (.D(_0046_),
    .CK(clknet_leaf_1_clk),
    .Q(\a_to_b_mem[12][1] ),
    .QN(_1178_));
 DFF_X1 \a_to_b_mem[12][2]$_DFFE_PP_  (.D(_0047_),
    .CK(clknet_leaf_1_clk),
    .Q(\a_to_b_mem[12][2] ),
    .QN(_1177_));
 DFF_X1 \a_to_b_mem[12][3]$_DFFE_PP_  (.D(_0048_),
    .CK(clknet_leaf_2_clk),
    .Q(\a_to_b_mem[12][3] ),
    .QN(_1176_));
 DFF_X1 \a_to_b_mem[12][4]$_DFFE_PP_  (.D(_0049_),
    .CK(clknet_leaf_5_clk),
    .Q(\a_to_b_mem[12][4] ),
    .QN(_1175_));
 DFF_X1 \a_to_b_mem[12][5]$_DFFE_PP_  (.D(_0050_),
    .CK(clknet_leaf_3_clk),
    .Q(\a_to_b_mem[12][5] ),
    .QN(_1174_));
 DFF_X1 \a_to_b_mem[12][6]$_DFFE_PP_  (.D(_0051_),
    .CK(clknet_leaf_1_clk),
    .Q(\a_to_b_mem[12][6] ),
    .QN(_1173_));
 DFF_X1 \a_to_b_mem[12][7]$_DFFE_PP_  (.D(_0052_),
    .CK(clknet_leaf_9_clk),
    .Q(\a_to_b_mem[12][7] ),
    .QN(_1172_));
 DFF_X1 \a_to_b_mem[13][0]$_DFFE_PP_  (.D(_0053_),
    .CK(clknet_leaf_4_clk),
    .Q(\a_to_b_mem[13][0] ),
    .QN(_1171_));
 DFF_X1 \a_to_b_mem[13][1]$_DFFE_PP_  (.D(_0054_),
    .CK(clknet_leaf_0_clk),
    .Q(\a_to_b_mem[13][1] ),
    .QN(_1170_));
 DFF_X1 \a_to_b_mem[13][2]$_DFFE_PP_  (.D(_0055_),
    .CK(clknet_leaf_8_clk),
    .Q(\a_to_b_mem[13][2] ),
    .QN(_1169_));
 DFF_X1 \a_to_b_mem[13][3]$_DFFE_PP_  (.D(_0056_),
    .CK(clknet_leaf_2_clk),
    .Q(\a_to_b_mem[13][3] ),
    .QN(_1168_));
 DFF_X1 \a_to_b_mem[13][4]$_DFFE_PP_  (.D(_0057_),
    .CK(clknet_leaf_4_clk),
    .Q(\a_to_b_mem[13][4] ),
    .QN(_1167_));
 DFF_X1 \a_to_b_mem[13][5]$_DFFE_PP_  (.D(_0058_),
    .CK(clknet_leaf_3_clk),
    .Q(\a_to_b_mem[13][5] ),
    .QN(_1166_));
 DFF_X1 \a_to_b_mem[13][6]$_DFFE_PP_  (.D(_0059_),
    .CK(clknet_leaf_0_clk),
    .Q(\a_to_b_mem[13][6] ),
    .QN(_1165_));
 DFF_X1 \a_to_b_mem[13][7]$_DFFE_PP_  (.D(_0060_),
    .CK(clknet_leaf_8_clk),
    .Q(\a_to_b_mem[13][7] ),
    .QN(_1164_));
 DFF_X1 \a_to_b_mem[14][0]$_DFFE_PP_  (.D(_0061_),
    .CK(clknet_leaf_5_clk),
    .Q(\a_to_b_mem[14][0] ),
    .QN(_1163_));
 DFF_X1 \a_to_b_mem[14][1]$_DFFE_PP_  (.D(_0062_),
    .CK(clknet_leaf_1_clk),
    .Q(\a_to_b_mem[14][1] ),
    .QN(_1162_));
 DFF_X1 \a_to_b_mem[14][2]$_DFFE_PP_  (.D(_0063_),
    .CK(clknet_leaf_1_clk),
    .Q(\a_to_b_mem[14][2] ),
    .QN(_1161_));
 DFF_X1 \a_to_b_mem[14][3]$_DFFE_PP_  (.D(_0064_),
    .CK(clknet_leaf_8_clk),
    .Q(\a_to_b_mem[14][3] ),
    .QN(_1160_));
 DFF_X1 \a_to_b_mem[14][4]$_DFFE_PP_  (.D(_0065_),
    .CK(clknet_leaf_5_clk),
    .Q(\a_to_b_mem[14][4] ),
    .QN(_1159_));
 DFF_X1 \a_to_b_mem[14][5]$_DFFE_PP_  (.D(_0066_),
    .CK(clknet_leaf_3_clk),
    .Q(\a_to_b_mem[14][5] ),
    .QN(_1158_));
 DFF_X1 \a_to_b_mem[14][6]$_DFFE_PP_  (.D(_0067_),
    .CK(clknet_leaf_2_clk),
    .Q(\a_to_b_mem[14][6] ),
    .QN(_1157_));
 DFF_X1 \a_to_b_mem[14][7]$_DFFE_PP_  (.D(_0068_),
    .CK(clknet_leaf_9_clk),
    .Q(\a_to_b_mem[14][7] ),
    .QN(_1156_));
 DFF_X1 \a_to_b_mem[15][0]$_DFFE_PP_  (.D(_0069_),
    .CK(clknet_leaf_5_clk),
    .Q(\a_to_b_mem[15][0] ),
    .QN(_1155_));
 DFF_X1 \a_to_b_mem[15][1]$_DFFE_PP_  (.D(_0070_),
    .CK(clknet_leaf_0_clk),
    .Q(\a_to_b_mem[15][1] ),
    .QN(_1154_));
 DFF_X1 \a_to_b_mem[15][2]$_DFFE_PP_  (.D(_0071_),
    .CK(clknet_leaf_1_clk),
    .Q(\a_to_b_mem[15][2] ),
    .QN(_1153_));
 DFF_X1 \a_to_b_mem[15][3]$_DFFE_PP_  (.D(_0072_),
    .CK(clknet_leaf_0_clk),
    .Q(\a_to_b_mem[15][3] ),
    .QN(_1152_));
 DFF_X1 \a_to_b_mem[15][4]$_DFFE_PP_  (.D(_0073_),
    .CK(clknet_leaf_4_clk),
    .Q(\a_to_b_mem[15][4] ),
    .QN(_1151_));
 DFF_X1 \a_to_b_mem[15][5]$_DFFE_PP_  (.D(_0074_),
    .CK(clknet_leaf_5_clk),
    .Q(\a_to_b_mem[15][5] ),
    .QN(_1150_));
 DFF_X1 \a_to_b_mem[15][6]$_DFFE_PP_  (.D(_0075_),
    .CK(clknet_leaf_0_clk),
    .Q(\a_to_b_mem[15][6] ),
    .QN(_1149_));
 DFF_X1 \a_to_b_mem[15][7]$_DFFE_PP_  (.D(_0076_),
    .CK(clknet_leaf_1_clk),
    .Q(\a_to_b_mem[15][7] ),
    .QN(_1148_));
 DFF_X1 \a_to_b_mem[1][0]$_DFFE_PP_  (.D(_0077_),
    .CK(clknet_leaf_18_clk),
    .Q(\a_to_b_mem[1][0] ),
    .QN(_1147_));
 DFF_X1 \a_to_b_mem[1][1]$_DFFE_PP_  (.D(_0078_),
    .CK(clknet_leaf_8_clk),
    .Q(\a_to_b_mem[1][1] ),
    .QN(_1146_));
 DFF_X1 \a_to_b_mem[1][2]$_DFFE_PP_  (.D(_0079_),
    .CK(clknet_leaf_8_clk),
    .Q(\a_to_b_mem[1][2] ),
    .QN(_1145_));
 DFF_X1 \a_to_b_mem[1][3]$_DFFE_PP_  (.D(_0080_),
    .CK(clknet_leaf_11_clk),
    .Q(\a_to_b_mem[1][3] ),
    .QN(_1144_));
 DFF_X1 \a_to_b_mem[1][4]$_DFFE_PP_  (.D(_0081_),
    .CK(clknet_leaf_7_clk),
    .Q(\a_to_b_mem[1][4] ),
    .QN(_1143_));
 DFF_X1 \a_to_b_mem[1][5]$_DFFE_PP_  (.D(_0082_),
    .CK(clknet_leaf_7_clk),
    .Q(\a_to_b_mem[1][5] ),
    .QN(_1142_));
 DFF_X1 \a_to_b_mem[1][6]$_DFFE_PP_  (.D(_0083_),
    .CK(clknet_leaf_11_clk),
    .Q(\a_to_b_mem[1][6] ),
    .QN(_1141_));
 DFF_X1 \a_to_b_mem[1][7]$_DFFE_PP_  (.D(_0084_),
    .CK(clknet_leaf_11_clk),
    .Q(\a_to_b_mem[1][7] ),
    .QN(_1140_));
 DFF_X1 \a_to_b_mem[2][0]$_DFFE_PP_  (.D(_0085_),
    .CK(clknet_leaf_6_clk),
    .Q(\a_to_b_mem[2][0] ),
    .QN(_1139_));
 DFF_X1 \a_to_b_mem[2][1]$_DFFE_PP_  (.D(_0086_),
    .CK(clknet_leaf_3_clk),
    .Q(\a_to_b_mem[2][1] ),
    .QN(_1138_));
 DFF_X1 \a_to_b_mem[2][2]$_DFFE_PP_  (.D(_0087_),
    .CK(clknet_leaf_2_clk),
    .Q(\a_to_b_mem[2][2] ),
    .QN(_1137_));
 DFF_X1 \a_to_b_mem[2][3]$_DFFE_PP_  (.D(_0088_),
    .CK(clknet_leaf_3_clk),
    .Q(\a_to_b_mem[2][3] ),
    .QN(_1136_));
 DFF_X1 \a_to_b_mem[2][4]$_DFFE_PP_  (.D(_0089_),
    .CK(clknet_leaf_4_clk),
    .Q(\a_to_b_mem[2][4] ),
    .QN(_1135_));
 DFF_X1 \a_to_b_mem[2][5]$_DFFE_PP_  (.D(_0090_),
    .CK(clknet_leaf_6_clk),
    .Q(\a_to_b_mem[2][5] ),
    .QN(_1134_));
 DFF_X1 \a_to_b_mem[2][6]$_DFFE_PP_  (.D(_0091_),
    .CK(clknet_leaf_0_clk),
    .Q(\a_to_b_mem[2][6] ),
    .QN(_1133_));
 DFF_X1 \a_to_b_mem[2][7]$_DFFE_PP_  (.D(_0092_),
    .CK(clknet_leaf_7_clk),
    .Q(\a_to_b_mem[2][7] ),
    .QN(_1132_));
 DFF_X1 \a_to_b_mem[3][0]$_DFFE_PP_  (.D(_0093_),
    .CK(clknet_leaf_18_clk),
    .Q(\a_to_b_mem[3][0] ),
    .QN(_1131_));
 DFF_X1 \a_to_b_mem[3][1]$_DFFE_PP_  (.D(_0094_),
    .CK(clknet_leaf_8_clk),
    .Q(\a_to_b_mem[3][1] ),
    .QN(_1130_));
 DFF_X1 \a_to_b_mem[3][2]$_DFFE_PP_  (.D(_0095_),
    .CK(clknet_leaf_8_clk),
    .Q(\a_to_b_mem[3][2] ),
    .QN(_1129_));
 DFF_X1 \a_to_b_mem[3][3]$_DFFE_PP_  (.D(_0096_),
    .CK(clknet_leaf_11_clk),
    .Q(\a_to_b_mem[3][3] ),
    .QN(_1128_));
 DFF_X1 \a_to_b_mem[3][4]$_DFFE_PP_  (.D(_0097_),
    .CK(clknet_leaf_18_clk),
    .Q(\a_to_b_mem[3][4] ),
    .QN(_1127_));
 DFF_X1 \a_to_b_mem[3][5]$_DFFE_PP_  (.D(_0098_),
    .CK(clknet_leaf_7_clk),
    .Q(\a_to_b_mem[3][5] ),
    .QN(_1126_));
 DFF_X1 \a_to_b_mem[3][6]$_DFFE_PP_  (.D(_0099_),
    .CK(clknet_leaf_11_clk),
    .Q(\a_to_b_mem[3][6] ),
    .QN(_1125_));
 DFF_X1 \a_to_b_mem[3][7]$_DFFE_PP_  (.D(_0100_),
    .CK(clknet_leaf_7_clk),
    .Q(\a_to_b_mem[3][7] ),
    .QN(_1124_));
 DFF_X1 \a_to_b_mem[4][0]$_DFFE_PP_  (.D(_0101_),
    .CK(clknet_leaf_17_clk),
    .Q(\a_to_b_mem[4][0] ),
    .QN(_1123_));
 DFF_X1 \a_to_b_mem[4][1]$_DFFE_PP_  (.D(_0102_),
    .CK(clknet_leaf_10_clk),
    .Q(\a_to_b_mem[4][1] ),
    .QN(_1122_));
 DFF_X1 \a_to_b_mem[4][2]$_DFFE_PP_  (.D(_0103_),
    .CK(clknet_leaf_9_clk),
    .Q(\a_to_b_mem[4][2] ),
    .QN(_1121_));
 DFF_X1 \a_to_b_mem[4][3]$_DFFE_PP_  (.D(_0104_),
    .CK(clknet_leaf_14_clk),
    .Q(\a_to_b_mem[4][3] ),
    .QN(_1120_));
 DFF_X1 \a_to_b_mem[4][4]$_DFFE_PP_  (.D(_0105_),
    .CK(clknet_leaf_16_clk),
    .Q(\a_to_b_mem[4][4] ),
    .QN(_1119_));
 DFF_X1 \a_to_b_mem[4][5]$_DFFE_PP_  (.D(_0106_),
    .CK(clknet_leaf_14_clk),
    .Q(\a_to_b_mem[4][5] ),
    .QN(_1118_));
 DFF_X1 \a_to_b_mem[4][6]$_DFFE_PP_  (.D(_0107_),
    .CK(clknet_leaf_13_clk),
    .Q(\a_to_b_mem[4][6] ),
    .QN(_1117_));
 DFF_X1 \a_to_b_mem[4][7]$_DFFE_PP_  (.D(_0108_),
    .CK(clknet_leaf_12_clk),
    .Q(\a_to_b_mem[4][7] ),
    .QN(_1116_));
 DFF_X1 \a_to_b_mem[5][0]$_DFFE_PP_  (.D(_0109_),
    .CK(clknet_leaf_17_clk),
    .Q(\a_to_b_mem[5][0] ),
    .QN(_1115_));
 DFF_X1 \a_to_b_mem[5][1]$_DFFE_PP_  (.D(_0110_),
    .CK(clknet_leaf_12_clk),
    .Q(\a_to_b_mem[5][1] ),
    .QN(_1114_));
 DFF_X1 \a_to_b_mem[5][2]$_DFFE_PP_  (.D(_0111_),
    .CK(clknet_leaf_9_clk),
    .Q(\a_to_b_mem[5][2] ),
    .QN(_1113_));
 DFF_X1 \a_to_b_mem[5][3]$_DFFE_PP_  (.D(_0112_),
    .CK(clknet_leaf_14_clk),
    .Q(\a_to_b_mem[5][3] ),
    .QN(_1112_));
 DFF_X1 \a_to_b_mem[5][4]$_DFFE_PP_  (.D(_0113_),
    .CK(clknet_leaf_17_clk),
    .Q(\a_to_b_mem[5][4] ),
    .QN(_1111_));
 DFF_X1 \a_to_b_mem[5][5]$_DFFE_PP_  (.D(_0114_),
    .CK(clknet_leaf_14_clk),
    .Q(\a_to_b_mem[5][5] ),
    .QN(_1110_));
 DFF_X1 \a_to_b_mem[5][6]$_DFFE_PP_  (.D(_0115_),
    .CK(clknet_leaf_13_clk),
    .Q(\a_to_b_mem[5][6] ),
    .QN(_1109_));
 DFF_X1 \a_to_b_mem[5][7]$_DFFE_PP_  (.D(_0116_),
    .CK(clknet_leaf_12_clk),
    .Q(\a_to_b_mem[5][7] ),
    .QN(_1108_));
 DFF_X1 \a_to_b_mem[6][0]$_DFFE_PP_  (.D(_0117_),
    .CK(clknet_leaf_16_clk),
    .Q(\a_to_b_mem[6][0] ),
    .QN(_1107_));
 DFF_X1 \a_to_b_mem[6][1]$_DFFE_PP_  (.D(_0118_),
    .CK(clknet_leaf_10_clk),
    .Q(\a_to_b_mem[6][1] ),
    .QN(_1106_));
 DFF_X1 \a_to_b_mem[6][2]$_DFFE_PP_  (.D(_0119_),
    .CK(clknet_leaf_9_clk),
    .Q(\a_to_b_mem[6][2] ),
    .QN(_1105_));
 DFF_X1 \a_to_b_mem[6][3]$_DFFE_PP_  (.D(_0120_),
    .CK(clknet_leaf_15_clk),
    .Q(\a_to_b_mem[6][3] ),
    .QN(_1104_));
 DFF_X1 \a_to_b_mem[6][4]$_DFFE_PP_  (.D(_0121_),
    .CK(clknet_leaf_16_clk),
    .Q(\a_to_b_mem[6][4] ),
    .QN(_1103_));
 DFF_X1 \a_to_b_mem[6][5]$_DFFE_PP_  (.D(_0122_),
    .CK(clknet_leaf_14_clk),
    .Q(\a_to_b_mem[6][5] ),
    .QN(_1102_));
 DFF_X1 \a_to_b_mem[6][6]$_DFFE_PP_  (.D(_0123_),
    .CK(clknet_leaf_13_clk),
    .Q(\a_to_b_mem[6][6] ),
    .QN(_1101_));
 DFF_X1 \a_to_b_mem[6][7]$_DFFE_PP_  (.D(_0124_),
    .CK(clknet_leaf_12_clk),
    .Q(\a_to_b_mem[6][7] ),
    .QN(_1100_));
 DFF_X1 \a_to_b_mem[7][0]$_DFFE_PP_  (.D(_0125_),
    .CK(clknet_leaf_17_clk),
    .Q(\a_to_b_mem[7][0] ),
    .QN(_1099_));
 DFF_X1 \a_to_b_mem[7][1]$_DFFE_PP_  (.D(_0126_),
    .CK(clknet_leaf_12_clk),
    .Q(\a_to_b_mem[7][1] ),
    .QN(_1098_));
 DFF_X1 \a_to_b_mem[7][2]$_DFFE_PP_  (.D(_0127_),
    .CK(clknet_leaf_9_clk),
    .Q(\a_to_b_mem[7][2] ),
    .QN(_1097_));
 DFF_X1 \a_to_b_mem[7][3]$_DFFE_PP_  (.D(_0128_),
    .CK(clknet_leaf_14_clk),
    .Q(\a_to_b_mem[7][3] ),
    .QN(_1096_));
 DFF_X1 \a_to_b_mem[7][4]$_DFFE_PP_  (.D(_0129_),
    .CK(clknet_leaf_17_clk),
    .Q(\a_to_b_mem[7][4] ),
    .QN(_1095_));
 DFF_X1 \a_to_b_mem[7][5]$_DFFE_PP_  (.D(_0130_),
    .CK(clknet_leaf_14_clk),
    .Q(\a_to_b_mem[7][5] ),
    .QN(_1094_));
 DFF_X1 \a_to_b_mem[7][6]$_DFFE_PP_  (.D(_0131_),
    .CK(clknet_leaf_13_clk),
    .Q(\a_to_b_mem[7][6] ),
    .QN(_1093_));
 DFF_X1 \a_to_b_mem[7][7]$_DFFE_PP_  (.D(_0132_),
    .CK(clknet_leaf_13_clk),
    .Q(\a_to_b_mem[7][7] ),
    .QN(_1092_));
 DFF_X1 \a_to_b_mem[8][0]$_DFFE_PP_  (.D(_0133_),
    .CK(clknet_leaf_18_clk),
    .Q(\a_to_b_mem[8][0] ),
    .QN(_1091_));
 DFF_X1 \a_to_b_mem[8][1]$_DFFE_PP_  (.D(_0134_),
    .CK(clknet_leaf_10_clk),
    .Q(\a_to_b_mem[8][1] ),
    .QN(_1090_));
 DFF_X1 \a_to_b_mem[8][2]$_DFFE_PP_  (.D(_0135_),
    .CK(clknet_leaf_9_clk),
    .Q(\a_to_b_mem[8][2] ),
    .QN(_1089_));
 DFF_X1 \a_to_b_mem[8][3]$_DFFE_PP_  (.D(_0136_),
    .CK(clknet_leaf_15_clk),
    .Q(\a_to_b_mem[8][3] ),
    .QN(_1088_));
 DFF_X1 \a_to_b_mem[8][4]$_DFFE_PP_  (.D(_0137_),
    .CK(clknet_leaf_16_clk),
    .Q(\a_to_b_mem[8][4] ),
    .QN(_1087_));
 DFF_X1 \a_to_b_mem[8][5]$_DFFE_PP_  (.D(_0138_),
    .CK(clknet_leaf_16_clk),
    .Q(\a_to_b_mem[8][5] ),
    .QN(_1086_));
 DFF_X1 \a_to_b_mem[8][6]$_DFFE_PP_  (.D(_0139_),
    .CK(clknet_leaf_14_clk),
    .Q(\a_to_b_mem[8][6] ),
    .QN(_1085_));
 DFF_X1 \a_to_b_mem[8][7]$_DFFE_PP_  (.D(_0140_),
    .CK(clknet_leaf_13_clk),
    .Q(\a_to_b_mem[8][7] ),
    .QN(_1084_));
 DFF_X1 \a_to_b_mem[9][0]$_DFFE_PP_  (.D(_0141_),
    .CK(clknet_leaf_17_clk),
    .Q(\a_to_b_mem[9][0] ),
    .QN(_1083_));
 DFF_X1 \a_to_b_mem[9][1]$_DFFE_PP_  (.D(_0142_),
    .CK(clknet_leaf_10_clk),
    .Q(\a_to_b_mem[9][1] ),
    .QN(_1082_));
 DFF_X1 \a_to_b_mem[9][2]$_DFFE_PP_  (.D(_0143_),
    .CK(clknet_leaf_10_clk),
    .Q(\a_to_b_mem[9][2] ),
    .QN(_1081_));
 DFF_X1 \a_to_b_mem[9][3]$_DFFE_PP_  (.D(_0144_),
    .CK(clknet_leaf_15_clk),
    .Q(\a_to_b_mem[9][3] ),
    .QN(_1080_));
 DFF_X1 \a_to_b_mem[9][4]$_DFFE_PP_  (.D(_0145_),
    .CK(clknet_leaf_16_clk),
    .Q(\a_to_b_mem[9][4] ),
    .QN(_1079_));
 DFF_X1 \a_to_b_mem[9][5]$_DFFE_PP_  (.D(_0146_),
    .CK(clknet_leaf_15_clk),
    .Q(\a_to_b_mem[9][5] ),
    .QN(_1078_));
 DFF_X1 \a_to_b_mem[9][6]$_DFFE_PP_  (.D(_0147_),
    .CK(clknet_leaf_13_clk),
    .Q(\a_to_b_mem[9][6] ),
    .QN(_1077_));
 DFF_X1 \a_to_b_mem[9][7]$_DFFE_PP_  (.D(_0148_),
    .CK(clknet_leaf_12_clk),
    .Q(\a_to_b_mem[9][7] ),
    .QN(_1076_));
 DFF_X2 \a_wr_ptr[0]$_SDFFE_PN0P_  (.D(_0149_),
    .CK(clknet_leaf_40_clk),
    .Q(\a_wr_ptr[0] ),
    .QN(_0000_));
 DFF_X2 \a_wr_ptr[1]$_SDFFE_PN0P_  (.D(_0150_),
    .CK(clknet_leaf_40_clk),
    .Q(\a_wr_ptr[1] ),
    .QN(_1245_));
 DFF_X2 \a_wr_ptr[2]$_SDFFE_PN0P_  (.D(_0151_),
    .CK(clknet_leaf_6_clk),
    .Q(\a_wr_ptr[2] ),
    .QN(_1075_));
 DFF_X1 \a_wr_ptr[3]$_SDFFE_PN0P_  (.D(_0152_),
    .CK(clknet_leaf_19_clk),
    .Q(\a_wr_ptr[3] ),
    .QN(_1074_));
 DFF_X1 \a_wr_ptr[4]$_SDFFE_PN0P_  (.D(_0153_),
    .CK(clknet_leaf_40_clk),
    .Q(\a_wr_ptr[4] ),
    .QN(_1073_));
 DFF_X2 \b_rd_data_reg[0]$_SDFFE_PN0P_  (.D(_0154_),
    .CK(clknet_leaf_40_clk),
    .Q(net22),
    .QN(_1072_));
 DFF_X2 \b_rd_data_reg[1]$_SDFFE_PN0P_  (.D(_0155_),
    .CK(clknet_leaf_40_clk),
    .Q(net23),
    .QN(_1071_));
 DFF_X2 \b_rd_data_reg[2]$_SDFFE_PN0P_  (.D(_0156_),
    .CK(clknet_leaf_3_clk),
    .Q(net24),
    .QN(_1070_));
 DFF_X2 \b_rd_data_reg[3]$_SDFFE_PN0P_  (.D(_0157_),
    .CK(clknet_leaf_41_clk),
    .Q(net25),
    .QN(_1069_));
 DFF_X2 \b_rd_data_reg[4]$_SDFFE_PN0P_  (.D(_0158_),
    .CK(clknet_leaf_4_clk),
    .Q(net26),
    .QN(_1068_));
 DFF_X2 \b_rd_data_reg[5]$_SDFFE_PN0P_  (.D(_0159_),
    .CK(clknet_leaf_4_clk),
    .Q(net27),
    .QN(_1067_));
 DFF_X2 \b_rd_data_reg[6]$_SDFFE_PN0P_  (.D(_0160_),
    .CK(clknet_leaf_4_clk),
    .Q(net28),
    .QN(_1066_));
 DFF_X2 \b_rd_data_reg[7]$_SDFFE_PN0P_  (.D(_0161_),
    .CK(clknet_leaf_3_clk),
    .Q(net29),
    .QN(_1065_));
 DFF_X2 \b_rd_ptr[0]$_SDFFE_PN0P_  (.D(_0162_),
    .CK(clknet_leaf_6_clk),
    .Q(\b_rd_ptr[0] ),
    .QN(_0002_));
 DFF_X1 \b_rd_ptr[1]$_SDFFE_PN0P_  (.D(_0163_),
    .CK(clknet_leaf_6_clk),
    .Q(\b_rd_ptr[1] ),
    .QN(_1213_));
 DFF_X1 \b_rd_ptr[2]$_SDFFE_PN0P_  (.D(_0164_),
    .CK(clknet_leaf_19_clk),
    .Q(\b_rd_ptr[2] ),
    .QN(_1229_));
 DFF_X1 \b_rd_ptr[3]$_SDFFE_PN0P_  (.D(_0165_),
    .CK(clknet_leaf_19_clk),
    .Q(\b_rd_ptr[3] ),
    .QN(_1224_));
 DFF_X1 \b_rd_ptr[4]$_SDFFE_PN0P_  (.D(_0166_),
    .CK(clknet_leaf_40_clk),
    .Q(\b_rd_ptr[4] ),
    .QN(_1064_));
 DFF_X1 \b_to_a_mem[0][0]$_DFFE_PP_  (.D(_0167_),
    .CK(clknet_leaf_37_clk),
    .Q(\b_to_a_mem[0][0] ),
    .QN(_1063_));
 DFF_X1 \b_to_a_mem[0][1]$_DFFE_PP_  (.D(_0168_),
    .CK(clknet_leaf_33_clk),
    .Q(\b_to_a_mem[0][1] ),
    .QN(_1062_));
 DFF_X1 \b_to_a_mem[0][2]$_DFFE_PP_  (.D(_0169_),
    .CK(clknet_leaf_33_clk),
    .Q(\b_to_a_mem[0][2] ),
    .QN(_1061_));
 DFF_X1 \b_to_a_mem[0][3]$_DFFE_PP_  (.D(_0170_),
    .CK(clknet_leaf_32_clk),
    .Q(\b_to_a_mem[0][3] ),
    .QN(_1060_));
 DFF_X1 \b_to_a_mem[0][4]$_DFFE_PP_  (.D(_0171_),
    .CK(clknet_leaf_36_clk),
    .Q(\b_to_a_mem[0][4] ),
    .QN(_1059_));
 DFF_X1 \b_to_a_mem[0][5]$_DFFE_PP_  (.D(_0172_),
    .CK(clknet_leaf_36_clk),
    .Q(\b_to_a_mem[0][5] ),
    .QN(_1058_));
 DFF_X1 \b_to_a_mem[0][6]$_DFFE_PP_  (.D(_0173_),
    .CK(clknet_leaf_36_clk),
    .Q(\b_to_a_mem[0][6] ),
    .QN(_1057_));
 DFF_X1 \b_to_a_mem[0][7]$_DFFE_PP_  (.D(_0174_),
    .CK(clknet_leaf_35_clk),
    .Q(\b_to_a_mem[0][7] ),
    .QN(_1056_));
 DFF_X1 \b_to_a_mem[10][0]$_DFFE_PP_  (.D(_0175_),
    .CK(clknet_leaf_26_clk),
    .Q(\b_to_a_mem[10][0] ),
    .QN(_1055_));
 DFF_X1 \b_to_a_mem[10][1]$_DFFE_PP_  (.D(_0176_),
    .CK(clknet_leaf_31_clk),
    .Q(\b_to_a_mem[10][1] ),
    .QN(_1054_));
 DFF_X1 \b_to_a_mem[10][2]$_DFFE_PP_  (.D(_0177_),
    .CK(clknet_leaf_31_clk),
    .Q(\b_to_a_mem[10][2] ),
    .QN(_1053_));
 DFF_X1 \b_to_a_mem[10][3]$_DFFE_PP_  (.D(_0178_),
    .CK(clknet_leaf_29_clk),
    .Q(\b_to_a_mem[10][3] ),
    .QN(_1052_));
 DFF_X1 \b_to_a_mem[10][4]$_DFFE_PP_  (.D(_0179_),
    .CK(clknet_leaf_24_clk),
    .Q(\b_to_a_mem[10][4] ),
    .QN(_1051_));
 DFF_X1 \b_to_a_mem[10][5]$_DFFE_PP_  (.D(_0180_),
    .CK(clknet_leaf_24_clk),
    .Q(\b_to_a_mem[10][5] ),
    .QN(_1050_));
 DFF_X1 \b_to_a_mem[10][6]$_DFFE_PP_  (.D(_0181_),
    .CK(clknet_leaf_23_clk),
    .Q(\b_to_a_mem[10][6] ),
    .QN(_1049_));
 DFF_X1 \b_to_a_mem[10][7]$_DFFE_PP_  (.D(_0182_),
    .CK(clknet_leaf_22_clk),
    .Q(\b_to_a_mem[10][7] ),
    .QN(_1048_));
 DFF_X1 \b_to_a_mem[11][0]$_DFFE_PP_  (.D(_0183_),
    .CK(clknet_leaf_25_clk),
    .Q(\b_to_a_mem[11][0] ),
    .QN(_1047_));
 DFF_X1 \b_to_a_mem[11][1]$_DFFE_PP_  (.D(_0184_),
    .CK(clknet_leaf_30_clk),
    .Q(\b_to_a_mem[11][1] ),
    .QN(_1046_));
 DFF_X1 \b_to_a_mem[11][2]$_DFFE_PP_  (.D(_0185_),
    .CK(clknet_leaf_30_clk),
    .Q(\b_to_a_mem[11][2] ),
    .QN(_1045_));
 DFF_X1 \b_to_a_mem[11][3]$_DFFE_PP_  (.D(_0186_),
    .CK(clknet_leaf_29_clk),
    .Q(\b_to_a_mem[11][3] ),
    .QN(_1044_));
 DFF_X1 \b_to_a_mem[11][4]$_DFFE_PP_  (.D(_0187_),
    .CK(clknet_leaf_25_clk),
    .Q(\b_to_a_mem[11][4] ),
    .QN(_1043_));
 DFF_X1 \b_to_a_mem[11][5]$_DFFE_PP_  (.D(_0188_),
    .CK(clknet_leaf_25_clk),
    .Q(\b_to_a_mem[11][5] ),
    .QN(_1042_));
 DFF_X1 \b_to_a_mem[11][6]$_DFFE_PP_  (.D(_0189_),
    .CK(clknet_leaf_22_clk),
    .Q(\b_to_a_mem[11][6] ),
    .QN(_1041_));
 DFF_X1 \b_to_a_mem[11][7]$_DFFE_PP_  (.D(_0190_),
    .CK(clknet_leaf_21_clk),
    .Q(\b_to_a_mem[11][7] ),
    .QN(_1040_));
 DFF_X1 \b_to_a_mem[12][0]$_DFFE_PP_  (.D(_0191_),
    .CK(clknet_leaf_38_clk),
    .Q(\b_to_a_mem[12][0] ),
    .QN(_1039_));
 DFF_X1 \b_to_a_mem[12][1]$_DFFE_PP_  (.D(_0192_),
    .CK(clknet_leaf_32_clk),
    .Q(\b_to_a_mem[12][1] ),
    .QN(_1038_));
 DFF_X1 \b_to_a_mem[12][2]$_DFFE_PP_  (.D(_0193_),
    .CK(clknet_leaf_33_clk),
    .Q(\b_to_a_mem[12][2] ),
    .QN(_1037_));
 DFF_X1 \b_to_a_mem[12][3]$_DFFE_PP_  (.D(_0194_),
    .CK(clknet_leaf_32_clk),
    .Q(\b_to_a_mem[12][3] ),
    .QN(_1036_));
 DFF_X1 \b_to_a_mem[12][4]$_DFFE_PP_  (.D(_0195_),
    .CK(clknet_leaf_38_clk),
    .Q(\b_to_a_mem[12][4] ),
    .QN(_1035_));
 DFF_X1 \b_to_a_mem[12][5]$_DFFE_PP_  (.D(_0196_),
    .CK(clknet_leaf_27_clk),
    .Q(\b_to_a_mem[12][5] ),
    .QN(_1034_));
 DFF_X1 \b_to_a_mem[12][6]$_DFFE_PP_  (.D(_0197_),
    .CK(clknet_leaf_27_clk),
    .Q(\b_to_a_mem[12][6] ),
    .QN(_1033_));
 DFF_X1 \b_to_a_mem[12][7]$_DFFE_PP_  (.D(_0198_),
    .CK(clknet_leaf_35_clk),
    .Q(\b_to_a_mem[12][7] ),
    .QN(_1032_));
 DFF_X1 \b_to_a_mem[13][0]$_DFFE_PP_  (.D(_0199_),
    .CK(clknet_leaf_38_clk),
    .Q(\b_to_a_mem[13][0] ),
    .QN(_1031_));
 DFF_X1 \b_to_a_mem[13][1]$_DFFE_PP_  (.D(_0200_),
    .CK(clknet_leaf_34_clk),
    .Q(\b_to_a_mem[13][1] ),
    .QN(_1030_));
 DFF_X1 \b_to_a_mem[13][2]$_DFFE_PP_  (.D(_0201_),
    .CK(clknet_leaf_34_clk),
    .Q(\b_to_a_mem[13][2] ),
    .QN(_1029_));
 DFF_X1 \b_to_a_mem[13][3]$_DFFE_PP_  (.D(_0202_),
    .CK(clknet_leaf_35_clk),
    .Q(\b_to_a_mem[13][3] ),
    .QN(_1028_));
 DFF_X1 \b_to_a_mem[13][4]$_DFFE_PP_  (.D(_0203_),
    .CK(clknet_leaf_35_clk),
    .Q(\b_to_a_mem[13][4] ),
    .QN(_1027_));
 DFF_X1 \b_to_a_mem[13][5]$_DFFE_PP_  (.D(_0204_),
    .CK(clknet_leaf_36_clk),
    .Q(\b_to_a_mem[13][5] ),
    .QN(_1026_));
 DFF_X1 \b_to_a_mem[13][6]$_DFFE_PP_  (.D(_0205_),
    .CK(clknet_leaf_34_clk),
    .Q(\b_to_a_mem[13][6] ),
    .QN(_1025_));
 DFF_X1 \b_to_a_mem[13][7]$_DFFE_PP_  (.D(_0206_),
    .CK(clknet_leaf_31_clk),
    .Q(\b_to_a_mem[13][7] ),
    .QN(_1024_));
 DFF_X1 \b_to_a_mem[14][0]$_DFFE_PP_  (.D(_0207_),
    .CK(clknet_leaf_27_clk),
    .Q(\b_to_a_mem[14][0] ),
    .QN(_1023_));
 DFF_X1 \b_to_a_mem[14][1]$_DFFE_PP_  (.D(_0208_),
    .CK(clknet_leaf_32_clk),
    .Q(\b_to_a_mem[14][1] ),
    .QN(_1022_));
 DFF_X1 \b_to_a_mem[14][2]$_DFFE_PP_  (.D(_0209_),
    .CK(clknet_leaf_33_clk),
    .Q(\b_to_a_mem[14][2] ),
    .QN(_1021_));
 DFF_X1 \b_to_a_mem[14][3]$_DFFE_PP_  (.D(_0210_),
    .CK(clknet_leaf_32_clk),
    .Q(\b_to_a_mem[14][3] ),
    .QN(_1020_));
 DFF_X1 \b_to_a_mem[14][4]$_DFFE_PP_  (.D(_0211_),
    .CK(clknet_leaf_38_clk),
    .Q(\b_to_a_mem[14][4] ),
    .QN(_1019_));
 DFF_X1 \b_to_a_mem[14][5]$_DFFE_PP_  (.D(_0212_),
    .CK(clknet_leaf_27_clk),
    .Q(\b_to_a_mem[14][5] ),
    .QN(_1018_));
 DFF_X1 \b_to_a_mem[14][6]$_DFFE_PP_  (.D(_0213_),
    .CK(clknet_leaf_27_clk),
    .Q(\b_to_a_mem[14][6] ),
    .QN(_1017_));
 DFF_X1 \b_to_a_mem[14][7]$_DFFE_PP_  (.D(_0214_),
    .CK(clknet_leaf_35_clk),
    .Q(\b_to_a_mem[14][7] ),
    .QN(_1016_));
 DFF_X1 \b_to_a_mem[15][0]$_DFFE_PP_  (.D(_0215_),
    .CK(clknet_leaf_38_clk),
    .Q(\b_to_a_mem[15][0] ),
    .QN(_1015_));
 DFF_X1 \b_to_a_mem[15][1]$_DFFE_PP_  (.D(_0216_),
    .CK(clknet_leaf_34_clk),
    .Q(\b_to_a_mem[15][1] ),
    .QN(_1014_));
 DFF_X1 \b_to_a_mem[15][2]$_DFFE_PP_  (.D(_0217_),
    .CK(clknet_leaf_33_clk),
    .Q(\b_to_a_mem[15][2] ),
    .QN(_1013_));
 DFF_X1 \b_to_a_mem[15][3]$_DFFE_PP_  (.D(_0218_),
    .CK(clknet_leaf_35_clk),
    .Q(\b_to_a_mem[15][3] ),
    .QN(_1012_));
 DFF_X1 \b_to_a_mem[15][4]$_DFFE_PP_  (.D(_0219_),
    .CK(clknet_leaf_35_clk),
    .Q(\b_to_a_mem[15][4] ),
    .QN(_1011_));
 DFF_X1 \b_to_a_mem[15][5]$_DFFE_PP_  (.D(_0220_),
    .CK(clknet_leaf_36_clk),
    .Q(\b_to_a_mem[15][5] ),
    .QN(_1010_));
 DFF_X1 \b_to_a_mem[15][6]$_DFFE_PP_  (.D(_0221_),
    .CK(clknet_leaf_34_clk),
    .Q(\b_to_a_mem[15][6] ),
    .QN(_1009_));
 DFF_X1 \b_to_a_mem[15][7]$_DFFE_PP_  (.D(_0222_),
    .CK(clknet_leaf_31_clk),
    .Q(\b_to_a_mem[15][7] ),
    .QN(_1008_));
 DFF_X1 \b_to_a_mem[1][0]$_DFFE_PP_  (.D(_0223_),
    .CK(clknet_leaf_26_clk),
    .Q(\b_to_a_mem[1][0] ),
    .QN(_1007_));
 DFF_X1 \b_to_a_mem[1][1]$_DFFE_PP_  (.D(_0224_),
    .CK(clknet_leaf_32_clk),
    .Q(\b_to_a_mem[1][1] ),
    .QN(_1006_));
 DFF_X1 \b_to_a_mem[1][2]$_DFFE_PP_  (.D(_0225_),
    .CK(clknet_leaf_31_clk),
    .Q(\b_to_a_mem[1][2] ),
    .QN(_1005_));
 DFF_X1 \b_to_a_mem[1][3]$_DFFE_PP_  (.D(_0226_),
    .CK(clknet_leaf_28_clk),
    .Q(\b_to_a_mem[1][3] ),
    .QN(_1004_));
 DFF_X1 \b_to_a_mem[1][4]$_DFFE_PP_  (.D(_0227_),
    .CK(clknet_leaf_26_clk),
    .Q(\b_to_a_mem[1][4] ),
    .QN(_1003_));
 DFF_X1 \b_to_a_mem[1][5]$_DFFE_PP_  (.D(_0228_),
    .CK(clknet_leaf_26_clk),
    .Q(\b_to_a_mem[1][5] ),
    .QN(_1002_));
 DFF_X1 \b_to_a_mem[1][6]$_DFFE_PP_  (.D(_0229_),
    .CK(clknet_leaf_28_clk),
    .Q(\b_to_a_mem[1][6] ),
    .QN(_1001_));
 DFF_X1 \b_to_a_mem[1][7]$_DFFE_PP_  (.D(_0230_),
    .CK(clknet_leaf_28_clk),
    .Q(\b_to_a_mem[1][7] ),
    .QN(_1000_));
 DFF_X1 \b_to_a_mem[2][0]$_DFFE_PP_  (.D(_0231_),
    .CK(clknet_leaf_36_clk),
    .Q(\b_to_a_mem[2][0] ),
    .QN(_0999_));
 DFF_X1 \b_to_a_mem[2][1]$_DFFE_PP_  (.D(_0232_),
    .CK(clknet_leaf_33_clk),
    .Q(\b_to_a_mem[2][1] ),
    .QN(_0998_));
 DFF_X1 \b_to_a_mem[2][2]$_DFFE_PP_  (.D(_0233_),
    .CK(clknet_leaf_33_clk),
    .Q(\b_to_a_mem[2][2] ),
    .QN(_0997_));
 DFF_X1 \b_to_a_mem[2][3]$_DFFE_PP_  (.D(_0234_),
    .CK(clknet_leaf_32_clk),
    .Q(\b_to_a_mem[2][3] ),
    .QN(_0996_));
 DFF_X1 \b_to_a_mem[2][4]$_DFFE_PP_  (.D(_0235_),
    .CK(clknet_leaf_35_clk),
    .Q(\b_to_a_mem[2][4] ),
    .QN(_0995_));
 DFF_X1 \b_to_a_mem[2][5]$_DFFE_PP_  (.D(_0236_),
    .CK(clknet_leaf_36_clk),
    .Q(\b_to_a_mem[2][5] ),
    .QN(_0994_));
 DFF_X1 \b_to_a_mem[2][6]$_DFFE_PP_  (.D(_0237_),
    .CK(clknet_leaf_34_clk),
    .Q(\b_to_a_mem[2][6] ),
    .QN(_0993_));
 DFF_X1 \b_to_a_mem[2][7]$_DFFE_PP_  (.D(_0238_),
    .CK(clknet_leaf_34_clk),
    .Q(\b_to_a_mem[2][7] ),
    .QN(_0992_));
 DFF_X1 \b_to_a_mem[3][0]$_DFFE_PP_  (.D(_0239_),
    .CK(clknet_leaf_26_clk),
    .Q(\b_to_a_mem[3][0] ),
    .QN(_0991_));
 DFF_X1 \b_to_a_mem[3][1]$_DFFE_PP_  (.D(_0240_),
    .CK(clknet_leaf_32_clk),
    .Q(\b_to_a_mem[3][1] ),
    .QN(_0990_));
 DFF_X1 \b_to_a_mem[3][2]$_DFFE_PP_  (.D(_0241_),
    .CK(clknet_leaf_31_clk),
    .Q(\b_to_a_mem[3][2] ),
    .QN(_0989_));
 DFF_X1 \b_to_a_mem[3][3]$_DFFE_PP_  (.D(_0242_),
    .CK(clknet_leaf_28_clk),
    .Q(\b_to_a_mem[3][3] ),
    .QN(_0988_));
 DFF_X1 \b_to_a_mem[3][4]$_DFFE_PP_  (.D(_0243_),
    .CK(clknet_leaf_25_clk),
    .Q(\b_to_a_mem[3][4] ),
    .QN(_0987_));
 DFF_X1 \b_to_a_mem[3][5]$_DFFE_PP_  (.D(_0244_),
    .CK(clknet_leaf_26_clk),
    .Q(\b_to_a_mem[3][5] ),
    .QN(_0986_));
 DFF_X1 \b_to_a_mem[3][6]$_DFFE_PP_  (.D(_0245_),
    .CK(clknet_leaf_28_clk),
    .Q(\b_to_a_mem[3][6] ),
    .QN(_0985_));
 DFF_X1 \b_to_a_mem[3][7]$_DFFE_PP_  (.D(_0246_),
    .CK(clknet_leaf_22_clk),
    .Q(\b_to_a_mem[3][7] ),
    .QN(_0984_));
 DFF_X1 \b_to_a_mem[4][0]$_DFFE_PP_  (.D(_0247_),
    .CK(clknet_leaf_25_clk),
    .Q(\b_to_a_mem[4][0] ),
    .QN(_0983_));
 DFF_X1 \b_to_a_mem[4][1]$_DFFE_PP_  (.D(_0248_),
    .CK(clknet_leaf_29_clk),
    .Q(\b_to_a_mem[4][1] ),
    .QN(_0982_));
 DFF_X1 \b_to_a_mem[4][2]$_DFFE_PP_  (.D(_0249_),
    .CK(clknet_leaf_30_clk),
    .Q(\b_to_a_mem[4][2] ),
    .QN(_0981_));
 DFF_X1 \b_to_a_mem[4][3]$_DFFE_PP_  (.D(_0250_),
    .CK(clknet_leaf_29_clk),
    .Q(\b_to_a_mem[4][3] ),
    .QN(_0980_));
 DFF_X1 \b_to_a_mem[4][4]$_DFFE_PP_  (.D(_0251_),
    .CK(clknet_leaf_21_clk),
    .Q(\b_to_a_mem[4][4] ),
    .QN(_0979_));
 DFF_X1 \b_to_a_mem[4][5]$_DFFE_PP_  (.D(_0252_),
    .CK(clknet_leaf_20_clk),
    .Q(\b_to_a_mem[4][5] ),
    .QN(_0978_));
 DFF_X1 \b_to_a_mem[4][6]$_DFFE_PP_  (.D(_0253_),
    .CK(clknet_leaf_20_clk),
    .Q(\b_to_a_mem[4][6] ),
    .QN(_0977_));
 DFF_X1 \b_to_a_mem[4][7]$_DFFE_PP_  (.D(_0254_),
    .CK(clknet_leaf_21_clk),
    .Q(\b_to_a_mem[4][7] ),
    .QN(_0976_));
 DFF_X1 \b_to_a_mem[5][0]$_DFFE_PP_  (.D(_0255_),
    .CK(clknet_leaf_24_clk),
    .Q(\b_to_a_mem[5][0] ),
    .QN(_0975_));
 DFF_X1 \b_to_a_mem[5][1]$_DFFE_PP_  (.D(_0256_),
    .CK(clknet_leaf_22_clk),
    .Q(\b_to_a_mem[5][1] ),
    .QN(_0974_));
 DFF_X1 \b_to_a_mem[5][2]$_DFFE_PP_  (.D(_0257_),
    .CK(clknet_leaf_28_clk),
    .Q(\b_to_a_mem[5][2] ),
    .QN(_0973_));
 DFF_X1 \b_to_a_mem[5][3]$_DFFE_PP_  (.D(_0258_),
    .CK(clknet_leaf_22_clk),
    .Q(\b_to_a_mem[5][3] ),
    .QN(_0972_));
 DFF_X1 \b_to_a_mem[5][4]$_DFFE_PP_  (.D(_0259_),
    .CK(clknet_leaf_23_clk),
    .Q(\b_to_a_mem[5][4] ),
    .QN(_0971_));
 DFF_X1 \b_to_a_mem[5][5]$_DFFE_PP_  (.D(_0260_),
    .CK(clknet_leaf_24_clk),
    .Q(\b_to_a_mem[5][5] ),
    .QN(_0970_));
 DFF_X1 \b_to_a_mem[5][6]$_DFFE_PP_  (.D(_0261_),
    .CK(clknet_leaf_23_clk),
    .Q(\b_to_a_mem[5][6] ),
    .QN(_0969_));
 DFF_X1 \b_to_a_mem[5][7]$_DFFE_PP_  (.D(_0262_),
    .CK(clknet_leaf_22_clk),
    .Q(\b_to_a_mem[5][7] ),
    .QN(_0968_));
 DFF_X1 \b_to_a_mem[6][0]$_DFFE_PP_  (.D(_0263_),
    .CK(clknet_leaf_19_clk),
    .Q(\b_to_a_mem[6][0] ),
    .QN(_0967_));
 DFF_X1 \b_to_a_mem[6][1]$_DFFE_PP_  (.D(_0264_),
    .CK(clknet_leaf_30_clk),
    .Q(\b_to_a_mem[6][1] ),
    .QN(_0966_));
 DFF_X1 \b_to_a_mem[6][2]$_DFFE_PP_  (.D(_0265_),
    .CK(clknet_leaf_30_clk),
    .Q(\b_to_a_mem[6][2] ),
    .QN(_0965_));
 DFF_X1 \b_to_a_mem[6][3]$_DFFE_PP_  (.D(_0266_),
    .CK(clknet_leaf_29_clk),
    .Q(\b_to_a_mem[6][3] ),
    .QN(_0964_));
 DFF_X1 \b_to_a_mem[6][4]$_DFFE_PP_  (.D(_0267_),
    .CK(clknet_leaf_20_clk),
    .Q(\b_to_a_mem[6][4] ),
    .QN(_0963_));
 DFF_X1 \b_to_a_mem[6][5]$_DFFE_PP_  (.D(_0268_),
    .CK(clknet_leaf_20_clk),
    .Q(\b_to_a_mem[6][5] ),
    .QN(_0962_));
 DFF_X1 \b_to_a_mem[6][6]$_DFFE_PP_  (.D(_0269_),
    .CK(clknet_leaf_20_clk),
    .Q(\b_to_a_mem[6][6] ),
    .QN(_0961_));
 DFF_X1 \b_to_a_mem[6][7]$_DFFE_PP_  (.D(_0270_),
    .CK(clknet_leaf_21_clk),
    .Q(\b_to_a_mem[6][7] ),
    .QN(_0960_));
 DFF_X1 \b_to_a_mem[7][0]$_DFFE_PP_  (.D(_0271_),
    .CK(clknet_leaf_19_clk),
    .Q(\b_to_a_mem[7][0] ),
    .QN(_0959_));
 DFF_X1 \b_to_a_mem[7][1]$_DFFE_PP_  (.D(_0272_),
    .CK(clknet_leaf_28_clk),
    .Q(\b_to_a_mem[7][1] ),
    .QN(_0958_));
 DFF_X1 \b_to_a_mem[7][2]$_DFFE_PP_  (.D(_0273_),
    .CK(clknet_leaf_29_clk),
    .Q(\b_to_a_mem[7][2] ),
    .QN(_0957_));
 DFF_X1 \b_to_a_mem[7][3]$_DFFE_PP_  (.D(_0274_),
    .CK(clknet_leaf_21_clk),
    .Q(\b_to_a_mem[7][3] ),
    .QN(_0956_));
 DFF_X1 \b_to_a_mem[7][4]$_DFFE_PP_  (.D(_0275_),
    .CK(clknet_leaf_23_clk),
    .Q(\b_to_a_mem[7][4] ),
    .QN(_0955_));
 DFF_X1 \b_to_a_mem[7][5]$_DFFE_PP_  (.D(_0276_),
    .CK(clknet_leaf_23_clk),
    .Q(\b_to_a_mem[7][5] ),
    .QN(_0954_));
 DFF_X1 \b_to_a_mem[7][6]$_DFFE_PP_  (.D(_0277_),
    .CK(clknet_leaf_23_clk),
    .Q(\b_to_a_mem[7][6] ),
    .QN(_0953_));
 DFF_X1 \b_to_a_mem[7][7]$_DFFE_PP_  (.D(_0278_),
    .CK(clknet_leaf_20_clk),
    .Q(\b_to_a_mem[7][7] ),
    .QN(_0952_));
 DFF_X1 \b_to_a_mem[8][0]$_DFFE_PP_  (.D(_0279_),
    .CK(clknet_leaf_25_clk),
    .Q(\b_to_a_mem[8][0] ),
    .QN(_0951_));
 DFF_X1 \b_to_a_mem[8][1]$_DFFE_PP_  (.D(_0280_),
    .CK(clknet_leaf_29_clk),
    .Q(\b_to_a_mem[8][1] ),
    .QN(_0950_));
 DFF_X1 \b_to_a_mem[8][2]$_DFFE_PP_  (.D(_0281_),
    .CK(clknet_leaf_31_clk),
    .Q(\b_to_a_mem[8][2] ),
    .QN(_0949_));
 DFF_X1 \b_to_a_mem[8][3]$_DFFE_PP_  (.D(_0282_),
    .CK(clknet_leaf_29_clk),
    .Q(\b_to_a_mem[8][3] ),
    .QN(_0948_));
 DFF_X1 \b_to_a_mem[8][4]$_DFFE_PP_  (.D(_0283_),
    .CK(clknet_leaf_24_clk),
    .Q(\b_to_a_mem[8][4] ),
    .QN(_0947_));
 DFF_X1 \b_to_a_mem[8][5]$_DFFE_PP_  (.D(_0284_),
    .CK(clknet_leaf_24_clk),
    .Q(\b_to_a_mem[8][5] ),
    .QN(_0946_));
 DFF_X1 \b_to_a_mem[8][6]$_DFFE_PP_  (.D(_0285_),
    .CK(clknet_leaf_23_clk),
    .Q(\b_to_a_mem[8][6] ),
    .QN(_0945_));
 DFF_X1 \b_to_a_mem[8][7]$_DFFE_PP_  (.D(_0286_),
    .CK(clknet_leaf_20_clk),
    .Q(\b_to_a_mem[8][7] ),
    .QN(_0944_));
 DFF_X1 \b_to_a_mem[9][0]$_DFFE_PP_  (.D(_0287_),
    .CK(clknet_leaf_25_clk),
    .Q(\b_to_a_mem[9][0] ),
    .QN(_0943_));
 DFF_X1 \b_to_a_mem[9][1]$_DFFE_PP_  (.D(_0288_),
    .CK(clknet_leaf_30_clk),
    .Q(\b_to_a_mem[9][1] ),
    .QN(_0942_));
 DFF_X1 \b_to_a_mem[9][2]$_DFFE_PP_  (.D(_0289_),
    .CK(clknet_leaf_30_clk),
    .Q(\b_to_a_mem[9][2] ),
    .QN(_0941_));
 DFF_X1 \b_to_a_mem[9][3]$_DFFE_PP_  (.D(_0290_),
    .CK(clknet_leaf_21_clk),
    .Q(\b_to_a_mem[9][3] ),
    .QN(_0940_));
 DFF_X1 \b_to_a_mem[9][4]$_DFFE_PP_  (.D(_0291_),
    .CK(clknet_leaf_24_clk),
    .Q(\b_to_a_mem[9][4] ),
    .QN(_0939_));
 DFF_X1 \b_to_a_mem[9][5]$_DFFE_PP_  (.D(_0292_),
    .CK(clknet_leaf_25_clk),
    .Q(\b_to_a_mem[9][5] ),
    .QN(_0938_));
 DFF_X1 \b_to_a_mem[9][6]$_DFFE_PP_  (.D(_0293_),
    .CK(clknet_leaf_22_clk),
    .Q(\b_to_a_mem[9][6] ),
    .QN(_0937_));
 DFF_X1 \b_to_a_mem[9][7]$_DFFE_PP_  (.D(_0294_),
    .CK(clknet_leaf_21_clk),
    .Q(\b_to_a_mem[9][7] ),
    .QN(_0936_));
 DFF_X2 \b_wr_ptr[0]$_SDFFE_PN0P_  (.D(_0295_),
    .CK(clknet_leaf_37_clk),
    .Q(\b_wr_ptr[0] ),
    .QN(_0004_));
 DFF_X2 \b_wr_ptr[1]$_SDFFE_PN0P_  (.D(_0296_),
    .CK(clknet_leaf_37_clk),
    .Q(\b_wr_ptr[1] ),
    .QN(_1236_));
 DFF_X2 \b_wr_ptr[2]$_SDFFE_PN0P_  (.D(_0297_),
    .CK(clknet_leaf_37_clk),
    .Q(\b_wr_ptr[2] ),
    .QN(_0935_));
 DFF_X1 \b_wr_ptr[3]$_SDFFE_PN0P_  (.D(_0298_),
    .CK(clknet_leaf_41_clk),
    .Q(\b_wr_ptr[3] ),
    .QN(_0934_));
 DFF_X1 \b_wr_ptr[4]$_SDFFE_PN0P_  (.D(_0299_),
    .CK(clknet_leaf_41_clk),
    .Q(\b_wr_ptr[4] ),
    .QN(_0933_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Right_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Right_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Right_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Right_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Right_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Right_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Right_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Right_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Right_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Right_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Right_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Right_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Right_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Right_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Right_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Right_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Right_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Right_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Right_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Right_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Right_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Right_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Right_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Right_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Right_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Right_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Right_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Right_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Right_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Right_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Right_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Right_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Right_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Right_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Right_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Right_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Right_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Right_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Right_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Right_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Right_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Right_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Right_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Right_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Right_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Right_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Right_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Right_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Right_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Right_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Right_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Right_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Right_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Right_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Right_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Right_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Right_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Right_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Right_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Right_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Right_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Right_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Right_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Right_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Right_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Right_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Right_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Right_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Right_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Right_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Right_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Right_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Right_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Right_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Right_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Right_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Right_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Right_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Right_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Right_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Right_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Right_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Right_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_238_Right_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_239_Right_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_240_Right_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_241_Right_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_242_Right_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_243_Right_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_244_Right_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_245_Right_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_246_Right_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_247_Right_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_248_Right_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_249_Right_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_250_Right_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_251_Right_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_252_Right_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_253_Right_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_254_Right_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_255_Right_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_256_Right_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_257_Right_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_258_Right_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_259_Right_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_260_Right_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_261_Right_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_262_Right_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_263_Right_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_264_Right_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_265_Right_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_266_Right_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_267_Right_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_268_Right_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_269_Right_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_270_Right_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_271_Right_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_272_Right_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_273_Right_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_274_Right_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_275_Right_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_276_Right_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_277_Right_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_278_Right_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_279_Right_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_280_Right_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_281_Right_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_282_Right_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_283_Right_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_284_Right_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_285_Right_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_286_Right_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_287_Right_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_288_Right_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_289_Right_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_290_Right_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_291_Right_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_292_Right_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_293_Right_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_294_Right_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_295_Right_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_296_Right_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_297_Right_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_298_Right_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_299_Right_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_300_Right_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_301_Right_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_302_Right_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_303_Right_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_304_Right_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_305_Right_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_306_Right_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_307_Right_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_308_Right_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_309_Right_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_310_Right_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_311_Right_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_312_Right_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_313_Right_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_314_Right_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_315_Right_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_316_Right_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_317_Right_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_318_Right_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_319_Right_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_320_Right_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_321_Right_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_322_Right_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_323_Right_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_324_Right_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_325_Right_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_326_Right_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_327_Right_327 ();
 TAPCELL_X1 PHY_EDGE_ROW_328_Right_328 ();
 TAPCELL_X1 PHY_EDGE_ROW_329_Right_329 ();
 TAPCELL_X1 PHY_EDGE_ROW_330_Right_330 ();
 TAPCELL_X1 PHY_EDGE_ROW_331_Right_331 ();
 TAPCELL_X1 PHY_EDGE_ROW_332_Right_332 ();
 TAPCELL_X1 PHY_EDGE_ROW_333_Right_333 ();
 TAPCELL_X1 PHY_EDGE_ROW_334_Right_334 ();
 TAPCELL_X1 PHY_EDGE_ROW_335_Right_335 ();
 TAPCELL_X1 PHY_EDGE_ROW_336_Right_336 ();
 TAPCELL_X1 PHY_EDGE_ROW_337_Right_337 ();
 TAPCELL_X1 PHY_EDGE_ROW_338_Right_338 ();
 TAPCELL_X1 PHY_EDGE_ROW_339_Right_339 ();
 TAPCELL_X1 PHY_EDGE_ROW_340_Right_340 ();
 TAPCELL_X1 PHY_EDGE_ROW_341_Right_341 ();
 TAPCELL_X1 PHY_EDGE_ROW_342_Right_342 ();
 TAPCELL_X1 PHY_EDGE_ROW_343_Right_343 ();
 TAPCELL_X1 PHY_EDGE_ROW_344_Right_344 ();
 TAPCELL_X1 PHY_EDGE_ROW_345_Right_345 ();
 TAPCELL_X1 PHY_EDGE_ROW_346_Right_346 ();
 TAPCELL_X1 PHY_EDGE_ROW_347_Right_347 ();
 TAPCELL_X1 PHY_EDGE_ROW_348_Right_348 ();
 TAPCELL_X1 PHY_EDGE_ROW_349_Right_349 ();
 TAPCELL_X1 PHY_EDGE_ROW_350_Right_350 ();
 TAPCELL_X1 PHY_EDGE_ROW_351_Right_351 ();
 TAPCELL_X1 PHY_EDGE_ROW_352_Right_352 ();
 TAPCELL_X1 PHY_EDGE_ROW_353_Right_353 ();
 TAPCELL_X1 PHY_EDGE_ROW_354_Right_354 ();
 TAPCELL_X1 PHY_EDGE_ROW_355_Right_355 ();
 TAPCELL_X1 PHY_EDGE_ROW_356_Right_356 ();
 TAPCELL_X1 PHY_EDGE_ROW_357_Right_357 ();
 TAPCELL_X1 PHY_EDGE_ROW_358_Right_358 ();
 TAPCELL_X1 PHY_EDGE_ROW_359_Right_359 ();
 TAPCELL_X1 PHY_EDGE_ROW_360_Right_360 ();
 TAPCELL_X1 PHY_EDGE_ROW_361_Right_361 ();
 TAPCELL_X1 PHY_EDGE_ROW_362_Right_362 ();
 TAPCELL_X1 PHY_EDGE_ROW_363_Right_363 ();
 TAPCELL_X1 PHY_EDGE_ROW_364_Right_364 ();
 TAPCELL_X1 PHY_EDGE_ROW_365_Right_365 ();
 TAPCELL_X1 PHY_EDGE_ROW_366_Right_366 ();
 TAPCELL_X1 PHY_EDGE_ROW_367_Right_367 ();
 TAPCELL_X1 PHY_EDGE_ROW_368_Right_368 ();
 TAPCELL_X1 PHY_EDGE_ROW_369_Right_369 ();
 TAPCELL_X1 PHY_EDGE_ROW_370_Right_370 ();
 TAPCELL_X1 PHY_EDGE_ROW_371_Right_371 ();
 TAPCELL_X1 PHY_EDGE_ROW_372_Right_372 ();
 TAPCELL_X1 PHY_EDGE_ROW_373_Right_373 ();
 TAPCELL_X1 PHY_EDGE_ROW_374_Right_374 ();
 TAPCELL_X1 PHY_EDGE_ROW_375_Right_375 ();
 TAPCELL_X1 PHY_EDGE_ROW_376_Right_376 ();
 TAPCELL_X1 PHY_EDGE_ROW_377_Right_377 ();
 TAPCELL_X1 PHY_EDGE_ROW_378_Right_378 ();
 TAPCELL_X1 PHY_EDGE_ROW_379_Right_379 ();
 TAPCELL_X1 PHY_EDGE_ROW_380_Right_380 ();
 TAPCELL_X1 PHY_EDGE_ROW_381_Right_381 ();
 TAPCELL_X1 PHY_EDGE_ROW_382_Right_382 ();
 TAPCELL_X1 PHY_EDGE_ROW_383_Right_383 ();
 TAPCELL_X1 PHY_EDGE_ROW_384_Right_384 ();
 TAPCELL_X1 PHY_EDGE_ROW_385_Right_385 ();
 TAPCELL_X1 PHY_EDGE_ROW_386_Right_386 ();
 TAPCELL_X1 PHY_EDGE_ROW_387_Right_387 ();
 TAPCELL_X1 PHY_EDGE_ROW_388_Right_388 ();
 TAPCELL_X1 PHY_EDGE_ROW_389_Right_389 ();
 TAPCELL_X1 PHY_EDGE_ROW_390_Right_390 ();
 TAPCELL_X1 PHY_EDGE_ROW_391_Right_391 ();
 TAPCELL_X1 PHY_EDGE_ROW_392_Right_392 ();
 TAPCELL_X1 PHY_EDGE_ROW_393_Right_393 ();
 TAPCELL_X1 PHY_EDGE_ROW_394_Right_394 ();
 TAPCELL_X1 PHY_EDGE_ROW_395_Right_395 ();
 TAPCELL_X1 PHY_EDGE_ROW_396_Right_396 ();
 TAPCELL_X1 PHY_EDGE_ROW_397_Right_397 ();
 TAPCELL_X1 PHY_EDGE_ROW_398_Right_398 ();
 TAPCELL_X1 PHY_EDGE_ROW_399_Right_399 ();
 TAPCELL_X1 PHY_EDGE_ROW_400_Right_400 ();
 TAPCELL_X1 PHY_EDGE_ROW_401_Right_401 ();
 TAPCELL_X1 PHY_EDGE_ROW_402_Right_402 ();
 TAPCELL_X1 PHY_EDGE_ROW_403_Right_403 ();
 TAPCELL_X1 PHY_EDGE_ROW_404_Right_404 ();
 TAPCELL_X1 PHY_EDGE_ROW_405_Right_405 ();
 TAPCELL_X1 PHY_EDGE_ROW_406_Right_406 ();
 TAPCELL_X1 PHY_EDGE_ROW_407_Right_407 ();
 TAPCELL_X1 PHY_EDGE_ROW_408_Right_408 ();
 TAPCELL_X1 PHY_EDGE_ROW_409_Right_409 ();
 TAPCELL_X1 PHY_EDGE_ROW_410_Right_410 ();
 TAPCELL_X1 PHY_EDGE_ROW_411_Right_411 ();
 TAPCELL_X1 PHY_EDGE_ROW_412_Right_412 ();
 TAPCELL_X1 PHY_EDGE_ROW_413_Right_413 ();
 TAPCELL_X1 PHY_EDGE_ROW_414_Right_414 ();
 TAPCELL_X1 PHY_EDGE_ROW_415_Right_415 ();
 TAPCELL_X1 PHY_EDGE_ROW_416_Right_416 ();
 TAPCELL_X1 PHY_EDGE_ROW_417_Right_417 ();
 TAPCELL_X1 PHY_EDGE_ROW_418_Right_418 ();
 TAPCELL_X1 PHY_EDGE_ROW_419_Right_419 ();
 TAPCELL_X1 PHY_EDGE_ROW_420_Right_420 ();
 TAPCELL_X1 PHY_EDGE_ROW_421_Right_421 ();
 TAPCELL_X1 PHY_EDGE_ROW_422_Right_422 ();
 TAPCELL_X1 PHY_EDGE_ROW_423_Right_423 ();
 TAPCELL_X1 PHY_EDGE_ROW_424_Right_424 ();
 TAPCELL_X1 PHY_EDGE_ROW_425_Right_425 ();
 TAPCELL_X1 PHY_EDGE_ROW_426_Right_426 ();
 TAPCELL_X1 PHY_EDGE_ROW_427_Right_427 ();
 TAPCELL_X1 PHY_EDGE_ROW_428_Right_428 ();
 TAPCELL_X1 PHY_EDGE_ROW_429_Right_429 ();
 TAPCELL_X1 PHY_EDGE_ROW_430_Right_430 ();
 TAPCELL_X1 PHY_EDGE_ROW_431_Right_431 ();
 TAPCELL_X1 PHY_EDGE_ROW_432_Right_432 ();
 TAPCELL_X1 PHY_EDGE_ROW_433_Right_433 ();
 TAPCELL_X1 PHY_EDGE_ROW_434_Right_434 ();
 TAPCELL_X1 PHY_EDGE_ROW_435_Right_435 ();
 TAPCELL_X1 PHY_EDGE_ROW_436_Right_436 ();
 TAPCELL_X1 PHY_EDGE_ROW_437_Right_437 ();
 TAPCELL_X1 PHY_EDGE_ROW_438_Right_438 ();
 TAPCELL_X1 PHY_EDGE_ROW_439_Right_439 ();
 TAPCELL_X1 PHY_EDGE_ROW_440_Right_440 ();
 TAPCELL_X1 PHY_EDGE_ROW_441_Right_441 ();
 TAPCELL_X1 PHY_EDGE_ROW_442_Right_442 ();
 TAPCELL_X1 PHY_EDGE_ROW_443_Right_443 ();
 TAPCELL_X1 PHY_EDGE_ROW_444_Right_444 ();
 TAPCELL_X1 PHY_EDGE_ROW_445_Right_445 ();
 TAPCELL_X1 PHY_EDGE_ROW_446_Right_446 ();
 TAPCELL_X1 PHY_EDGE_ROW_447_Right_447 ();
 TAPCELL_X1 PHY_EDGE_ROW_448_Right_448 ();
 TAPCELL_X1 PHY_EDGE_ROW_449_Right_449 ();
 TAPCELL_X1 PHY_EDGE_ROW_450_Right_450 ();
 TAPCELL_X1 PHY_EDGE_ROW_451_Right_451 ();
 TAPCELL_X1 PHY_EDGE_ROW_452_Right_452 ();
 TAPCELL_X1 PHY_EDGE_ROW_453_Right_453 ();
 TAPCELL_X1 PHY_EDGE_ROW_454_Right_454 ();
 TAPCELL_X1 PHY_EDGE_ROW_455_Right_455 ();
 TAPCELL_X1 PHY_EDGE_ROW_456_Right_456 ();
 TAPCELL_X1 PHY_EDGE_ROW_457_Right_457 ();
 TAPCELL_X1 PHY_EDGE_ROW_458_Right_458 ();
 TAPCELL_X1 PHY_EDGE_ROW_459_Right_459 ();
 TAPCELL_X1 PHY_EDGE_ROW_460_Right_460 ();
 TAPCELL_X1 PHY_EDGE_ROW_461_Right_461 ();
 TAPCELL_X1 PHY_EDGE_ROW_462_Right_462 ();
 TAPCELL_X1 PHY_EDGE_ROW_463_Right_463 ();
 TAPCELL_X1 PHY_EDGE_ROW_464_Right_464 ();
 TAPCELL_X1 PHY_EDGE_ROW_465_Right_465 ();
 TAPCELL_X1 PHY_EDGE_ROW_466_Right_466 ();
 TAPCELL_X1 PHY_EDGE_ROW_467_Right_467 ();
 TAPCELL_X1 PHY_EDGE_ROW_468_Right_468 ();
 TAPCELL_X1 PHY_EDGE_ROW_469_Right_469 ();
 TAPCELL_X1 PHY_EDGE_ROW_470_Right_470 ();
 TAPCELL_X1 PHY_EDGE_ROW_471_Right_471 ();
 TAPCELL_X1 PHY_EDGE_ROW_472_Right_472 ();
 TAPCELL_X1 PHY_EDGE_ROW_473_Right_473 ();
 TAPCELL_X1 PHY_EDGE_ROW_474_Right_474 ();
 TAPCELL_X1 PHY_EDGE_ROW_475_Right_475 ();
 TAPCELL_X1 PHY_EDGE_ROW_476_Right_476 ();
 TAPCELL_X1 PHY_EDGE_ROW_477_Right_477 ();
 TAPCELL_X1 PHY_EDGE_ROW_478_Right_478 ();
 TAPCELL_X1 PHY_EDGE_ROW_479_Right_479 ();
 TAPCELL_X1 PHY_EDGE_ROW_480_Right_480 ();
 TAPCELL_X1 PHY_EDGE_ROW_481_Right_481 ();
 TAPCELL_X1 PHY_EDGE_ROW_482_Right_482 ();
 TAPCELL_X1 PHY_EDGE_ROW_483_Right_483 ();
 TAPCELL_X1 PHY_EDGE_ROW_484_Right_484 ();
 TAPCELL_X1 PHY_EDGE_ROW_485_Right_485 ();
 TAPCELL_X1 PHY_EDGE_ROW_486_Right_486 ();
 TAPCELL_X1 PHY_EDGE_ROW_487_Right_487 ();
 TAPCELL_X1 PHY_EDGE_ROW_488_Right_488 ();
 TAPCELL_X1 PHY_EDGE_ROW_489_Right_489 ();
 TAPCELL_X1 PHY_EDGE_ROW_490_Right_490 ();
 TAPCELL_X1 PHY_EDGE_ROW_491_Right_491 ();
 TAPCELL_X1 PHY_EDGE_ROW_492_Right_492 ();
 TAPCELL_X1 PHY_EDGE_ROW_493_Right_493 ();
 TAPCELL_X1 PHY_EDGE_ROW_494_Right_494 ();
 TAPCELL_X1 PHY_EDGE_ROW_495_Right_495 ();
 TAPCELL_X1 PHY_EDGE_ROW_496_Right_496 ();
 TAPCELL_X1 PHY_EDGE_ROW_497_Right_497 ();
 TAPCELL_X1 PHY_EDGE_ROW_498_Right_498 ();
 TAPCELL_X1 PHY_EDGE_ROW_499_Right_499 ();
 TAPCELL_X1 PHY_EDGE_ROW_500_Right_500 ();
 TAPCELL_X1 PHY_EDGE_ROW_501_Right_501 ();
 TAPCELL_X1 PHY_EDGE_ROW_502_Right_502 ();
 TAPCELL_X1 PHY_EDGE_ROW_503_Right_503 ();
 TAPCELL_X1 PHY_EDGE_ROW_504_Right_504 ();
 TAPCELL_X1 PHY_EDGE_ROW_505_Right_505 ();
 TAPCELL_X1 PHY_EDGE_ROW_506_Right_506 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_507 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_508 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_509 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_510 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_511 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_512 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_513 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_514 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_515 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_516 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_517 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_518 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_519 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_520 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_521 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_522 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_523 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_524 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_525 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_526 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_527 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_528 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_529 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_530 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_531 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_532 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_533 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_534 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_535 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_536 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_537 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_538 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_539 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_540 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_541 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_542 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_543 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_544 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_545 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_546 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_547 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_548 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_549 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_550 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_551 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_552 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_553 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_554 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_555 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_556 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_557 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_558 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_559 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_560 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_561 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_562 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_563 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_564 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_565 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_566 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_567 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_568 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_569 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_570 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_571 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_572 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_573 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_574 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_575 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_576 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_577 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_578 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_579 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_580 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_581 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_582 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_583 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_584 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_585 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_586 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_587 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_588 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_589 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_590 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_591 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_592 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_593 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_594 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_595 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_596 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_597 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_598 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_599 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_600 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_601 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_602 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_603 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_604 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_605 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_606 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_607 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_608 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_609 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_610 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_611 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_612 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_613 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_614 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_615 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_616 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Left_617 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Left_618 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Left_619 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Left_620 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Left_621 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Left_622 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Left_623 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_624 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_625 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_626 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_627 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_628 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_629 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_630 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_631 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_632 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_633 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_634 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_635 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_636 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_637 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_638 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_639 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Left_640 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Left_641 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Left_642 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Left_643 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Left_644 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Left_645 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Left_646 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Left_647 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Left_648 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Left_649 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Left_650 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Left_651 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Left_652 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Left_653 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Left_654 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Left_655 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Left_656 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Left_657 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Left_658 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Left_659 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Left_660 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Left_661 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Left_662 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Left_663 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Left_664 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Left_665 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Left_666 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Left_667 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Left_668 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Left_669 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Left_670 ();
 TAPCELL_X1 PHY_EDGE_ROW_164_Left_671 ();
 TAPCELL_X1 PHY_EDGE_ROW_165_Left_672 ();
 TAPCELL_X1 PHY_EDGE_ROW_166_Left_673 ();
 TAPCELL_X1 PHY_EDGE_ROW_167_Left_674 ();
 TAPCELL_X1 PHY_EDGE_ROW_168_Left_675 ();
 TAPCELL_X1 PHY_EDGE_ROW_169_Left_676 ();
 TAPCELL_X1 PHY_EDGE_ROW_170_Left_677 ();
 TAPCELL_X1 PHY_EDGE_ROW_171_Left_678 ();
 TAPCELL_X1 PHY_EDGE_ROW_172_Left_679 ();
 TAPCELL_X1 PHY_EDGE_ROW_173_Left_680 ();
 TAPCELL_X1 PHY_EDGE_ROW_174_Left_681 ();
 TAPCELL_X1 PHY_EDGE_ROW_175_Left_682 ();
 TAPCELL_X1 PHY_EDGE_ROW_176_Left_683 ();
 TAPCELL_X1 PHY_EDGE_ROW_177_Left_684 ();
 TAPCELL_X1 PHY_EDGE_ROW_178_Left_685 ();
 TAPCELL_X1 PHY_EDGE_ROW_179_Left_686 ();
 TAPCELL_X1 PHY_EDGE_ROW_180_Left_687 ();
 TAPCELL_X1 PHY_EDGE_ROW_181_Left_688 ();
 TAPCELL_X1 PHY_EDGE_ROW_182_Left_689 ();
 TAPCELL_X1 PHY_EDGE_ROW_183_Left_690 ();
 TAPCELL_X1 PHY_EDGE_ROW_184_Left_691 ();
 TAPCELL_X1 PHY_EDGE_ROW_185_Left_692 ();
 TAPCELL_X1 PHY_EDGE_ROW_186_Left_693 ();
 TAPCELL_X1 PHY_EDGE_ROW_187_Left_694 ();
 TAPCELL_X1 PHY_EDGE_ROW_188_Left_695 ();
 TAPCELL_X1 PHY_EDGE_ROW_189_Left_696 ();
 TAPCELL_X1 PHY_EDGE_ROW_190_Left_697 ();
 TAPCELL_X1 PHY_EDGE_ROW_191_Left_698 ();
 TAPCELL_X1 PHY_EDGE_ROW_192_Left_699 ();
 TAPCELL_X1 PHY_EDGE_ROW_193_Left_700 ();
 TAPCELL_X1 PHY_EDGE_ROW_194_Left_701 ();
 TAPCELL_X1 PHY_EDGE_ROW_195_Left_702 ();
 TAPCELL_X1 PHY_EDGE_ROW_196_Left_703 ();
 TAPCELL_X1 PHY_EDGE_ROW_197_Left_704 ();
 TAPCELL_X1 PHY_EDGE_ROW_198_Left_705 ();
 TAPCELL_X1 PHY_EDGE_ROW_199_Left_706 ();
 TAPCELL_X1 PHY_EDGE_ROW_200_Left_707 ();
 TAPCELL_X1 PHY_EDGE_ROW_201_Left_708 ();
 TAPCELL_X1 PHY_EDGE_ROW_202_Left_709 ();
 TAPCELL_X1 PHY_EDGE_ROW_203_Left_710 ();
 TAPCELL_X1 PHY_EDGE_ROW_204_Left_711 ();
 TAPCELL_X1 PHY_EDGE_ROW_205_Left_712 ();
 TAPCELL_X1 PHY_EDGE_ROW_206_Left_713 ();
 TAPCELL_X1 PHY_EDGE_ROW_207_Left_714 ();
 TAPCELL_X1 PHY_EDGE_ROW_208_Left_715 ();
 TAPCELL_X1 PHY_EDGE_ROW_209_Left_716 ();
 TAPCELL_X1 PHY_EDGE_ROW_210_Left_717 ();
 TAPCELL_X1 PHY_EDGE_ROW_211_Left_718 ();
 TAPCELL_X1 PHY_EDGE_ROW_212_Left_719 ();
 TAPCELL_X1 PHY_EDGE_ROW_213_Left_720 ();
 TAPCELL_X1 PHY_EDGE_ROW_214_Left_721 ();
 TAPCELL_X1 PHY_EDGE_ROW_215_Left_722 ();
 TAPCELL_X1 PHY_EDGE_ROW_216_Left_723 ();
 TAPCELL_X1 PHY_EDGE_ROW_217_Left_724 ();
 TAPCELL_X1 PHY_EDGE_ROW_218_Left_725 ();
 TAPCELL_X1 PHY_EDGE_ROW_219_Left_726 ();
 TAPCELL_X1 PHY_EDGE_ROW_220_Left_727 ();
 TAPCELL_X1 PHY_EDGE_ROW_221_Left_728 ();
 TAPCELL_X1 PHY_EDGE_ROW_222_Left_729 ();
 TAPCELL_X1 PHY_EDGE_ROW_223_Left_730 ();
 TAPCELL_X1 PHY_EDGE_ROW_224_Left_731 ();
 TAPCELL_X1 PHY_EDGE_ROW_225_Left_732 ();
 TAPCELL_X1 PHY_EDGE_ROW_226_Left_733 ();
 TAPCELL_X1 PHY_EDGE_ROW_227_Left_734 ();
 TAPCELL_X1 PHY_EDGE_ROW_228_Left_735 ();
 TAPCELL_X1 PHY_EDGE_ROW_229_Left_736 ();
 TAPCELL_X1 PHY_EDGE_ROW_230_Left_737 ();
 TAPCELL_X1 PHY_EDGE_ROW_231_Left_738 ();
 TAPCELL_X1 PHY_EDGE_ROW_232_Left_739 ();
 TAPCELL_X1 PHY_EDGE_ROW_233_Left_740 ();
 TAPCELL_X1 PHY_EDGE_ROW_234_Left_741 ();
 TAPCELL_X1 PHY_EDGE_ROW_235_Left_742 ();
 TAPCELL_X1 PHY_EDGE_ROW_236_Left_743 ();
 TAPCELL_X1 PHY_EDGE_ROW_237_Left_744 ();
 TAPCELL_X1 PHY_EDGE_ROW_238_Left_745 ();
 TAPCELL_X1 PHY_EDGE_ROW_239_Left_746 ();
 TAPCELL_X1 PHY_EDGE_ROW_240_Left_747 ();
 TAPCELL_X1 PHY_EDGE_ROW_241_Left_748 ();
 TAPCELL_X1 PHY_EDGE_ROW_242_Left_749 ();
 TAPCELL_X1 PHY_EDGE_ROW_243_Left_750 ();
 TAPCELL_X1 PHY_EDGE_ROW_244_Left_751 ();
 TAPCELL_X1 PHY_EDGE_ROW_245_Left_752 ();
 TAPCELL_X1 PHY_EDGE_ROW_246_Left_753 ();
 TAPCELL_X1 PHY_EDGE_ROW_247_Left_754 ();
 TAPCELL_X1 PHY_EDGE_ROW_248_Left_755 ();
 TAPCELL_X1 PHY_EDGE_ROW_249_Left_756 ();
 TAPCELL_X1 PHY_EDGE_ROW_250_Left_757 ();
 TAPCELL_X1 PHY_EDGE_ROW_251_Left_758 ();
 TAPCELL_X1 PHY_EDGE_ROW_252_Left_759 ();
 TAPCELL_X1 PHY_EDGE_ROW_253_Left_760 ();
 TAPCELL_X1 PHY_EDGE_ROW_254_Left_761 ();
 TAPCELL_X1 PHY_EDGE_ROW_255_Left_762 ();
 TAPCELL_X1 PHY_EDGE_ROW_256_Left_763 ();
 TAPCELL_X1 PHY_EDGE_ROW_257_Left_764 ();
 TAPCELL_X1 PHY_EDGE_ROW_258_Left_765 ();
 TAPCELL_X1 PHY_EDGE_ROW_259_Left_766 ();
 TAPCELL_X1 PHY_EDGE_ROW_260_Left_767 ();
 TAPCELL_X1 PHY_EDGE_ROW_261_Left_768 ();
 TAPCELL_X1 PHY_EDGE_ROW_262_Left_769 ();
 TAPCELL_X1 PHY_EDGE_ROW_263_Left_770 ();
 TAPCELL_X1 PHY_EDGE_ROW_264_Left_771 ();
 TAPCELL_X1 PHY_EDGE_ROW_265_Left_772 ();
 TAPCELL_X1 PHY_EDGE_ROW_266_Left_773 ();
 TAPCELL_X1 PHY_EDGE_ROW_267_Left_774 ();
 TAPCELL_X1 PHY_EDGE_ROW_268_Left_775 ();
 TAPCELL_X1 PHY_EDGE_ROW_269_Left_776 ();
 TAPCELL_X1 PHY_EDGE_ROW_270_Left_777 ();
 TAPCELL_X1 PHY_EDGE_ROW_271_Left_778 ();
 TAPCELL_X1 PHY_EDGE_ROW_272_Left_779 ();
 TAPCELL_X1 PHY_EDGE_ROW_273_Left_780 ();
 TAPCELL_X1 PHY_EDGE_ROW_274_Left_781 ();
 TAPCELL_X1 PHY_EDGE_ROW_275_Left_782 ();
 TAPCELL_X1 PHY_EDGE_ROW_276_Left_783 ();
 TAPCELL_X1 PHY_EDGE_ROW_277_Left_784 ();
 TAPCELL_X1 PHY_EDGE_ROW_278_Left_785 ();
 TAPCELL_X1 PHY_EDGE_ROW_279_Left_786 ();
 TAPCELL_X1 PHY_EDGE_ROW_280_Left_787 ();
 TAPCELL_X1 PHY_EDGE_ROW_281_Left_788 ();
 TAPCELL_X1 PHY_EDGE_ROW_282_Left_789 ();
 TAPCELL_X1 PHY_EDGE_ROW_283_Left_790 ();
 TAPCELL_X1 PHY_EDGE_ROW_284_Left_791 ();
 TAPCELL_X1 PHY_EDGE_ROW_285_Left_792 ();
 TAPCELL_X1 PHY_EDGE_ROW_286_Left_793 ();
 TAPCELL_X1 PHY_EDGE_ROW_287_Left_794 ();
 TAPCELL_X1 PHY_EDGE_ROW_288_Left_795 ();
 TAPCELL_X1 PHY_EDGE_ROW_289_Left_796 ();
 TAPCELL_X1 PHY_EDGE_ROW_290_Left_797 ();
 TAPCELL_X1 PHY_EDGE_ROW_291_Left_798 ();
 TAPCELL_X1 PHY_EDGE_ROW_292_Left_799 ();
 TAPCELL_X1 PHY_EDGE_ROW_293_Left_800 ();
 TAPCELL_X1 PHY_EDGE_ROW_294_Left_801 ();
 TAPCELL_X1 PHY_EDGE_ROW_295_Left_802 ();
 TAPCELL_X1 PHY_EDGE_ROW_296_Left_803 ();
 TAPCELL_X1 PHY_EDGE_ROW_297_Left_804 ();
 TAPCELL_X1 PHY_EDGE_ROW_298_Left_805 ();
 TAPCELL_X1 PHY_EDGE_ROW_299_Left_806 ();
 TAPCELL_X1 PHY_EDGE_ROW_300_Left_807 ();
 TAPCELL_X1 PHY_EDGE_ROW_301_Left_808 ();
 TAPCELL_X1 PHY_EDGE_ROW_302_Left_809 ();
 TAPCELL_X1 PHY_EDGE_ROW_303_Left_810 ();
 TAPCELL_X1 PHY_EDGE_ROW_304_Left_811 ();
 TAPCELL_X1 PHY_EDGE_ROW_305_Left_812 ();
 TAPCELL_X1 PHY_EDGE_ROW_306_Left_813 ();
 TAPCELL_X1 PHY_EDGE_ROW_307_Left_814 ();
 TAPCELL_X1 PHY_EDGE_ROW_308_Left_815 ();
 TAPCELL_X1 PHY_EDGE_ROW_309_Left_816 ();
 TAPCELL_X1 PHY_EDGE_ROW_310_Left_817 ();
 TAPCELL_X1 PHY_EDGE_ROW_311_Left_818 ();
 TAPCELL_X1 PHY_EDGE_ROW_312_Left_819 ();
 TAPCELL_X1 PHY_EDGE_ROW_313_Left_820 ();
 TAPCELL_X1 PHY_EDGE_ROW_314_Left_821 ();
 TAPCELL_X1 PHY_EDGE_ROW_315_Left_822 ();
 TAPCELL_X1 PHY_EDGE_ROW_316_Left_823 ();
 TAPCELL_X1 PHY_EDGE_ROW_317_Left_824 ();
 TAPCELL_X1 PHY_EDGE_ROW_318_Left_825 ();
 TAPCELL_X1 PHY_EDGE_ROW_319_Left_826 ();
 TAPCELL_X1 PHY_EDGE_ROW_320_Left_827 ();
 TAPCELL_X1 PHY_EDGE_ROW_321_Left_828 ();
 TAPCELL_X1 PHY_EDGE_ROW_322_Left_829 ();
 TAPCELL_X1 PHY_EDGE_ROW_323_Left_830 ();
 TAPCELL_X1 PHY_EDGE_ROW_324_Left_831 ();
 TAPCELL_X1 PHY_EDGE_ROW_325_Left_832 ();
 TAPCELL_X1 PHY_EDGE_ROW_326_Left_833 ();
 TAPCELL_X1 PHY_EDGE_ROW_327_Left_834 ();
 TAPCELL_X1 PHY_EDGE_ROW_328_Left_835 ();
 TAPCELL_X1 PHY_EDGE_ROW_329_Left_836 ();
 TAPCELL_X1 PHY_EDGE_ROW_330_Left_837 ();
 TAPCELL_X1 PHY_EDGE_ROW_331_Left_838 ();
 TAPCELL_X1 PHY_EDGE_ROW_332_Left_839 ();
 TAPCELL_X1 PHY_EDGE_ROW_333_Left_840 ();
 TAPCELL_X1 PHY_EDGE_ROW_334_Left_841 ();
 TAPCELL_X1 PHY_EDGE_ROW_335_Left_842 ();
 TAPCELL_X1 PHY_EDGE_ROW_336_Left_843 ();
 TAPCELL_X1 PHY_EDGE_ROW_337_Left_844 ();
 TAPCELL_X1 PHY_EDGE_ROW_338_Left_845 ();
 TAPCELL_X1 PHY_EDGE_ROW_339_Left_846 ();
 TAPCELL_X1 PHY_EDGE_ROW_340_Left_847 ();
 TAPCELL_X1 PHY_EDGE_ROW_341_Left_848 ();
 TAPCELL_X1 PHY_EDGE_ROW_342_Left_849 ();
 TAPCELL_X1 PHY_EDGE_ROW_343_Left_850 ();
 TAPCELL_X1 PHY_EDGE_ROW_344_Left_851 ();
 TAPCELL_X1 PHY_EDGE_ROW_345_Left_852 ();
 TAPCELL_X1 PHY_EDGE_ROW_346_Left_853 ();
 TAPCELL_X1 PHY_EDGE_ROW_347_Left_854 ();
 TAPCELL_X1 PHY_EDGE_ROW_348_Left_855 ();
 TAPCELL_X1 PHY_EDGE_ROW_349_Left_856 ();
 TAPCELL_X1 PHY_EDGE_ROW_350_Left_857 ();
 TAPCELL_X1 PHY_EDGE_ROW_351_Left_858 ();
 TAPCELL_X1 PHY_EDGE_ROW_352_Left_859 ();
 TAPCELL_X1 PHY_EDGE_ROW_353_Left_860 ();
 TAPCELL_X1 PHY_EDGE_ROW_354_Left_861 ();
 TAPCELL_X1 PHY_EDGE_ROW_355_Left_862 ();
 TAPCELL_X1 PHY_EDGE_ROW_356_Left_863 ();
 TAPCELL_X1 PHY_EDGE_ROW_357_Left_864 ();
 TAPCELL_X1 PHY_EDGE_ROW_358_Left_865 ();
 TAPCELL_X1 PHY_EDGE_ROW_359_Left_866 ();
 TAPCELL_X1 PHY_EDGE_ROW_360_Left_867 ();
 TAPCELL_X1 PHY_EDGE_ROW_361_Left_868 ();
 TAPCELL_X1 PHY_EDGE_ROW_362_Left_869 ();
 TAPCELL_X1 PHY_EDGE_ROW_363_Left_870 ();
 TAPCELL_X1 PHY_EDGE_ROW_364_Left_871 ();
 TAPCELL_X1 PHY_EDGE_ROW_365_Left_872 ();
 TAPCELL_X1 PHY_EDGE_ROW_366_Left_873 ();
 TAPCELL_X1 PHY_EDGE_ROW_367_Left_874 ();
 TAPCELL_X1 PHY_EDGE_ROW_368_Left_875 ();
 TAPCELL_X1 PHY_EDGE_ROW_369_Left_876 ();
 TAPCELL_X1 PHY_EDGE_ROW_370_Left_877 ();
 TAPCELL_X1 PHY_EDGE_ROW_371_Left_878 ();
 TAPCELL_X1 PHY_EDGE_ROW_372_Left_879 ();
 TAPCELL_X1 PHY_EDGE_ROW_373_Left_880 ();
 TAPCELL_X1 PHY_EDGE_ROW_374_Left_881 ();
 TAPCELL_X1 PHY_EDGE_ROW_375_Left_882 ();
 TAPCELL_X1 PHY_EDGE_ROW_376_Left_883 ();
 TAPCELL_X1 PHY_EDGE_ROW_377_Left_884 ();
 TAPCELL_X1 PHY_EDGE_ROW_378_Left_885 ();
 TAPCELL_X1 PHY_EDGE_ROW_379_Left_886 ();
 TAPCELL_X1 PHY_EDGE_ROW_380_Left_887 ();
 TAPCELL_X1 PHY_EDGE_ROW_381_Left_888 ();
 TAPCELL_X1 PHY_EDGE_ROW_382_Left_889 ();
 TAPCELL_X1 PHY_EDGE_ROW_383_Left_890 ();
 TAPCELL_X1 PHY_EDGE_ROW_384_Left_891 ();
 TAPCELL_X1 PHY_EDGE_ROW_385_Left_892 ();
 TAPCELL_X1 PHY_EDGE_ROW_386_Left_893 ();
 TAPCELL_X1 PHY_EDGE_ROW_387_Left_894 ();
 TAPCELL_X1 PHY_EDGE_ROW_388_Left_895 ();
 TAPCELL_X1 PHY_EDGE_ROW_389_Left_896 ();
 TAPCELL_X1 PHY_EDGE_ROW_390_Left_897 ();
 TAPCELL_X1 PHY_EDGE_ROW_391_Left_898 ();
 TAPCELL_X1 PHY_EDGE_ROW_392_Left_899 ();
 TAPCELL_X1 PHY_EDGE_ROW_393_Left_900 ();
 TAPCELL_X1 PHY_EDGE_ROW_394_Left_901 ();
 TAPCELL_X1 PHY_EDGE_ROW_395_Left_902 ();
 TAPCELL_X1 PHY_EDGE_ROW_396_Left_903 ();
 TAPCELL_X1 PHY_EDGE_ROW_397_Left_904 ();
 TAPCELL_X1 PHY_EDGE_ROW_398_Left_905 ();
 TAPCELL_X1 PHY_EDGE_ROW_399_Left_906 ();
 TAPCELL_X1 PHY_EDGE_ROW_400_Left_907 ();
 TAPCELL_X1 PHY_EDGE_ROW_401_Left_908 ();
 TAPCELL_X1 PHY_EDGE_ROW_402_Left_909 ();
 TAPCELL_X1 PHY_EDGE_ROW_403_Left_910 ();
 TAPCELL_X1 PHY_EDGE_ROW_404_Left_911 ();
 TAPCELL_X1 PHY_EDGE_ROW_405_Left_912 ();
 TAPCELL_X1 PHY_EDGE_ROW_406_Left_913 ();
 TAPCELL_X1 PHY_EDGE_ROW_407_Left_914 ();
 TAPCELL_X1 PHY_EDGE_ROW_408_Left_915 ();
 TAPCELL_X1 PHY_EDGE_ROW_409_Left_916 ();
 TAPCELL_X1 PHY_EDGE_ROW_410_Left_917 ();
 TAPCELL_X1 PHY_EDGE_ROW_411_Left_918 ();
 TAPCELL_X1 PHY_EDGE_ROW_412_Left_919 ();
 TAPCELL_X1 PHY_EDGE_ROW_413_Left_920 ();
 TAPCELL_X1 PHY_EDGE_ROW_414_Left_921 ();
 TAPCELL_X1 PHY_EDGE_ROW_415_Left_922 ();
 TAPCELL_X1 PHY_EDGE_ROW_416_Left_923 ();
 TAPCELL_X1 PHY_EDGE_ROW_417_Left_924 ();
 TAPCELL_X1 PHY_EDGE_ROW_418_Left_925 ();
 TAPCELL_X1 PHY_EDGE_ROW_419_Left_926 ();
 TAPCELL_X1 PHY_EDGE_ROW_420_Left_927 ();
 TAPCELL_X1 PHY_EDGE_ROW_421_Left_928 ();
 TAPCELL_X1 PHY_EDGE_ROW_422_Left_929 ();
 TAPCELL_X1 PHY_EDGE_ROW_423_Left_930 ();
 TAPCELL_X1 PHY_EDGE_ROW_424_Left_931 ();
 TAPCELL_X1 PHY_EDGE_ROW_425_Left_932 ();
 TAPCELL_X1 PHY_EDGE_ROW_426_Left_933 ();
 TAPCELL_X1 PHY_EDGE_ROW_427_Left_934 ();
 TAPCELL_X1 PHY_EDGE_ROW_428_Left_935 ();
 TAPCELL_X1 PHY_EDGE_ROW_429_Left_936 ();
 TAPCELL_X1 PHY_EDGE_ROW_430_Left_937 ();
 TAPCELL_X1 PHY_EDGE_ROW_431_Left_938 ();
 TAPCELL_X1 PHY_EDGE_ROW_432_Left_939 ();
 TAPCELL_X1 PHY_EDGE_ROW_433_Left_940 ();
 TAPCELL_X1 PHY_EDGE_ROW_434_Left_941 ();
 TAPCELL_X1 PHY_EDGE_ROW_435_Left_942 ();
 TAPCELL_X1 PHY_EDGE_ROW_436_Left_943 ();
 TAPCELL_X1 PHY_EDGE_ROW_437_Left_944 ();
 TAPCELL_X1 PHY_EDGE_ROW_438_Left_945 ();
 TAPCELL_X1 PHY_EDGE_ROW_439_Left_946 ();
 TAPCELL_X1 PHY_EDGE_ROW_440_Left_947 ();
 TAPCELL_X1 PHY_EDGE_ROW_441_Left_948 ();
 TAPCELL_X1 PHY_EDGE_ROW_442_Left_949 ();
 TAPCELL_X1 PHY_EDGE_ROW_443_Left_950 ();
 TAPCELL_X1 PHY_EDGE_ROW_444_Left_951 ();
 TAPCELL_X1 PHY_EDGE_ROW_445_Left_952 ();
 TAPCELL_X1 PHY_EDGE_ROW_446_Left_953 ();
 TAPCELL_X1 PHY_EDGE_ROW_447_Left_954 ();
 TAPCELL_X1 PHY_EDGE_ROW_448_Left_955 ();
 TAPCELL_X1 PHY_EDGE_ROW_449_Left_956 ();
 TAPCELL_X1 PHY_EDGE_ROW_450_Left_957 ();
 TAPCELL_X1 PHY_EDGE_ROW_451_Left_958 ();
 TAPCELL_X1 PHY_EDGE_ROW_452_Left_959 ();
 TAPCELL_X1 PHY_EDGE_ROW_453_Left_960 ();
 TAPCELL_X1 PHY_EDGE_ROW_454_Left_961 ();
 TAPCELL_X1 PHY_EDGE_ROW_455_Left_962 ();
 TAPCELL_X1 PHY_EDGE_ROW_456_Left_963 ();
 TAPCELL_X1 PHY_EDGE_ROW_457_Left_964 ();
 TAPCELL_X1 PHY_EDGE_ROW_458_Left_965 ();
 TAPCELL_X1 PHY_EDGE_ROW_459_Left_966 ();
 TAPCELL_X1 PHY_EDGE_ROW_460_Left_967 ();
 TAPCELL_X1 PHY_EDGE_ROW_461_Left_968 ();
 TAPCELL_X1 PHY_EDGE_ROW_462_Left_969 ();
 TAPCELL_X1 PHY_EDGE_ROW_463_Left_970 ();
 TAPCELL_X1 PHY_EDGE_ROW_464_Left_971 ();
 TAPCELL_X1 PHY_EDGE_ROW_465_Left_972 ();
 TAPCELL_X1 PHY_EDGE_ROW_466_Left_973 ();
 TAPCELL_X1 PHY_EDGE_ROW_467_Left_974 ();
 TAPCELL_X1 PHY_EDGE_ROW_468_Left_975 ();
 TAPCELL_X1 PHY_EDGE_ROW_469_Left_976 ();
 TAPCELL_X1 PHY_EDGE_ROW_470_Left_977 ();
 TAPCELL_X1 PHY_EDGE_ROW_471_Left_978 ();
 TAPCELL_X1 PHY_EDGE_ROW_472_Left_979 ();
 TAPCELL_X1 PHY_EDGE_ROW_473_Left_980 ();
 TAPCELL_X1 PHY_EDGE_ROW_474_Left_981 ();
 TAPCELL_X1 PHY_EDGE_ROW_475_Left_982 ();
 TAPCELL_X1 PHY_EDGE_ROW_476_Left_983 ();
 TAPCELL_X1 PHY_EDGE_ROW_477_Left_984 ();
 TAPCELL_X1 PHY_EDGE_ROW_478_Left_985 ();
 TAPCELL_X1 PHY_EDGE_ROW_479_Left_986 ();
 TAPCELL_X1 PHY_EDGE_ROW_480_Left_987 ();
 TAPCELL_X1 PHY_EDGE_ROW_481_Left_988 ();
 TAPCELL_X1 PHY_EDGE_ROW_482_Left_989 ();
 TAPCELL_X1 PHY_EDGE_ROW_483_Left_990 ();
 TAPCELL_X1 PHY_EDGE_ROW_484_Left_991 ();
 TAPCELL_X1 PHY_EDGE_ROW_485_Left_992 ();
 TAPCELL_X1 PHY_EDGE_ROW_486_Left_993 ();
 TAPCELL_X1 PHY_EDGE_ROW_487_Left_994 ();
 TAPCELL_X1 PHY_EDGE_ROW_488_Left_995 ();
 TAPCELL_X1 PHY_EDGE_ROW_489_Left_996 ();
 TAPCELL_X1 PHY_EDGE_ROW_490_Left_997 ();
 TAPCELL_X1 PHY_EDGE_ROW_491_Left_998 ();
 TAPCELL_X1 PHY_EDGE_ROW_492_Left_999 ();
 TAPCELL_X1 PHY_EDGE_ROW_493_Left_1000 ();
 TAPCELL_X1 PHY_EDGE_ROW_494_Left_1001 ();
 TAPCELL_X1 PHY_EDGE_ROW_495_Left_1002 ();
 TAPCELL_X1 PHY_EDGE_ROW_496_Left_1003 ();
 TAPCELL_X1 PHY_EDGE_ROW_497_Left_1004 ();
 TAPCELL_X1 PHY_EDGE_ROW_498_Left_1005 ();
 TAPCELL_X1 PHY_EDGE_ROW_499_Left_1006 ();
 TAPCELL_X1 PHY_EDGE_ROW_500_Left_1007 ();
 TAPCELL_X1 PHY_EDGE_ROW_501_Left_1008 ();
 TAPCELL_X1 PHY_EDGE_ROW_502_Left_1009 ();
 TAPCELL_X1 PHY_EDGE_ROW_503_Left_1010 ();
 TAPCELL_X1 PHY_EDGE_ROW_504_Left_1011 ();
 TAPCELL_X1 PHY_EDGE_ROW_505_Left_1012 ();
 TAPCELL_X1 PHY_EDGE_ROW_506_Left_1013 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_1014 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_1015 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_1016 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_1017 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_1018 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_1019 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_1_1020 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_1021 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_1022 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_1023 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_1024 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_3_1025 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_1026 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_1027 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_1028 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_1029 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_5_1030 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_1031 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_1032 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_1033 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_1034 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_7_1035 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_1036 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_1037 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_1038 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_1039 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_9_1040 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_1041 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_1042 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_1043 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_1044 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_11_1045 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_1046 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_1047 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_1048 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_1049 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_13_1050 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_1051 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_1052 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_1053 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_1054 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_15_1055 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_1056 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_1057 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_1058 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_1059 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_17_1060 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_1061 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_1062 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_1063 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_1064 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_19_1065 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_1066 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_1067 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_1068 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_1069 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_21_1070 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_1071 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_1072 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_1073 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_1074 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_23_1075 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_1076 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_1077 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_1078 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_1079 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_25_1080 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_1081 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_1082 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_1083 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_1084 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_27_1085 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_1086 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_1087 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_1088 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_1089 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_29_1090 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_1091 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_1092 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_1093 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_1094 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_31_1095 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_1096 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_1097 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_1098 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_1099 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_33_1100 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_1101 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_1102 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_1103 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_1104 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_35_1105 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_1106 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_1107 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_1108 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_1109 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_37_1110 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_1111 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_1112 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_1113 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_1114 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_39_1115 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_1116 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_1117 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_1118 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_1119 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_41_1120 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_1121 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_1122 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_1123 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_1124 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_43_1125 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_1126 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_1127 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_1128 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_1129 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_45_1130 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_1131 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_1132 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_1133 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_1134 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_47_1135 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_1136 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_1137 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_1138 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_1139 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_49_1140 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_1141 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_1142 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_1143 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_1144 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_51_1145 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_1146 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_1147 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_1148 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_1149 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_53_1150 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_1151 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_1152 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_1153 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_1154 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_55_1155 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_1156 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_1157 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_1158 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_57_1159 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_57_1160 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_1161 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_1162 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_1163 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_59_1164 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_59_1165 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_1166 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_1167 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_1168 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_61_1169 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_61_1170 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_1171 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_1172 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_1173 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_63_1174 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_63_1175 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_1176 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_1177 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_1178 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_1179 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_65_1180 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_1181 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_1182 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_1183 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_67_1184 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_67_1185 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_1186 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_1187 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_1188 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_1189 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_69_1190 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_1191 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_1192 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_1193 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_1194 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_71_1195 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_1196 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_1197 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_1198 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_73_1199 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_73_1200 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_1201 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_1202 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_1203 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_75_1204 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_75_1205 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_1206 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_1207 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_1208 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_77_1209 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_77_1210 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_1211 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_1212 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_1213 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_79_1214 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_79_1215 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_1216 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_1217 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_1218 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_81_1219 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_81_1220 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_1221 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_1222 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_1223 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_83_1224 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_83_1225 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_1226 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_1227 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_1228 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_85_1229 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_85_1230 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_1231 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_1232 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_1233 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_87_1234 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_87_1235 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_1236 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_1237 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_1238 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_89_1239 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_89_1240 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_1241 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_1242 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_1243 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_91_1244 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_91_1245 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_1246 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_1247 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_1248 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_93_1249 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_93_1250 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_1251 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_1252 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_1253 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_95_1254 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_95_1255 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_1256 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_1257 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_1258 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_97_1259 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_97_1260 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_1261 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_1262 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_1263 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_99_1264 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_99_1265 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_1266 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_1267 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_1268 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_101_1269 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_101_1270 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_1271 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_1272 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_1273 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_103_1274 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_103_1275 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_1276 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_1277 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_1278 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_105_1279 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_105_1280 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_1281 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_1282 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_1283 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_107_1284 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_107_1285 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_1286 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_1287 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_1288 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_109_1289 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_109_1290 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_1291 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_1292 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_1293 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_111_1294 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_111_1295 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_1296 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_1297 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_1298 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_113_1299 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_113_1300 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_1301 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_1302 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_1303 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_115_1304 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_115_1305 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_1306 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_1307 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_1308 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_117_1309 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_117_1310 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_1311 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_1312 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_1313 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_119_1314 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_119_1315 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_1316 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_1317 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_1318 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_121_1319 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_121_1320 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_1321 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_1322 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_1323 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_123_1324 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_123_1325 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_1326 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_1327 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_1328 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_125_1329 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_125_1330 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_1331 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_1332 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_1333 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_127_1334 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_127_1335 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_1336 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_1337 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_1338 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_129_1339 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_129_1340 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_1341 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_1342 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_1343 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_131_1344 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_131_1345 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_1346 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_1347 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_1348 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_133_1349 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_133_1350 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_1351 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_1352 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_1353 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_135_1354 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_135_1355 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_1356 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_1357 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_1358 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_137_1359 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_137_1360 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_1361 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_1362 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_1363 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_139_1364 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_139_1365 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_1366 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_1367 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_1368 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_141_1369 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_141_1370 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_1371 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_1372 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_1373 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_143_1374 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_143_1375 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_1376 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_1377 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_1378 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_145_1379 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_145_1380 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_1381 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_1382 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_1383 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_147_1384 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_147_1385 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_1386 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_1387 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_1388 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_149_1389 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_149_1390 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_1391 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_1392 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_1393 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_151_1394 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_151_1395 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_1396 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_1397 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_1398 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_153_1399 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_153_1400 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_1401 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_1402 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_1403 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_155_1404 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_155_1405 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_1406 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_1407 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_1408 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_157_1409 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_157_1410 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_1411 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_1412 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_1413 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_159_1414 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_159_1415 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_1416 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_1417 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_1418 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_161_1419 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_161_1420 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_1421 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_1422 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_1423 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_163_1424 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_163_1425 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_1426 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_1427 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_164_1428 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_165_1429 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_165_1430 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_1431 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_1432 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_166_1433 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_167_1434 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_167_1435 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_1436 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_1437 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_168_1438 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_169_1439 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_169_1440 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_1441 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_1442 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_170_1443 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_171_1444 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_171_1445 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_1446 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_1447 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_172_1448 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_173_1449 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_173_1450 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_1451 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_1452 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_174_1453 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_175_1454 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_175_1455 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_1456 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_1457 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_176_1458 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_177_1459 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_177_1460 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_1461 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_1462 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_178_1463 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_179_1464 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_179_1465 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_180_1466 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_180_1467 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_180_1468 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_181_1469 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_181_1470 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_182_1471 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_182_1472 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_182_1473 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_183_1474 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_183_1475 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_184_1476 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_184_1477 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_184_1478 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_185_1479 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_185_1480 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_186_1481 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_186_1482 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_186_1483 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_187_1484 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_187_1485 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_188_1486 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_188_1487 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_188_1488 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_189_1489 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_189_1490 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_190_1491 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_190_1492 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_190_1493 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_191_1494 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_191_1495 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_192_1496 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_192_1497 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_192_1498 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_193_1499 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_193_1500 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_194_1501 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_194_1502 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_194_1503 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_195_1504 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_195_1505 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_196_1506 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_196_1507 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_196_1508 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_197_1509 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_197_1510 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_198_1511 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_198_1512 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_198_1513 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_199_1514 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_199_1515 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_200_1516 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_200_1517 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_200_1518 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_201_1519 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_201_1520 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_202_1521 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_202_1522 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_202_1523 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_203_1524 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_203_1525 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_204_1526 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_204_1527 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_204_1528 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_205_1529 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_205_1530 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_206_1531 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_206_1532 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_206_1533 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_207_1534 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_207_1535 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_1536 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_1537 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_208_1538 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_209_1539 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_209_1540 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_1541 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_1542 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_210_1543 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_211_1544 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_211_1545 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_1546 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_1547 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_212_1548 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_213_1549 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_213_1550 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_1551 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_1552 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_214_1553 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_215_1554 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_215_1555 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_1556 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_1557 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_216_1558 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_217_1559 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_217_1560 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_1561 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_1562 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_218_1563 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_219_1564 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_219_1565 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_1566 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_1567 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_220_1568 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_221_1569 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_221_1570 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_1571 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_1572 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_222_1573 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_223_1574 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_223_1575 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_1576 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_1577 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_224_1578 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_225_1579 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_225_1580 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_1581 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_1582 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_226_1583 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_227_1584 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_227_1585 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_1586 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_1587 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_228_1588 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_229_1589 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_229_1590 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_230_1591 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_230_1592 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_230_1593 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_231_1594 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_231_1595 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_232_1596 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_232_1597 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_232_1598 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_233_1599 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_233_1600 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_234_1601 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_234_1602 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_234_1603 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_235_1604 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_235_1605 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_236_1606 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_236_1607 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_236_1608 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_237_1609 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_237_1610 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_238_1611 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_238_1612 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_238_1613 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_239_1614 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_239_1615 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_240_1616 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_240_1617 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_240_1618 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_241_1619 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_241_1620 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_242_1621 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_242_1622 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_242_1623 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_243_1624 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_243_1625 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_244_1626 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_244_1627 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_244_1628 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_245_1629 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_245_1630 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_246_1631 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_246_1632 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_246_1633 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_247_1634 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_247_1635 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_248_1636 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_248_1637 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_248_1638 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_249_1639 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_249_1640 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_250_1641 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_250_1642 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_250_1643 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_251_1644 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_251_1645 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_252_1646 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_252_1647 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_252_1648 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_253_1649 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_253_1650 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_254_1651 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_254_1652 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_254_1653 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_255_1654 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_255_1655 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_256_1656 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_256_1657 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_256_1658 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_257_1659 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_257_1660 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_258_1661 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_258_1662 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_258_1663 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_259_1664 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_259_1665 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_260_1666 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_260_1667 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_260_1668 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_261_1669 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_261_1670 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_262_1671 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_262_1672 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_262_1673 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_263_1674 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_263_1675 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_264_1676 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_264_1677 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_264_1678 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_265_1679 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_265_1680 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_266_1681 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_266_1682 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_266_1683 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_267_1684 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_267_1685 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_268_1686 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_268_1687 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_268_1688 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_269_1689 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_269_1690 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_270_1691 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_270_1692 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_270_1693 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_271_1694 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_271_1695 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_272_1696 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_272_1697 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_272_1698 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_273_1699 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_273_1700 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_274_1701 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_274_1702 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_274_1703 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_275_1704 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_275_1705 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_276_1706 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_276_1707 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_276_1708 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_277_1709 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_277_1710 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_278_1711 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_278_1712 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_278_1713 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_279_1714 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_279_1715 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_280_1716 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_280_1717 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_280_1718 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_281_1719 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_281_1720 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_282_1721 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_282_1722 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_282_1723 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_283_1724 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_283_1725 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_284_1726 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_284_1727 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_284_1728 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_285_1729 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_285_1730 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_286_1731 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_286_1732 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_286_1733 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_287_1734 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_287_1735 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_288_1736 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_288_1737 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_288_1738 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_289_1739 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_289_1740 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_290_1741 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_290_1742 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_290_1743 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_291_1744 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_291_1745 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_292_1746 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_292_1747 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_292_1748 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_293_1749 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_293_1750 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_294_1751 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_294_1752 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_294_1753 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_295_1754 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_295_1755 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_296_1756 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_296_1757 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_296_1758 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_297_1759 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_297_1760 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_298_1761 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_298_1762 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_298_1763 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_299_1764 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_299_1765 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_300_1766 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_300_1767 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_300_1768 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_301_1769 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_301_1770 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_302_1771 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_302_1772 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_302_1773 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_303_1774 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_303_1775 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_304_1776 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_304_1777 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_304_1778 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_305_1779 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_305_1780 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_306_1781 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_306_1782 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_306_1783 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_307_1784 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_307_1785 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_308_1786 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_308_1787 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_308_1788 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_309_1789 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_309_1790 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_310_1791 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_310_1792 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_310_1793 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_311_1794 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_311_1795 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_312_1796 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_312_1797 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_312_1798 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_313_1799 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_313_1800 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_314_1801 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_314_1802 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_314_1803 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_315_1804 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_315_1805 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_316_1806 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_316_1807 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_316_1808 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_317_1809 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_317_1810 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_318_1811 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_318_1812 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_318_1813 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_319_1814 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_319_1815 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_320_1816 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_320_1817 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_320_1818 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_321_1819 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_321_1820 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_322_1821 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_322_1822 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_322_1823 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_323_1824 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_323_1825 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_324_1826 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_324_1827 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_324_1828 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_325_1829 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_325_1830 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_326_1831 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_326_1832 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_326_1833 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_327_1834 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_327_1835 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_328_1836 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_328_1837 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_328_1838 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_329_1839 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_329_1840 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_330_1841 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_330_1842 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_330_1843 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_331_1844 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_331_1845 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_332_1846 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_332_1847 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_332_1848 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_333_1849 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_333_1850 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_334_1851 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_334_1852 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_334_1853 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_335_1854 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_335_1855 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_336_1856 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_336_1857 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_336_1858 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_337_1859 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_337_1860 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_338_1861 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_338_1862 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_338_1863 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_339_1864 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_339_1865 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_340_1866 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_340_1867 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_340_1868 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_341_1869 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_341_1870 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_342_1871 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_342_1872 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_342_1873 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_343_1874 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_343_1875 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_344_1876 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_344_1877 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_344_1878 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_345_1879 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_345_1880 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_346_1881 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_346_1882 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_346_1883 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_347_1884 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_347_1885 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_348_1886 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_348_1887 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_348_1888 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_349_1889 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_349_1890 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_350_1891 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_350_1892 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_350_1893 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_351_1894 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_351_1895 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_352_1896 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_352_1897 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_352_1898 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_353_1899 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_353_1900 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_354_1901 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_354_1902 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_354_1903 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_355_1904 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_355_1905 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_356_1906 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_356_1907 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_356_1908 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_357_1909 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_357_1910 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_358_1911 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_358_1912 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_358_1913 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_359_1914 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_359_1915 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_360_1916 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_360_1917 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_360_1918 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_361_1919 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_361_1920 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_362_1921 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_362_1922 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_362_1923 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_363_1924 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_363_1925 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_364_1926 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_364_1927 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_364_1928 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_365_1929 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_365_1930 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_366_1931 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_366_1932 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_366_1933 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_367_1934 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_367_1935 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_368_1936 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_368_1937 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_368_1938 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_369_1939 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_369_1940 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_370_1941 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_370_1942 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_370_1943 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_371_1944 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_371_1945 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_372_1946 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_372_1947 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_372_1948 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_373_1949 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_373_1950 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_374_1951 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_374_1952 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_374_1953 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_375_1954 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_375_1955 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_376_1956 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_376_1957 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_376_1958 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_377_1959 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_377_1960 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_378_1961 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_378_1962 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_378_1963 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_379_1964 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_379_1965 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_380_1966 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_380_1967 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_380_1968 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_381_1969 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_381_1970 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_382_1971 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_382_1972 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_382_1973 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_383_1974 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_383_1975 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_384_1976 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_384_1977 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_384_1978 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_385_1979 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_385_1980 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_386_1981 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_386_1982 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_386_1983 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_387_1984 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_387_1985 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_388_1986 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_388_1987 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_388_1988 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_389_1989 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_389_1990 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_390_1991 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_390_1992 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_390_1993 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_391_1994 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_391_1995 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_392_1996 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_392_1997 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_392_1998 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_393_1999 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_393_2000 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_394_2001 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_394_2002 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_394_2003 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_395_2004 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_395_2005 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_396_2006 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_396_2007 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_396_2008 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_397_2009 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_397_2010 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_398_2011 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_398_2012 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_398_2013 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_399_2014 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_399_2015 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_400_2016 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_400_2017 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_400_2018 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_401_2019 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_401_2020 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_402_2021 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_402_2022 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_402_2023 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_403_2024 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_403_2025 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_404_2026 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_404_2027 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_404_2028 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_405_2029 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_405_2030 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_406_2031 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_406_2032 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_406_2033 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_407_2034 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_407_2035 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_408_2036 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_408_2037 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_408_2038 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_409_2039 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_409_2040 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_410_2041 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_410_2042 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_410_2043 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_411_2044 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_411_2045 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_412_2046 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_412_2047 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_412_2048 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_413_2049 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_413_2050 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_414_2051 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_414_2052 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_414_2053 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_415_2054 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_415_2055 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_416_2056 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_416_2057 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_416_2058 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_417_2059 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_417_2060 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_418_2061 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_418_2062 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_418_2063 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_419_2064 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_419_2065 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_420_2066 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_420_2067 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_420_2068 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_421_2069 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_421_2070 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_422_2071 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_422_2072 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_422_2073 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_423_2074 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_423_2075 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_424_2076 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_424_2077 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_424_2078 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_425_2079 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_425_2080 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_426_2081 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_426_2082 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_426_2083 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_427_2084 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_427_2085 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_428_2086 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_428_2087 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_428_2088 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_429_2089 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_429_2090 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_430_2091 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_430_2092 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_430_2093 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_431_2094 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_431_2095 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_432_2096 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_432_2097 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_432_2098 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_433_2099 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_433_2100 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_434_2101 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_434_2102 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_434_2103 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_435_2104 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_435_2105 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_436_2106 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_436_2107 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_436_2108 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_437_2109 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_437_2110 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_438_2111 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_438_2112 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_438_2113 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_439_2114 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_439_2115 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_440_2116 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_440_2117 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_440_2118 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_441_2119 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_441_2120 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_442_2121 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_442_2122 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_442_2123 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_443_2124 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_443_2125 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_444_2126 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_444_2127 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_444_2128 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_445_2129 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_445_2130 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_446_2131 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_446_2132 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_446_2133 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_447_2134 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_447_2135 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_448_2136 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_448_2137 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_448_2138 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_449_2139 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_449_2140 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_450_2141 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_450_2142 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_450_2143 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_451_2144 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_451_2145 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_452_2146 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_452_2147 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_452_2148 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_453_2149 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_453_2150 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_454_2151 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_454_2152 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_454_2153 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_455_2154 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_455_2155 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_456_2156 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_456_2157 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_456_2158 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_457_2159 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_457_2160 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_458_2161 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_458_2162 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_458_2163 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_459_2164 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_459_2165 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_460_2166 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_460_2167 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_460_2168 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_461_2169 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_461_2170 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_462_2171 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_462_2172 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_462_2173 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_463_2174 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_463_2175 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_464_2176 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_464_2177 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_464_2178 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_465_2179 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_465_2180 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_466_2181 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_466_2182 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_466_2183 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_467_2184 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_467_2185 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_468_2186 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_468_2187 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_468_2188 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_469_2189 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_469_2190 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_470_2191 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_470_2192 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_470_2193 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_471_2194 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_471_2195 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_472_2196 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_472_2197 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_472_2198 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_473_2199 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_473_2200 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_474_2201 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_474_2202 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_474_2203 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_475_2204 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_475_2205 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_476_2206 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_476_2207 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_476_2208 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_477_2209 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_477_2210 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_478_2211 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_478_2212 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_478_2213 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_479_2214 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_479_2215 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_480_2216 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_480_2217 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_480_2218 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_481_2219 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_481_2220 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_482_2221 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_482_2222 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_482_2223 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_483_2224 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_483_2225 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_484_2226 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_484_2227 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_484_2228 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_485_2229 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_485_2230 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_486_2231 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_486_2232 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_486_2233 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_487_2234 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_487_2235 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_488_2236 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_488_2237 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_488_2238 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_489_2239 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_489_2240 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_490_2241 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_490_2242 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_490_2243 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_491_2244 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_491_2245 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_492_2246 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_492_2247 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_492_2248 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_493_2249 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_493_2250 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_494_2251 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_494_2252 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_494_2253 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_495_2254 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_495_2255 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_496_2256 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_496_2257 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_496_2258 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_497_2259 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_497_2260 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_498_2261 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_498_2262 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_498_2263 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_499_2264 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_499_2265 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_500_2266 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_500_2267 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_500_2268 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_501_2269 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_501_2270 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_502_2271 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_502_2272 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_502_2273 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_503_2274 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_503_2275 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_504_2276 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_504_2277 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_504_2278 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_505_2279 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_505_2280 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_506_2281 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_506_2282 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_506_2283 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_506_2284 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_506_2285 ();
 BUF_X1 output1 (.A(net1),
    .Z(a_almost_empty));
 BUF_X1 output2 (.A(net2),
    .Z(a_almost_full));
 BUF_X1 output3 (.A(net3),
    .Z(a_empty));
 BUF_X1 output4 (.A(net4),
    .Z(a_full));
 BUF_X1 output5 (.A(net5),
    .Z(a_rd_data[0]));
 BUF_X1 output6 (.A(net6),
    .Z(a_rd_data[1]));
 BUF_X1 output7 (.A(net7),
    .Z(a_rd_data[2]));
 BUF_X1 output8 (.A(net8),
    .Z(a_rd_data[3]));
 BUF_X1 output9 (.A(net9),
    .Z(a_rd_data[4]));
 BUF_X1 output10 (.A(net10),
    .Z(a_rd_data[5]));
 BUF_X1 output11 (.A(net11),
    .Z(a_rd_data[6]));
 BUF_X1 output12 (.A(net12),
    .Z(a_rd_data[7]));
 BUF_X1 output13 (.A(net13),
    .Z(a_to_b_count[0]));
 BUF_X1 output14 (.A(net40),
    .Z(a_to_b_count[1]));
 BUF_X1 output15 (.A(net41),
    .Z(a_to_b_count[2]));
 BUF_X1 output16 (.A(net16),
    .Z(a_to_b_count[3]));
 BUF_X1 output17 (.A(_0795_),
    .Z(a_to_b_count[4]));
 BUF_X1 output18 (.A(net18),
    .Z(b_almost_empty));
 BUF_X1 output19 (.A(net19),
    .Z(b_almost_full));
 BUF_X1 output20 (.A(net20),
    .Z(b_empty));
 BUF_X1 output21 (.A(net21),
    .Z(b_full));
 BUF_X1 output22 (.A(net22),
    .Z(b_rd_data[0]));
 BUF_X1 output23 (.A(net23),
    .Z(b_rd_data[1]));
 BUF_X1 output24 (.A(net24),
    .Z(b_rd_data[2]));
 BUF_X1 output25 (.A(net25),
    .Z(b_rd_data[3]));
 BUF_X1 output26 (.A(net26),
    .Z(b_rd_data[4]));
 BUF_X1 output27 (.A(net27),
    .Z(b_rd_data[5]));
 BUF_X1 output28 (.A(net28),
    .Z(b_rd_data[6]));
 BUF_X1 output29 (.A(net29),
    .Z(b_rd_data[7]));
 BUF_X1 output30 (.A(net30),
    .Z(b_to_a_count[0]));
 BUF_X1 output31 (.A(net35),
    .Z(b_to_a_count[1]));
 BUF_X1 output32 (.A(net39),
    .Z(b_to_a_count[2]));
 BUF_X1 output33 (.A(net33),
    .Z(b_to_a_count[3]));
 BUF_X1 output34 (.A(net34),
    .Z(b_to_a_count[4]));
 CLKBUF_X3 clkbuf_leaf_0_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_0_clk));
 CLKBUF_X3 clkbuf_leaf_1_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_1_clk));
 CLKBUF_X3 clkbuf_leaf_2_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_2_clk));
 CLKBUF_X3 clkbuf_leaf_3_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_3_clk));
 CLKBUF_X3 clkbuf_leaf_4_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_4_clk));
 CLKBUF_X3 clkbuf_leaf_5_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_5_clk));
 CLKBUF_X3 clkbuf_leaf_6_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_6_clk));
 CLKBUF_X3 clkbuf_leaf_7_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_7_clk));
 CLKBUF_X3 clkbuf_leaf_8_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_8_clk));
 CLKBUF_X3 clkbuf_leaf_9_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_9_clk));
 CLKBUF_X3 clkbuf_leaf_10_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_10_clk));
 CLKBUF_X3 clkbuf_leaf_11_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_11_clk));
 CLKBUF_X3 clkbuf_leaf_12_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_12_clk));
 CLKBUF_X3 clkbuf_leaf_13_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_13_clk));
 CLKBUF_X3 clkbuf_leaf_14_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_14_clk));
 CLKBUF_X3 clkbuf_leaf_15_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_15_clk));
 CLKBUF_X3 clkbuf_leaf_16_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_16_clk));
 CLKBUF_X3 clkbuf_leaf_17_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_17_clk));
 CLKBUF_X3 clkbuf_leaf_18_clk (.A(clknet_2_1__leaf_clk),
    .Z(clknet_leaf_18_clk));
 CLKBUF_X3 clkbuf_leaf_19_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_19_clk));
 CLKBUF_X3 clkbuf_leaf_20_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_20_clk));
 CLKBUF_X3 clkbuf_leaf_21_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_21_clk));
 CLKBUF_X3 clkbuf_leaf_22_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_22_clk));
 CLKBUF_X3 clkbuf_leaf_23_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_23_clk));
 CLKBUF_X3 clkbuf_leaf_24_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_24_clk));
 CLKBUF_X3 clkbuf_leaf_25_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_25_clk));
 CLKBUF_X3 clkbuf_leaf_26_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_26_clk));
 CLKBUF_X3 clkbuf_leaf_27_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_27_clk));
 CLKBUF_X3 clkbuf_leaf_28_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_28_clk));
 CLKBUF_X3 clkbuf_leaf_29_clk (.A(clknet_2_3__leaf_clk),
    .Z(clknet_leaf_29_clk));
 CLKBUF_X3 clkbuf_leaf_30_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_30_clk));
 CLKBUF_X3 clkbuf_leaf_31_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_31_clk));
 CLKBUF_X3 clkbuf_leaf_32_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_32_clk));
 CLKBUF_X3 clkbuf_leaf_33_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_33_clk));
 CLKBUF_X3 clkbuf_leaf_34_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_34_clk));
 CLKBUF_X3 clkbuf_leaf_35_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_35_clk));
 CLKBUF_X3 clkbuf_leaf_36_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_36_clk));
 CLKBUF_X3 clkbuf_leaf_37_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_37_clk));
 CLKBUF_X3 clkbuf_leaf_38_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_38_clk));
 CLKBUF_X3 clkbuf_leaf_39_clk (.A(clknet_2_2__leaf_clk),
    .Z(clknet_leaf_39_clk));
 CLKBUF_X3 clkbuf_leaf_40_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_40_clk));
 CLKBUF_X3 clkbuf_leaf_41_clk (.A(clknet_2_0__leaf_clk),
    .Z(clknet_leaf_41_clk));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 CLKBUF_X3 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 CLKBUF_X3 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 CLKBUF_X3 clkload0 (.A(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkload1 (.A(clknet_2_3__leaf_clk));
 CLKBUF_X1 clkload2 (.A(clknet_leaf_0_clk));
 CLKBUF_X1 clkload3 (.A(clknet_leaf_1_clk));
 CLKBUF_X1 clkload4 (.A(clknet_leaf_2_clk));
 CLKBUF_X1 clkload5 (.A(clknet_leaf_4_clk));
 INV_X1 clkload6 (.A(clknet_leaf_5_clk));
 INV_X1 clkload7 (.A(clknet_leaf_6_clk));
 CLKBUF_X1 clkload8 (.A(clknet_leaf_8_clk));
 INV_X1 clkload9 (.A(clknet_leaf_40_clk));
 INV_X2 clkload10 (.A(clknet_leaf_41_clk));
 INV_X2 clkload11 (.A(clknet_leaf_7_clk));
 INV_X1 clkload12 (.A(clknet_leaf_9_clk));
 INV_X1 clkload13 (.A(clknet_leaf_10_clk));
 CLKBUF_X1 clkload14 (.A(clknet_leaf_11_clk));
 INV_X1 clkload15 (.A(clknet_leaf_13_clk));
 CLKBUF_X1 clkload16 (.A(clknet_leaf_14_clk));
 INV_X1 clkload17 (.A(clknet_leaf_15_clk));
 CLKBUF_X1 clkload18 (.A(clknet_leaf_16_clk));
 INV_X2 clkload19 (.A(clknet_leaf_17_clk));
 INV_X1 clkload20 (.A(clknet_leaf_18_clk));
 INV_X1 clkload21 (.A(clknet_leaf_27_clk));
 CLKBUF_X1 clkload22 (.A(clknet_leaf_30_clk));
 CLKBUF_X1 clkload23 (.A(clknet_leaf_31_clk));
 CLKBUF_X1 clkload24 (.A(clknet_leaf_33_clk));
 CLKBUF_X1 clkload25 (.A(clknet_leaf_34_clk));
 CLKBUF_X1 clkload26 (.A(clknet_leaf_36_clk));
 INV_X1 clkload27 (.A(clknet_leaf_37_clk));
 INV_X1 clkload28 (.A(clknet_leaf_38_clk));
 CLKBUF_X1 clkload29 (.A(clknet_leaf_39_clk));
 INV_X2 clkload30 (.A(clknet_leaf_19_clk));
 CLKBUF_X1 clkload31 (.A(clknet_leaf_20_clk));
 CLKBUF_X1 clkload32 (.A(clknet_leaf_21_clk));
 CLKBUF_X1 clkload33 (.A(clknet_leaf_22_clk));
 CLKBUF_X1 clkload34 (.A(clknet_leaf_23_clk));
 CLKBUF_X1 clkload35 (.A(clknet_leaf_24_clk));
 CLKBUF_X1 clkload36 (.A(clknet_leaf_26_clk));
 CLKBUF_X1 clkload37 (.A(clknet_leaf_28_clk));
 BUF_X1 rebuffer1 (.A(net31),
    .Z(net35));
 BUF_X1 rebuffer2 (.A(_0806_),
    .Z(net36));
 BUF_X1 rebuffer3 (.A(_0794_),
    .Z(net37));
 BUF_X2 rebuffer4 (.A(_1218_),
    .Z(net38));
 BUF_X1 rebuffer5 (.A(net32),
    .Z(net39));
 BUF_X1 rebuffer7 (.A(net15),
    .Z(net41));
 BUF_X1 rebuffer8 (.A(_0794_),
    .Z(net43));
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X32 FILLER_0_257 ();
 FILLCELL_X32 FILLER_0_289 ();
 FILLCELL_X32 FILLER_0_321 ();
 FILLCELL_X32 FILLER_0_353 ();
 FILLCELL_X32 FILLER_0_385 ();
 FILLCELL_X32 FILLER_0_417 ();
 FILLCELL_X32 FILLER_0_449 ();
 FILLCELL_X32 FILLER_0_481 ();
 FILLCELL_X32 FILLER_0_513 ();
 FILLCELL_X32 FILLER_0_545 ();
 FILLCELL_X32 FILLER_0_577 ();
 FILLCELL_X16 FILLER_0_609 ();
 FILLCELL_X4 FILLER_0_625 ();
 FILLCELL_X2 FILLER_0_629 ();
 FILLCELL_X32 FILLER_0_632 ();
 FILLCELL_X32 FILLER_0_664 ();
 FILLCELL_X32 FILLER_0_696 ();
 FILLCELL_X32 FILLER_0_728 ();
 FILLCELL_X32 FILLER_0_760 ();
 FILLCELL_X32 FILLER_0_792 ();
 FILLCELL_X32 FILLER_0_824 ();
 FILLCELL_X32 FILLER_0_856 ();
 FILLCELL_X32 FILLER_0_888 ();
 FILLCELL_X32 FILLER_0_920 ();
 FILLCELL_X32 FILLER_0_952 ();
 FILLCELL_X32 FILLER_0_984 ();
 FILLCELL_X32 FILLER_0_1016 ();
 FILLCELL_X32 FILLER_0_1048 ();
 FILLCELL_X32 FILLER_0_1080 ();
 FILLCELL_X32 FILLER_0_1112 ();
 FILLCELL_X32 FILLER_0_1144 ();
 FILLCELL_X32 FILLER_0_1176 ();
 FILLCELL_X32 FILLER_0_1208 ();
 FILLCELL_X16 FILLER_0_1240 ();
 FILLCELL_X4 FILLER_0_1256 ();
 FILLCELL_X2 FILLER_0_1260 ();
 FILLCELL_X32 FILLER_0_1263 ();
 FILLCELL_X32 FILLER_0_1295 ();
 FILLCELL_X32 FILLER_0_1327 ();
 FILLCELL_X32 FILLER_0_1359 ();
 FILLCELL_X32 FILLER_0_1391 ();
 FILLCELL_X32 FILLER_0_1423 ();
 FILLCELL_X32 FILLER_0_1455 ();
 FILLCELL_X32 FILLER_0_1487 ();
 FILLCELL_X32 FILLER_0_1519 ();
 FILLCELL_X32 FILLER_0_1551 ();
 FILLCELL_X32 FILLER_0_1583 ();
 FILLCELL_X32 FILLER_0_1615 ();
 FILLCELL_X32 FILLER_0_1647 ();
 FILLCELL_X32 FILLER_0_1679 ();
 FILLCELL_X32 FILLER_0_1711 ();
 FILLCELL_X32 FILLER_0_1743 ();
 FILLCELL_X32 FILLER_0_1775 ();
 FILLCELL_X32 FILLER_0_1807 ();
 FILLCELL_X32 FILLER_0_1839 ();
 FILLCELL_X4 FILLER_0_1871 ();
 FILLCELL_X2 FILLER_0_1875 ();
 FILLCELL_X1 FILLER_0_1877 ();
 FILLCELL_X4 FILLER_0_1887 ();
 FILLCELL_X2 FILLER_0_1891 ();
 FILLCELL_X4 FILLER_0_1894 ();
 FILLCELL_X1 FILLER_0_1898 ();
 FILLCELL_X2 FILLER_0_1902 ();
 FILLCELL_X1 FILLER_0_1904 ();
 FILLCELL_X16 FILLER_0_1908 ();
 FILLCELL_X4 FILLER_0_1924 ();
 FILLCELL_X2 FILLER_0_1928 ();
 FILLCELL_X16 FILLER_0_1933 ();
 FILLCELL_X8 FILLER_0_1949 ();
 FILLCELL_X2 FILLER_0_1957 ();
 FILLCELL_X1 FILLER_0_1959 ();
 FILLCELL_X4 FILLER_0_1963 ();
 FILLCELL_X32 FILLER_0_1970 ();
 FILLCELL_X8 FILLER_0_2002 ();
 FILLCELL_X1 FILLER_0_2010 ();
 FILLCELL_X32 FILLER_0_2014 ();
 FILLCELL_X32 FILLER_0_2046 ();
 FILLCELL_X32 FILLER_0_2078 ();
 FILLCELL_X32 FILLER_0_2110 ();
 FILLCELL_X32 FILLER_0_2142 ();
 FILLCELL_X32 FILLER_0_2174 ();
 FILLCELL_X32 FILLER_0_2206 ();
 FILLCELL_X32 FILLER_0_2238 ();
 FILLCELL_X32 FILLER_0_2270 ();
 FILLCELL_X32 FILLER_0_2302 ();
 FILLCELL_X32 FILLER_0_2334 ();
 FILLCELL_X32 FILLER_0_2366 ();
 FILLCELL_X32 FILLER_0_2398 ();
 FILLCELL_X32 FILLER_0_2430 ();
 FILLCELL_X32 FILLER_0_2462 ();
 FILLCELL_X16 FILLER_0_2494 ();
 FILLCELL_X8 FILLER_0_2510 ();
 FILLCELL_X4 FILLER_0_2518 ();
 FILLCELL_X2 FILLER_0_2522 ();
 FILLCELL_X32 FILLER_0_2525 ();
 FILLCELL_X32 FILLER_0_2557 ();
 FILLCELL_X32 FILLER_0_2589 ();
 FILLCELL_X32 FILLER_0_2621 ();
 FILLCELL_X32 FILLER_0_2653 ();
 FILLCELL_X32 FILLER_0_2685 ();
 FILLCELL_X32 FILLER_0_2717 ();
 FILLCELL_X32 FILLER_0_2749 ();
 FILLCELL_X32 FILLER_0_2781 ();
 FILLCELL_X32 FILLER_0_2813 ();
 FILLCELL_X32 FILLER_0_2845 ();
 FILLCELL_X32 FILLER_0_2877 ();
 FILLCELL_X32 FILLER_0_2909 ();
 FILLCELL_X32 FILLER_0_2941 ();
 FILLCELL_X32 FILLER_0_2973 ();
 FILLCELL_X32 FILLER_0_3005 ();
 FILLCELL_X32 FILLER_0_3037 ();
 FILLCELL_X32 FILLER_0_3069 ();
 FILLCELL_X32 FILLER_0_3101 ();
 FILLCELL_X16 FILLER_0_3133 ();
 FILLCELL_X4 FILLER_0_3149 ();
 FILLCELL_X2 FILLER_0_3153 ();
 FILLCELL_X32 FILLER_0_3156 ();
 FILLCELL_X32 FILLER_0_3188 ();
 FILLCELL_X32 FILLER_0_3220 ();
 FILLCELL_X32 FILLER_0_3252 ();
 FILLCELL_X32 FILLER_0_3284 ();
 FILLCELL_X32 FILLER_0_3316 ();
 FILLCELL_X32 FILLER_0_3348 ();
 FILLCELL_X32 FILLER_0_3380 ();
 FILLCELL_X32 FILLER_0_3412 ();
 FILLCELL_X32 FILLER_0_3444 ();
 FILLCELL_X32 FILLER_0_3476 ();
 FILLCELL_X32 FILLER_0_3508 ();
 FILLCELL_X32 FILLER_0_3540 ();
 FILLCELL_X32 FILLER_0_3572 ();
 FILLCELL_X32 FILLER_0_3604 ();
 FILLCELL_X32 FILLER_0_3636 ();
 FILLCELL_X32 FILLER_0_3668 ();
 FILLCELL_X32 FILLER_0_3700 ();
 FILLCELL_X4 FILLER_0_3732 ();
 FILLCELL_X2 FILLER_0_3736 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X32 FILLER_1_321 ();
 FILLCELL_X32 FILLER_1_353 ();
 FILLCELL_X32 FILLER_1_385 ();
 FILLCELL_X32 FILLER_1_417 ();
 FILLCELL_X32 FILLER_1_449 ();
 FILLCELL_X32 FILLER_1_481 ();
 FILLCELL_X32 FILLER_1_513 ();
 FILLCELL_X32 FILLER_1_545 ();
 FILLCELL_X32 FILLER_1_577 ();
 FILLCELL_X32 FILLER_1_609 ();
 FILLCELL_X32 FILLER_1_641 ();
 FILLCELL_X32 FILLER_1_673 ();
 FILLCELL_X32 FILLER_1_705 ();
 FILLCELL_X32 FILLER_1_737 ();
 FILLCELL_X32 FILLER_1_769 ();
 FILLCELL_X32 FILLER_1_801 ();
 FILLCELL_X32 FILLER_1_833 ();
 FILLCELL_X32 FILLER_1_865 ();
 FILLCELL_X32 FILLER_1_897 ();
 FILLCELL_X32 FILLER_1_929 ();
 FILLCELL_X32 FILLER_1_961 ();
 FILLCELL_X32 FILLER_1_993 ();
 FILLCELL_X32 FILLER_1_1025 ();
 FILLCELL_X32 FILLER_1_1057 ();
 FILLCELL_X32 FILLER_1_1089 ();
 FILLCELL_X32 FILLER_1_1121 ();
 FILLCELL_X32 FILLER_1_1153 ();
 FILLCELL_X32 FILLER_1_1185 ();
 FILLCELL_X32 FILLER_1_1217 ();
 FILLCELL_X8 FILLER_1_1249 ();
 FILLCELL_X4 FILLER_1_1257 ();
 FILLCELL_X2 FILLER_1_1261 ();
 FILLCELL_X32 FILLER_1_1264 ();
 FILLCELL_X32 FILLER_1_1296 ();
 FILLCELL_X32 FILLER_1_1328 ();
 FILLCELL_X32 FILLER_1_1360 ();
 FILLCELL_X32 FILLER_1_1392 ();
 FILLCELL_X32 FILLER_1_1424 ();
 FILLCELL_X32 FILLER_1_1456 ();
 FILLCELL_X32 FILLER_1_1488 ();
 FILLCELL_X32 FILLER_1_1520 ();
 FILLCELL_X32 FILLER_1_1552 ();
 FILLCELL_X32 FILLER_1_1584 ();
 FILLCELL_X32 FILLER_1_1616 ();
 FILLCELL_X32 FILLER_1_1648 ();
 FILLCELL_X32 FILLER_1_1680 ();
 FILLCELL_X32 FILLER_1_1712 ();
 FILLCELL_X32 FILLER_1_1744 ();
 FILLCELL_X32 FILLER_1_1776 ();
 FILLCELL_X32 FILLER_1_1808 ();
 FILLCELL_X32 FILLER_1_1840 ();
 FILLCELL_X16 FILLER_1_1872 ();
 FILLCELL_X8 FILLER_1_1888 ();
 FILLCELL_X1 FILLER_1_1896 ();
 FILLCELL_X8 FILLER_1_1903 ();
 FILLCELL_X4 FILLER_1_1911 ();
 FILLCELL_X32 FILLER_1_1918 ();
 FILLCELL_X1 FILLER_1_1950 ();
 FILLCELL_X32 FILLER_1_1954 ();
 FILLCELL_X32 FILLER_1_1986 ();
 FILLCELL_X32 FILLER_1_2018 ();
 FILLCELL_X32 FILLER_1_2050 ();
 FILLCELL_X32 FILLER_1_2082 ();
 FILLCELL_X32 FILLER_1_2114 ();
 FILLCELL_X32 FILLER_1_2146 ();
 FILLCELL_X32 FILLER_1_2178 ();
 FILLCELL_X32 FILLER_1_2210 ();
 FILLCELL_X32 FILLER_1_2242 ();
 FILLCELL_X32 FILLER_1_2274 ();
 FILLCELL_X32 FILLER_1_2306 ();
 FILLCELL_X32 FILLER_1_2338 ();
 FILLCELL_X32 FILLER_1_2370 ();
 FILLCELL_X32 FILLER_1_2402 ();
 FILLCELL_X32 FILLER_1_2434 ();
 FILLCELL_X32 FILLER_1_2466 ();
 FILLCELL_X16 FILLER_1_2498 ();
 FILLCELL_X8 FILLER_1_2514 ();
 FILLCELL_X4 FILLER_1_2522 ();
 FILLCELL_X32 FILLER_1_2527 ();
 FILLCELL_X32 FILLER_1_2559 ();
 FILLCELL_X32 FILLER_1_2591 ();
 FILLCELL_X32 FILLER_1_2623 ();
 FILLCELL_X32 FILLER_1_2655 ();
 FILLCELL_X32 FILLER_1_2687 ();
 FILLCELL_X32 FILLER_1_2719 ();
 FILLCELL_X32 FILLER_1_2751 ();
 FILLCELL_X32 FILLER_1_2783 ();
 FILLCELL_X32 FILLER_1_2815 ();
 FILLCELL_X32 FILLER_1_2847 ();
 FILLCELL_X32 FILLER_1_2879 ();
 FILLCELL_X32 FILLER_1_2911 ();
 FILLCELL_X32 FILLER_1_2943 ();
 FILLCELL_X32 FILLER_1_2975 ();
 FILLCELL_X32 FILLER_1_3007 ();
 FILLCELL_X32 FILLER_1_3039 ();
 FILLCELL_X32 FILLER_1_3071 ();
 FILLCELL_X32 FILLER_1_3103 ();
 FILLCELL_X32 FILLER_1_3135 ();
 FILLCELL_X32 FILLER_1_3167 ();
 FILLCELL_X32 FILLER_1_3199 ();
 FILLCELL_X32 FILLER_1_3231 ();
 FILLCELL_X32 FILLER_1_3263 ();
 FILLCELL_X32 FILLER_1_3295 ();
 FILLCELL_X32 FILLER_1_3327 ();
 FILLCELL_X32 FILLER_1_3359 ();
 FILLCELL_X32 FILLER_1_3391 ();
 FILLCELL_X32 FILLER_1_3423 ();
 FILLCELL_X32 FILLER_1_3455 ();
 FILLCELL_X32 FILLER_1_3487 ();
 FILLCELL_X32 FILLER_1_3519 ();
 FILLCELL_X32 FILLER_1_3551 ();
 FILLCELL_X32 FILLER_1_3583 ();
 FILLCELL_X32 FILLER_1_3615 ();
 FILLCELL_X32 FILLER_1_3647 ();
 FILLCELL_X32 FILLER_1_3679 ();
 FILLCELL_X16 FILLER_1_3711 ();
 FILLCELL_X8 FILLER_1_3727 ();
 FILLCELL_X2 FILLER_1_3735 ();
 FILLCELL_X1 FILLER_1_3737 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X32 FILLER_2_385 ();
 FILLCELL_X32 FILLER_2_417 ();
 FILLCELL_X32 FILLER_2_449 ();
 FILLCELL_X32 FILLER_2_481 ();
 FILLCELL_X32 FILLER_2_513 ();
 FILLCELL_X32 FILLER_2_545 ();
 FILLCELL_X32 FILLER_2_577 ();
 FILLCELL_X16 FILLER_2_609 ();
 FILLCELL_X4 FILLER_2_625 ();
 FILLCELL_X2 FILLER_2_629 ();
 FILLCELL_X32 FILLER_2_632 ();
 FILLCELL_X32 FILLER_2_664 ();
 FILLCELL_X32 FILLER_2_696 ();
 FILLCELL_X32 FILLER_2_728 ();
 FILLCELL_X32 FILLER_2_760 ();
 FILLCELL_X32 FILLER_2_792 ();
 FILLCELL_X32 FILLER_2_824 ();
 FILLCELL_X32 FILLER_2_856 ();
 FILLCELL_X32 FILLER_2_888 ();
 FILLCELL_X32 FILLER_2_920 ();
 FILLCELL_X32 FILLER_2_952 ();
 FILLCELL_X32 FILLER_2_984 ();
 FILLCELL_X32 FILLER_2_1016 ();
 FILLCELL_X32 FILLER_2_1048 ();
 FILLCELL_X32 FILLER_2_1080 ();
 FILLCELL_X32 FILLER_2_1112 ();
 FILLCELL_X32 FILLER_2_1144 ();
 FILLCELL_X32 FILLER_2_1176 ();
 FILLCELL_X32 FILLER_2_1208 ();
 FILLCELL_X32 FILLER_2_1240 ();
 FILLCELL_X32 FILLER_2_1272 ();
 FILLCELL_X32 FILLER_2_1304 ();
 FILLCELL_X32 FILLER_2_1336 ();
 FILLCELL_X32 FILLER_2_1368 ();
 FILLCELL_X32 FILLER_2_1400 ();
 FILLCELL_X32 FILLER_2_1432 ();
 FILLCELL_X32 FILLER_2_1464 ();
 FILLCELL_X32 FILLER_2_1496 ();
 FILLCELL_X32 FILLER_2_1528 ();
 FILLCELL_X32 FILLER_2_1560 ();
 FILLCELL_X32 FILLER_2_1592 ();
 FILLCELL_X32 FILLER_2_1624 ();
 FILLCELL_X32 FILLER_2_1656 ();
 FILLCELL_X32 FILLER_2_1688 ();
 FILLCELL_X32 FILLER_2_1720 ();
 FILLCELL_X32 FILLER_2_1752 ();
 FILLCELL_X32 FILLER_2_1784 ();
 FILLCELL_X32 FILLER_2_1816 ();
 FILLCELL_X32 FILLER_2_1848 ();
 FILLCELL_X8 FILLER_2_1880 ();
 FILLCELL_X4 FILLER_2_1888 ();
 FILLCELL_X2 FILLER_2_1892 ();
 FILLCELL_X32 FILLER_2_1895 ();
 FILLCELL_X32 FILLER_2_1927 ();
 FILLCELL_X32 FILLER_2_1959 ();
 FILLCELL_X32 FILLER_2_1991 ();
 FILLCELL_X32 FILLER_2_2023 ();
 FILLCELL_X32 FILLER_2_2055 ();
 FILLCELL_X32 FILLER_2_2087 ();
 FILLCELL_X32 FILLER_2_2119 ();
 FILLCELL_X32 FILLER_2_2151 ();
 FILLCELL_X32 FILLER_2_2183 ();
 FILLCELL_X32 FILLER_2_2215 ();
 FILLCELL_X32 FILLER_2_2247 ();
 FILLCELL_X32 FILLER_2_2279 ();
 FILLCELL_X32 FILLER_2_2311 ();
 FILLCELL_X32 FILLER_2_2343 ();
 FILLCELL_X32 FILLER_2_2375 ();
 FILLCELL_X32 FILLER_2_2407 ();
 FILLCELL_X32 FILLER_2_2439 ();
 FILLCELL_X32 FILLER_2_2471 ();
 FILLCELL_X32 FILLER_2_2503 ();
 FILLCELL_X32 FILLER_2_2535 ();
 FILLCELL_X32 FILLER_2_2567 ();
 FILLCELL_X32 FILLER_2_2599 ();
 FILLCELL_X32 FILLER_2_2631 ();
 FILLCELL_X32 FILLER_2_2663 ();
 FILLCELL_X32 FILLER_2_2695 ();
 FILLCELL_X32 FILLER_2_2727 ();
 FILLCELL_X32 FILLER_2_2759 ();
 FILLCELL_X32 FILLER_2_2791 ();
 FILLCELL_X32 FILLER_2_2823 ();
 FILLCELL_X32 FILLER_2_2855 ();
 FILLCELL_X32 FILLER_2_2887 ();
 FILLCELL_X32 FILLER_2_2919 ();
 FILLCELL_X32 FILLER_2_2951 ();
 FILLCELL_X32 FILLER_2_2983 ();
 FILLCELL_X32 FILLER_2_3015 ();
 FILLCELL_X32 FILLER_2_3047 ();
 FILLCELL_X32 FILLER_2_3079 ();
 FILLCELL_X32 FILLER_2_3111 ();
 FILLCELL_X8 FILLER_2_3143 ();
 FILLCELL_X4 FILLER_2_3151 ();
 FILLCELL_X2 FILLER_2_3155 ();
 FILLCELL_X32 FILLER_2_3158 ();
 FILLCELL_X32 FILLER_2_3190 ();
 FILLCELL_X32 FILLER_2_3222 ();
 FILLCELL_X32 FILLER_2_3254 ();
 FILLCELL_X32 FILLER_2_3286 ();
 FILLCELL_X32 FILLER_2_3318 ();
 FILLCELL_X32 FILLER_2_3350 ();
 FILLCELL_X32 FILLER_2_3382 ();
 FILLCELL_X32 FILLER_2_3414 ();
 FILLCELL_X32 FILLER_2_3446 ();
 FILLCELL_X32 FILLER_2_3478 ();
 FILLCELL_X32 FILLER_2_3510 ();
 FILLCELL_X32 FILLER_2_3542 ();
 FILLCELL_X32 FILLER_2_3574 ();
 FILLCELL_X32 FILLER_2_3606 ();
 FILLCELL_X32 FILLER_2_3638 ();
 FILLCELL_X32 FILLER_2_3670 ();
 FILLCELL_X32 FILLER_2_3702 ();
 FILLCELL_X4 FILLER_2_3734 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X32 FILLER_3_385 ();
 FILLCELL_X32 FILLER_3_417 ();
 FILLCELL_X32 FILLER_3_449 ();
 FILLCELL_X32 FILLER_3_481 ();
 FILLCELL_X32 FILLER_3_513 ();
 FILLCELL_X32 FILLER_3_545 ();
 FILLCELL_X32 FILLER_3_577 ();
 FILLCELL_X32 FILLER_3_609 ();
 FILLCELL_X32 FILLER_3_641 ();
 FILLCELL_X32 FILLER_3_673 ();
 FILLCELL_X32 FILLER_3_705 ();
 FILLCELL_X32 FILLER_3_737 ();
 FILLCELL_X32 FILLER_3_769 ();
 FILLCELL_X32 FILLER_3_801 ();
 FILLCELL_X32 FILLER_3_833 ();
 FILLCELL_X32 FILLER_3_865 ();
 FILLCELL_X32 FILLER_3_897 ();
 FILLCELL_X32 FILLER_3_929 ();
 FILLCELL_X32 FILLER_3_961 ();
 FILLCELL_X32 FILLER_3_993 ();
 FILLCELL_X32 FILLER_3_1025 ();
 FILLCELL_X32 FILLER_3_1057 ();
 FILLCELL_X32 FILLER_3_1089 ();
 FILLCELL_X32 FILLER_3_1121 ();
 FILLCELL_X32 FILLER_3_1153 ();
 FILLCELL_X32 FILLER_3_1185 ();
 FILLCELL_X32 FILLER_3_1217 ();
 FILLCELL_X8 FILLER_3_1249 ();
 FILLCELL_X4 FILLER_3_1257 ();
 FILLCELL_X2 FILLER_3_1261 ();
 FILLCELL_X32 FILLER_3_1264 ();
 FILLCELL_X32 FILLER_3_1296 ();
 FILLCELL_X32 FILLER_3_1328 ();
 FILLCELL_X32 FILLER_3_1360 ();
 FILLCELL_X32 FILLER_3_1392 ();
 FILLCELL_X32 FILLER_3_1424 ();
 FILLCELL_X32 FILLER_3_1456 ();
 FILLCELL_X32 FILLER_3_1488 ();
 FILLCELL_X32 FILLER_3_1520 ();
 FILLCELL_X32 FILLER_3_1552 ();
 FILLCELL_X32 FILLER_3_1584 ();
 FILLCELL_X32 FILLER_3_1616 ();
 FILLCELL_X32 FILLER_3_1648 ();
 FILLCELL_X32 FILLER_3_1680 ();
 FILLCELL_X32 FILLER_3_1712 ();
 FILLCELL_X32 FILLER_3_1744 ();
 FILLCELL_X32 FILLER_3_1776 ();
 FILLCELL_X32 FILLER_3_1808 ();
 FILLCELL_X32 FILLER_3_1840 ();
 FILLCELL_X32 FILLER_3_1872 ();
 FILLCELL_X32 FILLER_3_1904 ();
 FILLCELL_X32 FILLER_3_1936 ();
 FILLCELL_X32 FILLER_3_1968 ();
 FILLCELL_X32 FILLER_3_2000 ();
 FILLCELL_X32 FILLER_3_2032 ();
 FILLCELL_X32 FILLER_3_2064 ();
 FILLCELL_X32 FILLER_3_2096 ();
 FILLCELL_X32 FILLER_3_2128 ();
 FILLCELL_X32 FILLER_3_2160 ();
 FILLCELL_X32 FILLER_3_2192 ();
 FILLCELL_X32 FILLER_3_2224 ();
 FILLCELL_X32 FILLER_3_2256 ();
 FILLCELL_X32 FILLER_3_2288 ();
 FILLCELL_X32 FILLER_3_2320 ();
 FILLCELL_X32 FILLER_3_2352 ();
 FILLCELL_X32 FILLER_3_2384 ();
 FILLCELL_X32 FILLER_3_2416 ();
 FILLCELL_X32 FILLER_3_2448 ();
 FILLCELL_X32 FILLER_3_2480 ();
 FILLCELL_X8 FILLER_3_2512 ();
 FILLCELL_X4 FILLER_3_2520 ();
 FILLCELL_X2 FILLER_3_2524 ();
 FILLCELL_X32 FILLER_3_2527 ();
 FILLCELL_X32 FILLER_3_2559 ();
 FILLCELL_X32 FILLER_3_2591 ();
 FILLCELL_X32 FILLER_3_2623 ();
 FILLCELL_X32 FILLER_3_2655 ();
 FILLCELL_X32 FILLER_3_2687 ();
 FILLCELL_X32 FILLER_3_2719 ();
 FILLCELL_X32 FILLER_3_2751 ();
 FILLCELL_X32 FILLER_3_2783 ();
 FILLCELL_X32 FILLER_3_2815 ();
 FILLCELL_X32 FILLER_3_2847 ();
 FILLCELL_X32 FILLER_3_2879 ();
 FILLCELL_X32 FILLER_3_2911 ();
 FILLCELL_X32 FILLER_3_2943 ();
 FILLCELL_X32 FILLER_3_2975 ();
 FILLCELL_X32 FILLER_3_3007 ();
 FILLCELL_X32 FILLER_3_3039 ();
 FILLCELL_X32 FILLER_3_3071 ();
 FILLCELL_X32 FILLER_3_3103 ();
 FILLCELL_X32 FILLER_3_3135 ();
 FILLCELL_X32 FILLER_3_3167 ();
 FILLCELL_X32 FILLER_3_3199 ();
 FILLCELL_X32 FILLER_3_3231 ();
 FILLCELL_X32 FILLER_3_3263 ();
 FILLCELL_X32 FILLER_3_3295 ();
 FILLCELL_X32 FILLER_3_3327 ();
 FILLCELL_X32 FILLER_3_3359 ();
 FILLCELL_X32 FILLER_3_3391 ();
 FILLCELL_X32 FILLER_3_3423 ();
 FILLCELL_X32 FILLER_3_3455 ();
 FILLCELL_X32 FILLER_3_3487 ();
 FILLCELL_X32 FILLER_3_3519 ();
 FILLCELL_X32 FILLER_3_3551 ();
 FILLCELL_X32 FILLER_3_3583 ();
 FILLCELL_X32 FILLER_3_3615 ();
 FILLCELL_X32 FILLER_3_3647 ();
 FILLCELL_X32 FILLER_3_3679 ();
 FILLCELL_X16 FILLER_3_3711 ();
 FILLCELL_X8 FILLER_3_3727 ();
 FILLCELL_X2 FILLER_3_3735 ();
 FILLCELL_X1 FILLER_3_3737 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X32 FILLER_4_353 ();
 FILLCELL_X32 FILLER_4_385 ();
 FILLCELL_X32 FILLER_4_417 ();
 FILLCELL_X32 FILLER_4_449 ();
 FILLCELL_X32 FILLER_4_481 ();
 FILLCELL_X32 FILLER_4_513 ();
 FILLCELL_X32 FILLER_4_545 ();
 FILLCELL_X32 FILLER_4_577 ();
 FILLCELL_X16 FILLER_4_609 ();
 FILLCELL_X4 FILLER_4_625 ();
 FILLCELL_X2 FILLER_4_629 ();
 FILLCELL_X32 FILLER_4_632 ();
 FILLCELL_X32 FILLER_4_664 ();
 FILLCELL_X32 FILLER_4_696 ();
 FILLCELL_X32 FILLER_4_728 ();
 FILLCELL_X32 FILLER_4_760 ();
 FILLCELL_X32 FILLER_4_792 ();
 FILLCELL_X32 FILLER_4_824 ();
 FILLCELL_X32 FILLER_4_856 ();
 FILLCELL_X32 FILLER_4_888 ();
 FILLCELL_X32 FILLER_4_920 ();
 FILLCELL_X32 FILLER_4_952 ();
 FILLCELL_X32 FILLER_4_984 ();
 FILLCELL_X32 FILLER_4_1016 ();
 FILLCELL_X32 FILLER_4_1048 ();
 FILLCELL_X32 FILLER_4_1080 ();
 FILLCELL_X32 FILLER_4_1112 ();
 FILLCELL_X32 FILLER_4_1144 ();
 FILLCELL_X32 FILLER_4_1176 ();
 FILLCELL_X32 FILLER_4_1208 ();
 FILLCELL_X32 FILLER_4_1240 ();
 FILLCELL_X32 FILLER_4_1272 ();
 FILLCELL_X32 FILLER_4_1304 ();
 FILLCELL_X32 FILLER_4_1336 ();
 FILLCELL_X32 FILLER_4_1368 ();
 FILLCELL_X32 FILLER_4_1400 ();
 FILLCELL_X32 FILLER_4_1432 ();
 FILLCELL_X32 FILLER_4_1464 ();
 FILLCELL_X32 FILLER_4_1496 ();
 FILLCELL_X32 FILLER_4_1528 ();
 FILLCELL_X32 FILLER_4_1560 ();
 FILLCELL_X32 FILLER_4_1592 ();
 FILLCELL_X32 FILLER_4_1624 ();
 FILLCELL_X32 FILLER_4_1656 ();
 FILLCELL_X32 FILLER_4_1688 ();
 FILLCELL_X32 FILLER_4_1720 ();
 FILLCELL_X32 FILLER_4_1752 ();
 FILLCELL_X32 FILLER_4_1784 ();
 FILLCELL_X32 FILLER_4_1816 ();
 FILLCELL_X32 FILLER_4_1848 ();
 FILLCELL_X8 FILLER_4_1880 ();
 FILLCELL_X4 FILLER_4_1888 ();
 FILLCELL_X2 FILLER_4_1892 ();
 FILLCELL_X32 FILLER_4_1895 ();
 FILLCELL_X32 FILLER_4_1927 ();
 FILLCELL_X32 FILLER_4_1959 ();
 FILLCELL_X32 FILLER_4_1991 ();
 FILLCELL_X32 FILLER_4_2023 ();
 FILLCELL_X32 FILLER_4_2055 ();
 FILLCELL_X32 FILLER_4_2087 ();
 FILLCELL_X32 FILLER_4_2119 ();
 FILLCELL_X32 FILLER_4_2151 ();
 FILLCELL_X32 FILLER_4_2183 ();
 FILLCELL_X32 FILLER_4_2215 ();
 FILLCELL_X32 FILLER_4_2247 ();
 FILLCELL_X32 FILLER_4_2279 ();
 FILLCELL_X32 FILLER_4_2311 ();
 FILLCELL_X32 FILLER_4_2343 ();
 FILLCELL_X32 FILLER_4_2375 ();
 FILLCELL_X32 FILLER_4_2407 ();
 FILLCELL_X32 FILLER_4_2439 ();
 FILLCELL_X32 FILLER_4_2471 ();
 FILLCELL_X32 FILLER_4_2503 ();
 FILLCELL_X32 FILLER_4_2535 ();
 FILLCELL_X32 FILLER_4_2567 ();
 FILLCELL_X32 FILLER_4_2599 ();
 FILLCELL_X32 FILLER_4_2631 ();
 FILLCELL_X32 FILLER_4_2663 ();
 FILLCELL_X32 FILLER_4_2695 ();
 FILLCELL_X32 FILLER_4_2727 ();
 FILLCELL_X32 FILLER_4_2759 ();
 FILLCELL_X32 FILLER_4_2791 ();
 FILLCELL_X32 FILLER_4_2823 ();
 FILLCELL_X32 FILLER_4_2855 ();
 FILLCELL_X32 FILLER_4_2887 ();
 FILLCELL_X32 FILLER_4_2919 ();
 FILLCELL_X32 FILLER_4_2951 ();
 FILLCELL_X32 FILLER_4_2983 ();
 FILLCELL_X32 FILLER_4_3015 ();
 FILLCELL_X32 FILLER_4_3047 ();
 FILLCELL_X32 FILLER_4_3079 ();
 FILLCELL_X32 FILLER_4_3111 ();
 FILLCELL_X8 FILLER_4_3143 ();
 FILLCELL_X4 FILLER_4_3151 ();
 FILLCELL_X2 FILLER_4_3155 ();
 FILLCELL_X32 FILLER_4_3158 ();
 FILLCELL_X32 FILLER_4_3190 ();
 FILLCELL_X32 FILLER_4_3222 ();
 FILLCELL_X32 FILLER_4_3254 ();
 FILLCELL_X32 FILLER_4_3286 ();
 FILLCELL_X32 FILLER_4_3318 ();
 FILLCELL_X32 FILLER_4_3350 ();
 FILLCELL_X32 FILLER_4_3382 ();
 FILLCELL_X32 FILLER_4_3414 ();
 FILLCELL_X32 FILLER_4_3446 ();
 FILLCELL_X32 FILLER_4_3478 ();
 FILLCELL_X32 FILLER_4_3510 ();
 FILLCELL_X32 FILLER_4_3542 ();
 FILLCELL_X32 FILLER_4_3574 ();
 FILLCELL_X32 FILLER_4_3606 ();
 FILLCELL_X32 FILLER_4_3638 ();
 FILLCELL_X32 FILLER_4_3670 ();
 FILLCELL_X32 FILLER_4_3702 ();
 FILLCELL_X4 FILLER_4_3734 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X32 FILLER_5_353 ();
 FILLCELL_X32 FILLER_5_385 ();
 FILLCELL_X32 FILLER_5_417 ();
 FILLCELL_X32 FILLER_5_449 ();
 FILLCELL_X32 FILLER_5_481 ();
 FILLCELL_X32 FILLER_5_513 ();
 FILLCELL_X32 FILLER_5_545 ();
 FILLCELL_X32 FILLER_5_577 ();
 FILLCELL_X32 FILLER_5_609 ();
 FILLCELL_X32 FILLER_5_641 ();
 FILLCELL_X32 FILLER_5_673 ();
 FILLCELL_X32 FILLER_5_705 ();
 FILLCELL_X32 FILLER_5_737 ();
 FILLCELL_X32 FILLER_5_769 ();
 FILLCELL_X32 FILLER_5_801 ();
 FILLCELL_X32 FILLER_5_833 ();
 FILLCELL_X32 FILLER_5_865 ();
 FILLCELL_X32 FILLER_5_897 ();
 FILLCELL_X32 FILLER_5_929 ();
 FILLCELL_X32 FILLER_5_961 ();
 FILLCELL_X32 FILLER_5_993 ();
 FILLCELL_X32 FILLER_5_1025 ();
 FILLCELL_X32 FILLER_5_1057 ();
 FILLCELL_X32 FILLER_5_1089 ();
 FILLCELL_X32 FILLER_5_1121 ();
 FILLCELL_X32 FILLER_5_1153 ();
 FILLCELL_X32 FILLER_5_1185 ();
 FILLCELL_X32 FILLER_5_1217 ();
 FILLCELL_X8 FILLER_5_1249 ();
 FILLCELL_X4 FILLER_5_1257 ();
 FILLCELL_X2 FILLER_5_1261 ();
 FILLCELL_X32 FILLER_5_1264 ();
 FILLCELL_X32 FILLER_5_1296 ();
 FILLCELL_X32 FILLER_5_1328 ();
 FILLCELL_X32 FILLER_5_1360 ();
 FILLCELL_X32 FILLER_5_1392 ();
 FILLCELL_X32 FILLER_5_1424 ();
 FILLCELL_X32 FILLER_5_1456 ();
 FILLCELL_X32 FILLER_5_1488 ();
 FILLCELL_X32 FILLER_5_1520 ();
 FILLCELL_X32 FILLER_5_1552 ();
 FILLCELL_X32 FILLER_5_1584 ();
 FILLCELL_X32 FILLER_5_1616 ();
 FILLCELL_X32 FILLER_5_1648 ();
 FILLCELL_X32 FILLER_5_1680 ();
 FILLCELL_X32 FILLER_5_1712 ();
 FILLCELL_X32 FILLER_5_1744 ();
 FILLCELL_X32 FILLER_5_1776 ();
 FILLCELL_X32 FILLER_5_1808 ();
 FILLCELL_X32 FILLER_5_1840 ();
 FILLCELL_X32 FILLER_5_1872 ();
 FILLCELL_X32 FILLER_5_1904 ();
 FILLCELL_X32 FILLER_5_1936 ();
 FILLCELL_X32 FILLER_5_1968 ();
 FILLCELL_X32 FILLER_5_2000 ();
 FILLCELL_X32 FILLER_5_2032 ();
 FILLCELL_X32 FILLER_5_2064 ();
 FILLCELL_X32 FILLER_5_2096 ();
 FILLCELL_X32 FILLER_5_2128 ();
 FILLCELL_X32 FILLER_5_2160 ();
 FILLCELL_X32 FILLER_5_2192 ();
 FILLCELL_X32 FILLER_5_2224 ();
 FILLCELL_X32 FILLER_5_2256 ();
 FILLCELL_X32 FILLER_5_2288 ();
 FILLCELL_X32 FILLER_5_2320 ();
 FILLCELL_X32 FILLER_5_2352 ();
 FILLCELL_X32 FILLER_5_2384 ();
 FILLCELL_X32 FILLER_5_2416 ();
 FILLCELL_X32 FILLER_5_2448 ();
 FILLCELL_X32 FILLER_5_2480 ();
 FILLCELL_X8 FILLER_5_2512 ();
 FILLCELL_X4 FILLER_5_2520 ();
 FILLCELL_X2 FILLER_5_2524 ();
 FILLCELL_X32 FILLER_5_2527 ();
 FILLCELL_X32 FILLER_5_2559 ();
 FILLCELL_X32 FILLER_5_2591 ();
 FILLCELL_X32 FILLER_5_2623 ();
 FILLCELL_X32 FILLER_5_2655 ();
 FILLCELL_X32 FILLER_5_2687 ();
 FILLCELL_X32 FILLER_5_2719 ();
 FILLCELL_X32 FILLER_5_2751 ();
 FILLCELL_X32 FILLER_5_2783 ();
 FILLCELL_X32 FILLER_5_2815 ();
 FILLCELL_X32 FILLER_5_2847 ();
 FILLCELL_X32 FILLER_5_2879 ();
 FILLCELL_X32 FILLER_5_2911 ();
 FILLCELL_X32 FILLER_5_2943 ();
 FILLCELL_X32 FILLER_5_2975 ();
 FILLCELL_X32 FILLER_5_3007 ();
 FILLCELL_X32 FILLER_5_3039 ();
 FILLCELL_X32 FILLER_5_3071 ();
 FILLCELL_X32 FILLER_5_3103 ();
 FILLCELL_X32 FILLER_5_3135 ();
 FILLCELL_X32 FILLER_5_3167 ();
 FILLCELL_X32 FILLER_5_3199 ();
 FILLCELL_X32 FILLER_5_3231 ();
 FILLCELL_X32 FILLER_5_3263 ();
 FILLCELL_X32 FILLER_5_3295 ();
 FILLCELL_X32 FILLER_5_3327 ();
 FILLCELL_X32 FILLER_5_3359 ();
 FILLCELL_X32 FILLER_5_3391 ();
 FILLCELL_X32 FILLER_5_3423 ();
 FILLCELL_X32 FILLER_5_3455 ();
 FILLCELL_X32 FILLER_5_3487 ();
 FILLCELL_X32 FILLER_5_3519 ();
 FILLCELL_X32 FILLER_5_3551 ();
 FILLCELL_X32 FILLER_5_3583 ();
 FILLCELL_X32 FILLER_5_3615 ();
 FILLCELL_X32 FILLER_5_3647 ();
 FILLCELL_X32 FILLER_5_3679 ();
 FILLCELL_X16 FILLER_5_3711 ();
 FILLCELL_X8 FILLER_5_3727 ();
 FILLCELL_X2 FILLER_5_3735 ();
 FILLCELL_X1 FILLER_5_3737 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X32 FILLER_6_321 ();
 FILLCELL_X32 FILLER_6_353 ();
 FILLCELL_X32 FILLER_6_385 ();
 FILLCELL_X32 FILLER_6_417 ();
 FILLCELL_X32 FILLER_6_449 ();
 FILLCELL_X32 FILLER_6_481 ();
 FILLCELL_X32 FILLER_6_513 ();
 FILLCELL_X32 FILLER_6_545 ();
 FILLCELL_X32 FILLER_6_577 ();
 FILLCELL_X16 FILLER_6_609 ();
 FILLCELL_X4 FILLER_6_625 ();
 FILLCELL_X2 FILLER_6_629 ();
 FILLCELL_X32 FILLER_6_632 ();
 FILLCELL_X32 FILLER_6_664 ();
 FILLCELL_X32 FILLER_6_696 ();
 FILLCELL_X32 FILLER_6_728 ();
 FILLCELL_X32 FILLER_6_760 ();
 FILLCELL_X32 FILLER_6_792 ();
 FILLCELL_X32 FILLER_6_824 ();
 FILLCELL_X32 FILLER_6_856 ();
 FILLCELL_X32 FILLER_6_888 ();
 FILLCELL_X32 FILLER_6_920 ();
 FILLCELL_X32 FILLER_6_952 ();
 FILLCELL_X32 FILLER_6_984 ();
 FILLCELL_X32 FILLER_6_1016 ();
 FILLCELL_X32 FILLER_6_1048 ();
 FILLCELL_X32 FILLER_6_1080 ();
 FILLCELL_X32 FILLER_6_1112 ();
 FILLCELL_X32 FILLER_6_1144 ();
 FILLCELL_X32 FILLER_6_1176 ();
 FILLCELL_X32 FILLER_6_1208 ();
 FILLCELL_X32 FILLER_6_1240 ();
 FILLCELL_X32 FILLER_6_1272 ();
 FILLCELL_X32 FILLER_6_1304 ();
 FILLCELL_X32 FILLER_6_1336 ();
 FILLCELL_X32 FILLER_6_1368 ();
 FILLCELL_X32 FILLER_6_1400 ();
 FILLCELL_X32 FILLER_6_1432 ();
 FILLCELL_X32 FILLER_6_1464 ();
 FILLCELL_X32 FILLER_6_1496 ();
 FILLCELL_X32 FILLER_6_1528 ();
 FILLCELL_X32 FILLER_6_1560 ();
 FILLCELL_X32 FILLER_6_1592 ();
 FILLCELL_X32 FILLER_6_1624 ();
 FILLCELL_X32 FILLER_6_1656 ();
 FILLCELL_X32 FILLER_6_1688 ();
 FILLCELL_X32 FILLER_6_1720 ();
 FILLCELL_X32 FILLER_6_1752 ();
 FILLCELL_X32 FILLER_6_1784 ();
 FILLCELL_X32 FILLER_6_1816 ();
 FILLCELL_X32 FILLER_6_1848 ();
 FILLCELL_X8 FILLER_6_1880 ();
 FILLCELL_X4 FILLER_6_1888 ();
 FILLCELL_X2 FILLER_6_1892 ();
 FILLCELL_X32 FILLER_6_1895 ();
 FILLCELL_X32 FILLER_6_1927 ();
 FILLCELL_X32 FILLER_6_1959 ();
 FILLCELL_X32 FILLER_6_1991 ();
 FILLCELL_X32 FILLER_6_2023 ();
 FILLCELL_X32 FILLER_6_2055 ();
 FILLCELL_X32 FILLER_6_2087 ();
 FILLCELL_X32 FILLER_6_2119 ();
 FILLCELL_X32 FILLER_6_2151 ();
 FILLCELL_X32 FILLER_6_2183 ();
 FILLCELL_X32 FILLER_6_2215 ();
 FILLCELL_X32 FILLER_6_2247 ();
 FILLCELL_X32 FILLER_6_2279 ();
 FILLCELL_X32 FILLER_6_2311 ();
 FILLCELL_X32 FILLER_6_2343 ();
 FILLCELL_X32 FILLER_6_2375 ();
 FILLCELL_X32 FILLER_6_2407 ();
 FILLCELL_X32 FILLER_6_2439 ();
 FILLCELL_X32 FILLER_6_2471 ();
 FILLCELL_X32 FILLER_6_2503 ();
 FILLCELL_X32 FILLER_6_2535 ();
 FILLCELL_X32 FILLER_6_2567 ();
 FILLCELL_X32 FILLER_6_2599 ();
 FILLCELL_X32 FILLER_6_2631 ();
 FILLCELL_X32 FILLER_6_2663 ();
 FILLCELL_X32 FILLER_6_2695 ();
 FILLCELL_X32 FILLER_6_2727 ();
 FILLCELL_X32 FILLER_6_2759 ();
 FILLCELL_X32 FILLER_6_2791 ();
 FILLCELL_X32 FILLER_6_2823 ();
 FILLCELL_X32 FILLER_6_2855 ();
 FILLCELL_X32 FILLER_6_2887 ();
 FILLCELL_X32 FILLER_6_2919 ();
 FILLCELL_X32 FILLER_6_2951 ();
 FILLCELL_X32 FILLER_6_2983 ();
 FILLCELL_X32 FILLER_6_3015 ();
 FILLCELL_X32 FILLER_6_3047 ();
 FILLCELL_X32 FILLER_6_3079 ();
 FILLCELL_X32 FILLER_6_3111 ();
 FILLCELL_X8 FILLER_6_3143 ();
 FILLCELL_X4 FILLER_6_3151 ();
 FILLCELL_X2 FILLER_6_3155 ();
 FILLCELL_X32 FILLER_6_3158 ();
 FILLCELL_X32 FILLER_6_3190 ();
 FILLCELL_X32 FILLER_6_3222 ();
 FILLCELL_X32 FILLER_6_3254 ();
 FILLCELL_X32 FILLER_6_3286 ();
 FILLCELL_X32 FILLER_6_3318 ();
 FILLCELL_X32 FILLER_6_3350 ();
 FILLCELL_X32 FILLER_6_3382 ();
 FILLCELL_X32 FILLER_6_3414 ();
 FILLCELL_X32 FILLER_6_3446 ();
 FILLCELL_X32 FILLER_6_3478 ();
 FILLCELL_X32 FILLER_6_3510 ();
 FILLCELL_X32 FILLER_6_3542 ();
 FILLCELL_X32 FILLER_6_3574 ();
 FILLCELL_X32 FILLER_6_3606 ();
 FILLCELL_X32 FILLER_6_3638 ();
 FILLCELL_X32 FILLER_6_3670 ();
 FILLCELL_X32 FILLER_6_3702 ();
 FILLCELL_X4 FILLER_6_3734 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X32 FILLER_7_321 ();
 FILLCELL_X32 FILLER_7_353 ();
 FILLCELL_X32 FILLER_7_385 ();
 FILLCELL_X32 FILLER_7_417 ();
 FILLCELL_X32 FILLER_7_449 ();
 FILLCELL_X32 FILLER_7_481 ();
 FILLCELL_X32 FILLER_7_513 ();
 FILLCELL_X32 FILLER_7_545 ();
 FILLCELL_X32 FILLER_7_577 ();
 FILLCELL_X32 FILLER_7_609 ();
 FILLCELL_X32 FILLER_7_641 ();
 FILLCELL_X32 FILLER_7_673 ();
 FILLCELL_X32 FILLER_7_705 ();
 FILLCELL_X32 FILLER_7_737 ();
 FILLCELL_X32 FILLER_7_769 ();
 FILLCELL_X32 FILLER_7_801 ();
 FILLCELL_X32 FILLER_7_833 ();
 FILLCELL_X32 FILLER_7_865 ();
 FILLCELL_X32 FILLER_7_897 ();
 FILLCELL_X32 FILLER_7_929 ();
 FILLCELL_X32 FILLER_7_961 ();
 FILLCELL_X32 FILLER_7_993 ();
 FILLCELL_X32 FILLER_7_1025 ();
 FILLCELL_X32 FILLER_7_1057 ();
 FILLCELL_X32 FILLER_7_1089 ();
 FILLCELL_X32 FILLER_7_1121 ();
 FILLCELL_X32 FILLER_7_1153 ();
 FILLCELL_X32 FILLER_7_1185 ();
 FILLCELL_X32 FILLER_7_1217 ();
 FILLCELL_X8 FILLER_7_1249 ();
 FILLCELL_X4 FILLER_7_1257 ();
 FILLCELL_X2 FILLER_7_1261 ();
 FILLCELL_X32 FILLER_7_1264 ();
 FILLCELL_X32 FILLER_7_1296 ();
 FILLCELL_X32 FILLER_7_1328 ();
 FILLCELL_X32 FILLER_7_1360 ();
 FILLCELL_X32 FILLER_7_1392 ();
 FILLCELL_X32 FILLER_7_1424 ();
 FILLCELL_X32 FILLER_7_1456 ();
 FILLCELL_X32 FILLER_7_1488 ();
 FILLCELL_X32 FILLER_7_1520 ();
 FILLCELL_X32 FILLER_7_1552 ();
 FILLCELL_X32 FILLER_7_1584 ();
 FILLCELL_X32 FILLER_7_1616 ();
 FILLCELL_X32 FILLER_7_1648 ();
 FILLCELL_X32 FILLER_7_1680 ();
 FILLCELL_X32 FILLER_7_1712 ();
 FILLCELL_X32 FILLER_7_1744 ();
 FILLCELL_X32 FILLER_7_1776 ();
 FILLCELL_X32 FILLER_7_1808 ();
 FILLCELL_X32 FILLER_7_1840 ();
 FILLCELL_X32 FILLER_7_1872 ();
 FILLCELL_X32 FILLER_7_1904 ();
 FILLCELL_X32 FILLER_7_1936 ();
 FILLCELL_X32 FILLER_7_1968 ();
 FILLCELL_X32 FILLER_7_2000 ();
 FILLCELL_X32 FILLER_7_2032 ();
 FILLCELL_X32 FILLER_7_2064 ();
 FILLCELL_X32 FILLER_7_2096 ();
 FILLCELL_X32 FILLER_7_2128 ();
 FILLCELL_X32 FILLER_7_2160 ();
 FILLCELL_X32 FILLER_7_2192 ();
 FILLCELL_X32 FILLER_7_2224 ();
 FILLCELL_X32 FILLER_7_2256 ();
 FILLCELL_X32 FILLER_7_2288 ();
 FILLCELL_X32 FILLER_7_2320 ();
 FILLCELL_X32 FILLER_7_2352 ();
 FILLCELL_X32 FILLER_7_2384 ();
 FILLCELL_X32 FILLER_7_2416 ();
 FILLCELL_X32 FILLER_7_2448 ();
 FILLCELL_X32 FILLER_7_2480 ();
 FILLCELL_X8 FILLER_7_2512 ();
 FILLCELL_X4 FILLER_7_2520 ();
 FILLCELL_X2 FILLER_7_2524 ();
 FILLCELL_X32 FILLER_7_2527 ();
 FILLCELL_X32 FILLER_7_2559 ();
 FILLCELL_X32 FILLER_7_2591 ();
 FILLCELL_X32 FILLER_7_2623 ();
 FILLCELL_X32 FILLER_7_2655 ();
 FILLCELL_X32 FILLER_7_2687 ();
 FILLCELL_X32 FILLER_7_2719 ();
 FILLCELL_X32 FILLER_7_2751 ();
 FILLCELL_X32 FILLER_7_2783 ();
 FILLCELL_X32 FILLER_7_2815 ();
 FILLCELL_X32 FILLER_7_2847 ();
 FILLCELL_X32 FILLER_7_2879 ();
 FILLCELL_X32 FILLER_7_2911 ();
 FILLCELL_X32 FILLER_7_2943 ();
 FILLCELL_X32 FILLER_7_2975 ();
 FILLCELL_X32 FILLER_7_3007 ();
 FILLCELL_X32 FILLER_7_3039 ();
 FILLCELL_X32 FILLER_7_3071 ();
 FILLCELL_X32 FILLER_7_3103 ();
 FILLCELL_X32 FILLER_7_3135 ();
 FILLCELL_X32 FILLER_7_3167 ();
 FILLCELL_X32 FILLER_7_3199 ();
 FILLCELL_X32 FILLER_7_3231 ();
 FILLCELL_X32 FILLER_7_3263 ();
 FILLCELL_X32 FILLER_7_3295 ();
 FILLCELL_X32 FILLER_7_3327 ();
 FILLCELL_X32 FILLER_7_3359 ();
 FILLCELL_X32 FILLER_7_3391 ();
 FILLCELL_X32 FILLER_7_3423 ();
 FILLCELL_X32 FILLER_7_3455 ();
 FILLCELL_X32 FILLER_7_3487 ();
 FILLCELL_X32 FILLER_7_3519 ();
 FILLCELL_X32 FILLER_7_3551 ();
 FILLCELL_X32 FILLER_7_3583 ();
 FILLCELL_X32 FILLER_7_3615 ();
 FILLCELL_X32 FILLER_7_3647 ();
 FILLCELL_X32 FILLER_7_3679 ();
 FILLCELL_X16 FILLER_7_3711 ();
 FILLCELL_X8 FILLER_7_3727 ();
 FILLCELL_X2 FILLER_7_3735 ();
 FILLCELL_X1 FILLER_7_3737 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X32 FILLER_8_321 ();
 FILLCELL_X32 FILLER_8_353 ();
 FILLCELL_X32 FILLER_8_385 ();
 FILLCELL_X32 FILLER_8_417 ();
 FILLCELL_X32 FILLER_8_449 ();
 FILLCELL_X32 FILLER_8_481 ();
 FILLCELL_X32 FILLER_8_513 ();
 FILLCELL_X32 FILLER_8_545 ();
 FILLCELL_X32 FILLER_8_577 ();
 FILLCELL_X16 FILLER_8_609 ();
 FILLCELL_X4 FILLER_8_625 ();
 FILLCELL_X2 FILLER_8_629 ();
 FILLCELL_X32 FILLER_8_632 ();
 FILLCELL_X32 FILLER_8_664 ();
 FILLCELL_X32 FILLER_8_696 ();
 FILLCELL_X32 FILLER_8_728 ();
 FILLCELL_X32 FILLER_8_760 ();
 FILLCELL_X32 FILLER_8_792 ();
 FILLCELL_X32 FILLER_8_824 ();
 FILLCELL_X32 FILLER_8_856 ();
 FILLCELL_X32 FILLER_8_888 ();
 FILLCELL_X32 FILLER_8_920 ();
 FILLCELL_X32 FILLER_8_952 ();
 FILLCELL_X32 FILLER_8_984 ();
 FILLCELL_X32 FILLER_8_1016 ();
 FILLCELL_X32 FILLER_8_1048 ();
 FILLCELL_X32 FILLER_8_1080 ();
 FILLCELL_X32 FILLER_8_1112 ();
 FILLCELL_X32 FILLER_8_1144 ();
 FILLCELL_X32 FILLER_8_1176 ();
 FILLCELL_X32 FILLER_8_1208 ();
 FILLCELL_X32 FILLER_8_1240 ();
 FILLCELL_X32 FILLER_8_1272 ();
 FILLCELL_X32 FILLER_8_1304 ();
 FILLCELL_X32 FILLER_8_1336 ();
 FILLCELL_X32 FILLER_8_1368 ();
 FILLCELL_X32 FILLER_8_1400 ();
 FILLCELL_X32 FILLER_8_1432 ();
 FILLCELL_X32 FILLER_8_1464 ();
 FILLCELL_X32 FILLER_8_1496 ();
 FILLCELL_X32 FILLER_8_1528 ();
 FILLCELL_X32 FILLER_8_1560 ();
 FILLCELL_X32 FILLER_8_1592 ();
 FILLCELL_X32 FILLER_8_1624 ();
 FILLCELL_X32 FILLER_8_1656 ();
 FILLCELL_X32 FILLER_8_1688 ();
 FILLCELL_X32 FILLER_8_1720 ();
 FILLCELL_X32 FILLER_8_1752 ();
 FILLCELL_X32 FILLER_8_1784 ();
 FILLCELL_X32 FILLER_8_1816 ();
 FILLCELL_X32 FILLER_8_1848 ();
 FILLCELL_X8 FILLER_8_1880 ();
 FILLCELL_X4 FILLER_8_1888 ();
 FILLCELL_X2 FILLER_8_1892 ();
 FILLCELL_X32 FILLER_8_1895 ();
 FILLCELL_X32 FILLER_8_1927 ();
 FILLCELL_X32 FILLER_8_1959 ();
 FILLCELL_X32 FILLER_8_1991 ();
 FILLCELL_X32 FILLER_8_2023 ();
 FILLCELL_X32 FILLER_8_2055 ();
 FILLCELL_X32 FILLER_8_2087 ();
 FILLCELL_X32 FILLER_8_2119 ();
 FILLCELL_X32 FILLER_8_2151 ();
 FILLCELL_X32 FILLER_8_2183 ();
 FILLCELL_X32 FILLER_8_2215 ();
 FILLCELL_X32 FILLER_8_2247 ();
 FILLCELL_X32 FILLER_8_2279 ();
 FILLCELL_X32 FILLER_8_2311 ();
 FILLCELL_X32 FILLER_8_2343 ();
 FILLCELL_X32 FILLER_8_2375 ();
 FILLCELL_X32 FILLER_8_2407 ();
 FILLCELL_X32 FILLER_8_2439 ();
 FILLCELL_X32 FILLER_8_2471 ();
 FILLCELL_X32 FILLER_8_2503 ();
 FILLCELL_X32 FILLER_8_2535 ();
 FILLCELL_X32 FILLER_8_2567 ();
 FILLCELL_X32 FILLER_8_2599 ();
 FILLCELL_X32 FILLER_8_2631 ();
 FILLCELL_X32 FILLER_8_2663 ();
 FILLCELL_X32 FILLER_8_2695 ();
 FILLCELL_X32 FILLER_8_2727 ();
 FILLCELL_X32 FILLER_8_2759 ();
 FILLCELL_X32 FILLER_8_2791 ();
 FILLCELL_X32 FILLER_8_2823 ();
 FILLCELL_X32 FILLER_8_2855 ();
 FILLCELL_X32 FILLER_8_2887 ();
 FILLCELL_X32 FILLER_8_2919 ();
 FILLCELL_X32 FILLER_8_2951 ();
 FILLCELL_X32 FILLER_8_2983 ();
 FILLCELL_X32 FILLER_8_3015 ();
 FILLCELL_X32 FILLER_8_3047 ();
 FILLCELL_X32 FILLER_8_3079 ();
 FILLCELL_X32 FILLER_8_3111 ();
 FILLCELL_X8 FILLER_8_3143 ();
 FILLCELL_X4 FILLER_8_3151 ();
 FILLCELL_X2 FILLER_8_3155 ();
 FILLCELL_X32 FILLER_8_3158 ();
 FILLCELL_X32 FILLER_8_3190 ();
 FILLCELL_X32 FILLER_8_3222 ();
 FILLCELL_X32 FILLER_8_3254 ();
 FILLCELL_X32 FILLER_8_3286 ();
 FILLCELL_X32 FILLER_8_3318 ();
 FILLCELL_X32 FILLER_8_3350 ();
 FILLCELL_X32 FILLER_8_3382 ();
 FILLCELL_X32 FILLER_8_3414 ();
 FILLCELL_X32 FILLER_8_3446 ();
 FILLCELL_X32 FILLER_8_3478 ();
 FILLCELL_X32 FILLER_8_3510 ();
 FILLCELL_X32 FILLER_8_3542 ();
 FILLCELL_X32 FILLER_8_3574 ();
 FILLCELL_X32 FILLER_8_3606 ();
 FILLCELL_X32 FILLER_8_3638 ();
 FILLCELL_X32 FILLER_8_3670 ();
 FILLCELL_X32 FILLER_8_3702 ();
 FILLCELL_X4 FILLER_8_3734 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X32 FILLER_9_353 ();
 FILLCELL_X32 FILLER_9_385 ();
 FILLCELL_X32 FILLER_9_417 ();
 FILLCELL_X32 FILLER_9_449 ();
 FILLCELL_X32 FILLER_9_481 ();
 FILLCELL_X32 FILLER_9_513 ();
 FILLCELL_X32 FILLER_9_545 ();
 FILLCELL_X32 FILLER_9_577 ();
 FILLCELL_X32 FILLER_9_609 ();
 FILLCELL_X32 FILLER_9_641 ();
 FILLCELL_X32 FILLER_9_673 ();
 FILLCELL_X32 FILLER_9_705 ();
 FILLCELL_X32 FILLER_9_737 ();
 FILLCELL_X32 FILLER_9_769 ();
 FILLCELL_X32 FILLER_9_801 ();
 FILLCELL_X32 FILLER_9_833 ();
 FILLCELL_X32 FILLER_9_865 ();
 FILLCELL_X32 FILLER_9_897 ();
 FILLCELL_X32 FILLER_9_929 ();
 FILLCELL_X32 FILLER_9_961 ();
 FILLCELL_X32 FILLER_9_993 ();
 FILLCELL_X32 FILLER_9_1025 ();
 FILLCELL_X32 FILLER_9_1057 ();
 FILLCELL_X32 FILLER_9_1089 ();
 FILLCELL_X32 FILLER_9_1121 ();
 FILLCELL_X32 FILLER_9_1153 ();
 FILLCELL_X32 FILLER_9_1185 ();
 FILLCELL_X32 FILLER_9_1217 ();
 FILLCELL_X8 FILLER_9_1249 ();
 FILLCELL_X4 FILLER_9_1257 ();
 FILLCELL_X2 FILLER_9_1261 ();
 FILLCELL_X32 FILLER_9_1264 ();
 FILLCELL_X32 FILLER_9_1296 ();
 FILLCELL_X32 FILLER_9_1328 ();
 FILLCELL_X32 FILLER_9_1360 ();
 FILLCELL_X32 FILLER_9_1392 ();
 FILLCELL_X32 FILLER_9_1424 ();
 FILLCELL_X32 FILLER_9_1456 ();
 FILLCELL_X32 FILLER_9_1488 ();
 FILLCELL_X32 FILLER_9_1520 ();
 FILLCELL_X32 FILLER_9_1552 ();
 FILLCELL_X32 FILLER_9_1584 ();
 FILLCELL_X32 FILLER_9_1616 ();
 FILLCELL_X32 FILLER_9_1648 ();
 FILLCELL_X32 FILLER_9_1680 ();
 FILLCELL_X32 FILLER_9_1712 ();
 FILLCELL_X32 FILLER_9_1744 ();
 FILLCELL_X32 FILLER_9_1776 ();
 FILLCELL_X32 FILLER_9_1808 ();
 FILLCELL_X32 FILLER_9_1840 ();
 FILLCELL_X32 FILLER_9_1872 ();
 FILLCELL_X32 FILLER_9_1904 ();
 FILLCELL_X32 FILLER_9_1936 ();
 FILLCELL_X32 FILLER_9_1968 ();
 FILLCELL_X32 FILLER_9_2000 ();
 FILLCELL_X32 FILLER_9_2032 ();
 FILLCELL_X32 FILLER_9_2064 ();
 FILLCELL_X32 FILLER_9_2096 ();
 FILLCELL_X32 FILLER_9_2128 ();
 FILLCELL_X32 FILLER_9_2160 ();
 FILLCELL_X32 FILLER_9_2192 ();
 FILLCELL_X32 FILLER_9_2224 ();
 FILLCELL_X32 FILLER_9_2256 ();
 FILLCELL_X32 FILLER_9_2288 ();
 FILLCELL_X32 FILLER_9_2320 ();
 FILLCELL_X32 FILLER_9_2352 ();
 FILLCELL_X32 FILLER_9_2384 ();
 FILLCELL_X32 FILLER_9_2416 ();
 FILLCELL_X32 FILLER_9_2448 ();
 FILLCELL_X32 FILLER_9_2480 ();
 FILLCELL_X8 FILLER_9_2512 ();
 FILLCELL_X4 FILLER_9_2520 ();
 FILLCELL_X2 FILLER_9_2524 ();
 FILLCELL_X32 FILLER_9_2527 ();
 FILLCELL_X32 FILLER_9_2559 ();
 FILLCELL_X32 FILLER_9_2591 ();
 FILLCELL_X32 FILLER_9_2623 ();
 FILLCELL_X32 FILLER_9_2655 ();
 FILLCELL_X32 FILLER_9_2687 ();
 FILLCELL_X32 FILLER_9_2719 ();
 FILLCELL_X32 FILLER_9_2751 ();
 FILLCELL_X32 FILLER_9_2783 ();
 FILLCELL_X32 FILLER_9_2815 ();
 FILLCELL_X32 FILLER_9_2847 ();
 FILLCELL_X32 FILLER_9_2879 ();
 FILLCELL_X32 FILLER_9_2911 ();
 FILLCELL_X32 FILLER_9_2943 ();
 FILLCELL_X32 FILLER_9_2975 ();
 FILLCELL_X32 FILLER_9_3007 ();
 FILLCELL_X32 FILLER_9_3039 ();
 FILLCELL_X32 FILLER_9_3071 ();
 FILLCELL_X32 FILLER_9_3103 ();
 FILLCELL_X32 FILLER_9_3135 ();
 FILLCELL_X32 FILLER_9_3167 ();
 FILLCELL_X32 FILLER_9_3199 ();
 FILLCELL_X32 FILLER_9_3231 ();
 FILLCELL_X32 FILLER_9_3263 ();
 FILLCELL_X32 FILLER_9_3295 ();
 FILLCELL_X32 FILLER_9_3327 ();
 FILLCELL_X32 FILLER_9_3359 ();
 FILLCELL_X32 FILLER_9_3391 ();
 FILLCELL_X32 FILLER_9_3423 ();
 FILLCELL_X32 FILLER_9_3455 ();
 FILLCELL_X32 FILLER_9_3487 ();
 FILLCELL_X32 FILLER_9_3519 ();
 FILLCELL_X32 FILLER_9_3551 ();
 FILLCELL_X32 FILLER_9_3583 ();
 FILLCELL_X32 FILLER_9_3615 ();
 FILLCELL_X32 FILLER_9_3647 ();
 FILLCELL_X32 FILLER_9_3679 ();
 FILLCELL_X16 FILLER_9_3711 ();
 FILLCELL_X8 FILLER_9_3727 ();
 FILLCELL_X2 FILLER_9_3735 ();
 FILLCELL_X1 FILLER_9_3737 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X32 FILLER_10_353 ();
 FILLCELL_X32 FILLER_10_385 ();
 FILLCELL_X32 FILLER_10_417 ();
 FILLCELL_X32 FILLER_10_449 ();
 FILLCELL_X32 FILLER_10_481 ();
 FILLCELL_X32 FILLER_10_513 ();
 FILLCELL_X32 FILLER_10_545 ();
 FILLCELL_X32 FILLER_10_577 ();
 FILLCELL_X16 FILLER_10_609 ();
 FILLCELL_X4 FILLER_10_625 ();
 FILLCELL_X2 FILLER_10_629 ();
 FILLCELL_X32 FILLER_10_632 ();
 FILLCELL_X32 FILLER_10_664 ();
 FILLCELL_X32 FILLER_10_696 ();
 FILLCELL_X32 FILLER_10_728 ();
 FILLCELL_X32 FILLER_10_760 ();
 FILLCELL_X32 FILLER_10_792 ();
 FILLCELL_X32 FILLER_10_824 ();
 FILLCELL_X32 FILLER_10_856 ();
 FILLCELL_X32 FILLER_10_888 ();
 FILLCELL_X32 FILLER_10_920 ();
 FILLCELL_X32 FILLER_10_952 ();
 FILLCELL_X32 FILLER_10_984 ();
 FILLCELL_X32 FILLER_10_1016 ();
 FILLCELL_X32 FILLER_10_1048 ();
 FILLCELL_X32 FILLER_10_1080 ();
 FILLCELL_X32 FILLER_10_1112 ();
 FILLCELL_X32 FILLER_10_1144 ();
 FILLCELL_X32 FILLER_10_1176 ();
 FILLCELL_X32 FILLER_10_1208 ();
 FILLCELL_X32 FILLER_10_1240 ();
 FILLCELL_X32 FILLER_10_1272 ();
 FILLCELL_X32 FILLER_10_1304 ();
 FILLCELL_X32 FILLER_10_1336 ();
 FILLCELL_X32 FILLER_10_1368 ();
 FILLCELL_X32 FILLER_10_1400 ();
 FILLCELL_X32 FILLER_10_1432 ();
 FILLCELL_X32 FILLER_10_1464 ();
 FILLCELL_X32 FILLER_10_1496 ();
 FILLCELL_X32 FILLER_10_1528 ();
 FILLCELL_X32 FILLER_10_1560 ();
 FILLCELL_X32 FILLER_10_1592 ();
 FILLCELL_X32 FILLER_10_1624 ();
 FILLCELL_X32 FILLER_10_1656 ();
 FILLCELL_X32 FILLER_10_1688 ();
 FILLCELL_X32 FILLER_10_1720 ();
 FILLCELL_X32 FILLER_10_1752 ();
 FILLCELL_X32 FILLER_10_1784 ();
 FILLCELL_X32 FILLER_10_1816 ();
 FILLCELL_X32 FILLER_10_1848 ();
 FILLCELL_X8 FILLER_10_1880 ();
 FILLCELL_X4 FILLER_10_1888 ();
 FILLCELL_X2 FILLER_10_1892 ();
 FILLCELL_X32 FILLER_10_1895 ();
 FILLCELL_X32 FILLER_10_1927 ();
 FILLCELL_X32 FILLER_10_1959 ();
 FILLCELL_X32 FILLER_10_1991 ();
 FILLCELL_X32 FILLER_10_2023 ();
 FILLCELL_X32 FILLER_10_2055 ();
 FILLCELL_X32 FILLER_10_2087 ();
 FILLCELL_X32 FILLER_10_2119 ();
 FILLCELL_X32 FILLER_10_2151 ();
 FILLCELL_X32 FILLER_10_2183 ();
 FILLCELL_X32 FILLER_10_2215 ();
 FILLCELL_X32 FILLER_10_2247 ();
 FILLCELL_X32 FILLER_10_2279 ();
 FILLCELL_X32 FILLER_10_2311 ();
 FILLCELL_X32 FILLER_10_2343 ();
 FILLCELL_X32 FILLER_10_2375 ();
 FILLCELL_X32 FILLER_10_2407 ();
 FILLCELL_X32 FILLER_10_2439 ();
 FILLCELL_X32 FILLER_10_2471 ();
 FILLCELL_X32 FILLER_10_2503 ();
 FILLCELL_X32 FILLER_10_2535 ();
 FILLCELL_X32 FILLER_10_2567 ();
 FILLCELL_X32 FILLER_10_2599 ();
 FILLCELL_X32 FILLER_10_2631 ();
 FILLCELL_X32 FILLER_10_2663 ();
 FILLCELL_X32 FILLER_10_2695 ();
 FILLCELL_X32 FILLER_10_2727 ();
 FILLCELL_X32 FILLER_10_2759 ();
 FILLCELL_X32 FILLER_10_2791 ();
 FILLCELL_X32 FILLER_10_2823 ();
 FILLCELL_X32 FILLER_10_2855 ();
 FILLCELL_X32 FILLER_10_2887 ();
 FILLCELL_X32 FILLER_10_2919 ();
 FILLCELL_X32 FILLER_10_2951 ();
 FILLCELL_X32 FILLER_10_2983 ();
 FILLCELL_X32 FILLER_10_3015 ();
 FILLCELL_X32 FILLER_10_3047 ();
 FILLCELL_X32 FILLER_10_3079 ();
 FILLCELL_X32 FILLER_10_3111 ();
 FILLCELL_X8 FILLER_10_3143 ();
 FILLCELL_X4 FILLER_10_3151 ();
 FILLCELL_X2 FILLER_10_3155 ();
 FILLCELL_X32 FILLER_10_3158 ();
 FILLCELL_X32 FILLER_10_3190 ();
 FILLCELL_X32 FILLER_10_3222 ();
 FILLCELL_X32 FILLER_10_3254 ();
 FILLCELL_X32 FILLER_10_3286 ();
 FILLCELL_X32 FILLER_10_3318 ();
 FILLCELL_X32 FILLER_10_3350 ();
 FILLCELL_X32 FILLER_10_3382 ();
 FILLCELL_X32 FILLER_10_3414 ();
 FILLCELL_X32 FILLER_10_3446 ();
 FILLCELL_X32 FILLER_10_3478 ();
 FILLCELL_X32 FILLER_10_3510 ();
 FILLCELL_X32 FILLER_10_3542 ();
 FILLCELL_X32 FILLER_10_3574 ();
 FILLCELL_X32 FILLER_10_3606 ();
 FILLCELL_X32 FILLER_10_3638 ();
 FILLCELL_X32 FILLER_10_3670 ();
 FILLCELL_X32 FILLER_10_3702 ();
 FILLCELL_X4 FILLER_10_3734 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X32 FILLER_11_321 ();
 FILLCELL_X32 FILLER_11_353 ();
 FILLCELL_X32 FILLER_11_385 ();
 FILLCELL_X32 FILLER_11_417 ();
 FILLCELL_X32 FILLER_11_449 ();
 FILLCELL_X32 FILLER_11_481 ();
 FILLCELL_X32 FILLER_11_513 ();
 FILLCELL_X32 FILLER_11_545 ();
 FILLCELL_X32 FILLER_11_577 ();
 FILLCELL_X32 FILLER_11_609 ();
 FILLCELL_X32 FILLER_11_641 ();
 FILLCELL_X32 FILLER_11_673 ();
 FILLCELL_X32 FILLER_11_705 ();
 FILLCELL_X32 FILLER_11_737 ();
 FILLCELL_X32 FILLER_11_769 ();
 FILLCELL_X32 FILLER_11_801 ();
 FILLCELL_X32 FILLER_11_833 ();
 FILLCELL_X32 FILLER_11_865 ();
 FILLCELL_X32 FILLER_11_897 ();
 FILLCELL_X32 FILLER_11_929 ();
 FILLCELL_X32 FILLER_11_961 ();
 FILLCELL_X32 FILLER_11_993 ();
 FILLCELL_X32 FILLER_11_1025 ();
 FILLCELL_X32 FILLER_11_1057 ();
 FILLCELL_X32 FILLER_11_1089 ();
 FILLCELL_X32 FILLER_11_1121 ();
 FILLCELL_X32 FILLER_11_1153 ();
 FILLCELL_X32 FILLER_11_1185 ();
 FILLCELL_X32 FILLER_11_1217 ();
 FILLCELL_X8 FILLER_11_1249 ();
 FILLCELL_X4 FILLER_11_1257 ();
 FILLCELL_X2 FILLER_11_1261 ();
 FILLCELL_X32 FILLER_11_1264 ();
 FILLCELL_X32 FILLER_11_1296 ();
 FILLCELL_X32 FILLER_11_1328 ();
 FILLCELL_X32 FILLER_11_1360 ();
 FILLCELL_X32 FILLER_11_1392 ();
 FILLCELL_X32 FILLER_11_1424 ();
 FILLCELL_X32 FILLER_11_1456 ();
 FILLCELL_X32 FILLER_11_1488 ();
 FILLCELL_X32 FILLER_11_1520 ();
 FILLCELL_X32 FILLER_11_1552 ();
 FILLCELL_X32 FILLER_11_1584 ();
 FILLCELL_X32 FILLER_11_1616 ();
 FILLCELL_X32 FILLER_11_1648 ();
 FILLCELL_X32 FILLER_11_1680 ();
 FILLCELL_X32 FILLER_11_1712 ();
 FILLCELL_X32 FILLER_11_1744 ();
 FILLCELL_X32 FILLER_11_1776 ();
 FILLCELL_X32 FILLER_11_1808 ();
 FILLCELL_X32 FILLER_11_1840 ();
 FILLCELL_X32 FILLER_11_1872 ();
 FILLCELL_X32 FILLER_11_1904 ();
 FILLCELL_X32 FILLER_11_1936 ();
 FILLCELL_X32 FILLER_11_1968 ();
 FILLCELL_X32 FILLER_11_2000 ();
 FILLCELL_X32 FILLER_11_2032 ();
 FILLCELL_X32 FILLER_11_2064 ();
 FILLCELL_X32 FILLER_11_2096 ();
 FILLCELL_X32 FILLER_11_2128 ();
 FILLCELL_X32 FILLER_11_2160 ();
 FILLCELL_X32 FILLER_11_2192 ();
 FILLCELL_X32 FILLER_11_2224 ();
 FILLCELL_X32 FILLER_11_2256 ();
 FILLCELL_X32 FILLER_11_2288 ();
 FILLCELL_X32 FILLER_11_2320 ();
 FILLCELL_X32 FILLER_11_2352 ();
 FILLCELL_X32 FILLER_11_2384 ();
 FILLCELL_X32 FILLER_11_2416 ();
 FILLCELL_X32 FILLER_11_2448 ();
 FILLCELL_X32 FILLER_11_2480 ();
 FILLCELL_X8 FILLER_11_2512 ();
 FILLCELL_X4 FILLER_11_2520 ();
 FILLCELL_X2 FILLER_11_2524 ();
 FILLCELL_X32 FILLER_11_2527 ();
 FILLCELL_X32 FILLER_11_2559 ();
 FILLCELL_X32 FILLER_11_2591 ();
 FILLCELL_X32 FILLER_11_2623 ();
 FILLCELL_X32 FILLER_11_2655 ();
 FILLCELL_X32 FILLER_11_2687 ();
 FILLCELL_X32 FILLER_11_2719 ();
 FILLCELL_X32 FILLER_11_2751 ();
 FILLCELL_X32 FILLER_11_2783 ();
 FILLCELL_X32 FILLER_11_2815 ();
 FILLCELL_X32 FILLER_11_2847 ();
 FILLCELL_X32 FILLER_11_2879 ();
 FILLCELL_X32 FILLER_11_2911 ();
 FILLCELL_X32 FILLER_11_2943 ();
 FILLCELL_X32 FILLER_11_2975 ();
 FILLCELL_X32 FILLER_11_3007 ();
 FILLCELL_X32 FILLER_11_3039 ();
 FILLCELL_X32 FILLER_11_3071 ();
 FILLCELL_X32 FILLER_11_3103 ();
 FILLCELL_X32 FILLER_11_3135 ();
 FILLCELL_X32 FILLER_11_3167 ();
 FILLCELL_X32 FILLER_11_3199 ();
 FILLCELL_X32 FILLER_11_3231 ();
 FILLCELL_X32 FILLER_11_3263 ();
 FILLCELL_X32 FILLER_11_3295 ();
 FILLCELL_X32 FILLER_11_3327 ();
 FILLCELL_X32 FILLER_11_3359 ();
 FILLCELL_X32 FILLER_11_3391 ();
 FILLCELL_X32 FILLER_11_3423 ();
 FILLCELL_X32 FILLER_11_3455 ();
 FILLCELL_X32 FILLER_11_3487 ();
 FILLCELL_X32 FILLER_11_3519 ();
 FILLCELL_X32 FILLER_11_3551 ();
 FILLCELL_X32 FILLER_11_3583 ();
 FILLCELL_X32 FILLER_11_3615 ();
 FILLCELL_X32 FILLER_11_3647 ();
 FILLCELL_X32 FILLER_11_3679 ();
 FILLCELL_X16 FILLER_11_3711 ();
 FILLCELL_X8 FILLER_11_3727 ();
 FILLCELL_X2 FILLER_11_3735 ();
 FILLCELL_X1 FILLER_11_3737 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X32 FILLER_12_321 ();
 FILLCELL_X32 FILLER_12_353 ();
 FILLCELL_X32 FILLER_12_385 ();
 FILLCELL_X32 FILLER_12_417 ();
 FILLCELL_X32 FILLER_12_449 ();
 FILLCELL_X32 FILLER_12_481 ();
 FILLCELL_X32 FILLER_12_513 ();
 FILLCELL_X32 FILLER_12_545 ();
 FILLCELL_X32 FILLER_12_577 ();
 FILLCELL_X16 FILLER_12_609 ();
 FILLCELL_X4 FILLER_12_625 ();
 FILLCELL_X2 FILLER_12_629 ();
 FILLCELL_X32 FILLER_12_632 ();
 FILLCELL_X32 FILLER_12_664 ();
 FILLCELL_X32 FILLER_12_696 ();
 FILLCELL_X32 FILLER_12_728 ();
 FILLCELL_X32 FILLER_12_760 ();
 FILLCELL_X32 FILLER_12_792 ();
 FILLCELL_X32 FILLER_12_824 ();
 FILLCELL_X32 FILLER_12_856 ();
 FILLCELL_X32 FILLER_12_888 ();
 FILLCELL_X32 FILLER_12_920 ();
 FILLCELL_X32 FILLER_12_952 ();
 FILLCELL_X32 FILLER_12_984 ();
 FILLCELL_X32 FILLER_12_1016 ();
 FILLCELL_X32 FILLER_12_1048 ();
 FILLCELL_X32 FILLER_12_1080 ();
 FILLCELL_X32 FILLER_12_1112 ();
 FILLCELL_X32 FILLER_12_1144 ();
 FILLCELL_X32 FILLER_12_1176 ();
 FILLCELL_X32 FILLER_12_1208 ();
 FILLCELL_X32 FILLER_12_1240 ();
 FILLCELL_X32 FILLER_12_1272 ();
 FILLCELL_X32 FILLER_12_1304 ();
 FILLCELL_X32 FILLER_12_1336 ();
 FILLCELL_X32 FILLER_12_1368 ();
 FILLCELL_X32 FILLER_12_1400 ();
 FILLCELL_X32 FILLER_12_1432 ();
 FILLCELL_X32 FILLER_12_1464 ();
 FILLCELL_X32 FILLER_12_1496 ();
 FILLCELL_X32 FILLER_12_1528 ();
 FILLCELL_X32 FILLER_12_1560 ();
 FILLCELL_X32 FILLER_12_1592 ();
 FILLCELL_X32 FILLER_12_1624 ();
 FILLCELL_X32 FILLER_12_1656 ();
 FILLCELL_X32 FILLER_12_1688 ();
 FILLCELL_X32 FILLER_12_1720 ();
 FILLCELL_X32 FILLER_12_1752 ();
 FILLCELL_X32 FILLER_12_1784 ();
 FILLCELL_X32 FILLER_12_1816 ();
 FILLCELL_X32 FILLER_12_1848 ();
 FILLCELL_X8 FILLER_12_1880 ();
 FILLCELL_X4 FILLER_12_1888 ();
 FILLCELL_X2 FILLER_12_1892 ();
 FILLCELL_X32 FILLER_12_1895 ();
 FILLCELL_X32 FILLER_12_1927 ();
 FILLCELL_X32 FILLER_12_1959 ();
 FILLCELL_X32 FILLER_12_1991 ();
 FILLCELL_X32 FILLER_12_2023 ();
 FILLCELL_X32 FILLER_12_2055 ();
 FILLCELL_X32 FILLER_12_2087 ();
 FILLCELL_X32 FILLER_12_2119 ();
 FILLCELL_X32 FILLER_12_2151 ();
 FILLCELL_X32 FILLER_12_2183 ();
 FILLCELL_X32 FILLER_12_2215 ();
 FILLCELL_X32 FILLER_12_2247 ();
 FILLCELL_X32 FILLER_12_2279 ();
 FILLCELL_X32 FILLER_12_2311 ();
 FILLCELL_X32 FILLER_12_2343 ();
 FILLCELL_X32 FILLER_12_2375 ();
 FILLCELL_X32 FILLER_12_2407 ();
 FILLCELL_X32 FILLER_12_2439 ();
 FILLCELL_X32 FILLER_12_2471 ();
 FILLCELL_X32 FILLER_12_2503 ();
 FILLCELL_X32 FILLER_12_2535 ();
 FILLCELL_X32 FILLER_12_2567 ();
 FILLCELL_X32 FILLER_12_2599 ();
 FILLCELL_X32 FILLER_12_2631 ();
 FILLCELL_X32 FILLER_12_2663 ();
 FILLCELL_X32 FILLER_12_2695 ();
 FILLCELL_X32 FILLER_12_2727 ();
 FILLCELL_X32 FILLER_12_2759 ();
 FILLCELL_X32 FILLER_12_2791 ();
 FILLCELL_X32 FILLER_12_2823 ();
 FILLCELL_X32 FILLER_12_2855 ();
 FILLCELL_X32 FILLER_12_2887 ();
 FILLCELL_X32 FILLER_12_2919 ();
 FILLCELL_X32 FILLER_12_2951 ();
 FILLCELL_X32 FILLER_12_2983 ();
 FILLCELL_X32 FILLER_12_3015 ();
 FILLCELL_X32 FILLER_12_3047 ();
 FILLCELL_X32 FILLER_12_3079 ();
 FILLCELL_X32 FILLER_12_3111 ();
 FILLCELL_X8 FILLER_12_3143 ();
 FILLCELL_X4 FILLER_12_3151 ();
 FILLCELL_X2 FILLER_12_3155 ();
 FILLCELL_X32 FILLER_12_3158 ();
 FILLCELL_X32 FILLER_12_3190 ();
 FILLCELL_X32 FILLER_12_3222 ();
 FILLCELL_X32 FILLER_12_3254 ();
 FILLCELL_X32 FILLER_12_3286 ();
 FILLCELL_X32 FILLER_12_3318 ();
 FILLCELL_X32 FILLER_12_3350 ();
 FILLCELL_X32 FILLER_12_3382 ();
 FILLCELL_X32 FILLER_12_3414 ();
 FILLCELL_X32 FILLER_12_3446 ();
 FILLCELL_X32 FILLER_12_3478 ();
 FILLCELL_X32 FILLER_12_3510 ();
 FILLCELL_X32 FILLER_12_3542 ();
 FILLCELL_X32 FILLER_12_3574 ();
 FILLCELL_X32 FILLER_12_3606 ();
 FILLCELL_X32 FILLER_12_3638 ();
 FILLCELL_X32 FILLER_12_3670 ();
 FILLCELL_X32 FILLER_12_3702 ();
 FILLCELL_X4 FILLER_12_3734 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X32 FILLER_13_321 ();
 FILLCELL_X32 FILLER_13_353 ();
 FILLCELL_X32 FILLER_13_385 ();
 FILLCELL_X32 FILLER_13_417 ();
 FILLCELL_X32 FILLER_13_449 ();
 FILLCELL_X32 FILLER_13_481 ();
 FILLCELL_X32 FILLER_13_513 ();
 FILLCELL_X32 FILLER_13_545 ();
 FILLCELL_X32 FILLER_13_577 ();
 FILLCELL_X32 FILLER_13_609 ();
 FILLCELL_X32 FILLER_13_641 ();
 FILLCELL_X32 FILLER_13_673 ();
 FILLCELL_X32 FILLER_13_705 ();
 FILLCELL_X32 FILLER_13_737 ();
 FILLCELL_X32 FILLER_13_769 ();
 FILLCELL_X32 FILLER_13_801 ();
 FILLCELL_X32 FILLER_13_833 ();
 FILLCELL_X32 FILLER_13_865 ();
 FILLCELL_X32 FILLER_13_897 ();
 FILLCELL_X32 FILLER_13_929 ();
 FILLCELL_X32 FILLER_13_961 ();
 FILLCELL_X32 FILLER_13_993 ();
 FILLCELL_X32 FILLER_13_1025 ();
 FILLCELL_X32 FILLER_13_1057 ();
 FILLCELL_X32 FILLER_13_1089 ();
 FILLCELL_X32 FILLER_13_1121 ();
 FILLCELL_X32 FILLER_13_1153 ();
 FILLCELL_X32 FILLER_13_1185 ();
 FILLCELL_X32 FILLER_13_1217 ();
 FILLCELL_X8 FILLER_13_1249 ();
 FILLCELL_X4 FILLER_13_1257 ();
 FILLCELL_X2 FILLER_13_1261 ();
 FILLCELL_X32 FILLER_13_1264 ();
 FILLCELL_X32 FILLER_13_1296 ();
 FILLCELL_X32 FILLER_13_1328 ();
 FILLCELL_X32 FILLER_13_1360 ();
 FILLCELL_X32 FILLER_13_1392 ();
 FILLCELL_X32 FILLER_13_1424 ();
 FILLCELL_X32 FILLER_13_1456 ();
 FILLCELL_X32 FILLER_13_1488 ();
 FILLCELL_X32 FILLER_13_1520 ();
 FILLCELL_X32 FILLER_13_1552 ();
 FILLCELL_X32 FILLER_13_1584 ();
 FILLCELL_X32 FILLER_13_1616 ();
 FILLCELL_X32 FILLER_13_1648 ();
 FILLCELL_X32 FILLER_13_1680 ();
 FILLCELL_X32 FILLER_13_1712 ();
 FILLCELL_X32 FILLER_13_1744 ();
 FILLCELL_X32 FILLER_13_1776 ();
 FILLCELL_X32 FILLER_13_1808 ();
 FILLCELL_X32 FILLER_13_1840 ();
 FILLCELL_X32 FILLER_13_1872 ();
 FILLCELL_X32 FILLER_13_1904 ();
 FILLCELL_X32 FILLER_13_1936 ();
 FILLCELL_X32 FILLER_13_1968 ();
 FILLCELL_X32 FILLER_13_2000 ();
 FILLCELL_X32 FILLER_13_2032 ();
 FILLCELL_X32 FILLER_13_2064 ();
 FILLCELL_X32 FILLER_13_2096 ();
 FILLCELL_X32 FILLER_13_2128 ();
 FILLCELL_X32 FILLER_13_2160 ();
 FILLCELL_X32 FILLER_13_2192 ();
 FILLCELL_X32 FILLER_13_2224 ();
 FILLCELL_X32 FILLER_13_2256 ();
 FILLCELL_X32 FILLER_13_2288 ();
 FILLCELL_X32 FILLER_13_2320 ();
 FILLCELL_X32 FILLER_13_2352 ();
 FILLCELL_X32 FILLER_13_2384 ();
 FILLCELL_X32 FILLER_13_2416 ();
 FILLCELL_X32 FILLER_13_2448 ();
 FILLCELL_X32 FILLER_13_2480 ();
 FILLCELL_X8 FILLER_13_2512 ();
 FILLCELL_X4 FILLER_13_2520 ();
 FILLCELL_X2 FILLER_13_2524 ();
 FILLCELL_X32 FILLER_13_2527 ();
 FILLCELL_X32 FILLER_13_2559 ();
 FILLCELL_X32 FILLER_13_2591 ();
 FILLCELL_X32 FILLER_13_2623 ();
 FILLCELL_X32 FILLER_13_2655 ();
 FILLCELL_X32 FILLER_13_2687 ();
 FILLCELL_X32 FILLER_13_2719 ();
 FILLCELL_X32 FILLER_13_2751 ();
 FILLCELL_X32 FILLER_13_2783 ();
 FILLCELL_X32 FILLER_13_2815 ();
 FILLCELL_X32 FILLER_13_2847 ();
 FILLCELL_X32 FILLER_13_2879 ();
 FILLCELL_X32 FILLER_13_2911 ();
 FILLCELL_X32 FILLER_13_2943 ();
 FILLCELL_X32 FILLER_13_2975 ();
 FILLCELL_X32 FILLER_13_3007 ();
 FILLCELL_X32 FILLER_13_3039 ();
 FILLCELL_X32 FILLER_13_3071 ();
 FILLCELL_X32 FILLER_13_3103 ();
 FILLCELL_X32 FILLER_13_3135 ();
 FILLCELL_X32 FILLER_13_3167 ();
 FILLCELL_X32 FILLER_13_3199 ();
 FILLCELL_X32 FILLER_13_3231 ();
 FILLCELL_X32 FILLER_13_3263 ();
 FILLCELL_X32 FILLER_13_3295 ();
 FILLCELL_X32 FILLER_13_3327 ();
 FILLCELL_X32 FILLER_13_3359 ();
 FILLCELL_X32 FILLER_13_3391 ();
 FILLCELL_X32 FILLER_13_3423 ();
 FILLCELL_X32 FILLER_13_3455 ();
 FILLCELL_X32 FILLER_13_3487 ();
 FILLCELL_X32 FILLER_13_3519 ();
 FILLCELL_X32 FILLER_13_3551 ();
 FILLCELL_X32 FILLER_13_3583 ();
 FILLCELL_X32 FILLER_13_3615 ();
 FILLCELL_X32 FILLER_13_3647 ();
 FILLCELL_X32 FILLER_13_3679 ();
 FILLCELL_X16 FILLER_13_3711 ();
 FILLCELL_X8 FILLER_13_3727 ();
 FILLCELL_X2 FILLER_13_3735 ();
 FILLCELL_X1 FILLER_13_3737 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X32 FILLER_14_321 ();
 FILLCELL_X32 FILLER_14_353 ();
 FILLCELL_X32 FILLER_14_385 ();
 FILLCELL_X32 FILLER_14_417 ();
 FILLCELL_X32 FILLER_14_449 ();
 FILLCELL_X32 FILLER_14_481 ();
 FILLCELL_X32 FILLER_14_513 ();
 FILLCELL_X32 FILLER_14_545 ();
 FILLCELL_X32 FILLER_14_577 ();
 FILLCELL_X16 FILLER_14_609 ();
 FILLCELL_X4 FILLER_14_625 ();
 FILLCELL_X2 FILLER_14_629 ();
 FILLCELL_X32 FILLER_14_632 ();
 FILLCELL_X32 FILLER_14_664 ();
 FILLCELL_X32 FILLER_14_696 ();
 FILLCELL_X32 FILLER_14_728 ();
 FILLCELL_X32 FILLER_14_760 ();
 FILLCELL_X32 FILLER_14_792 ();
 FILLCELL_X32 FILLER_14_824 ();
 FILLCELL_X32 FILLER_14_856 ();
 FILLCELL_X32 FILLER_14_888 ();
 FILLCELL_X32 FILLER_14_920 ();
 FILLCELL_X32 FILLER_14_952 ();
 FILLCELL_X32 FILLER_14_984 ();
 FILLCELL_X32 FILLER_14_1016 ();
 FILLCELL_X32 FILLER_14_1048 ();
 FILLCELL_X32 FILLER_14_1080 ();
 FILLCELL_X32 FILLER_14_1112 ();
 FILLCELL_X32 FILLER_14_1144 ();
 FILLCELL_X32 FILLER_14_1176 ();
 FILLCELL_X32 FILLER_14_1208 ();
 FILLCELL_X32 FILLER_14_1240 ();
 FILLCELL_X32 FILLER_14_1272 ();
 FILLCELL_X32 FILLER_14_1304 ();
 FILLCELL_X32 FILLER_14_1336 ();
 FILLCELL_X32 FILLER_14_1368 ();
 FILLCELL_X32 FILLER_14_1400 ();
 FILLCELL_X32 FILLER_14_1432 ();
 FILLCELL_X32 FILLER_14_1464 ();
 FILLCELL_X32 FILLER_14_1496 ();
 FILLCELL_X32 FILLER_14_1528 ();
 FILLCELL_X32 FILLER_14_1560 ();
 FILLCELL_X32 FILLER_14_1592 ();
 FILLCELL_X32 FILLER_14_1624 ();
 FILLCELL_X32 FILLER_14_1656 ();
 FILLCELL_X32 FILLER_14_1688 ();
 FILLCELL_X32 FILLER_14_1720 ();
 FILLCELL_X32 FILLER_14_1752 ();
 FILLCELL_X32 FILLER_14_1784 ();
 FILLCELL_X32 FILLER_14_1816 ();
 FILLCELL_X32 FILLER_14_1848 ();
 FILLCELL_X8 FILLER_14_1880 ();
 FILLCELL_X4 FILLER_14_1888 ();
 FILLCELL_X2 FILLER_14_1892 ();
 FILLCELL_X32 FILLER_14_1895 ();
 FILLCELL_X32 FILLER_14_1927 ();
 FILLCELL_X32 FILLER_14_1959 ();
 FILLCELL_X32 FILLER_14_1991 ();
 FILLCELL_X32 FILLER_14_2023 ();
 FILLCELL_X32 FILLER_14_2055 ();
 FILLCELL_X32 FILLER_14_2087 ();
 FILLCELL_X32 FILLER_14_2119 ();
 FILLCELL_X32 FILLER_14_2151 ();
 FILLCELL_X32 FILLER_14_2183 ();
 FILLCELL_X32 FILLER_14_2215 ();
 FILLCELL_X32 FILLER_14_2247 ();
 FILLCELL_X32 FILLER_14_2279 ();
 FILLCELL_X32 FILLER_14_2311 ();
 FILLCELL_X32 FILLER_14_2343 ();
 FILLCELL_X32 FILLER_14_2375 ();
 FILLCELL_X32 FILLER_14_2407 ();
 FILLCELL_X32 FILLER_14_2439 ();
 FILLCELL_X32 FILLER_14_2471 ();
 FILLCELL_X32 FILLER_14_2503 ();
 FILLCELL_X32 FILLER_14_2535 ();
 FILLCELL_X32 FILLER_14_2567 ();
 FILLCELL_X32 FILLER_14_2599 ();
 FILLCELL_X32 FILLER_14_2631 ();
 FILLCELL_X32 FILLER_14_2663 ();
 FILLCELL_X32 FILLER_14_2695 ();
 FILLCELL_X32 FILLER_14_2727 ();
 FILLCELL_X32 FILLER_14_2759 ();
 FILLCELL_X32 FILLER_14_2791 ();
 FILLCELL_X32 FILLER_14_2823 ();
 FILLCELL_X32 FILLER_14_2855 ();
 FILLCELL_X32 FILLER_14_2887 ();
 FILLCELL_X32 FILLER_14_2919 ();
 FILLCELL_X32 FILLER_14_2951 ();
 FILLCELL_X32 FILLER_14_2983 ();
 FILLCELL_X32 FILLER_14_3015 ();
 FILLCELL_X32 FILLER_14_3047 ();
 FILLCELL_X32 FILLER_14_3079 ();
 FILLCELL_X32 FILLER_14_3111 ();
 FILLCELL_X8 FILLER_14_3143 ();
 FILLCELL_X4 FILLER_14_3151 ();
 FILLCELL_X2 FILLER_14_3155 ();
 FILLCELL_X32 FILLER_14_3158 ();
 FILLCELL_X32 FILLER_14_3190 ();
 FILLCELL_X32 FILLER_14_3222 ();
 FILLCELL_X32 FILLER_14_3254 ();
 FILLCELL_X32 FILLER_14_3286 ();
 FILLCELL_X32 FILLER_14_3318 ();
 FILLCELL_X32 FILLER_14_3350 ();
 FILLCELL_X32 FILLER_14_3382 ();
 FILLCELL_X32 FILLER_14_3414 ();
 FILLCELL_X32 FILLER_14_3446 ();
 FILLCELL_X32 FILLER_14_3478 ();
 FILLCELL_X32 FILLER_14_3510 ();
 FILLCELL_X32 FILLER_14_3542 ();
 FILLCELL_X32 FILLER_14_3574 ();
 FILLCELL_X32 FILLER_14_3606 ();
 FILLCELL_X32 FILLER_14_3638 ();
 FILLCELL_X32 FILLER_14_3670 ();
 FILLCELL_X32 FILLER_14_3702 ();
 FILLCELL_X4 FILLER_14_3734 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X32 FILLER_15_289 ();
 FILLCELL_X32 FILLER_15_321 ();
 FILLCELL_X32 FILLER_15_353 ();
 FILLCELL_X32 FILLER_15_385 ();
 FILLCELL_X32 FILLER_15_417 ();
 FILLCELL_X32 FILLER_15_449 ();
 FILLCELL_X32 FILLER_15_481 ();
 FILLCELL_X32 FILLER_15_513 ();
 FILLCELL_X32 FILLER_15_545 ();
 FILLCELL_X32 FILLER_15_577 ();
 FILLCELL_X32 FILLER_15_609 ();
 FILLCELL_X32 FILLER_15_641 ();
 FILLCELL_X32 FILLER_15_673 ();
 FILLCELL_X32 FILLER_15_705 ();
 FILLCELL_X32 FILLER_15_737 ();
 FILLCELL_X32 FILLER_15_769 ();
 FILLCELL_X32 FILLER_15_801 ();
 FILLCELL_X32 FILLER_15_833 ();
 FILLCELL_X32 FILLER_15_865 ();
 FILLCELL_X32 FILLER_15_897 ();
 FILLCELL_X32 FILLER_15_929 ();
 FILLCELL_X32 FILLER_15_961 ();
 FILLCELL_X32 FILLER_15_993 ();
 FILLCELL_X32 FILLER_15_1025 ();
 FILLCELL_X32 FILLER_15_1057 ();
 FILLCELL_X32 FILLER_15_1089 ();
 FILLCELL_X32 FILLER_15_1121 ();
 FILLCELL_X32 FILLER_15_1153 ();
 FILLCELL_X32 FILLER_15_1185 ();
 FILLCELL_X32 FILLER_15_1217 ();
 FILLCELL_X8 FILLER_15_1249 ();
 FILLCELL_X4 FILLER_15_1257 ();
 FILLCELL_X2 FILLER_15_1261 ();
 FILLCELL_X32 FILLER_15_1264 ();
 FILLCELL_X32 FILLER_15_1296 ();
 FILLCELL_X32 FILLER_15_1328 ();
 FILLCELL_X32 FILLER_15_1360 ();
 FILLCELL_X32 FILLER_15_1392 ();
 FILLCELL_X32 FILLER_15_1424 ();
 FILLCELL_X32 FILLER_15_1456 ();
 FILLCELL_X32 FILLER_15_1488 ();
 FILLCELL_X32 FILLER_15_1520 ();
 FILLCELL_X32 FILLER_15_1552 ();
 FILLCELL_X32 FILLER_15_1584 ();
 FILLCELL_X32 FILLER_15_1616 ();
 FILLCELL_X32 FILLER_15_1648 ();
 FILLCELL_X32 FILLER_15_1680 ();
 FILLCELL_X32 FILLER_15_1712 ();
 FILLCELL_X32 FILLER_15_1744 ();
 FILLCELL_X32 FILLER_15_1776 ();
 FILLCELL_X32 FILLER_15_1808 ();
 FILLCELL_X32 FILLER_15_1840 ();
 FILLCELL_X32 FILLER_15_1872 ();
 FILLCELL_X32 FILLER_15_1904 ();
 FILLCELL_X32 FILLER_15_1936 ();
 FILLCELL_X32 FILLER_15_1968 ();
 FILLCELL_X32 FILLER_15_2000 ();
 FILLCELL_X32 FILLER_15_2032 ();
 FILLCELL_X32 FILLER_15_2064 ();
 FILLCELL_X32 FILLER_15_2096 ();
 FILLCELL_X32 FILLER_15_2128 ();
 FILLCELL_X32 FILLER_15_2160 ();
 FILLCELL_X32 FILLER_15_2192 ();
 FILLCELL_X32 FILLER_15_2224 ();
 FILLCELL_X32 FILLER_15_2256 ();
 FILLCELL_X32 FILLER_15_2288 ();
 FILLCELL_X32 FILLER_15_2320 ();
 FILLCELL_X32 FILLER_15_2352 ();
 FILLCELL_X32 FILLER_15_2384 ();
 FILLCELL_X32 FILLER_15_2416 ();
 FILLCELL_X32 FILLER_15_2448 ();
 FILLCELL_X32 FILLER_15_2480 ();
 FILLCELL_X8 FILLER_15_2512 ();
 FILLCELL_X4 FILLER_15_2520 ();
 FILLCELL_X2 FILLER_15_2524 ();
 FILLCELL_X32 FILLER_15_2527 ();
 FILLCELL_X32 FILLER_15_2559 ();
 FILLCELL_X32 FILLER_15_2591 ();
 FILLCELL_X32 FILLER_15_2623 ();
 FILLCELL_X32 FILLER_15_2655 ();
 FILLCELL_X32 FILLER_15_2687 ();
 FILLCELL_X32 FILLER_15_2719 ();
 FILLCELL_X32 FILLER_15_2751 ();
 FILLCELL_X32 FILLER_15_2783 ();
 FILLCELL_X32 FILLER_15_2815 ();
 FILLCELL_X32 FILLER_15_2847 ();
 FILLCELL_X32 FILLER_15_2879 ();
 FILLCELL_X32 FILLER_15_2911 ();
 FILLCELL_X32 FILLER_15_2943 ();
 FILLCELL_X32 FILLER_15_2975 ();
 FILLCELL_X32 FILLER_15_3007 ();
 FILLCELL_X32 FILLER_15_3039 ();
 FILLCELL_X32 FILLER_15_3071 ();
 FILLCELL_X32 FILLER_15_3103 ();
 FILLCELL_X32 FILLER_15_3135 ();
 FILLCELL_X32 FILLER_15_3167 ();
 FILLCELL_X32 FILLER_15_3199 ();
 FILLCELL_X32 FILLER_15_3231 ();
 FILLCELL_X32 FILLER_15_3263 ();
 FILLCELL_X32 FILLER_15_3295 ();
 FILLCELL_X32 FILLER_15_3327 ();
 FILLCELL_X32 FILLER_15_3359 ();
 FILLCELL_X32 FILLER_15_3391 ();
 FILLCELL_X32 FILLER_15_3423 ();
 FILLCELL_X32 FILLER_15_3455 ();
 FILLCELL_X32 FILLER_15_3487 ();
 FILLCELL_X32 FILLER_15_3519 ();
 FILLCELL_X32 FILLER_15_3551 ();
 FILLCELL_X32 FILLER_15_3583 ();
 FILLCELL_X32 FILLER_15_3615 ();
 FILLCELL_X32 FILLER_15_3647 ();
 FILLCELL_X32 FILLER_15_3679 ();
 FILLCELL_X16 FILLER_15_3711 ();
 FILLCELL_X8 FILLER_15_3727 ();
 FILLCELL_X2 FILLER_15_3735 ();
 FILLCELL_X1 FILLER_15_3737 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X32 FILLER_16_289 ();
 FILLCELL_X32 FILLER_16_321 ();
 FILLCELL_X32 FILLER_16_353 ();
 FILLCELL_X32 FILLER_16_385 ();
 FILLCELL_X32 FILLER_16_417 ();
 FILLCELL_X32 FILLER_16_449 ();
 FILLCELL_X32 FILLER_16_481 ();
 FILLCELL_X32 FILLER_16_513 ();
 FILLCELL_X32 FILLER_16_545 ();
 FILLCELL_X32 FILLER_16_577 ();
 FILLCELL_X16 FILLER_16_609 ();
 FILLCELL_X4 FILLER_16_625 ();
 FILLCELL_X2 FILLER_16_629 ();
 FILLCELL_X32 FILLER_16_632 ();
 FILLCELL_X32 FILLER_16_664 ();
 FILLCELL_X32 FILLER_16_696 ();
 FILLCELL_X32 FILLER_16_728 ();
 FILLCELL_X32 FILLER_16_760 ();
 FILLCELL_X32 FILLER_16_792 ();
 FILLCELL_X32 FILLER_16_824 ();
 FILLCELL_X32 FILLER_16_856 ();
 FILLCELL_X32 FILLER_16_888 ();
 FILLCELL_X32 FILLER_16_920 ();
 FILLCELL_X32 FILLER_16_952 ();
 FILLCELL_X32 FILLER_16_984 ();
 FILLCELL_X32 FILLER_16_1016 ();
 FILLCELL_X32 FILLER_16_1048 ();
 FILLCELL_X32 FILLER_16_1080 ();
 FILLCELL_X32 FILLER_16_1112 ();
 FILLCELL_X32 FILLER_16_1144 ();
 FILLCELL_X32 FILLER_16_1176 ();
 FILLCELL_X32 FILLER_16_1208 ();
 FILLCELL_X32 FILLER_16_1240 ();
 FILLCELL_X32 FILLER_16_1272 ();
 FILLCELL_X32 FILLER_16_1304 ();
 FILLCELL_X32 FILLER_16_1336 ();
 FILLCELL_X32 FILLER_16_1368 ();
 FILLCELL_X32 FILLER_16_1400 ();
 FILLCELL_X32 FILLER_16_1432 ();
 FILLCELL_X32 FILLER_16_1464 ();
 FILLCELL_X32 FILLER_16_1496 ();
 FILLCELL_X32 FILLER_16_1528 ();
 FILLCELL_X32 FILLER_16_1560 ();
 FILLCELL_X32 FILLER_16_1592 ();
 FILLCELL_X32 FILLER_16_1624 ();
 FILLCELL_X32 FILLER_16_1656 ();
 FILLCELL_X32 FILLER_16_1688 ();
 FILLCELL_X32 FILLER_16_1720 ();
 FILLCELL_X32 FILLER_16_1752 ();
 FILLCELL_X32 FILLER_16_1784 ();
 FILLCELL_X32 FILLER_16_1816 ();
 FILLCELL_X32 FILLER_16_1848 ();
 FILLCELL_X8 FILLER_16_1880 ();
 FILLCELL_X4 FILLER_16_1888 ();
 FILLCELL_X2 FILLER_16_1892 ();
 FILLCELL_X32 FILLER_16_1895 ();
 FILLCELL_X32 FILLER_16_1927 ();
 FILLCELL_X32 FILLER_16_1959 ();
 FILLCELL_X32 FILLER_16_1991 ();
 FILLCELL_X32 FILLER_16_2023 ();
 FILLCELL_X32 FILLER_16_2055 ();
 FILLCELL_X32 FILLER_16_2087 ();
 FILLCELL_X32 FILLER_16_2119 ();
 FILLCELL_X32 FILLER_16_2151 ();
 FILLCELL_X32 FILLER_16_2183 ();
 FILLCELL_X32 FILLER_16_2215 ();
 FILLCELL_X32 FILLER_16_2247 ();
 FILLCELL_X32 FILLER_16_2279 ();
 FILLCELL_X32 FILLER_16_2311 ();
 FILLCELL_X32 FILLER_16_2343 ();
 FILLCELL_X32 FILLER_16_2375 ();
 FILLCELL_X32 FILLER_16_2407 ();
 FILLCELL_X32 FILLER_16_2439 ();
 FILLCELL_X32 FILLER_16_2471 ();
 FILLCELL_X32 FILLER_16_2503 ();
 FILLCELL_X32 FILLER_16_2535 ();
 FILLCELL_X32 FILLER_16_2567 ();
 FILLCELL_X32 FILLER_16_2599 ();
 FILLCELL_X32 FILLER_16_2631 ();
 FILLCELL_X32 FILLER_16_2663 ();
 FILLCELL_X32 FILLER_16_2695 ();
 FILLCELL_X32 FILLER_16_2727 ();
 FILLCELL_X32 FILLER_16_2759 ();
 FILLCELL_X32 FILLER_16_2791 ();
 FILLCELL_X32 FILLER_16_2823 ();
 FILLCELL_X32 FILLER_16_2855 ();
 FILLCELL_X32 FILLER_16_2887 ();
 FILLCELL_X32 FILLER_16_2919 ();
 FILLCELL_X32 FILLER_16_2951 ();
 FILLCELL_X32 FILLER_16_2983 ();
 FILLCELL_X32 FILLER_16_3015 ();
 FILLCELL_X32 FILLER_16_3047 ();
 FILLCELL_X32 FILLER_16_3079 ();
 FILLCELL_X32 FILLER_16_3111 ();
 FILLCELL_X8 FILLER_16_3143 ();
 FILLCELL_X4 FILLER_16_3151 ();
 FILLCELL_X2 FILLER_16_3155 ();
 FILLCELL_X32 FILLER_16_3158 ();
 FILLCELL_X32 FILLER_16_3190 ();
 FILLCELL_X32 FILLER_16_3222 ();
 FILLCELL_X32 FILLER_16_3254 ();
 FILLCELL_X32 FILLER_16_3286 ();
 FILLCELL_X32 FILLER_16_3318 ();
 FILLCELL_X32 FILLER_16_3350 ();
 FILLCELL_X32 FILLER_16_3382 ();
 FILLCELL_X32 FILLER_16_3414 ();
 FILLCELL_X32 FILLER_16_3446 ();
 FILLCELL_X32 FILLER_16_3478 ();
 FILLCELL_X32 FILLER_16_3510 ();
 FILLCELL_X32 FILLER_16_3542 ();
 FILLCELL_X32 FILLER_16_3574 ();
 FILLCELL_X32 FILLER_16_3606 ();
 FILLCELL_X32 FILLER_16_3638 ();
 FILLCELL_X32 FILLER_16_3670 ();
 FILLCELL_X32 FILLER_16_3702 ();
 FILLCELL_X4 FILLER_16_3734 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X32 FILLER_17_289 ();
 FILLCELL_X32 FILLER_17_321 ();
 FILLCELL_X32 FILLER_17_353 ();
 FILLCELL_X32 FILLER_17_385 ();
 FILLCELL_X32 FILLER_17_417 ();
 FILLCELL_X32 FILLER_17_449 ();
 FILLCELL_X32 FILLER_17_481 ();
 FILLCELL_X32 FILLER_17_513 ();
 FILLCELL_X32 FILLER_17_545 ();
 FILLCELL_X32 FILLER_17_577 ();
 FILLCELL_X32 FILLER_17_609 ();
 FILLCELL_X32 FILLER_17_641 ();
 FILLCELL_X32 FILLER_17_673 ();
 FILLCELL_X32 FILLER_17_705 ();
 FILLCELL_X32 FILLER_17_737 ();
 FILLCELL_X32 FILLER_17_769 ();
 FILLCELL_X32 FILLER_17_801 ();
 FILLCELL_X32 FILLER_17_833 ();
 FILLCELL_X32 FILLER_17_865 ();
 FILLCELL_X32 FILLER_17_897 ();
 FILLCELL_X32 FILLER_17_929 ();
 FILLCELL_X32 FILLER_17_961 ();
 FILLCELL_X32 FILLER_17_993 ();
 FILLCELL_X32 FILLER_17_1025 ();
 FILLCELL_X32 FILLER_17_1057 ();
 FILLCELL_X32 FILLER_17_1089 ();
 FILLCELL_X32 FILLER_17_1121 ();
 FILLCELL_X32 FILLER_17_1153 ();
 FILLCELL_X32 FILLER_17_1185 ();
 FILLCELL_X32 FILLER_17_1217 ();
 FILLCELL_X8 FILLER_17_1249 ();
 FILLCELL_X4 FILLER_17_1257 ();
 FILLCELL_X2 FILLER_17_1261 ();
 FILLCELL_X32 FILLER_17_1264 ();
 FILLCELL_X32 FILLER_17_1296 ();
 FILLCELL_X32 FILLER_17_1328 ();
 FILLCELL_X32 FILLER_17_1360 ();
 FILLCELL_X32 FILLER_17_1392 ();
 FILLCELL_X32 FILLER_17_1424 ();
 FILLCELL_X32 FILLER_17_1456 ();
 FILLCELL_X32 FILLER_17_1488 ();
 FILLCELL_X32 FILLER_17_1520 ();
 FILLCELL_X32 FILLER_17_1552 ();
 FILLCELL_X32 FILLER_17_1584 ();
 FILLCELL_X32 FILLER_17_1616 ();
 FILLCELL_X32 FILLER_17_1648 ();
 FILLCELL_X32 FILLER_17_1680 ();
 FILLCELL_X32 FILLER_17_1712 ();
 FILLCELL_X32 FILLER_17_1744 ();
 FILLCELL_X32 FILLER_17_1776 ();
 FILLCELL_X32 FILLER_17_1808 ();
 FILLCELL_X32 FILLER_17_1840 ();
 FILLCELL_X32 FILLER_17_1872 ();
 FILLCELL_X32 FILLER_17_1904 ();
 FILLCELL_X32 FILLER_17_1936 ();
 FILLCELL_X32 FILLER_17_1968 ();
 FILLCELL_X32 FILLER_17_2000 ();
 FILLCELL_X32 FILLER_17_2032 ();
 FILLCELL_X32 FILLER_17_2064 ();
 FILLCELL_X32 FILLER_17_2096 ();
 FILLCELL_X32 FILLER_17_2128 ();
 FILLCELL_X32 FILLER_17_2160 ();
 FILLCELL_X32 FILLER_17_2192 ();
 FILLCELL_X32 FILLER_17_2224 ();
 FILLCELL_X32 FILLER_17_2256 ();
 FILLCELL_X32 FILLER_17_2288 ();
 FILLCELL_X32 FILLER_17_2320 ();
 FILLCELL_X32 FILLER_17_2352 ();
 FILLCELL_X32 FILLER_17_2384 ();
 FILLCELL_X32 FILLER_17_2416 ();
 FILLCELL_X32 FILLER_17_2448 ();
 FILLCELL_X32 FILLER_17_2480 ();
 FILLCELL_X8 FILLER_17_2512 ();
 FILLCELL_X4 FILLER_17_2520 ();
 FILLCELL_X2 FILLER_17_2524 ();
 FILLCELL_X32 FILLER_17_2527 ();
 FILLCELL_X32 FILLER_17_2559 ();
 FILLCELL_X32 FILLER_17_2591 ();
 FILLCELL_X32 FILLER_17_2623 ();
 FILLCELL_X32 FILLER_17_2655 ();
 FILLCELL_X32 FILLER_17_2687 ();
 FILLCELL_X32 FILLER_17_2719 ();
 FILLCELL_X32 FILLER_17_2751 ();
 FILLCELL_X32 FILLER_17_2783 ();
 FILLCELL_X32 FILLER_17_2815 ();
 FILLCELL_X32 FILLER_17_2847 ();
 FILLCELL_X32 FILLER_17_2879 ();
 FILLCELL_X32 FILLER_17_2911 ();
 FILLCELL_X32 FILLER_17_2943 ();
 FILLCELL_X32 FILLER_17_2975 ();
 FILLCELL_X32 FILLER_17_3007 ();
 FILLCELL_X32 FILLER_17_3039 ();
 FILLCELL_X32 FILLER_17_3071 ();
 FILLCELL_X32 FILLER_17_3103 ();
 FILLCELL_X32 FILLER_17_3135 ();
 FILLCELL_X32 FILLER_17_3167 ();
 FILLCELL_X32 FILLER_17_3199 ();
 FILLCELL_X32 FILLER_17_3231 ();
 FILLCELL_X32 FILLER_17_3263 ();
 FILLCELL_X32 FILLER_17_3295 ();
 FILLCELL_X32 FILLER_17_3327 ();
 FILLCELL_X32 FILLER_17_3359 ();
 FILLCELL_X32 FILLER_17_3391 ();
 FILLCELL_X32 FILLER_17_3423 ();
 FILLCELL_X32 FILLER_17_3455 ();
 FILLCELL_X32 FILLER_17_3487 ();
 FILLCELL_X32 FILLER_17_3519 ();
 FILLCELL_X32 FILLER_17_3551 ();
 FILLCELL_X32 FILLER_17_3583 ();
 FILLCELL_X32 FILLER_17_3615 ();
 FILLCELL_X32 FILLER_17_3647 ();
 FILLCELL_X32 FILLER_17_3679 ();
 FILLCELL_X16 FILLER_17_3711 ();
 FILLCELL_X8 FILLER_17_3727 ();
 FILLCELL_X2 FILLER_17_3735 ();
 FILLCELL_X1 FILLER_17_3737 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_289 ();
 FILLCELL_X32 FILLER_18_321 ();
 FILLCELL_X32 FILLER_18_353 ();
 FILLCELL_X32 FILLER_18_385 ();
 FILLCELL_X32 FILLER_18_417 ();
 FILLCELL_X32 FILLER_18_449 ();
 FILLCELL_X32 FILLER_18_481 ();
 FILLCELL_X32 FILLER_18_513 ();
 FILLCELL_X32 FILLER_18_545 ();
 FILLCELL_X32 FILLER_18_577 ();
 FILLCELL_X16 FILLER_18_609 ();
 FILLCELL_X4 FILLER_18_625 ();
 FILLCELL_X2 FILLER_18_629 ();
 FILLCELL_X32 FILLER_18_632 ();
 FILLCELL_X32 FILLER_18_664 ();
 FILLCELL_X32 FILLER_18_696 ();
 FILLCELL_X32 FILLER_18_728 ();
 FILLCELL_X32 FILLER_18_760 ();
 FILLCELL_X32 FILLER_18_792 ();
 FILLCELL_X32 FILLER_18_824 ();
 FILLCELL_X32 FILLER_18_856 ();
 FILLCELL_X32 FILLER_18_888 ();
 FILLCELL_X32 FILLER_18_920 ();
 FILLCELL_X32 FILLER_18_952 ();
 FILLCELL_X32 FILLER_18_984 ();
 FILLCELL_X32 FILLER_18_1016 ();
 FILLCELL_X32 FILLER_18_1048 ();
 FILLCELL_X32 FILLER_18_1080 ();
 FILLCELL_X32 FILLER_18_1112 ();
 FILLCELL_X32 FILLER_18_1144 ();
 FILLCELL_X32 FILLER_18_1176 ();
 FILLCELL_X32 FILLER_18_1208 ();
 FILLCELL_X32 FILLER_18_1240 ();
 FILLCELL_X32 FILLER_18_1272 ();
 FILLCELL_X32 FILLER_18_1304 ();
 FILLCELL_X32 FILLER_18_1336 ();
 FILLCELL_X32 FILLER_18_1368 ();
 FILLCELL_X32 FILLER_18_1400 ();
 FILLCELL_X32 FILLER_18_1432 ();
 FILLCELL_X32 FILLER_18_1464 ();
 FILLCELL_X32 FILLER_18_1496 ();
 FILLCELL_X32 FILLER_18_1528 ();
 FILLCELL_X32 FILLER_18_1560 ();
 FILLCELL_X32 FILLER_18_1592 ();
 FILLCELL_X32 FILLER_18_1624 ();
 FILLCELL_X32 FILLER_18_1656 ();
 FILLCELL_X32 FILLER_18_1688 ();
 FILLCELL_X32 FILLER_18_1720 ();
 FILLCELL_X32 FILLER_18_1752 ();
 FILLCELL_X32 FILLER_18_1784 ();
 FILLCELL_X32 FILLER_18_1816 ();
 FILLCELL_X32 FILLER_18_1848 ();
 FILLCELL_X8 FILLER_18_1880 ();
 FILLCELL_X4 FILLER_18_1888 ();
 FILLCELL_X2 FILLER_18_1892 ();
 FILLCELL_X32 FILLER_18_1895 ();
 FILLCELL_X32 FILLER_18_1927 ();
 FILLCELL_X32 FILLER_18_1959 ();
 FILLCELL_X32 FILLER_18_1991 ();
 FILLCELL_X32 FILLER_18_2023 ();
 FILLCELL_X32 FILLER_18_2055 ();
 FILLCELL_X32 FILLER_18_2087 ();
 FILLCELL_X32 FILLER_18_2119 ();
 FILLCELL_X32 FILLER_18_2151 ();
 FILLCELL_X32 FILLER_18_2183 ();
 FILLCELL_X32 FILLER_18_2215 ();
 FILLCELL_X32 FILLER_18_2247 ();
 FILLCELL_X32 FILLER_18_2279 ();
 FILLCELL_X32 FILLER_18_2311 ();
 FILLCELL_X32 FILLER_18_2343 ();
 FILLCELL_X32 FILLER_18_2375 ();
 FILLCELL_X32 FILLER_18_2407 ();
 FILLCELL_X32 FILLER_18_2439 ();
 FILLCELL_X32 FILLER_18_2471 ();
 FILLCELL_X32 FILLER_18_2503 ();
 FILLCELL_X32 FILLER_18_2535 ();
 FILLCELL_X32 FILLER_18_2567 ();
 FILLCELL_X32 FILLER_18_2599 ();
 FILLCELL_X32 FILLER_18_2631 ();
 FILLCELL_X32 FILLER_18_2663 ();
 FILLCELL_X32 FILLER_18_2695 ();
 FILLCELL_X32 FILLER_18_2727 ();
 FILLCELL_X32 FILLER_18_2759 ();
 FILLCELL_X32 FILLER_18_2791 ();
 FILLCELL_X32 FILLER_18_2823 ();
 FILLCELL_X32 FILLER_18_2855 ();
 FILLCELL_X32 FILLER_18_2887 ();
 FILLCELL_X32 FILLER_18_2919 ();
 FILLCELL_X32 FILLER_18_2951 ();
 FILLCELL_X32 FILLER_18_2983 ();
 FILLCELL_X32 FILLER_18_3015 ();
 FILLCELL_X32 FILLER_18_3047 ();
 FILLCELL_X32 FILLER_18_3079 ();
 FILLCELL_X32 FILLER_18_3111 ();
 FILLCELL_X8 FILLER_18_3143 ();
 FILLCELL_X4 FILLER_18_3151 ();
 FILLCELL_X2 FILLER_18_3155 ();
 FILLCELL_X32 FILLER_18_3158 ();
 FILLCELL_X32 FILLER_18_3190 ();
 FILLCELL_X32 FILLER_18_3222 ();
 FILLCELL_X32 FILLER_18_3254 ();
 FILLCELL_X32 FILLER_18_3286 ();
 FILLCELL_X32 FILLER_18_3318 ();
 FILLCELL_X32 FILLER_18_3350 ();
 FILLCELL_X32 FILLER_18_3382 ();
 FILLCELL_X32 FILLER_18_3414 ();
 FILLCELL_X32 FILLER_18_3446 ();
 FILLCELL_X32 FILLER_18_3478 ();
 FILLCELL_X32 FILLER_18_3510 ();
 FILLCELL_X32 FILLER_18_3542 ();
 FILLCELL_X32 FILLER_18_3574 ();
 FILLCELL_X32 FILLER_18_3606 ();
 FILLCELL_X32 FILLER_18_3638 ();
 FILLCELL_X32 FILLER_18_3670 ();
 FILLCELL_X32 FILLER_18_3702 ();
 FILLCELL_X4 FILLER_18_3734 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X32 FILLER_19_257 ();
 FILLCELL_X32 FILLER_19_289 ();
 FILLCELL_X32 FILLER_19_321 ();
 FILLCELL_X32 FILLER_19_353 ();
 FILLCELL_X32 FILLER_19_385 ();
 FILLCELL_X32 FILLER_19_417 ();
 FILLCELL_X32 FILLER_19_449 ();
 FILLCELL_X32 FILLER_19_481 ();
 FILLCELL_X32 FILLER_19_513 ();
 FILLCELL_X32 FILLER_19_545 ();
 FILLCELL_X32 FILLER_19_577 ();
 FILLCELL_X32 FILLER_19_609 ();
 FILLCELL_X32 FILLER_19_641 ();
 FILLCELL_X32 FILLER_19_673 ();
 FILLCELL_X32 FILLER_19_705 ();
 FILLCELL_X32 FILLER_19_737 ();
 FILLCELL_X32 FILLER_19_769 ();
 FILLCELL_X32 FILLER_19_801 ();
 FILLCELL_X32 FILLER_19_833 ();
 FILLCELL_X32 FILLER_19_865 ();
 FILLCELL_X32 FILLER_19_897 ();
 FILLCELL_X32 FILLER_19_929 ();
 FILLCELL_X32 FILLER_19_961 ();
 FILLCELL_X32 FILLER_19_993 ();
 FILLCELL_X32 FILLER_19_1025 ();
 FILLCELL_X32 FILLER_19_1057 ();
 FILLCELL_X32 FILLER_19_1089 ();
 FILLCELL_X32 FILLER_19_1121 ();
 FILLCELL_X32 FILLER_19_1153 ();
 FILLCELL_X32 FILLER_19_1185 ();
 FILLCELL_X32 FILLER_19_1217 ();
 FILLCELL_X8 FILLER_19_1249 ();
 FILLCELL_X4 FILLER_19_1257 ();
 FILLCELL_X2 FILLER_19_1261 ();
 FILLCELL_X32 FILLER_19_1264 ();
 FILLCELL_X32 FILLER_19_1296 ();
 FILLCELL_X32 FILLER_19_1328 ();
 FILLCELL_X32 FILLER_19_1360 ();
 FILLCELL_X32 FILLER_19_1392 ();
 FILLCELL_X32 FILLER_19_1424 ();
 FILLCELL_X32 FILLER_19_1456 ();
 FILLCELL_X32 FILLER_19_1488 ();
 FILLCELL_X32 FILLER_19_1520 ();
 FILLCELL_X32 FILLER_19_1552 ();
 FILLCELL_X32 FILLER_19_1584 ();
 FILLCELL_X32 FILLER_19_1616 ();
 FILLCELL_X32 FILLER_19_1648 ();
 FILLCELL_X32 FILLER_19_1680 ();
 FILLCELL_X32 FILLER_19_1712 ();
 FILLCELL_X32 FILLER_19_1744 ();
 FILLCELL_X32 FILLER_19_1776 ();
 FILLCELL_X32 FILLER_19_1808 ();
 FILLCELL_X32 FILLER_19_1840 ();
 FILLCELL_X32 FILLER_19_1872 ();
 FILLCELL_X32 FILLER_19_1904 ();
 FILLCELL_X32 FILLER_19_1936 ();
 FILLCELL_X32 FILLER_19_1968 ();
 FILLCELL_X32 FILLER_19_2000 ();
 FILLCELL_X32 FILLER_19_2032 ();
 FILLCELL_X32 FILLER_19_2064 ();
 FILLCELL_X32 FILLER_19_2096 ();
 FILLCELL_X32 FILLER_19_2128 ();
 FILLCELL_X32 FILLER_19_2160 ();
 FILLCELL_X32 FILLER_19_2192 ();
 FILLCELL_X32 FILLER_19_2224 ();
 FILLCELL_X32 FILLER_19_2256 ();
 FILLCELL_X32 FILLER_19_2288 ();
 FILLCELL_X32 FILLER_19_2320 ();
 FILLCELL_X32 FILLER_19_2352 ();
 FILLCELL_X32 FILLER_19_2384 ();
 FILLCELL_X32 FILLER_19_2416 ();
 FILLCELL_X32 FILLER_19_2448 ();
 FILLCELL_X32 FILLER_19_2480 ();
 FILLCELL_X8 FILLER_19_2512 ();
 FILLCELL_X4 FILLER_19_2520 ();
 FILLCELL_X2 FILLER_19_2524 ();
 FILLCELL_X32 FILLER_19_2527 ();
 FILLCELL_X32 FILLER_19_2559 ();
 FILLCELL_X32 FILLER_19_2591 ();
 FILLCELL_X32 FILLER_19_2623 ();
 FILLCELL_X32 FILLER_19_2655 ();
 FILLCELL_X32 FILLER_19_2687 ();
 FILLCELL_X32 FILLER_19_2719 ();
 FILLCELL_X32 FILLER_19_2751 ();
 FILLCELL_X32 FILLER_19_2783 ();
 FILLCELL_X32 FILLER_19_2815 ();
 FILLCELL_X32 FILLER_19_2847 ();
 FILLCELL_X32 FILLER_19_2879 ();
 FILLCELL_X32 FILLER_19_2911 ();
 FILLCELL_X32 FILLER_19_2943 ();
 FILLCELL_X32 FILLER_19_2975 ();
 FILLCELL_X32 FILLER_19_3007 ();
 FILLCELL_X32 FILLER_19_3039 ();
 FILLCELL_X32 FILLER_19_3071 ();
 FILLCELL_X32 FILLER_19_3103 ();
 FILLCELL_X32 FILLER_19_3135 ();
 FILLCELL_X32 FILLER_19_3167 ();
 FILLCELL_X32 FILLER_19_3199 ();
 FILLCELL_X32 FILLER_19_3231 ();
 FILLCELL_X32 FILLER_19_3263 ();
 FILLCELL_X32 FILLER_19_3295 ();
 FILLCELL_X32 FILLER_19_3327 ();
 FILLCELL_X32 FILLER_19_3359 ();
 FILLCELL_X32 FILLER_19_3391 ();
 FILLCELL_X32 FILLER_19_3423 ();
 FILLCELL_X32 FILLER_19_3455 ();
 FILLCELL_X32 FILLER_19_3487 ();
 FILLCELL_X32 FILLER_19_3519 ();
 FILLCELL_X32 FILLER_19_3551 ();
 FILLCELL_X32 FILLER_19_3583 ();
 FILLCELL_X32 FILLER_19_3615 ();
 FILLCELL_X32 FILLER_19_3647 ();
 FILLCELL_X32 FILLER_19_3679 ();
 FILLCELL_X16 FILLER_19_3711 ();
 FILLCELL_X8 FILLER_19_3727 ();
 FILLCELL_X2 FILLER_19_3735 ();
 FILLCELL_X1 FILLER_19_3737 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X32 FILLER_20_225 ();
 FILLCELL_X32 FILLER_20_257 ();
 FILLCELL_X32 FILLER_20_289 ();
 FILLCELL_X32 FILLER_20_321 ();
 FILLCELL_X32 FILLER_20_353 ();
 FILLCELL_X32 FILLER_20_385 ();
 FILLCELL_X32 FILLER_20_417 ();
 FILLCELL_X32 FILLER_20_449 ();
 FILLCELL_X32 FILLER_20_481 ();
 FILLCELL_X32 FILLER_20_513 ();
 FILLCELL_X32 FILLER_20_545 ();
 FILLCELL_X32 FILLER_20_577 ();
 FILLCELL_X16 FILLER_20_609 ();
 FILLCELL_X4 FILLER_20_625 ();
 FILLCELL_X2 FILLER_20_629 ();
 FILLCELL_X32 FILLER_20_632 ();
 FILLCELL_X32 FILLER_20_664 ();
 FILLCELL_X32 FILLER_20_696 ();
 FILLCELL_X32 FILLER_20_728 ();
 FILLCELL_X32 FILLER_20_760 ();
 FILLCELL_X32 FILLER_20_792 ();
 FILLCELL_X32 FILLER_20_824 ();
 FILLCELL_X32 FILLER_20_856 ();
 FILLCELL_X32 FILLER_20_888 ();
 FILLCELL_X32 FILLER_20_920 ();
 FILLCELL_X32 FILLER_20_952 ();
 FILLCELL_X32 FILLER_20_984 ();
 FILLCELL_X32 FILLER_20_1016 ();
 FILLCELL_X32 FILLER_20_1048 ();
 FILLCELL_X32 FILLER_20_1080 ();
 FILLCELL_X32 FILLER_20_1112 ();
 FILLCELL_X32 FILLER_20_1144 ();
 FILLCELL_X32 FILLER_20_1176 ();
 FILLCELL_X32 FILLER_20_1208 ();
 FILLCELL_X32 FILLER_20_1240 ();
 FILLCELL_X32 FILLER_20_1272 ();
 FILLCELL_X32 FILLER_20_1304 ();
 FILLCELL_X32 FILLER_20_1336 ();
 FILLCELL_X32 FILLER_20_1368 ();
 FILLCELL_X32 FILLER_20_1400 ();
 FILLCELL_X32 FILLER_20_1432 ();
 FILLCELL_X32 FILLER_20_1464 ();
 FILLCELL_X32 FILLER_20_1496 ();
 FILLCELL_X32 FILLER_20_1528 ();
 FILLCELL_X32 FILLER_20_1560 ();
 FILLCELL_X32 FILLER_20_1592 ();
 FILLCELL_X32 FILLER_20_1624 ();
 FILLCELL_X32 FILLER_20_1656 ();
 FILLCELL_X32 FILLER_20_1688 ();
 FILLCELL_X32 FILLER_20_1720 ();
 FILLCELL_X32 FILLER_20_1752 ();
 FILLCELL_X32 FILLER_20_1784 ();
 FILLCELL_X32 FILLER_20_1816 ();
 FILLCELL_X32 FILLER_20_1848 ();
 FILLCELL_X8 FILLER_20_1880 ();
 FILLCELL_X4 FILLER_20_1888 ();
 FILLCELL_X2 FILLER_20_1892 ();
 FILLCELL_X32 FILLER_20_1895 ();
 FILLCELL_X32 FILLER_20_1927 ();
 FILLCELL_X32 FILLER_20_1959 ();
 FILLCELL_X32 FILLER_20_1991 ();
 FILLCELL_X32 FILLER_20_2023 ();
 FILLCELL_X32 FILLER_20_2055 ();
 FILLCELL_X32 FILLER_20_2087 ();
 FILLCELL_X32 FILLER_20_2119 ();
 FILLCELL_X32 FILLER_20_2151 ();
 FILLCELL_X32 FILLER_20_2183 ();
 FILLCELL_X32 FILLER_20_2215 ();
 FILLCELL_X32 FILLER_20_2247 ();
 FILLCELL_X32 FILLER_20_2279 ();
 FILLCELL_X32 FILLER_20_2311 ();
 FILLCELL_X32 FILLER_20_2343 ();
 FILLCELL_X32 FILLER_20_2375 ();
 FILLCELL_X32 FILLER_20_2407 ();
 FILLCELL_X32 FILLER_20_2439 ();
 FILLCELL_X32 FILLER_20_2471 ();
 FILLCELL_X32 FILLER_20_2503 ();
 FILLCELL_X32 FILLER_20_2535 ();
 FILLCELL_X32 FILLER_20_2567 ();
 FILLCELL_X32 FILLER_20_2599 ();
 FILLCELL_X32 FILLER_20_2631 ();
 FILLCELL_X32 FILLER_20_2663 ();
 FILLCELL_X32 FILLER_20_2695 ();
 FILLCELL_X32 FILLER_20_2727 ();
 FILLCELL_X32 FILLER_20_2759 ();
 FILLCELL_X32 FILLER_20_2791 ();
 FILLCELL_X32 FILLER_20_2823 ();
 FILLCELL_X32 FILLER_20_2855 ();
 FILLCELL_X32 FILLER_20_2887 ();
 FILLCELL_X32 FILLER_20_2919 ();
 FILLCELL_X32 FILLER_20_2951 ();
 FILLCELL_X32 FILLER_20_2983 ();
 FILLCELL_X32 FILLER_20_3015 ();
 FILLCELL_X32 FILLER_20_3047 ();
 FILLCELL_X32 FILLER_20_3079 ();
 FILLCELL_X32 FILLER_20_3111 ();
 FILLCELL_X8 FILLER_20_3143 ();
 FILLCELL_X4 FILLER_20_3151 ();
 FILLCELL_X2 FILLER_20_3155 ();
 FILLCELL_X32 FILLER_20_3158 ();
 FILLCELL_X32 FILLER_20_3190 ();
 FILLCELL_X32 FILLER_20_3222 ();
 FILLCELL_X32 FILLER_20_3254 ();
 FILLCELL_X32 FILLER_20_3286 ();
 FILLCELL_X32 FILLER_20_3318 ();
 FILLCELL_X32 FILLER_20_3350 ();
 FILLCELL_X32 FILLER_20_3382 ();
 FILLCELL_X32 FILLER_20_3414 ();
 FILLCELL_X32 FILLER_20_3446 ();
 FILLCELL_X32 FILLER_20_3478 ();
 FILLCELL_X32 FILLER_20_3510 ();
 FILLCELL_X32 FILLER_20_3542 ();
 FILLCELL_X32 FILLER_20_3574 ();
 FILLCELL_X32 FILLER_20_3606 ();
 FILLCELL_X32 FILLER_20_3638 ();
 FILLCELL_X32 FILLER_20_3670 ();
 FILLCELL_X32 FILLER_20_3702 ();
 FILLCELL_X4 FILLER_20_3734 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X32 FILLER_21_225 ();
 FILLCELL_X32 FILLER_21_257 ();
 FILLCELL_X32 FILLER_21_289 ();
 FILLCELL_X32 FILLER_21_321 ();
 FILLCELL_X32 FILLER_21_353 ();
 FILLCELL_X32 FILLER_21_385 ();
 FILLCELL_X32 FILLER_21_417 ();
 FILLCELL_X32 FILLER_21_449 ();
 FILLCELL_X32 FILLER_21_481 ();
 FILLCELL_X32 FILLER_21_513 ();
 FILLCELL_X32 FILLER_21_545 ();
 FILLCELL_X32 FILLER_21_577 ();
 FILLCELL_X32 FILLER_21_609 ();
 FILLCELL_X32 FILLER_21_641 ();
 FILLCELL_X32 FILLER_21_673 ();
 FILLCELL_X32 FILLER_21_705 ();
 FILLCELL_X32 FILLER_21_737 ();
 FILLCELL_X32 FILLER_21_769 ();
 FILLCELL_X32 FILLER_21_801 ();
 FILLCELL_X32 FILLER_21_833 ();
 FILLCELL_X32 FILLER_21_865 ();
 FILLCELL_X32 FILLER_21_897 ();
 FILLCELL_X32 FILLER_21_929 ();
 FILLCELL_X32 FILLER_21_961 ();
 FILLCELL_X32 FILLER_21_993 ();
 FILLCELL_X32 FILLER_21_1025 ();
 FILLCELL_X32 FILLER_21_1057 ();
 FILLCELL_X32 FILLER_21_1089 ();
 FILLCELL_X32 FILLER_21_1121 ();
 FILLCELL_X32 FILLER_21_1153 ();
 FILLCELL_X32 FILLER_21_1185 ();
 FILLCELL_X32 FILLER_21_1217 ();
 FILLCELL_X8 FILLER_21_1249 ();
 FILLCELL_X4 FILLER_21_1257 ();
 FILLCELL_X2 FILLER_21_1261 ();
 FILLCELL_X32 FILLER_21_1264 ();
 FILLCELL_X32 FILLER_21_1296 ();
 FILLCELL_X32 FILLER_21_1328 ();
 FILLCELL_X32 FILLER_21_1360 ();
 FILLCELL_X32 FILLER_21_1392 ();
 FILLCELL_X32 FILLER_21_1424 ();
 FILLCELL_X32 FILLER_21_1456 ();
 FILLCELL_X32 FILLER_21_1488 ();
 FILLCELL_X32 FILLER_21_1520 ();
 FILLCELL_X32 FILLER_21_1552 ();
 FILLCELL_X32 FILLER_21_1584 ();
 FILLCELL_X32 FILLER_21_1616 ();
 FILLCELL_X32 FILLER_21_1648 ();
 FILLCELL_X32 FILLER_21_1680 ();
 FILLCELL_X32 FILLER_21_1712 ();
 FILLCELL_X32 FILLER_21_1744 ();
 FILLCELL_X32 FILLER_21_1776 ();
 FILLCELL_X32 FILLER_21_1808 ();
 FILLCELL_X32 FILLER_21_1840 ();
 FILLCELL_X32 FILLER_21_1872 ();
 FILLCELL_X32 FILLER_21_1904 ();
 FILLCELL_X32 FILLER_21_1936 ();
 FILLCELL_X32 FILLER_21_1968 ();
 FILLCELL_X32 FILLER_21_2000 ();
 FILLCELL_X32 FILLER_21_2032 ();
 FILLCELL_X32 FILLER_21_2064 ();
 FILLCELL_X32 FILLER_21_2096 ();
 FILLCELL_X32 FILLER_21_2128 ();
 FILLCELL_X32 FILLER_21_2160 ();
 FILLCELL_X32 FILLER_21_2192 ();
 FILLCELL_X32 FILLER_21_2224 ();
 FILLCELL_X32 FILLER_21_2256 ();
 FILLCELL_X32 FILLER_21_2288 ();
 FILLCELL_X32 FILLER_21_2320 ();
 FILLCELL_X32 FILLER_21_2352 ();
 FILLCELL_X32 FILLER_21_2384 ();
 FILLCELL_X32 FILLER_21_2416 ();
 FILLCELL_X32 FILLER_21_2448 ();
 FILLCELL_X32 FILLER_21_2480 ();
 FILLCELL_X8 FILLER_21_2512 ();
 FILLCELL_X4 FILLER_21_2520 ();
 FILLCELL_X2 FILLER_21_2524 ();
 FILLCELL_X32 FILLER_21_2527 ();
 FILLCELL_X32 FILLER_21_2559 ();
 FILLCELL_X32 FILLER_21_2591 ();
 FILLCELL_X32 FILLER_21_2623 ();
 FILLCELL_X32 FILLER_21_2655 ();
 FILLCELL_X32 FILLER_21_2687 ();
 FILLCELL_X32 FILLER_21_2719 ();
 FILLCELL_X32 FILLER_21_2751 ();
 FILLCELL_X32 FILLER_21_2783 ();
 FILLCELL_X32 FILLER_21_2815 ();
 FILLCELL_X32 FILLER_21_2847 ();
 FILLCELL_X32 FILLER_21_2879 ();
 FILLCELL_X32 FILLER_21_2911 ();
 FILLCELL_X32 FILLER_21_2943 ();
 FILLCELL_X32 FILLER_21_2975 ();
 FILLCELL_X32 FILLER_21_3007 ();
 FILLCELL_X32 FILLER_21_3039 ();
 FILLCELL_X32 FILLER_21_3071 ();
 FILLCELL_X32 FILLER_21_3103 ();
 FILLCELL_X32 FILLER_21_3135 ();
 FILLCELL_X32 FILLER_21_3167 ();
 FILLCELL_X32 FILLER_21_3199 ();
 FILLCELL_X32 FILLER_21_3231 ();
 FILLCELL_X32 FILLER_21_3263 ();
 FILLCELL_X32 FILLER_21_3295 ();
 FILLCELL_X32 FILLER_21_3327 ();
 FILLCELL_X32 FILLER_21_3359 ();
 FILLCELL_X32 FILLER_21_3391 ();
 FILLCELL_X32 FILLER_21_3423 ();
 FILLCELL_X32 FILLER_21_3455 ();
 FILLCELL_X32 FILLER_21_3487 ();
 FILLCELL_X32 FILLER_21_3519 ();
 FILLCELL_X32 FILLER_21_3551 ();
 FILLCELL_X32 FILLER_21_3583 ();
 FILLCELL_X32 FILLER_21_3615 ();
 FILLCELL_X32 FILLER_21_3647 ();
 FILLCELL_X32 FILLER_21_3679 ();
 FILLCELL_X16 FILLER_21_3711 ();
 FILLCELL_X8 FILLER_21_3727 ();
 FILLCELL_X2 FILLER_21_3735 ();
 FILLCELL_X1 FILLER_21_3737 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X32 FILLER_22_225 ();
 FILLCELL_X32 FILLER_22_257 ();
 FILLCELL_X32 FILLER_22_289 ();
 FILLCELL_X32 FILLER_22_321 ();
 FILLCELL_X32 FILLER_22_353 ();
 FILLCELL_X32 FILLER_22_385 ();
 FILLCELL_X32 FILLER_22_417 ();
 FILLCELL_X32 FILLER_22_449 ();
 FILLCELL_X32 FILLER_22_481 ();
 FILLCELL_X32 FILLER_22_513 ();
 FILLCELL_X32 FILLER_22_545 ();
 FILLCELL_X32 FILLER_22_577 ();
 FILLCELL_X16 FILLER_22_609 ();
 FILLCELL_X4 FILLER_22_625 ();
 FILLCELL_X2 FILLER_22_629 ();
 FILLCELL_X32 FILLER_22_632 ();
 FILLCELL_X32 FILLER_22_664 ();
 FILLCELL_X32 FILLER_22_696 ();
 FILLCELL_X32 FILLER_22_728 ();
 FILLCELL_X32 FILLER_22_760 ();
 FILLCELL_X32 FILLER_22_792 ();
 FILLCELL_X32 FILLER_22_824 ();
 FILLCELL_X32 FILLER_22_856 ();
 FILLCELL_X32 FILLER_22_888 ();
 FILLCELL_X32 FILLER_22_920 ();
 FILLCELL_X32 FILLER_22_952 ();
 FILLCELL_X32 FILLER_22_984 ();
 FILLCELL_X32 FILLER_22_1016 ();
 FILLCELL_X32 FILLER_22_1048 ();
 FILLCELL_X32 FILLER_22_1080 ();
 FILLCELL_X32 FILLER_22_1112 ();
 FILLCELL_X32 FILLER_22_1144 ();
 FILLCELL_X32 FILLER_22_1176 ();
 FILLCELL_X32 FILLER_22_1208 ();
 FILLCELL_X32 FILLER_22_1240 ();
 FILLCELL_X32 FILLER_22_1272 ();
 FILLCELL_X32 FILLER_22_1304 ();
 FILLCELL_X32 FILLER_22_1336 ();
 FILLCELL_X32 FILLER_22_1368 ();
 FILLCELL_X32 FILLER_22_1400 ();
 FILLCELL_X32 FILLER_22_1432 ();
 FILLCELL_X32 FILLER_22_1464 ();
 FILLCELL_X32 FILLER_22_1496 ();
 FILLCELL_X32 FILLER_22_1528 ();
 FILLCELL_X32 FILLER_22_1560 ();
 FILLCELL_X32 FILLER_22_1592 ();
 FILLCELL_X32 FILLER_22_1624 ();
 FILLCELL_X32 FILLER_22_1656 ();
 FILLCELL_X32 FILLER_22_1688 ();
 FILLCELL_X32 FILLER_22_1720 ();
 FILLCELL_X32 FILLER_22_1752 ();
 FILLCELL_X32 FILLER_22_1784 ();
 FILLCELL_X32 FILLER_22_1816 ();
 FILLCELL_X32 FILLER_22_1848 ();
 FILLCELL_X8 FILLER_22_1880 ();
 FILLCELL_X4 FILLER_22_1888 ();
 FILLCELL_X2 FILLER_22_1892 ();
 FILLCELL_X32 FILLER_22_1895 ();
 FILLCELL_X32 FILLER_22_1927 ();
 FILLCELL_X32 FILLER_22_1959 ();
 FILLCELL_X32 FILLER_22_1991 ();
 FILLCELL_X32 FILLER_22_2023 ();
 FILLCELL_X32 FILLER_22_2055 ();
 FILLCELL_X32 FILLER_22_2087 ();
 FILLCELL_X32 FILLER_22_2119 ();
 FILLCELL_X32 FILLER_22_2151 ();
 FILLCELL_X32 FILLER_22_2183 ();
 FILLCELL_X32 FILLER_22_2215 ();
 FILLCELL_X32 FILLER_22_2247 ();
 FILLCELL_X32 FILLER_22_2279 ();
 FILLCELL_X32 FILLER_22_2311 ();
 FILLCELL_X32 FILLER_22_2343 ();
 FILLCELL_X32 FILLER_22_2375 ();
 FILLCELL_X32 FILLER_22_2407 ();
 FILLCELL_X32 FILLER_22_2439 ();
 FILLCELL_X32 FILLER_22_2471 ();
 FILLCELL_X32 FILLER_22_2503 ();
 FILLCELL_X32 FILLER_22_2535 ();
 FILLCELL_X32 FILLER_22_2567 ();
 FILLCELL_X32 FILLER_22_2599 ();
 FILLCELL_X32 FILLER_22_2631 ();
 FILLCELL_X32 FILLER_22_2663 ();
 FILLCELL_X32 FILLER_22_2695 ();
 FILLCELL_X32 FILLER_22_2727 ();
 FILLCELL_X32 FILLER_22_2759 ();
 FILLCELL_X32 FILLER_22_2791 ();
 FILLCELL_X32 FILLER_22_2823 ();
 FILLCELL_X32 FILLER_22_2855 ();
 FILLCELL_X32 FILLER_22_2887 ();
 FILLCELL_X32 FILLER_22_2919 ();
 FILLCELL_X32 FILLER_22_2951 ();
 FILLCELL_X32 FILLER_22_2983 ();
 FILLCELL_X32 FILLER_22_3015 ();
 FILLCELL_X32 FILLER_22_3047 ();
 FILLCELL_X32 FILLER_22_3079 ();
 FILLCELL_X32 FILLER_22_3111 ();
 FILLCELL_X8 FILLER_22_3143 ();
 FILLCELL_X4 FILLER_22_3151 ();
 FILLCELL_X2 FILLER_22_3155 ();
 FILLCELL_X32 FILLER_22_3158 ();
 FILLCELL_X32 FILLER_22_3190 ();
 FILLCELL_X32 FILLER_22_3222 ();
 FILLCELL_X32 FILLER_22_3254 ();
 FILLCELL_X32 FILLER_22_3286 ();
 FILLCELL_X32 FILLER_22_3318 ();
 FILLCELL_X32 FILLER_22_3350 ();
 FILLCELL_X32 FILLER_22_3382 ();
 FILLCELL_X32 FILLER_22_3414 ();
 FILLCELL_X32 FILLER_22_3446 ();
 FILLCELL_X32 FILLER_22_3478 ();
 FILLCELL_X32 FILLER_22_3510 ();
 FILLCELL_X32 FILLER_22_3542 ();
 FILLCELL_X32 FILLER_22_3574 ();
 FILLCELL_X32 FILLER_22_3606 ();
 FILLCELL_X32 FILLER_22_3638 ();
 FILLCELL_X32 FILLER_22_3670 ();
 FILLCELL_X32 FILLER_22_3702 ();
 FILLCELL_X4 FILLER_22_3734 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X32 FILLER_23_225 ();
 FILLCELL_X32 FILLER_23_257 ();
 FILLCELL_X32 FILLER_23_289 ();
 FILLCELL_X32 FILLER_23_321 ();
 FILLCELL_X32 FILLER_23_353 ();
 FILLCELL_X32 FILLER_23_385 ();
 FILLCELL_X32 FILLER_23_417 ();
 FILLCELL_X32 FILLER_23_449 ();
 FILLCELL_X32 FILLER_23_481 ();
 FILLCELL_X32 FILLER_23_513 ();
 FILLCELL_X32 FILLER_23_545 ();
 FILLCELL_X32 FILLER_23_577 ();
 FILLCELL_X32 FILLER_23_609 ();
 FILLCELL_X32 FILLER_23_641 ();
 FILLCELL_X32 FILLER_23_673 ();
 FILLCELL_X32 FILLER_23_705 ();
 FILLCELL_X32 FILLER_23_737 ();
 FILLCELL_X32 FILLER_23_769 ();
 FILLCELL_X32 FILLER_23_801 ();
 FILLCELL_X32 FILLER_23_833 ();
 FILLCELL_X32 FILLER_23_865 ();
 FILLCELL_X32 FILLER_23_897 ();
 FILLCELL_X32 FILLER_23_929 ();
 FILLCELL_X32 FILLER_23_961 ();
 FILLCELL_X32 FILLER_23_993 ();
 FILLCELL_X32 FILLER_23_1025 ();
 FILLCELL_X32 FILLER_23_1057 ();
 FILLCELL_X32 FILLER_23_1089 ();
 FILLCELL_X32 FILLER_23_1121 ();
 FILLCELL_X32 FILLER_23_1153 ();
 FILLCELL_X32 FILLER_23_1185 ();
 FILLCELL_X32 FILLER_23_1217 ();
 FILLCELL_X8 FILLER_23_1249 ();
 FILLCELL_X4 FILLER_23_1257 ();
 FILLCELL_X2 FILLER_23_1261 ();
 FILLCELL_X32 FILLER_23_1264 ();
 FILLCELL_X32 FILLER_23_1296 ();
 FILLCELL_X32 FILLER_23_1328 ();
 FILLCELL_X32 FILLER_23_1360 ();
 FILLCELL_X32 FILLER_23_1392 ();
 FILLCELL_X32 FILLER_23_1424 ();
 FILLCELL_X32 FILLER_23_1456 ();
 FILLCELL_X32 FILLER_23_1488 ();
 FILLCELL_X32 FILLER_23_1520 ();
 FILLCELL_X32 FILLER_23_1552 ();
 FILLCELL_X32 FILLER_23_1584 ();
 FILLCELL_X32 FILLER_23_1616 ();
 FILLCELL_X32 FILLER_23_1648 ();
 FILLCELL_X32 FILLER_23_1680 ();
 FILLCELL_X32 FILLER_23_1712 ();
 FILLCELL_X32 FILLER_23_1744 ();
 FILLCELL_X32 FILLER_23_1776 ();
 FILLCELL_X32 FILLER_23_1808 ();
 FILLCELL_X32 FILLER_23_1840 ();
 FILLCELL_X32 FILLER_23_1872 ();
 FILLCELL_X32 FILLER_23_1904 ();
 FILLCELL_X32 FILLER_23_1936 ();
 FILLCELL_X32 FILLER_23_1968 ();
 FILLCELL_X32 FILLER_23_2000 ();
 FILLCELL_X32 FILLER_23_2032 ();
 FILLCELL_X32 FILLER_23_2064 ();
 FILLCELL_X32 FILLER_23_2096 ();
 FILLCELL_X32 FILLER_23_2128 ();
 FILLCELL_X32 FILLER_23_2160 ();
 FILLCELL_X32 FILLER_23_2192 ();
 FILLCELL_X32 FILLER_23_2224 ();
 FILLCELL_X32 FILLER_23_2256 ();
 FILLCELL_X32 FILLER_23_2288 ();
 FILLCELL_X32 FILLER_23_2320 ();
 FILLCELL_X32 FILLER_23_2352 ();
 FILLCELL_X32 FILLER_23_2384 ();
 FILLCELL_X32 FILLER_23_2416 ();
 FILLCELL_X32 FILLER_23_2448 ();
 FILLCELL_X32 FILLER_23_2480 ();
 FILLCELL_X8 FILLER_23_2512 ();
 FILLCELL_X4 FILLER_23_2520 ();
 FILLCELL_X2 FILLER_23_2524 ();
 FILLCELL_X32 FILLER_23_2527 ();
 FILLCELL_X32 FILLER_23_2559 ();
 FILLCELL_X32 FILLER_23_2591 ();
 FILLCELL_X32 FILLER_23_2623 ();
 FILLCELL_X32 FILLER_23_2655 ();
 FILLCELL_X32 FILLER_23_2687 ();
 FILLCELL_X32 FILLER_23_2719 ();
 FILLCELL_X32 FILLER_23_2751 ();
 FILLCELL_X32 FILLER_23_2783 ();
 FILLCELL_X32 FILLER_23_2815 ();
 FILLCELL_X32 FILLER_23_2847 ();
 FILLCELL_X32 FILLER_23_2879 ();
 FILLCELL_X32 FILLER_23_2911 ();
 FILLCELL_X32 FILLER_23_2943 ();
 FILLCELL_X32 FILLER_23_2975 ();
 FILLCELL_X32 FILLER_23_3007 ();
 FILLCELL_X32 FILLER_23_3039 ();
 FILLCELL_X32 FILLER_23_3071 ();
 FILLCELL_X32 FILLER_23_3103 ();
 FILLCELL_X32 FILLER_23_3135 ();
 FILLCELL_X32 FILLER_23_3167 ();
 FILLCELL_X32 FILLER_23_3199 ();
 FILLCELL_X32 FILLER_23_3231 ();
 FILLCELL_X32 FILLER_23_3263 ();
 FILLCELL_X32 FILLER_23_3295 ();
 FILLCELL_X32 FILLER_23_3327 ();
 FILLCELL_X32 FILLER_23_3359 ();
 FILLCELL_X32 FILLER_23_3391 ();
 FILLCELL_X32 FILLER_23_3423 ();
 FILLCELL_X32 FILLER_23_3455 ();
 FILLCELL_X32 FILLER_23_3487 ();
 FILLCELL_X32 FILLER_23_3519 ();
 FILLCELL_X32 FILLER_23_3551 ();
 FILLCELL_X32 FILLER_23_3583 ();
 FILLCELL_X32 FILLER_23_3615 ();
 FILLCELL_X32 FILLER_23_3647 ();
 FILLCELL_X32 FILLER_23_3679 ();
 FILLCELL_X16 FILLER_23_3711 ();
 FILLCELL_X8 FILLER_23_3727 ();
 FILLCELL_X2 FILLER_23_3735 ();
 FILLCELL_X1 FILLER_23_3737 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X32 FILLER_24_225 ();
 FILLCELL_X32 FILLER_24_257 ();
 FILLCELL_X32 FILLER_24_289 ();
 FILLCELL_X32 FILLER_24_321 ();
 FILLCELL_X32 FILLER_24_353 ();
 FILLCELL_X32 FILLER_24_385 ();
 FILLCELL_X32 FILLER_24_417 ();
 FILLCELL_X32 FILLER_24_449 ();
 FILLCELL_X32 FILLER_24_481 ();
 FILLCELL_X32 FILLER_24_513 ();
 FILLCELL_X32 FILLER_24_545 ();
 FILLCELL_X32 FILLER_24_577 ();
 FILLCELL_X16 FILLER_24_609 ();
 FILLCELL_X4 FILLER_24_625 ();
 FILLCELL_X2 FILLER_24_629 ();
 FILLCELL_X32 FILLER_24_632 ();
 FILLCELL_X32 FILLER_24_664 ();
 FILLCELL_X32 FILLER_24_696 ();
 FILLCELL_X32 FILLER_24_728 ();
 FILLCELL_X32 FILLER_24_760 ();
 FILLCELL_X32 FILLER_24_792 ();
 FILLCELL_X32 FILLER_24_824 ();
 FILLCELL_X32 FILLER_24_856 ();
 FILLCELL_X32 FILLER_24_888 ();
 FILLCELL_X32 FILLER_24_920 ();
 FILLCELL_X32 FILLER_24_952 ();
 FILLCELL_X32 FILLER_24_984 ();
 FILLCELL_X32 FILLER_24_1016 ();
 FILLCELL_X32 FILLER_24_1048 ();
 FILLCELL_X32 FILLER_24_1080 ();
 FILLCELL_X32 FILLER_24_1112 ();
 FILLCELL_X32 FILLER_24_1144 ();
 FILLCELL_X32 FILLER_24_1176 ();
 FILLCELL_X32 FILLER_24_1208 ();
 FILLCELL_X32 FILLER_24_1240 ();
 FILLCELL_X32 FILLER_24_1272 ();
 FILLCELL_X32 FILLER_24_1304 ();
 FILLCELL_X32 FILLER_24_1336 ();
 FILLCELL_X32 FILLER_24_1368 ();
 FILLCELL_X32 FILLER_24_1400 ();
 FILLCELL_X32 FILLER_24_1432 ();
 FILLCELL_X32 FILLER_24_1464 ();
 FILLCELL_X32 FILLER_24_1496 ();
 FILLCELL_X32 FILLER_24_1528 ();
 FILLCELL_X32 FILLER_24_1560 ();
 FILLCELL_X32 FILLER_24_1592 ();
 FILLCELL_X32 FILLER_24_1624 ();
 FILLCELL_X32 FILLER_24_1656 ();
 FILLCELL_X32 FILLER_24_1688 ();
 FILLCELL_X32 FILLER_24_1720 ();
 FILLCELL_X32 FILLER_24_1752 ();
 FILLCELL_X32 FILLER_24_1784 ();
 FILLCELL_X32 FILLER_24_1816 ();
 FILLCELL_X32 FILLER_24_1848 ();
 FILLCELL_X8 FILLER_24_1880 ();
 FILLCELL_X4 FILLER_24_1888 ();
 FILLCELL_X2 FILLER_24_1892 ();
 FILLCELL_X32 FILLER_24_1895 ();
 FILLCELL_X32 FILLER_24_1927 ();
 FILLCELL_X32 FILLER_24_1959 ();
 FILLCELL_X32 FILLER_24_1991 ();
 FILLCELL_X32 FILLER_24_2023 ();
 FILLCELL_X32 FILLER_24_2055 ();
 FILLCELL_X32 FILLER_24_2087 ();
 FILLCELL_X32 FILLER_24_2119 ();
 FILLCELL_X32 FILLER_24_2151 ();
 FILLCELL_X32 FILLER_24_2183 ();
 FILLCELL_X32 FILLER_24_2215 ();
 FILLCELL_X32 FILLER_24_2247 ();
 FILLCELL_X32 FILLER_24_2279 ();
 FILLCELL_X32 FILLER_24_2311 ();
 FILLCELL_X32 FILLER_24_2343 ();
 FILLCELL_X32 FILLER_24_2375 ();
 FILLCELL_X32 FILLER_24_2407 ();
 FILLCELL_X32 FILLER_24_2439 ();
 FILLCELL_X32 FILLER_24_2471 ();
 FILLCELL_X32 FILLER_24_2503 ();
 FILLCELL_X32 FILLER_24_2535 ();
 FILLCELL_X32 FILLER_24_2567 ();
 FILLCELL_X32 FILLER_24_2599 ();
 FILLCELL_X32 FILLER_24_2631 ();
 FILLCELL_X32 FILLER_24_2663 ();
 FILLCELL_X32 FILLER_24_2695 ();
 FILLCELL_X32 FILLER_24_2727 ();
 FILLCELL_X32 FILLER_24_2759 ();
 FILLCELL_X32 FILLER_24_2791 ();
 FILLCELL_X32 FILLER_24_2823 ();
 FILLCELL_X32 FILLER_24_2855 ();
 FILLCELL_X32 FILLER_24_2887 ();
 FILLCELL_X32 FILLER_24_2919 ();
 FILLCELL_X32 FILLER_24_2951 ();
 FILLCELL_X32 FILLER_24_2983 ();
 FILLCELL_X32 FILLER_24_3015 ();
 FILLCELL_X32 FILLER_24_3047 ();
 FILLCELL_X32 FILLER_24_3079 ();
 FILLCELL_X32 FILLER_24_3111 ();
 FILLCELL_X8 FILLER_24_3143 ();
 FILLCELL_X4 FILLER_24_3151 ();
 FILLCELL_X2 FILLER_24_3155 ();
 FILLCELL_X32 FILLER_24_3158 ();
 FILLCELL_X32 FILLER_24_3190 ();
 FILLCELL_X32 FILLER_24_3222 ();
 FILLCELL_X32 FILLER_24_3254 ();
 FILLCELL_X32 FILLER_24_3286 ();
 FILLCELL_X32 FILLER_24_3318 ();
 FILLCELL_X32 FILLER_24_3350 ();
 FILLCELL_X32 FILLER_24_3382 ();
 FILLCELL_X32 FILLER_24_3414 ();
 FILLCELL_X32 FILLER_24_3446 ();
 FILLCELL_X32 FILLER_24_3478 ();
 FILLCELL_X32 FILLER_24_3510 ();
 FILLCELL_X32 FILLER_24_3542 ();
 FILLCELL_X32 FILLER_24_3574 ();
 FILLCELL_X32 FILLER_24_3606 ();
 FILLCELL_X32 FILLER_24_3638 ();
 FILLCELL_X32 FILLER_24_3670 ();
 FILLCELL_X32 FILLER_24_3702 ();
 FILLCELL_X4 FILLER_24_3734 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X32 FILLER_25_225 ();
 FILLCELL_X32 FILLER_25_257 ();
 FILLCELL_X32 FILLER_25_289 ();
 FILLCELL_X32 FILLER_25_321 ();
 FILLCELL_X32 FILLER_25_353 ();
 FILLCELL_X32 FILLER_25_385 ();
 FILLCELL_X32 FILLER_25_417 ();
 FILLCELL_X32 FILLER_25_449 ();
 FILLCELL_X32 FILLER_25_481 ();
 FILLCELL_X32 FILLER_25_513 ();
 FILLCELL_X32 FILLER_25_545 ();
 FILLCELL_X32 FILLER_25_577 ();
 FILLCELL_X32 FILLER_25_609 ();
 FILLCELL_X32 FILLER_25_641 ();
 FILLCELL_X32 FILLER_25_673 ();
 FILLCELL_X32 FILLER_25_705 ();
 FILLCELL_X32 FILLER_25_737 ();
 FILLCELL_X32 FILLER_25_769 ();
 FILLCELL_X32 FILLER_25_801 ();
 FILLCELL_X32 FILLER_25_833 ();
 FILLCELL_X32 FILLER_25_865 ();
 FILLCELL_X32 FILLER_25_897 ();
 FILLCELL_X32 FILLER_25_929 ();
 FILLCELL_X32 FILLER_25_961 ();
 FILLCELL_X32 FILLER_25_993 ();
 FILLCELL_X32 FILLER_25_1025 ();
 FILLCELL_X32 FILLER_25_1057 ();
 FILLCELL_X32 FILLER_25_1089 ();
 FILLCELL_X32 FILLER_25_1121 ();
 FILLCELL_X32 FILLER_25_1153 ();
 FILLCELL_X32 FILLER_25_1185 ();
 FILLCELL_X32 FILLER_25_1217 ();
 FILLCELL_X8 FILLER_25_1249 ();
 FILLCELL_X4 FILLER_25_1257 ();
 FILLCELL_X2 FILLER_25_1261 ();
 FILLCELL_X32 FILLER_25_1264 ();
 FILLCELL_X32 FILLER_25_1296 ();
 FILLCELL_X32 FILLER_25_1328 ();
 FILLCELL_X32 FILLER_25_1360 ();
 FILLCELL_X32 FILLER_25_1392 ();
 FILLCELL_X32 FILLER_25_1424 ();
 FILLCELL_X32 FILLER_25_1456 ();
 FILLCELL_X32 FILLER_25_1488 ();
 FILLCELL_X32 FILLER_25_1520 ();
 FILLCELL_X32 FILLER_25_1552 ();
 FILLCELL_X32 FILLER_25_1584 ();
 FILLCELL_X32 FILLER_25_1616 ();
 FILLCELL_X32 FILLER_25_1648 ();
 FILLCELL_X32 FILLER_25_1680 ();
 FILLCELL_X32 FILLER_25_1712 ();
 FILLCELL_X32 FILLER_25_1744 ();
 FILLCELL_X32 FILLER_25_1776 ();
 FILLCELL_X32 FILLER_25_1808 ();
 FILLCELL_X32 FILLER_25_1840 ();
 FILLCELL_X32 FILLER_25_1872 ();
 FILLCELL_X32 FILLER_25_1904 ();
 FILLCELL_X32 FILLER_25_1936 ();
 FILLCELL_X32 FILLER_25_1968 ();
 FILLCELL_X32 FILLER_25_2000 ();
 FILLCELL_X32 FILLER_25_2032 ();
 FILLCELL_X32 FILLER_25_2064 ();
 FILLCELL_X32 FILLER_25_2096 ();
 FILLCELL_X32 FILLER_25_2128 ();
 FILLCELL_X32 FILLER_25_2160 ();
 FILLCELL_X32 FILLER_25_2192 ();
 FILLCELL_X32 FILLER_25_2224 ();
 FILLCELL_X32 FILLER_25_2256 ();
 FILLCELL_X32 FILLER_25_2288 ();
 FILLCELL_X32 FILLER_25_2320 ();
 FILLCELL_X32 FILLER_25_2352 ();
 FILLCELL_X32 FILLER_25_2384 ();
 FILLCELL_X32 FILLER_25_2416 ();
 FILLCELL_X32 FILLER_25_2448 ();
 FILLCELL_X32 FILLER_25_2480 ();
 FILLCELL_X8 FILLER_25_2512 ();
 FILLCELL_X4 FILLER_25_2520 ();
 FILLCELL_X2 FILLER_25_2524 ();
 FILLCELL_X32 FILLER_25_2527 ();
 FILLCELL_X32 FILLER_25_2559 ();
 FILLCELL_X32 FILLER_25_2591 ();
 FILLCELL_X32 FILLER_25_2623 ();
 FILLCELL_X32 FILLER_25_2655 ();
 FILLCELL_X32 FILLER_25_2687 ();
 FILLCELL_X32 FILLER_25_2719 ();
 FILLCELL_X32 FILLER_25_2751 ();
 FILLCELL_X32 FILLER_25_2783 ();
 FILLCELL_X32 FILLER_25_2815 ();
 FILLCELL_X32 FILLER_25_2847 ();
 FILLCELL_X32 FILLER_25_2879 ();
 FILLCELL_X32 FILLER_25_2911 ();
 FILLCELL_X32 FILLER_25_2943 ();
 FILLCELL_X32 FILLER_25_2975 ();
 FILLCELL_X32 FILLER_25_3007 ();
 FILLCELL_X32 FILLER_25_3039 ();
 FILLCELL_X32 FILLER_25_3071 ();
 FILLCELL_X32 FILLER_25_3103 ();
 FILLCELL_X32 FILLER_25_3135 ();
 FILLCELL_X32 FILLER_25_3167 ();
 FILLCELL_X32 FILLER_25_3199 ();
 FILLCELL_X32 FILLER_25_3231 ();
 FILLCELL_X32 FILLER_25_3263 ();
 FILLCELL_X32 FILLER_25_3295 ();
 FILLCELL_X32 FILLER_25_3327 ();
 FILLCELL_X32 FILLER_25_3359 ();
 FILLCELL_X32 FILLER_25_3391 ();
 FILLCELL_X32 FILLER_25_3423 ();
 FILLCELL_X32 FILLER_25_3455 ();
 FILLCELL_X32 FILLER_25_3487 ();
 FILLCELL_X32 FILLER_25_3519 ();
 FILLCELL_X32 FILLER_25_3551 ();
 FILLCELL_X32 FILLER_25_3583 ();
 FILLCELL_X32 FILLER_25_3615 ();
 FILLCELL_X32 FILLER_25_3647 ();
 FILLCELL_X32 FILLER_25_3679 ();
 FILLCELL_X16 FILLER_25_3711 ();
 FILLCELL_X8 FILLER_25_3727 ();
 FILLCELL_X2 FILLER_25_3735 ();
 FILLCELL_X1 FILLER_25_3737 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X32 FILLER_26_225 ();
 FILLCELL_X32 FILLER_26_257 ();
 FILLCELL_X32 FILLER_26_289 ();
 FILLCELL_X32 FILLER_26_321 ();
 FILLCELL_X32 FILLER_26_353 ();
 FILLCELL_X32 FILLER_26_385 ();
 FILLCELL_X32 FILLER_26_417 ();
 FILLCELL_X32 FILLER_26_449 ();
 FILLCELL_X32 FILLER_26_481 ();
 FILLCELL_X32 FILLER_26_513 ();
 FILLCELL_X32 FILLER_26_545 ();
 FILLCELL_X32 FILLER_26_577 ();
 FILLCELL_X16 FILLER_26_609 ();
 FILLCELL_X4 FILLER_26_625 ();
 FILLCELL_X2 FILLER_26_629 ();
 FILLCELL_X32 FILLER_26_632 ();
 FILLCELL_X32 FILLER_26_664 ();
 FILLCELL_X32 FILLER_26_696 ();
 FILLCELL_X32 FILLER_26_728 ();
 FILLCELL_X32 FILLER_26_760 ();
 FILLCELL_X32 FILLER_26_792 ();
 FILLCELL_X32 FILLER_26_824 ();
 FILLCELL_X32 FILLER_26_856 ();
 FILLCELL_X32 FILLER_26_888 ();
 FILLCELL_X32 FILLER_26_920 ();
 FILLCELL_X32 FILLER_26_952 ();
 FILLCELL_X32 FILLER_26_984 ();
 FILLCELL_X32 FILLER_26_1016 ();
 FILLCELL_X32 FILLER_26_1048 ();
 FILLCELL_X32 FILLER_26_1080 ();
 FILLCELL_X32 FILLER_26_1112 ();
 FILLCELL_X32 FILLER_26_1144 ();
 FILLCELL_X32 FILLER_26_1176 ();
 FILLCELL_X32 FILLER_26_1208 ();
 FILLCELL_X32 FILLER_26_1240 ();
 FILLCELL_X32 FILLER_26_1272 ();
 FILLCELL_X32 FILLER_26_1304 ();
 FILLCELL_X32 FILLER_26_1336 ();
 FILLCELL_X32 FILLER_26_1368 ();
 FILLCELL_X32 FILLER_26_1400 ();
 FILLCELL_X32 FILLER_26_1432 ();
 FILLCELL_X32 FILLER_26_1464 ();
 FILLCELL_X32 FILLER_26_1496 ();
 FILLCELL_X32 FILLER_26_1528 ();
 FILLCELL_X32 FILLER_26_1560 ();
 FILLCELL_X32 FILLER_26_1592 ();
 FILLCELL_X32 FILLER_26_1624 ();
 FILLCELL_X32 FILLER_26_1656 ();
 FILLCELL_X32 FILLER_26_1688 ();
 FILLCELL_X32 FILLER_26_1720 ();
 FILLCELL_X32 FILLER_26_1752 ();
 FILLCELL_X32 FILLER_26_1784 ();
 FILLCELL_X32 FILLER_26_1816 ();
 FILLCELL_X32 FILLER_26_1848 ();
 FILLCELL_X8 FILLER_26_1880 ();
 FILLCELL_X4 FILLER_26_1888 ();
 FILLCELL_X2 FILLER_26_1892 ();
 FILLCELL_X32 FILLER_26_1895 ();
 FILLCELL_X32 FILLER_26_1927 ();
 FILLCELL_X32 FILLER_26_1959 ();
 FILLCELL_X32 FILLER_26_1991 ();
 FILLCELL_X32 FILLER_26_2023 ();
 FILLCELL_X32 FILLER_26_2055 ();
 FILLCELL_X32 FILLER_26_2087 ();
 FILLCELL_X32 FILLER_26_2119 ();
 FILLCELL_X32 FILLER_26_2151 ();
 FILLCELL_X32 FILLER_26_2183 ();
 FILLCELL_X32 FILLER_26_2215 ();
 FILLCELL_X32 FILLER_26_2247 ();
 FILLCELL_X32 FILLER_26_2279 ();
 FILLCELL_X32 FILLER_26_2311 ();
 FILLCELL_X32 FILLER_26_2343 ();
 FILLCELL_X32 FILLER_26_2375 ();
 FILLCELL_X32 FILLER_26_2407 ();
 FILLCELL_X32 FILLER_26_2439 ();
 FILLCELL_X32 FILLER_26_2471 ();
 FILLCELL_X32 FILLER_26_2503 ();
 FILLCELL_X32 FILLER_26_2535 ();
 FILLCELL_X32 FILLER_26_2567 ();
 FILLCELL_X32 FILLER_26_2599 ();
 FILLCELL_X32 FILLER_26_2631 ();
 FILLCELL_X32 FILLER_26_2663 ();
 FILLCELL_X32 FILLER_26_2695 ();
 FILLCELL_X32 FILLER_26_2727 ();
 FILLCELL_X32 FILLER_26_2759 ();
 FILLCELL_X32 FILLER_26_2791 ();
 FILLCELL_X32 FILLER_26_2823 ();
 FILLCELL_X32 FILLER_26_2855 ();
 FILLCELL_X32 FILLER_26_2887 ();
 FILLCELL_X32 FILLER_26_2919 ();
 FILLCELL_X32 FILLER_26_2951 ();
 FILLCELL_X32 FILLER_26_2983 ();
 FILLCELL_X32 FILLER_26_3015 ();
 FILLCELL_X32 FILLER_26_3047 ();
 FILLCELL_X32 FILLER_26_3079 ();
 FILLCELL_X32 FILLER_26_3111 ();
 FILLCELL_X8 FILLER_26_3143 ();
 FILLCELL_X4 FILLER_26_3151 ();
 FILLCELL_X2 FILLER_26_3155 ();
 FILLCELL_X32 FILLER_26_3158 ();
 FILLCELL_X32 FILLER_26_3190 ();
 FILLCELL_X32 FILLER_26_3222 ();
 FILLCELL_X32 FILLER_26_3254 ();
 FILLCELL_X32 FILLER_26_3286 ();
 FILLCELL_X32 FILLER_26_3318 ();
 FILLCELL_X32 FILLER_26_3350 ();
 FILLCELL_X32 FILLER_26_3382 ();
 FILLCELL_X32 FILLER_26_3414 ();
 FILLCELL_X32 FILLER_26_3446 ();
 FILLCELL_X32 FILLER_26_3478 ();
 FILLCELL_X32 FILLER_26_3510 ();
 FILLCELL_X32 FILLER_26_3542 ();
 FILLCELL_X32 FILLER_26_3574 ();
 FILLCELL_X32 FILLER_26_3606 ();
 FILLCELL_X32 FILLER_26_3638 ();
 FILLCELL_X32 FILLER_26_3670 ();
 FILLCELL_X32 FILLER_26_3702 ();
 FILLCELL_X4 FILLER_26_3734 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X32 FILLER_27_225 ();
 FILLCELL_X32 FILLER_27_257 ();
 FILLCELL_X32 FILLER_27_289 ();
 FILLCELL_X32 FILLER_27_321 ();
 FILLCELL_X32 FILLER_27_353 ();
 FILLCELL_X32 FILLER_27_385 ();
 FILLCELL_X32 FILLER_27_417 ();
 FILLCELL_X32 FILLER_27_449 ();
 FILLCELL_X32 FILLER_27_481 ();
 FILLCELL_X32 FILLER_27_513 ();
 FILLCELL_X32 FILLER_27_545 ();
 FILLCELL_X32 FILLER_27_577 ();
 FILLCELL_X32 FILLER_27_609 ();
 FILLCELL_X32 FILLER_27_641 ();
 FILLCELL_X32 FILLER_27_673 ();
 FILLCELL_X32 FILLER_27_705 ();
 FILLCELL_X32 FILLER_27_737 ();
 FILLCELL_X32 FILLER_27_769 ();
 FILLCELL_X32 FILLER_27_801 ();
 FILLCELL_X32 FILLER_27_833 ();
 FILLCELL_X32 FILLER_27_865 ();
 FILLCELL_X32 FILLER_27_897 ();
 FILLCELL_X32 FILLER_27_929 ();
 FILLCELL_X32 FILLER_27_961 ();
 FILLCELL_X32 FILLER_27_993 ();
 FILLCELL_X32 FILLER_27_1025 ();
 FILLCELL_X32 FILLER_27_1057 ();
 FILLCELL_X32 FILLER_27_1089 ();
 FILLCELL_X32 FILLER_27_1121 ();
 FILLCELL_X32 FILLER_27_1153 ();
 FILLCELL_X32 FILLER_27_1185 ();
 FILLCELL_X32 FILLER_27_1217 ();
 FILLCELL_X8 FILLER_27_1249 ();
 FILLCELL_X4 FILLER_27_1257 ();
 FILLCELL_X2 FILLER_27_1261 ();
 FILLCELL_X32 FILLER_27_1264 ();
 FILLCELL_X32 FILLER_27_1296 ();
 FILLCELL_X32 FILLER_27_1328 ();
 FILLCELL_X32 FILLER_27_1360 ();
 FILLCELL_X32 FILLER_27_1392 ();
 FILLCELL_X32 FILLER_27_1424 ();
 FILLCELL_X32 FILLER_27_1456 ();
 FILLCELL_X32 FILLER_27_1488 ();
 FILLCELL_X32 FILLER_27_1520 ();
 FILLCELL_X32 FILLER_27_1552 ();
 FILLCELL_X32 FILLER_27_1584 ();
 FILLCELL_X32 FILLER_27_1616 ();
 FILLCELL_X32 FILLER_27_1648 ();
 FILLCELL_X32 FILLER_27_1680 ();
 FILLCELL_X32 FILLER_27_1712 ();
 FILLCELL_X32 FILLER_27_1744 ();
 FILLCELL_X32 FILLER_27_1776 ();
 FILLCELL_X32 FILLER_27_1808 ();
 FILLCELL_X32 FILLER_27_1840 ();
 FILLCELL_X32 FILLER_27_1872 ();
 FILLCELL_X32 FILLER_27_1904 ();
 FILLCELL_X32 FILLER_27_1936 ();
 FILLCELL_X32 FILLER_27_1968 ();
 FILLCELL_X32 FILLER_27_2000 ();
 FILLCELL_X32 FILLER_27_2032 ();
 FILLCELL_X32 FILLER_27_2064 ();
 FILLCELL_X32 FILLER_27_2096 ();
 FILLCELL_X32 FILLER_27_2128 ();
 FILLCELL_X32 FILLER_27_2160 ();
 FILLCELL_X32 FILLER_27_2192 ();
 FILLCELL_X32 FILLER_27_2224 ();
 FILLCELL_X32 FILLER_27_2256 ();
 FILLCELL_X32 FILLER_27_2288 ();
 FILLCELL_X32 FILLER_27_2320 ();
 FILLCELL_X32 FILLER_27_2352 ();
 FILLCELL_X32 FILLER_27_2384 ();
 FILLCELL_X32 FILLER_27_2416 ();
 FILLCELL_X32 FILLER_27_2448 ();
 FILLCELL_X32 FILLER_27_2480 ();
 FILLCELL_X8 FILLER_27_2512 ();
 FILLCELL_X4 FILLER_27_2520 ();
 FILLCELL_X2 FILLER_27_2524 ();
 FILLCELL_X32 FILLER_27_2527 ();
 FILLCELL_X32 FILLER_27_2559 ();
 FILLCELL_X32 FILLER_27_2591 ();
 FILLCELL_X32 FILLER_27_2623 ();
 FILLCELL_X32 FILLER_27_2655 ();
 FILLCELL_X32 FILLER_27_2687 ();
 FILLCELL_X32 FILLER_27_2719 ();
 FILLCELL_X32 FILLER_27_2751 ();
 FILLCELL_X32 FILLER_27_2783 ();
 FILLCELL_X32 FILLER_27_2815 ();
 FILLCELL_X32 FILLER_27_2847 ();
 FILLCELL_X32 FILLER_27_2879 ();
 FILLCELL_X32 FILLER_27_2911 ();
 FILLCELL_X32 FILLER_27_2943 ();
 FILLCELL_X32 FILLER_27_2975 ();
 FILLCELL_X32 FILLER_27_3007 ();
 FILLCELL_X32 FILLER_27_3039 ();
 FILLCELL_X32 FILLER_27_3071 ();
 FILLCELL_X32 FILLER_27_3103 ();
 FILLCELL_X32 FILLER_27_3135 ();
 FILLCELL_X32 FILLER_27_3167 ();
 FILLCELL_X32 FILLER_27_3199 ();
 FILLCELL_X32 FILLER_27_3231 ();
 FILLCELL_X32 FILLER_27_3263 ();
 FILLCELL_X32 FILLER_27_3295 ();
 FILLCELL_X32 FILLER_27_3327 ();
 FILLCELL_X32 FILLER_27_3359 ();
 FILLCELL_X32 FILLER_27_3391 ();
 FILLCELL_X32 FILLER_27_3423 ();
 FILLCELL_X32 FILLER_27_3455 ();
 FILLCELL_X32 FILLER_27_3487 ();
 FILLCELL_X32 FILLER_27_3519 ();
 FILLCELL_X32 FILLER_27_3551 ();
 FILLCELL_X32 FILLER_27_3583 ();
 FILLCELL_X32 FILLER_27_3615 ();
 FILLCELL_X32 FILLER_27_3647 ();
 FILLCELL_X32 FILLER_27_3679 ();
 FILLCELL_X16 FILLER_27_3711 ();
 FILLCELL_X8 FILLER_27_3727 ();
 FILLCELL_X2 FILLER_27_3735 ();
 FILLCELL_X1 FILLER_27_3737 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X32 FILLER_28_257 ();
 FILLCELL_X32 FILLER_28_289 ();
 FILLCELL_X32 FILLER_28_321 ();
 FILLCELL_X32 FILLER_28_353 ();
 FILLCELL_X32 FILLER_28_385 ();
 FILLCELL_X32 FILLER_28_417 ();
 FILLCELL_X32 FILLER_28_449 ();
 FILLCELL_X32 FILLER_28_481 ();
 FILLCELL_X32 FILLER_28_513 ();
 FILLCELL_X32 FILLER_28_545 ();
 FILLCELL_X32 FILLER_28_577 ();
 FILLCELL_X16 FILLER_28_609 ();
 FILLCELL_X4 FILLER_28_625 ();
 FILLCELL_X2 FILLER_28_629 ();
 FILLCELL_X32 FILLER_28_632 ();
 FILLCELL_X32 FILLER_28_664 ();
 FILLCELL_X32 FILLER_28_696 ();
 FILLCELL_X32 FILLER_28_728 ();
 FILLCELL_X32 FILLER_28_760 ();
 FILLCELL_X32 FILLER_28_792 ();
 FILLCELL_X32 FILLER_28_824 ();
 FILLCELL_X32 FILLER_28_856 ();
 FILLCELL_X32 FILLER_28_888 ();
 FILLCELL_X32 FILLER_28_920 ();
 FILLCELL_X32 FILLER_28_952 ();
 FILLCELL_X32 FILLER_28_984 ();
 FILLCELL_X32 FILLER_28_1016 ();
 FILLCELL_X32 FILLER_28_1048 ();
 FILLCELL_X32 FILLER_28_1080 ();
 FILLCELL_X32 FILLER_28_1112 ();
 FILLCELL_X32 FILLER_28_1144 ();
 FILLCELL_X32 FILLER_28_1176 ();
 FILLCELL_X32 FILLER_28_1208 ();
 FILLCELL_X32 FILLER_28_1240 ();
 FILLCELL_X32 FILLER_28_1272 ();
 FILLCELL_X32 FILLER_28_1304 ();
 FILLCELL_X32 FILLER_28_1336 ();
 FILLCELL_X32 FILLER_28_1368 ();
 FILLCELL_X32 FILLER_28_1400 ();
 FILLCELL_X32 FILLER_28_1432 ();
 FILLCELL_X32 FILLER_28_1464 ();
 FILLCELL_X32 FILLER_28_1496 ();
 FILLCELL_X32 FILLER_28_1528 ();
 FILLCELL_X32 FILLER_28_1560 ();
 FILLCELL_X32 FILLER_28_1592 ();
 FILLCELL_X32 FILLER_28_1624 ();
 FILLCELL_X32 FILLER_28_1656 ();
 FILLCELL_X32 FILLER_28_1688 ();
 FILLCELL_X32 FILLER_28_1720 ();
 FILLCELL_X32 FILLER_28_1752 ();
 FILLCELL_X32 FILLER_28_1784 ();
 FILLCELL_X32 FILLER_28_1816 ();
 FILLCELL_X32 FILLER_28_1848 ();
 FILLCELL_X8 FILLER_28_1880 ();
 FILLCELL_X4 FILLER_28_1888 ();
 FILLCELL_X2 FILLER_28_1892 ();
 FILLCELL_X32 FILLER_28_1895 ();
 FILLCELL_X32 FILLER_28_1927 ();
 FILLCELL_X32 FILLER_28_1959 ();
 FILLCELL_X32 FILLER_28_1991 ();
 FILLCELL_X32 FILLER_28_2023 ();
 FILLCELL_X32 FILLER_28_2055 ();
 FILLCELL_X32 FILLER_28_2087 ();
 FILLCELL_X32 FILLER_28_2119 ();
 FILLCELL_X32 FILLER_28_2151 ();
 FILLCELL_X32 FILLER_28_2183 ();
 FILLCELL_X32 FILLER_28_2215 ();
 FILLCELL_X32 FILLER_28_2247 ();
 FILLCELL_X32 FILLER_28_2279 ();
 FILLCELL_X32 FILLER_28_2311 ();
 FILLCELL_X32 FILLER_28_2343 ();
 FILLCELL_X32 FILLER_28_2375 ();
 FILLCELL_X32 FILLER_28_2407 ();
 FILLCELL_X32 FILLER_28_2439 ();
 FILLCELL_X32 FILLER_28_2471 ();
 FILLCELL_X32 FILLER_28_2503 ();
 FILLCELL_X32 FILLER_28_2535 ();
 FILLCELL_X32 FILLER_28_2567 ();
 FILLCELL_X32 FILLER_28_2599 ();
 FILLCELL_X32 FILLER_28_2631 ();
 FILLCELL_X32 FILLER_28_2663 ();
 FILLCELL_X32 FILLER_28_2695 ();
 FILLCELL_X32 FILLER_28_2727 ();
 FILLCELL_X32 FILLER_28_2759 ();
 FILLCELL_X32 FILLER_28_2791 ();
 FILLCELL_X32 FILLER_28_2823 ();
 FILLCELL_X32 FILLER_28_2855 ();
 FILLCELL_X32 FILLER_28_2887 ();
 FILLCELL_X32 FILLER_28_2919 ();
 FILLCELL_X32 FILLER_28_2951 ();
 FILLCELL_X32 FILLER_28_2983 ();
 FILLCELL_X32 FILLER_28_3015 ();
 FILLCELL_X32 FILLER_28_3047 ();
 FILLCELL_X32 FILLER_28_3079 ();
 FILLCELL_X32 FILLER_28_3111 ();
 FILLCELL_X8 FILLER_28_3143 ();
 FILLCELL_X4 FILLER_28_3151 ();
 FILLCELL_X2 FILLER_28_3155 ();
 FILLCELL_X32 FILLER_28_3158 ();
 FILLCELL_X32 FILLER_28_3190 ();
 FILLCELL_X32 FILLER_28_3222 ();
 FILLCELL_X32 FILLER_28_3254 ();
 FILLCELL_X32 FILLER_28_3286 ();
 FILLCELL_X32 FILLER_28_3318 ();
 FILLCELL_X32 FILLER_28_3350 ();
 FILLCELL_X32 FILLER_28_3382 ();
 FILLCELL_X32 FILLER_28_3414 ();
 FILLCELL_X32 FILLER_28_3446 ();
 FILLCELL_X32 FILLER_28_3478 ();
 FILLCELL_X32 FILLER_28_3510 ();
 FILLCELL_X32 FILLER_28_3542 ();
 FILLCELL_X32 FILLER_28_3574 ();
 FILLCELL_X32 FILLER_28_3606 ();
 FILLCELL_X32 FILLER_28_3638 ();
 FILLCELL_X32 FILLER_28_3670 ();
 FILLCELL_X32 FILLER_28_3702 ();
 FILLCELL_X4 FILLER_28_3734 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X32 FILLER_29_257 ();
 FILLCELL_X32 FILLER_29_289 ();
 FILLCELL_X32 FILLER_29_321 ();
 FILLCELL_X32 FILLER_29_353 ();
 FILLCELL_X32 FILLER_29_385 ();
 FILLCELL_X32 FILLER_29_417 ();
 FILLCELL_X32 FILLER_29_449 ();
 FILLCELL_X32 FILLER_29_481 ();
 FILLCELL_X32 FILLER_29_513 ();
 FILLCELL_X32 FILLER_29_545 ();
 FILLCELL_X32 FILLER_29_577 ();
 FILLCELL_X32 FILLER_29_609 ();
 FILLCELL_X32 FILLER_29_641 ();
 FILLCELL_X32 FILLER_29_673 ();
 FILLCELL_X32 FILLER_29_705 ();
 FILLCELL_X32 FILLER_29_737 ();
 FILLCELL_X32 FILLER_29_769 ();
 FILLCELL_X32 FILLER_29_801 ();
 FILLCELL_X32 FILLER_29_833 ();
 FILLCELL_X32 FILLER_29_865 ();
 FILLCELL_X32 FILLER_29_897 ();
 FILLCELL_X32 FILLER_29_929 ();
 FILLCELL_X32 FILLER_29_961 ();
 FILLCELL_X32 FILLER_29_993 ();
 FILLCELL_X32 FILLER_29_1025 ();
 FILLCELL_X32 FILLER_29_1057 ();
 FILLCELL_X32 FILLER_29_1089 ();
 FILLCELL_X32 FILLER_29_1121 ();
 FILLCELL_X32 FILLER_29_1153 ();
 FILLCELL_X32 FILLER_29_1185 ();
 FILLCELL_X32 FILLER_29_1217 ();
 FILLCELL_X8 FILLER_29_1249 ();
 FILLCELL_X4 FILLER_29_1257 ();
 FILLCELL_X2 FILLER_29_1261 ();
 FILLCELL_X32 FILLER_29_1264 ();
 FILLCELL_X32 FILLER_29_1296 ();
 FILLCELL_X32 FILLER_29_1328 ();
 FILLCELL_X32 FILLER_29_1360 ();
 FILLCELL_X32 FILLER_29_1392 ();
 FILLCELL_X32 FILLER_29_1424 ();
 FILLCELL_X32 FILLER_29_1456 ();
 FILLCELL_X32 FILLER_29_1488 ();
 FILLCELL_X32 FILLER_29_1520 ();
 FILLCELL_X32 FILLER_29_1552 ();
 FILLCELL_X32 FILLER_29_1584 ();
 FILLCELL_X32 FILLER_29_1616 ();
 FILLCELL_X32 FILLER_29_1648 ();
 FILLCELL_X32 FILLER_29_1680 ();
 FILLCELL_X32 FILLER_29_1712 ();
 FILLCELL_X32 FILLER_29_1744 ();
 FILLCELL_X32 FILLER_29_1776 ();
 FILLCELL_X32 FILLER_29_1808 ();
 FILLCELL_X32 FILLER_29_1840 ();
 FILLCELL_X32 FILLER_29_1872 ();
 FILLCELL_X32 FILLER_29_1904 ();
 FILLCELL_X32 FILLER_29_1936 ();
 FILLCELL_X32 FILLER_29_1968 ();
 FILLCELL_X32 FILLER_29_2000 ();
 FILLCELL_X32 FILLER_29_2032 ();
 FILLCELL_X32 FILLER_29_2064 ();
 FILLCELL_X32 FILLER_29_2096 ();
 FILLCELL_X32 FILLER_29_2128 ();
 FILLCELL_X32 FILLER_29_2160 ();
 FILLCELL_X32 FILLER_29_2192 ();
 FILLCELL_X32 FILLER_29_2224 ();
 FILLCELL_X32 FILLER_29_2256 ();
 FILLCELL_X32 FILLER_29_2288 ();
 FILLCELL_X32 FILLER_29_2320 ();
 FILLCELL_X32 FILLER_29_2352 ();
 FILLCELL_X32 FILLER_29_2384 ();
 FILLCELL_X32 FILLER_29_2416 ();
 FILLCELL_X32 FILLER_29_2448 ();
 FILLCELL_X32 FILLER_29_2480 ();
 FILLCELL_X8 FILLER_29_2512 ();
 FILLCELL_X4 FILLER_29_2520 ();
 FILLCELL_X2 FILLER_29_2524 ();
 FILLCELL_X32 FILLER_29_2527 ();
 FILLCELL_X32 FILLER_29_2559 ();
 FILLCELL_X32 FILLER_29_2591 ();
 FILLCELL_X32 FILLER_29_2623 ();
 FILLCELL_X32 FILLER_29_2655 ();
 FILLCELL_X32 FILLER_29_2687 ();
 FILLCELL_X32 FILLER_29_2719 ();
 FILLCELL_X32 FILLER_29_2751 ();
 FILLCELL_X32 FILLER_29_2783 ();
 FILLCELL_X32 FILLER_29_2815 ();
 FILLCELL_X32 FILLER_29_2847 ();
 FILLCELL_X32 FILLER_29_2879 ();
 FILLCELL_X32 FILLER_29_2911 ();
 FILLCELL_X32 FILLER_29_2943 ();
 FILLCELL_X32 FILLER_29_2975 ();
 FILLCELL_X32 FILLER_29_3007 ();
 FILLCELL_X32 FILLER_29_3039 ();
 FILLCELL_X32 FILLER_29_3071 ();
 FILLCELL_X32 FILLER_29_3103 ();
 FILLCELL_X32 FILLER_29_3135 ();
 FILLCELL_X32 FILLER_29_3167 ();
 FILLCELL_X32 FILLER_29_3199 ();
 FILLCELL_X32 FILLER_29_3231 ();
 FILLCELL_X32 FILLER_29_3263 ();
 FILLCELL_X32 FILLER_29_3295 ();
 FILLCELL_X32 FILLER_29_3327 ();
 FILLCELL_X32 FILLER_29_3359 ();
 FILLCELL_X32 FILLER_29_3391 ();
 FILLCELL_X32 FILLER_29_3423 ();
 FILLCELL_X32 FILLER_29_3455 ();
 FILLCELL_X32 FILLER_29_3487 ();
 FILLCELL_X32 FILLER_29_3519 ();
 FILLCELL_X32 FILLER_29_3551 ();
 FILLCELL_X32 FILLER_29_3583 ();
 FILLCELL_X32 FILLER_29_3615 ();
 FILLCELL_X32 FILLER_29_3647 ();
 FILLCELL_X32 FILLER_29_3679 ();
 FILLCELL_X16 FILLER_29_3711 ();
 FILLCELL_X8 FILLER_29_3727 ();
 FILLCELL_X2 FILLER_29_3735 ();
 FILLCELL_X1 FILLER_29_3737 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X32 FILLER_30_257 ();
 FILLCELL_X32 FILLER_30_289 ();
 FILLCELL_X32 FILLER_30_321 ();
 FILLCELL_X32 FILLER_30_353 ();
 FILLCELL_X32 FILLER_30_385 ();
 FILLCELL_X32 FILLER_30_417 ();
 FILLCELL_X32 FILLER_30_449 ();
 FILLCELL_X32 FILLER_30_481 ();
 FILLCELL_X32 FILLER_30_513 ();
 FILLCELL_X32 FILLER_30_545 ();
 FILLCELL_X32 FILLER_30_577 ();
 FILLCELL_X16 FILLER_30_609 ();
 FILLCELL_X4 FILLER_30_625 ();
 FILLCELL_X2 FILLER_30_629 ();
 FILLCELL_X32 FILLER_30_632 ();
 FILLCELL_X32 FILLER_30_664 ();
 FILLCELL_X32 FILLER_30_696 ();
 FILLCELL_X32 FILLER_30_728 ();
 FILLCELL_X32 FILLER_30_760 ();
 FILLCELL_X32 FILLER_30_792 ();
 FILLCELL_X32 FILLER_30_824 ();
 FILLCELL_X32 FILLER_30_856 ();
 FILLCELL_X32 FILLER_30_888 ();
 FILLCELL_X32 FILLER_30_920 ();
 FILLCELL_X32 FILLER_30_952 ();
 FILLCELL_X32 FILLER_30_984 ();
 FILLCELL_X32 FILLER_30_1016 ();
 FILLCELL_X32 FILLER_30_1048 ();
 FILLCELL_X32 FILLER_30_1080 ();
 FILLCELL_X32 FILLER_30_1112 ();
 FILLCELL_X32 FILLER_30_1144 ();
 FILLCELL_X32 FILLER_30_1176 ();
 FILLCELL_X32 FILLER_30_1208 ();
 FILLCELL_X32 FILLER_30_1240 ();
 FILLCELL_X32 FILLER_30_1272 ();
 FILLCELL_X32 FILLER_30_1304 ();
 FILLCELL_X32 FILLER_30_1336 ();
 FILLCELL_X32 FILLER_30_1368 ();
 FILLCELL_X32 FILLER_30_1400 ();
 FILLCELL_X32 FILLER_30_1432 ();
 FILLCELL_X32 FILLER_30_1464 ();
 FILLCELL_X32 FILLER_30_1496 ();
 FILLCELL_X32 FILLER_30_1528 ();
 FILLCELL_X32 FILLER_30_1560 ();
 FILLCELL_X32 FILLER_30_1592 ();
 FILLCELL_X32 FILLER_30_1624 ();
 FILLCELL_X32 FILLER_30_1656 ();
 FILLCELL_X32 FILLER_30_1688 ();
 FILLCELL_X32 FILLER_30_1720 ();
 FILLCELL_X32 FILLER_30_1752 ();
 FILLCELL_X32 FILLER_30_1784 ();
 FILLCELL_X32 FILLER_30_1816 ();
 FILLCELL_X32 FILLER_30_1848 ();
 FILLCELL_X8 FILLER_30_1880 ();
 FILLCELL_X4 FILLER_30_1888 ();
 FILLCELL_X2 FILLER_30_1892 ();
 FILLCELL_X32 FILLER_30_1895 ();
 FILLCELL_X32 FILLER_30_1927 ();
 FILLCELL_X32 FILLER_30_1959 ();
 FILLCELL_X32 FILLER_30_1991 ();
 FILLCELL_X32 FILLER_30_2023 ();
 FILLCELL_X32 FILLER_30_2055 ();
 FILLCELL_X32 FILLER_30_2087 ();
 FILLCELL_X32 FILLER_30_2119 ();
 FILLCELL_X32 FILLER_30_2151 ();
 FILLCELL_X32 FILLER_30_2183 ();
 FILLCELL_X32 FILLER_30_2215 ();
 FILLCELL_X32 FILLER_30_2247 ();
 FILLCELL_X32 FILLER_30_2279 ();
 FILLCELL_X32 FILLER_30_2311 ();
 FILLCELL_X32 FILLER_30_2343 ();
 FILLCELL_X32 FILLER_30_2375 ();
 FILLCELL_X32 FILLER_30_2407 ();
 FILLCELL_X32 FILLER_30_2439 ();
 FILLCELL_X32 FILLER_30_2471 ();
 FILLCELL_X32 FILLER_30_2503 ();
 FILLCELL_X32 FILLER_30_2535 ();
 FILLCELL_X32 FILLER_30_2567 ();
 FILLCELL_X32 FILLER_30_2599 ();
 FILLCELL_X32 FILLER_30_2631 ();
 FILLCELL_X32 FILLER_30_2663 ();
 FILLCELL_X32 FILLER_30_2695 ();
 FILLCELL_X32 FILLER_30_2727 ();
 FILLCELL_X32 FILLER_30_2759 ();
 FILLCELL_X32 FILLER_30_2791 ();
 FILLCELL_X32 FILLER_30_2823 ();
 FILLCELL_X32 FILLER_30_2855 ();
 FILLCELL_X32 FILLER_30_2887 ();
 FILLCELL_X32 FILLER_30_2919 ();
 FILLCELL_X32 FILLER_30_2951 ();
 FILLCELL_X32 FILLER_30_2983 ();
 FILLCELL_X32 FILLER_30_3015 ();
 FILLCELL_X32 FILLER_30_3047 ();
 FILLCELL_X32 FILLER_30_3079 ();
 FILLCELL_X32 FILLER_30_3111 ();
 FILLCELL_X8 FILLER_30_3143 ();
 FILLCELL_X4 FILLER_30_3151 ();
 FILLCELL_X2 FILLER_30_3155 ();
 FILLCELL_X32 FILLER_30_3158 ();
 FILLCELL_X32 FILLER_30_3190 ();
 FILLCELL_X32 FILLER_30_3222 ();
 FILLCELL_X32 FILLER_30_3254 ();
 FILLCELL_X32 FILLER_30_3286 ();
 FILLCELL_X32 FILLER_30_3318 ();
 FILLCELL_X32 FILLER_30_3350 ();
 FILLCELL_X32 FILLER_30_3382 ();
 FILLCELL_X32 FILLER_30_3414 ();
 FILLCELL_X32 FILLER_30_3446 ();
 FILLCELL_X32 FILLER_30_3478 ();
 FILLCELL_X32 FILLER_30_3510 ();
 FILLCELL_X32 FILLER_30_3542 ();
 FILLCELL_X32 FILLER_30_3574 ();
 FILLCELL_X32 FILLER_30_3606 ();
 FILLCELL_X32 FILLER_30_3638 ();
 FILLCELL_X32 FILLER_30_3670 ();
 FILLCELL_X32 FILLER_30_3702 ();
 FILLCELL_X4 FILLER_30_3734 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X32 FILLER_31_257 ();
 FILLCELL_X32 FILLER_31_289 ();
 FILLCELL_X32 FILLER_31_321 ();
 FILLCELL_X32 FILLER_31_353 ();
 FILLCELL_X32 FILLER_31_385 ();
 FILLCELL_X32 FILLER_31_417 ();
 FILLCELL_X32 FILLER_31_449 ();
 FILLCELL_X32 FILLER_31_481 ();
 FILLCELL_X32 FILLER_31_513 ();
 FILLCELL_X32 FILLER_31_545 ();
 FILLCELL_X32 FILLER_31_577 ();
 FILLCELL_X32 FILLER_31_609 ();
 FILLCELL_X32 FILLER_31_641 ();
 FILLCELL_X32 FILLER_31_673 ();
 FILLCELL_X32 FILLER_31_705 ();
 FILLCELL_X32 FILLER_31_737 ();
 FILLCELL_X32 FILLER_31_769 ();
 FILLCELL_X32 FILLER_31_801 ();
 FILLCELL_X32 FILLER_31_833 ();
 FILLCELL_X32 FILLER_31_865 ();
 FILLCELL_X32 FILLER_31_897 ();
 FILLCELL_X32 FILLER_31_929 ();
 FILLCELL_X32 FILLER_31_961 ();
 FILLCELL_X32 FILLER_31_993 ();
 FILLCELL_X32 FILLER_31_1025 ();
 FILLCELL_X32 FILLER_31_1057 ();
 FILLCELL_X32 FILLER_31_1089 ();
 FILLCELL_X32 FILLER_31_1121 ();
 FILLCELL_X32 FILLER_31_1153 ();
 FILLCELL_X32 FILLER_31_1185 ();
 FILLCELL_X32 FILLER_31_1217 ();
 FILLCELL_X8 FILLER_31_1249 ();
 FILLCELL_X4 FILLER_31_1257 ();
 FILLCELL_X2 FILLER_31_1261 ();
 FILLCELL_X32 FILLER_31_1264 ();
 FILLCELL_X32 FILLER_31_1296 ();
 FILLCELL_X32 FILLER_31_1328 ();
 FILLCELL_X32 FILLER_31_1360 ();
 FILLCELL_X32 FILLER_31_1392 ();
 FILLCELL_X32 FILLER_31_1424 ();
 FILLCELL_X32 FILLER_31_1456 ();
 FILLCELL_X32 FILLER_31_1488 ();
 FILLCELL_X32 FILLER_31_1520 ();
 FILLCELL_X32 FILLER_31_1552 ();
 FILLCELL_X32 FILLER_31_1584 ();
 FILLCELL_X32 FILLER_31_1616 ();
 FILLCELL_X32 FILLER_31_1648 ();
 FILLCELL_X32 FILLER_31_1680 ();
 FILLCELL_X32 FILLER_31_1712 ();
 FILLCELL_X32 FILLER_31_1744 ();
 FILLCELL_X32 FILLER_31_1776 ();
 FILLCELL_X32 FILLER_31_1808 ();
 FILLCELL_X32 FILLER_31_1840 ();
 FILLCELL_X32 FILLER_31_1872 ();
 FILLCELL_X32 FILLER_31_1904 ();
 FILLCELL_X32 FILLER_31_1936 ();
 FILLCELL_X32 FILLER_31_1968 ();
 FILLCELL_X32 FILLER_31_2000 ();
 FILLCELL_X32 FILLER_31_2032 ();
 FILLCELL_X32 FILLER_31_2064 ();
 FILLCELL_X32 FILLER_31_2096 ();
 FILLCELL_X32 FILLER_31_2128 ();
 FILLCELL_X32 FILLER_31_2160 ();
 FILLCELL_X32 FILLER_31_2192 ();
 FILLCELL_X32 FILLER_31_2224 ();
 FILLCELL_X32 FILLER_31_2256 ();
 FILLCELL_X32 FILLER_31_2288 ();
 FILLCELL_X32 FILLER_31_2320 ();
 FILLCELL_X32 FILLER_31_2352 ();
 FILLCELL_X32 FILLER_31_2384 ();
 FILLCELL_X32 FILLER_31_2416 ();
 FILLCELL_X32 FILLER_31_2448 ();
 FILLCELL_X32 FILLER_31_2480 ();
 FILLCELL_X8 FILLER_31_2512 ();
 FILLCELL_X4 FILLER_31_2520 ();
 FILLCELL_X2 FILLER_31_2524 ();
 FILLCELL_X32 FILLER_31_2527 ();
 FILLCELL_X32 FILLER_31_2559 ();
 FILLCELL_X32 FILLER_31_2591 ();
 FILLCELL_X32 FILLER_31_2623 ();
 FILLCELL_X32 FILLER_31_2655 ();
 FILLCELL_X32 FILLER_31_2687 ();
 FILLCELL_X32 FILLER_31_2719 ();
 FILLCELL_X32 FILLER_31_2751 ();
 FILLCELL_X32 FILLER_31_2783 ();
 FILLCELL_X32 FILLER_31_2815 ();
 FILLCELL_X32 FILLER_31_2847 ();
 FILLCELL_X32 FILLER_31_2879 ();
 FILLCELL_X32 FILLER_31_2911 ();
 FILLCELL_X32 FILLER_31_2943 ();
 FILLCELL_X32 FILLER_31_2975 ();
 FILLCELL_X32 FILLER_31_3007 ();
 FILLCELL_X32 FILLER_31_3039 ();
 FILLCELL_X32 FILLER_31_3071 ();
 FILLCELL_X32 FILLER_31_3103 ();
 FILLCELL_X32 FILLER_31_3135 ();
 FILLCELL_X32 FILLER_31_3167 ();
 FILLCELL_X32 FILLER_31_3199 ();
 FILLCELL_X32 FILLER_31_3231 ();
 FILLCELL_X32 FILLER_31_3263 ();
 FILLCELL_X32 FILLER_31_3295 ();
 FILLCELL_X32 FILLER_31_3327 ();
 FILLCELL_X32 FILLER_31_3359 ();
 FILLCELL_X32 FILLER_31_3391 ();
 FILLCELL_X32 FILLER_31_3423 ();
 FILLCELL_X32 FILLER_31_3455 ();
 FILLCELL_X32 FILLER_31_3487 ();
 FILLCELL_X32 FILLER_31_3519 ();
 FILLCELL_X32 FILLER_31_3551 ();
 FILLCELL_X32 FILLER_31_3583 ();
 FILLCELL_X32 FILLER_31_3615 ();
 FILLCELL_X32 FILLER_31_3647 ();
 FILLCELL_X32 FILLER_31_3679 ();
 FILLCELL_X16 FILLER_31_3711 ();
 FILLCELL_X8 FILLER_31_3727 ();
 FILLCELL_X2 FILLER_31_3735 ();
 FILLCELL_X1 FILLER_31_3737 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X32 FILLER_32_289 ();
 FILLCELL_X32 FILLER_32_321 ();
 FILLCELL_X32 FILLER_32_353 ();
 FILLCELL_X32 FILLER_32_385 ();
 FILLCELL_X32 FILLER_32_417 ();
 FILLCELL_X32 FILLER_32_449 ();
 FILLCELL_X32 FILLER_32_481 ();
 FILLCELL_X32 FILLER_32_513 ();
 FILLCELL_X32 FILLER_32_545 ();
 FILLCELL_X32 FILLER_32_577 ();
 FILLCELL_X16 FILLER_32_609 ();
 FILLCELL_X4 FILLER_32_625 ();
 FILLCELL_X2 FILLER_32_629 ();
 FILLCELL_X32 FILLER_32_632 ();
 FILLCELL_X32 FILLER_32_664 ();
 FILLCELL_X32 FILLER_32_696 ();
 FILLCELL_X32 FILLER_32_728 ();
 FILLCELL_X32 FILLER_32_760 ();
 FILLCELL_X32 FILLER_32_792 ();
 FILLCELL_X32 FILLER_32_824 ();
 FILLCELL_X32 FILLER_32_856 ();
 FILLCELL_X32 FILLER_32_888 ();
 FILLCELL_X32 FILLER_32_920 ();
 FILLCELL_X32 FILLER_32_952 ();
 FILLCELL_X32 FILLER_32_984 ();
 FILLCELL_X32 FILLER_32_1016 ();
 FILLCELL_X32 FILLER_32_1048 ();
 FILLCELL_X32 FILLER_32_1080 ();
 FILLCELL_X32 FILLER_32_1112 ();
 FILLCELL_X32 FILLER_32_1144 ();
 FILLCELL_X32 FILLER_32_1176 ();
 FILLCELL_X32 FILLER_32_1208 ();
 FILLCELL_X32 FILLER_32_1240 ();
 FILLCELL_X32 FILLER_32_1272 ();
 FILLCELL_X32 FILLER_32_1304 ();
 FILLCELL_X32 FILLER_32_1336 ();
 FILLCELL_X32 FILLER_32_1368 ();
 FILLCELL_X32 FILLER_32_1400 ();
 FILLCELL_X32 FILLER_32_1432 ();
 FILLCELL_X32 FILLER_32_1464 ();
 FILLCELL_X32 FILLER_32_1496 ();
 FILLCELL_X32 FILLER_32_1528 ();
 FILLCELL_X32 FILLER_32_1560 ();
 FILLCELL_X32 FILLER_32_1592 ();
 FILLCELL_X32 FILLER_32_1624 ();
 FILLCELL_X32 FILLER_32_1656 ();
 FILLCELL_X32 FILLER_32_1688 ();
 FILLCELL_X32 FILLER_32_1720 ();
 FILLCELL_X32 FILLER_32_1752 ();
 FILLCELL_X32 FILLER_32_1784 ();
 FILLCELL_X32 FILLER_32_1816 ();
 FILLCELL_X32 FILLER_32_1848 ();
 FILLCELL_X8 FILLER_32_1880 ();
 FILLCELL_X4 FILLER_32_1888 ();
 FILLCELL_X2 FILLER_32_1892 ();
 FILLCELL_X32 FILLER_32_1895 ();
 FILLCELL_X32 FILLER_32_1927 ();
 FILLCELL_X32 FILLER_32_1959 ();
 FILLCELL_X32 FILLER_32_1991 ();
 FILLCELL_X32 FILLER_32_2023 ();
 FILLCELL_X32 FILLER_32_2055 ();
 FILLCELL_X32 FILLER_32_2087 ();
 FILLCELL_X32 FILLER_32_2119 ();
 FILLCELL_X32 FILLER_32_2151 ();
 FILLCELL_X32 FILLER_32_2183 ();
 FILLCELL_X32 FILLER_32_2215 ();
 FILLCELL_X32 FILLER_32_2247 ();
 FILLCELL_X32 FILLER_32_2279 ();
 FILLCELL_X32 FILLER_32_2311 ();
 FILLCELL_X32 FILLER_32_2343 ();
 FILLCELL_X32 FILLER_32_2375 ();
 FILLCELL_X32 FILLER_32_2407 ();
 FILLCELL_X32 FILLER_32_2439 ();
 FILLCELL_X32 FILLER_32_2471 ();
 FILLCELL_X32 FILLER_32_2503 ();
 FILLCELL_X32 FILLER_32_2535 ();
 FILLCELL_X32 FILLER_32_2567 ();
 FILLCELL_X32 FILLER_32_2599 ();
 FILLCELL_X32 FILLER_32_2631 ();
 FILLCELL_X32 FILLER_32_2663 ();
 FILLCELL_X32 FILLER_32_2695 ();
 FILLCELL_X32 FILLER_32_2727 ();
 FILLCELL_X32 FILLER_32_2759 ();
 FILLCELL_X32 FILLER_32_2791 ();
 FILLCELL_X32 FILLER_32_2823 ();
 FILLCELL_X32 FILLER_32_2855 ();
 FILLCELL_X32 FILLER_32_2887 ();
 FILLCELL_X32 FILLER_32_2919 ();
 FILLCELL_X32 FILLER_32_2951 ();
 FILLCELL_X32 FILLER_32_2983 ();
 FILLCELL_X32 FILLER_32_3015 ();
 FILLCELL_X32 FILLER_32_3047 ();
 FILLCELL_X32 FILLER_32_3079 ();
 FILLCELL_X32 FILLER_32_3111 ();
 FILLCELL_X8 FILLER_32_3143 ();
 FILLCELL_X4 FILLER_32_3151 ();
 FILLCELL_X2 FILLER_32_3155 ();
 FILLCELL_X32 FILLER_32_3158 ();
 FILLCELL_X32 FILLER_32_3190 ();
 FILLCELL_X32 FILLER_32_3222 ();
 FILLCELL_X32 FILLER_32_3254 ();
 FILLCELL_X32 FILLER_32_3286 ();
 FILLCELL_X32 FILLER_32_3318 ();
 FILLCELL_X32 FILLER_32_3350 ();
 FILLCELL_X32 FILLER_32_3382 ();
 FILLCELL_X32 FILLER_32_3414 ();
 FILLCELL_X32 FILLER_32_3446 ();
 FILLCELL_X32 FILLER_32_3478 ();
 FILLCELL_X32 FILLER_32_3510 ();
 FILLCELL_X32 FILLER_32_3542 ();
 FILLCELL_X32 FILLER_32_3574 ();
 FILLCELL_X32 FILLER_32_3606 ();
 FILLCELL_X32 FILLER_32_3638 ();
 FILLCELL_X32 FILLER_32_3670 ();
 FILLCELL_X32 FILLER_32_3702 ();
 FILLCELL_X4 FILLER_32_3734 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X32 FILLER_33_289 ();
 FILLCELL_X32 FILLER_33_321 ();
 FILLCELL_X32 FILLER_33_353 ();
 FILLCELL_X32 FILLER_33_385 ();
 FILLCELL_X32 FILLER_33_417 ();
 FILLCELL_X32 FILLER_33_449 ();
 FILLCELL_X32 FILLER_33_481 ();
 FILLCELL_X32 FILLER_33_513 ();
 FILLCELL_X32 FILLER_33_545 ();
 FILLCELL_X32 FILLER_33_577 ();
 FILLCELL_X32 FILLER_33_609 ();
 FILLCELL_X32 FILLER_33_641 ();
 FILLCELL_X32 FILLER_33_673 ();
 FILLCELL_X32 FILLER_33_705 ();
 FILLCELL_X32 FILLER_33_737 ();
 FILLCELL_X32 FILLER_33_769 ();
 FILLCELL_X32 FILLER_33_801 ();
 FILLCELL_X32 FILLER_33_833 ();
 FILLCELL_X32 FILLER_33_865 ();
 FILLCELL_X32 FILLER_33_897 ();
 FILLCELL_X32 FILLER_33_929 ();
 FILLCELL_X32 FILLER_33_961 ();
 FILLCELL_X32 FILLER_33_993 ();
 FILLCELL_X32 FILLER_33_1025 ();
 FILLCELL_X32 FILLER_33_1057 ();
 FILLCELL_X32 FILLER_33_1089 ();
 FILLCELL_X32 FILLER_33_1121 ();
 FILLCELL_X32 FILLER_33_1153 ();
 FILLCELL_X32 FILLER_33_1185 ();
 FILLCELL_X32 FILLER_33_1217 ();
 FILLCELL_X8 FILLER_33_1249 ();
 FILLCELL_X4 FILLER_33_1257 ();
 FILLCELL_X2 FILLER_33_1261 ();
 FILLCELL_X32 FILLER_33_1264 ();
 FILLCELL_X32 FILLER_33_1296 ();
 FILLCELL_X32 FILLER_33_1328 ();
 FILLCELL_X32 FILLER_33_1360 ();
 FILLCELL_X32 FILLER_33_1392 ();
 FILLCELL_X32 FILLER_33_1424 ();
 FILLCELL_X32 FILLER_33_1456 ();
 FILLCELL_X32 FILLER_33_1488 ();
 FILLCELL_X32 FILLER_33_1520 ();
 FILLCELL_X32 FILLER_33_1552 ();
 FILLCELL_X32 FILLER_33_1584 ();
 FILLCELL_X32 FILLER_33_1616 ();
 FILLCELL_X32 FILLER_33_1648 ();
 FILLCELL_X32 FILLER_33_1680 ();
 FILLCELL_X32 FILLER_33_1712 ();
 FILLCELL_X32 FILLER_33_1744 ();
 FILLCELL_X32 FILLER_33_1776 ();
 FILLCELL_X32 FILLER_33_1808 ();
 FILLCELL_X32 FILLER_33_1840 ();
 FILLCELL_X32 FILLER_33_1872 ();
 FILLCELL_X32 FILLER_33_1904 ();
 FILLCELL_X32 FILLER_33_1936 ();
 FILLCELL_X32 FILLER_33_1968 ();
 FILLCELL_X32 FILLER_33_2000 ();
 FILLCELL_X32 FILLER_33_2032 ();
 FILLCELL_X32 FILLER_33_2064 ();
 FILLCELL_X32 FILLER_33_2096 ();
 FILLCELL_X32 FILLER_33_2128 ();
 FILLCELL_X32 FILLER_33_2160 ();
 FILLCELL_X32 FILLER_33_2192 ();
 FILLCELL_X32 FILLER_33_2224 ();
 FILLCELL_X32 FILLER_33_2256 ();
 FILLCELL_X32 FILLER_33_2288 ();
 FILLCELL_X32 FILLER_33_2320 ();
 FILLCELL_X32 FILLER_33_2352 ();
 FILLCELL_X32 FILLER_33_2384 ();
 FILLCELL_X32 FILLER_33_2416 ();
 FILLCELL_X32 FILLER_33_2448 ();
 FILLCELL_X32 FILLER_33_2480 ();
 FILLCELL_X8 FILLER_33_2512 ();
 FILLCELL_X4 FILLER_33_2520 ();
 FILLCELL_X2 FILLER_33_2524 ();
 FILLCELL_X32 FILLER_33_2527 ();
 FILLCELL_X32 FILLER_33_2559 ();
 FILLCELL_X32 FILLER_33_2591 ();
 FILLCELL_X32 FILLER_33_2623 ();
 FILLCELL_X32 FILLER_33_2655 ();
 FILLCELL_X32 FILLER_33_2687 ();
 FILLCELL_X32 FILLER_33_2719 ();
 FILLCELL_X32 FILLER_33_2751 ();
 FILLCELL_X32 FILLER_33_2783 ();
 FILLCELL_X32 FILLER_33_2815 ();
 FILLCELL_X32 FILLER_33_2847 ();
 FILLCELL_X32 FILLER_33_2879 ();
 FILLCELL_X32 FILLER_33_2911 ();
 FILLCELL_X32 FILLER_33_2943 ();
 FILLCELL_X32 FILLER_33_2975 ();
 FILLCELL_X32 FILLER_33_3007 ();
 FILLCELL_X32 FILLER_33_3039 ();
 FILLCELL_X32 FILLER_33_3071 ();
 FILLCELL_X32 FILLER_33_3103 ();
 FILLCELL_X32 FILLER_33_3135 ();
 FILLCELL_X32 FILLER_33_3167 ();
 FILLCELL_X32 FILLER_33_3199 ();
 FILLCELL_X32 FILLER_33_3231 ();
 FILLCELL_X32 FILLER_33_3263 ();
 FILLCELL_X32 FILLER_33_3295 ();
 FILLCELL_X32 FILLER_33_3327 ();
 FILLCELL_X32 FILLER_33_3359 ();
 FILLCELL_X32 FILLER_33_3391 ();
 FILLCELL_X32 FILLER_33_3423 ();
 FILLCELL_X32 FILLER_33_3455 ();
 FILLCELL_X32 FILLER_33_3487 ();
 FILLCELL_X32 FILLER_33_3519 ();
 FILLCELL_X32 FILLER_33_3551 ();
 FILLCELL_X32 FILLER_33_3583 ();
 FILLCELL_X32 FILLER_33_3615 ();
 FILLCELL_X32 FILLER_33_3647 ();
 FILLCELL_X32 FILLER_33_3679 ();
 FILLCELL_X16 FILLER_33_3711 ();
 FILLCELL_X8 FILLER_33_3727 ();
 FILLCELL_X2 FILLER_33_3735 ();
 FILLCELL_X1 FILLER_33_3737 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X32 FILLER_34_257 ();
 FILLCELL_X32 FILLER_34_289 ();
 FILLCELL_X32 FILLER_34_321 ();
 FILLCELL_X32 FILLER_34_353 ();
 FILLCELL_X32 FILLER_34_385 ();
 FILLCELL_X32 FILLER_34_417 ();
 FILLCELL_X32 FILLER_34_449 ();
 FILLCELL_X32 FILLER_34_481 ();
 FILLCELL_X32 FILLER_34_513 ();
 FILLCELL_X32 FILLER_34_545 ();
 FILLCELL_X32 FILLER_34_577 ();
 FILLCELL_X16 FILLER_34_609 ();
 FILLCELL_X4 FILLER_34_625 ();
 FILLCELL_X2 FILLER_34_629 ();
 FILLCELL_X32 FILLER_34_632 ();
 FILLCELL_X32 FILLER_34_664 ();
 FILLCELL_X32 FILLER_34_696 ();
 FILLCELL_X32 FILLER_34_728 ();
 FILLCELL_X32 FILLER_34_760 ();
 FILLCELL_X32 FILLER_34_792 ();
 FILLCELL_X32 FILLER_34_824 ();
 FILLCELL_X32 FILLER_34_856 ();
 FILLCELL_X32 FILLER_34_888 ();
 FILLCELL_X32 FILLER_34_920 ();
 FILLCELL_X32 FILLER_34_952 ();
 FILLCELL_X32 FILLER_34_984 ();
 FILLCELL_X32 FILLER_34_1016 ();
 FILLCELL_X32 FILLER_34_1048 ();
 FILLCELL_X32 FILLER_34_1080 ();
 FILLCELL_X32 FILLER_34_1112 ();
 FILLCELL_X32 FILLER_34_1144 ();
 FILLCELL_X32 FILLER_34_1176 ();
 FILLCELL_X32 FILLER_34_1208 ();
 FILLCELL_X32 FILLER_34_1240 ();
 FILLCELL_X32 FILLER_34_1272 ();
 FILLCELL_X32 FILLER_34_1304 ();
 FILLCELL_X32 FILLER_34_1336 ();
 FILLCELL_X32 FILLER_34_1368 ();
 FILLCELL_X32 FILLER_34_1400 ();
 FILLCELL_X32 FILLER_34_1432 ();
 FILLCELL_X32 FILLER_34_1464 ();
 FILLCELL_X32 FILLER_34_1496 ();
 FILLCELL_X32 FILLER_34_1528 ();
 FILLCELL_X32 FILLER_34_1560 ();
 FILLCELL_X32 FILLER_34_1592 ();
 FILLCELL_X32 FILLER_34_1624 ();
 FILLCELL_X32 FILLER_34_1656 ();
 FILLCELL_X32 FILLER_34_1688 ();
 FILLCELL_X32 FILLER_34_1720 ();
 FILLCELL_X32 FILLER_34_1752 ();
 FILLCELL_X32 FILLER_34_1784 ();
 FILLCELL_X32 FILLER_34_1816 ();
 FILLCELL_X32 FILLER_34_1848 ();
 FILLCELL_X8 FILLER_34_1880 ();
 FILLCELL_X4 FILLER_34_1888 ();
 FILLCELL_X2 FILLER_34_1892 ();
 FILLCELL_X32 FILLER_34_1895 ();
 FILLCELL_X32 FILLER_34_1927 ();
 FILLCELL_X32 FILLER_34_1959 ();
 FILLCELL_X32 FILLER_34_1991 ();
 FILLCELL_X32 FILLER_34_2023 ();
 FILLCELL_X32 FILLER_34_2055 ();
 FILLCELL_X32 FILLER_34_2087 ();
 FILLCELL_X32 FILLER_34_2119 ();
 FILLCELL_X32 FILLER_34_2151 ();
 FILLCELL_X32 FILLER_34_2183 ();
 FILLCELL_X32 FILLER_34_2215 ();
 FILLCELL_X32 FILLER_34_2247 ();
 FILLCELL_X32 FILLER_34_2279 ();
 FILLCELL_X32 FILLER_34_2311 ();
 FILLCELL_X32 FILLER_34_2343 ();
 FILLCELL_X32 FILLER_34_2375 ();
 FILLCELL_X32 FILLER_34_2407 ();
 FILLCELL_X32 FILLER_34_2439 ();
 FILLCELL_X32 FILLER_34_2471 ();
 FILLCELL_X32 FILLER_34_2503 ();
 FILLCELL_X32 FILLER_34_2535 ();
 FILLCELL_X32 FILLER_34_2567 ();
 FILLCELL_X32 FILLER_34_2599 ();
 FILLCELL_X32 FILLER_34_2631 ();
 FILLCELL_X32 FILLER_34_2663 ();
 FILLCELL_X32 FILLER_34_2695 ();
 FILLCELL_X32 FILLER_34_2727 ();
 FILLCELL_X32 FILLER_34_2759 ();
 FILLCELL_X32 FILLER_34_2791 ();
 FILLCELL_X32 FILLER_34_2823 ();
 FILLCELL_X32 FILLER_34_2855 ();
 FILLCELL_X32 FILLER_34_2887 ();
 FILLCELL_X32 FILLER_34_2919 ();
 FILLCELL_X32 FILLER_34_2951 ();
 FILLCELL_X32 FILLER_34_2983 ();
 FILLCELL_X32 FILLER_34_3015 ();
 FILLCELL_X32 FILLER_34_3047 ();
 FILLCELL_X32 FILLER_34_3079 ();
 FILLCELL_X32 FILLER_34_3111 ();
 FILLCELL_X8 FILLER_34_3143 ();
 FILLCELL_X4 FILLER_34_3151 ();
 FILLCELL_X2 FILLER_34_3155 ();
 FILLCELL_X32 FILLER_34_3158 ();
 FILLCELL_X32 FILLER_34_3190 ();
 FILLCELL_X32 FILLER_34_3222 ();
 FILLCELL_X32 FILLER_34_3254 ();
 FILLCELL_X32 FILLER_34_3286 ();
 FILLCELL_X32 FILLER_34_3318 ();
 FILLCELL_X32 FILLER_34_3350 ();
 FILLCELL_X32 FILLER_34_3382 ();
 FILLCELL_X32 FILLER_34_3414 ();
 FILLCELL_X32 FILLER_34_3446 ();
 FILLCELL_X32 FILLER_34_3478 ();
 FILLCELL_X32 FILLER_34_3510 ();
 FILLCELL_X32 FILLER_34_3542 ();
 FILLCELL_X32 FILLER_34_3574 ();
 FILLCELL_X32 FILLER_34_3606 ();
 FILLCELL_X32 FILLER_34_3638 ();
 FILLCELL_X32 FILLER_34_3670 ();
 FILLCELL_X32 FILLER_34_3702 ();
 FILLCELL_X4 FILLER_34_3734 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X32 FILLER_35_289 ();
 FILLCELL_X32 FILLER_35_321 ();
 FILLCELL_X32 FILLER_35_353 ();
 FILLCELL_X32 FILLER_35_385 ();
 FILLCELL_X32 FILLER_35_417 ();
 FILLCELL_X32 FILLER_35_449 ();
 FILLCELL_X32 FILLER_35_481 ();
 FILLCELL_X32 FILLER_35_513 ();
 FILLCELL_X32 FILLER_35_545 ();
 FILLCELL_X32 FILLER_35_577 ();
 FILLCELL_X32 FILLER_35_609 ();
 FILLCELL_X32 FILLER_35_641 ();
 FILLCELL_X32 FILLER_35_673 ();
 FILLCELL_X32 FILLER_35_705 ();
 FILLCELL_X32 FILLER_35_737 ();
 FILLCELL_X32 FILLER_35_769 ();
 FILLCELL_X32 FILLER_35_801 ();
 FILLCELL_X32 FILLER_35_833 ();
 FILLCELL_X32 FILLER_35_865 ();
 FILLCELL_X32 FILLER_35_897 ();
 FILLCELL_X32 FILLER_35_929 ();
 FILLCELL_X32 FILLER_35_961 ();
 FILLCELL_X32 FILLER_35_993 ();
 FILLCELL_X32 FILLER_35_1025 ();
 FILLCELL_X32 FILLER_35_1057 ();
 FILLCELL_X32 FILLER_35_1089 ();
 FILLCELL_X32 FILLER_35_1121 ();
 FILLCELL_X32 FILLER_35_1153 ();
 FILLCELL_X32 FILLER_35_1185 ();
 FILLCELL_X32 FILLER_35_1217 ();
 FILLCELL_X8 FILLER_35_1249 ();
 FILLCELL_X4 FILLER_35_1257 ();
 FILLCELL_X2 FILLER_35_1261 ();
 FILLCELL_X32 FILLER_35_1264 ();
 FILLCELL_X32 FILLER_35_1296 ();
 FILLCELL_X32 FILLER_35_1328 ();
 FILLCELL_X32 FILLER_35_1360 ();
 FILLCELL_X32 FILLER_35_1392 ();
 FILLCELL_X32 FILLER_35_1424 ();
 FILLCELL_X32 FILLER_35_1456 ();
 FILLCELL_X32 FILLER_35_1488 ();
 FILLCELL_X32 FILLER_35_1520 ();
 FILLCELL_X32 FILLER_35_1552 ();
 FILLCELL_X32 FILLER_35_1584 ();
 FILLCELL_X32 FILLER_35_1616 ();
 FILLCELL_X32 FILLER_35_1648 ();
 FILLCELL_X32 FILLER_35_1680 ();
 FILLCELL_X32 FILLER_35_1712 ();
 FILLCELL_X32 FILLER_35_1744 ();
 FILLCELL_X32 FILLER_35_1776 ();
 FILLCELL_X32 FILLER_35_1808 ();
 FILLCELL_X32 FILLER_35_1840 ();
 FILLCELL_X32 FILLER_35_1872 ();
 FILLCELL_X32 FILLER_35_1904 ();
 FILLCELL_X32 FILLER_35_1936 ();
 FILLCELL_X32 FILLER_35_1968 ();
 FILLCELL_X32 FILLER_35_2000 ();
 FILLCELL_X32 FILLER_35_2032 ();
 FILLCELL_X32 FILLER_35_2064 ();
 FILLCELL_X32 FILLER_35_2096 ();
 FILLCELL_X32 FILLER_35_2128 ();
 FILLCELL_X32 FILLER_35_2160 ();
 FILLCELL_X32 FILLER_35_2192 ();
 FILLCELL_X32 FILLER_35_2224 ();
 FILLCELL_X32 FILLER_35_2256 ();
 FILLCELL_X32 FILLER_35_2288 ();
 FILLCELL_X32 FILLER_35_2320 ();
 FILLCELL_X32 FILLER_35_2352 ();
 FILLCELL_X32 FILLER_35_2384 ();
 FILLCELL_X32 FILLER_35_2416 ();
 FILLCELL_X32 FILLER_35_2448 ();
 FILLCELL_X32 FILLER_35_2480 ();
 FILLCELL_X8 FILLER_35_2512 ();
 FILLCELL_X4 FILLER_35_2520 ();
 FILLCELL_X2 FILLER_35_2524 ();
 FILLCELL_X32 FILLER_35_2527 ();
 FILLCELL_X32 FILLER_35_2559 ();
 FILLCELL_X32 FILLER_35_2591 ();
 FILLCELL_X32 FILLER_35_2623 ();
 FILLCELL_X32 FILLER_35_2655 ();
 FILLCELL_X32 FILLER_35_2687 ();
 FILLCELL_X32 FILLER_35_2719 ();
 FILLCELL_X32 FILLER_35_2751 ();
 FILLCELL_X32 FILLER_35_2783 ();
 FILLCELL_X32 FILLER_35_2815 ();
 FILLCELL_X32 FILLER_35_2847 ();
 FILLCELL_X32 FILLER_35_2879 ();
 FILLCELL_X32 FILLER_35_2911 ();
 FILLCELL_X32 FILLER_35_2943 ();
 FILLCELL_X32 FILLER_35_2975 ();
 FILLCELL_X32 FILLER_35_3007 ();
 FILLCELL_X32 FILLER_35_3039 ();
 FILLCELL_X32 FILLER_35_3071 ();
 FILLCELL_X32 FILLER_35_3103 ();
 FILLCELL_X32 FILLER_35_3135 ();
 FILLCELL_X32 FILLER_35_3167 ();
 FILLCELL_X32 FILLER_35_3199 ();
 FILLCELL_X32 FILLER_35_3231 ();
 FILLCELL_X32 FILLER_35_3263 ();
 FILLCELL_X32 FILLER_35_3295 ();
 FILLCELL_X32 FILLER_35_3327 ();
 FILLCELL_X32 FILLER_35_3359 ();
 FILLCELL_X32 FILLER_35_3391 ();
 FILLCELL_X32 FILLER_35_3423 ();
 FILLCELL_X32 FILLER_35_3455 ();
 FILLCELL_X32 FILLER_35_3487 ();
 FILLCELL_X32 FILLER_35_3519 ();
 FILLCELL_X32 FILLER_35_3551 ();
 FILLCELL_X32 FILLER_35_3583 ();
 FILLCELL_X32 FILLER_35_3615 ();
 FILLCELL_X32 FILLER_35_3647 ();
 FILLCELL_X32 FILLER_35_3679 ();
 FILLCELL_X16 FILLER_35_3711 ();
 FILLCELL_X8 FILLER_35_3727 ();
 FILLCELL_X2 FILLER_35_3735 ();
 FILLCELL_X1 FILLER_35_3737 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X32 FILLER_36_289 ();
 FILLCELL_X32 FILLER_36_321 ();
 FILLCELL_X32 FILLER_36_353 ();
 FILLCELL_X32 FILLER_36_385 ();
 FILLCELL_X32 FILLER_36_417 ();
 FILLCELL_X32 FILLER_36_449 ();
 FILLCELL_X32 FILLER_36_481 ();
 FILLCELL_X32 FILLER_36_513 ();
 FILLCELL_X32 FILLER_36_545 ();
 FILLCELL_X32 FILLER_36_577 ();
 FILLCELL_X16 FILLER_36_609 ();
 FILLCELL_X4 FILLER_36_625 ();
 FILLCELL_X2 FILLER_36_629 ();
 FILLCELL_X32 FILLER_36_632 ();
 FILLCELL_X32 FILLER_36_664 ();
 FILLCELL_X32 FILLER_36_696 ();
 FILLCELL_X32 FILLER_36_728 ();
 FILLCELL_X32 FILLER_36_760 ();
 FILLCELL_X32 FILLER_36_792 ();
 FILLCELL_X32 FILLER_36_824 ();
 FILLCELL_X32 FILLER_36_856 ();
 FILLCELL_X32 FILLER_36_888 ();
 FILLCELL_X32 FILLER_36_920 ();
 FILLCELL_X32 FILLER_36_952 ();
 FILLCELL_X32 FILLER_36_984 ();
 FILLCELL_X32 FILLER_36_1016 ();
 FILLCELL_X32 FILLER_36_1048 ();
 FILLCELL_X32 FILLER_36_1080 ();
 FILLCELL_X32 FILLER_36_1112 ();
 FILLCELL_X32 FILLER_36_1144 ();
 FILLCELL_X32 FILLER_36_1176 ();
 FILLCELL_X32 FILLER_36_1208 ();
 FILLCELL_X32 FILLER_36_1240 ();
 FILLCELL_X32 FILLER_36_1272 ();
 FILLCELL_X32 FILLER_36_1304 ();
 FILLCELL_X32 FILLER_36_1336 ();
 FILLCELL_X32 FILLER_36_1368 ();
 FILLCELL_X32 FILLER_36_1400 ();
 FILLCELL_X32 FILLER_36_1432 ();
 FILLCELL_X32 FILLER_36_1464 ();
 FILLCELL_X32 FILLER_36_1496 ();
 FILLCELL_X32 FILLER_36_1528 ();
 FILLCELL_X32 FILLER_36_1560 ();
 FILLCELL_X32 FILLER_36_1592 ();
 FILLCELL_X32 FILLER_36_1624 ();
 FILLCELL_X32 FILLER_36_1656 ();
 FILLCELL_X32 FILLER_36_1688 ();
 FILLCELL_X32 FILLER_36_1720 ();
 FILLCELL_X32 FILLER_36_1752 ();
 FILLCELL_X32 FILLER_36_1784 ();
 FILLCELL_X32 FILLER_36_1816 ();
 FILLCELL_X32 FILLER_36_1848 ();
 FILLCELL_X8 FILLER_36_1880 ();
 FILLCELL_X4 FILLER_36_1888 ();
 FILLCELL_X2 FILLER_36_1892 ();
 FILLCELL_X32 FILLER_36_1895 ();
 FILLCELL_X32 FILLER_36_1927 ();
 FILLCELL_X32 FILLER_36_1959 ();
 FILLCELL_X32 FILLER_36_1991 ();
 FILLCELL_X32 FILLER_36_2023 ();
 FILLCELL_X32 FILLER_36_2055 ();
 FILLCELL_X32 FILLER_36_2087 ();
 FILLCELL_X32 FILLER_36_2119 ();
 FILLCELL_X32 FILLER_36_2151 ();
 FILLCELL_X32 FILLER_36_2183 ();
 FILLCELL_X32 FILLER_36_2215 ();
 FILLCELL_X32 FILLER_36_2247 ();
 FILLCELL_X32 FILLER_36_2279 ();
 FILLCELL_X32 FILLER_36_2311 ();
 FILLCELL_X32 FILLER_36_2343 ();
 FILLCELL_X32 FILLER_36_2375 ();
 FILLCELL_X32 FILLER_36_2407 ();
 FILLCELL_X32 FILLER_36_2439 ();
 FILLCELL_X32 FILLER_36_2471 ();
 FILLCELL_X32 FILLER_36_2503 ();
 FILLCELL_X32 FILLER_36_2535 ();
 FILLCELL_X32 FILLER_36_2567 ();
 FILLCELL_X32 FILLER_36_2599 ();
 FILLCELL_X32 FILLER_36_2631 ();
 FILLCELL_X32 FILLER_36_2663 ();
 FILLCELL_X32 FILLER_36_2695 ();
 FILLCELL_X32 FILLER_36_2727 ();
 FILLCELL_X32 FILLER_36_2759 ();
 FILLCELL_X32 FILLER_36_2791 ();
 FILLCELL_X32 FILLER_36_2823 ();
 FILLCELL_X32 FILLER_36_2855 ();
 FILLCELL_X32 FILLER_36_2887 ();
 FILLCELL_X32 FILLER_36_2919 ();
 FILLCELL_X32 FILLER_36_2951 ();
 FILLCELL_X32 FILLER_36_2983 ();
 FILLCELL_X32 FILLER_36_3015 ();
 FILLCELL_X32 FILLER_36_3047 ();
 FILLCELL_X32 FILLER_36_3079 ();
 FILLCELL_X32 FILLER_36_3111 ();
 FILLCELL_X8 FILLER_36_3143 ();
 FILLCELL_X4 FILLER_36_3151 ();
 FILLCELL_X2 FILLER_36_3155 ();
 FILLCELL_X32 FILLER_36_3158 ();
 FILLCELL_X32 FILLER_36_3190 ();
 FILLCELL_X32 FILLER_36_3222 ();
 FILLCELL_X32 FILLER_36_3254 ();
 FILLCELL_X32 FILLER_36_3286 ();
 FILLCELL_X32 FILLER_36_3318 ();
 FILLCELL_X32 FILLER_36_3350 ();
 FILLCELL_X32 FILLER_36_3382 ();
 FILLCELL_X32 FILLER_36_3414 ();
 FILLCELL_X32 FILLER_36_3446 ();
 FILLCELL_X32 FILLER_36_3478 ();
 FILLCELL_X32 FILLER_36_3510 ();
 FILLCELL_X32 FILLER_36_3542 ();
 FILLCELL_X32 FILLER_36_3574 ();
 FILLCELL_X32 FILLER_36_3606 ();
 FILLCELL_X32 FILLER_36_3638 ();
 FILLCELL_X32 FILLER_36_3670 ();
 FILLCELL_X32 FILLER_36_3702 ();
 FILLCELL_X4 FILLER_36_3734 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X32 FILLER_37_289 ();
 FILLCELL_X32 FILLER_37_321 ();
 FILLCELL_X32 FILLER_37_353 ();
 FILLCELL_X32 FILLER_37_385 ();
 FILLCELL_X32 FILLER_37_417 ();
 FILLCELL_X32 FILLER_37_449 ();
 FILLCELL_X32 FILLER_37_481 ();
 FILLCELL_X32 FILLER_37_513 ();
 FILLCELL_X32 FILLER_37_545 ();
 FILLCELL_X32 FILLER_37_577 ();
 FILLCELL_X32 FILLER_37_609 ();
 FILLCELL_X32 FILLER_37_641 ();
 FILLCELL_X32 FILLER_37_673 ();
 FILLCELL_X32 FILLER_37_705 ();
 FILLCELL_X32 FILLER_37_737 ();
 FILLCELL_X32 FILLER_37_769 ();
 FILLCELL_X32 FILLER_37_801 ();
 FILLCELL_X32 FILLER_37_833 ();
 FILLCELL_X32 FILLER_37_865 ();
 FILLCELL_X32 FILLER_37_897 ();
 FILLCELL_X32 FILLER_37_929 ();
 FILLCELL_X32 FILLER_37_961 ();
 FILLCELL_X32 FILLER_37_993 ();
 FILLCELL_X32 FILLER_37_1025 ();
 FILLCELL_X32 FILLER_37_1057 ();
 FILLCELL_X32 FILLER_37_1089 ();
 FILLCELL_X32 FILLER_37_1121 ();
 FILLCELL_X32 FILLER_37_1153 ();
 FILLCELL_X32 FILLER_37_1185 ();
 FILLCELL_X32 FILLER_37_1217 ();
 FILLCELL_X8 FILLER_37_1249 ();
 FILLCELL_X4 FILLER_37_1257 ();
 FILLCELL_X2 FILLER_37_1261 ();
 FILLCELL_X32 FILLER_37_1264 ();
 FILLCELL_X32 FILLER_37_1296 ();
 FILLCELL_X32 FILLER_37_1328 ();
 FILLCELL_X32 FILLER_37_1360 ();
 FILLCELL_X32 FILLER_37_1392 ();
 FILLCELL_X32 FILLER_37_1424 ();
 FILLCELL_X32 FILLER_37_1456 ();
 FILLCELL_X32 FILLER_37_1488 ();
 FILLCELL_X32 FILLER_37_1520 ();
 FILLCELL_X32 FILLER_37_1552 ();
 FILLCELL_X32 FILLER_37_1584 ();
 FILLCELL_X32 FILLER_37_1616 ();
 FILLCELL_X32 FILLER_37_1648 ();
 FILLCELL_X32 FILLER_37_1680 ();
 FILLCELL_X32 FILLER_37_1712 ();
 FILLCELL_X32 FILLER_37_1744 ();
 FILLCELL_X32 FILLER_37_1776 ();
 FILLCELL_X32 FILLER_37_1808 ();
 FILLCELL_X32 FILLER_37_1840 ();
 FILLCELL_X32 FILLER_37_1872 ();
 FILLCELL_X32 FILLER_37_1904 ();
 FILLCELL_X32 FILLER_37_1936 ();
 FILLCELL_X32 FILLER_37_1968 ();
 FILLCELL_X32 FILLER_37_2000 ();
 FILLCELL_X32 FILLER_37_2032 ();
 FILLCELL_X32 FILLER_37_2064 ();
 FILLCELL_X32 FILLER_37_2096 ();
 FILLCELL_X32 FILLER_37_2128 ();
 FILLCELL_X32 FILLER_37_2160 ();
 FILLCELL_X32 FILLER_37_2192 ();
 FILLCELL_X32 FILLER_37_2224 ();
 FILLCELL_X32 FILLER_37_2256 ();
 FILLCELL_X32 FILLER_37_2288 ();
 FILLCELL_X32 FILLER_37_2320 ();
 FILLCELL_X32 FILLER_37_2352 ();
 FILLCELL_X32 FILLER_37_2384 ();
 FILLCELL_X32 FILLER_37_2416 ();
 FILLCELL_X32 FILLER_37_2448 ();
 FILLCELL_X32 FILLER_37_2480 ();
 FILLCELL_X8 FILLER_37_2512 ();
 FILLCELL_X4 FILLER_37_2520 ();
 FILLCELL_X2 FILLER_37_2524 ();
 FILLCELL_X32 FILLER_37_2527 ();
 FILLCELL_X32 FILLER_37_2559 ();
 FILLCELL_X32 FILLER_37_2591 ();
 FILLCELL_X32 FILLER_37_2623 ();
 FILLCELL_X32 FILLER_37_2655 ();
 FILLCELL_X32 FILLER_37_2687 ();
 FILLCELL_X32 FILLER_37_2719 ();
 FILLCELL_X32 FILLER_37_2751 ();
 FILLCELL_X32 FILLER_37_2783 ();
 FILLCELL_X32 FILLER_37_2815 ();
 FILLCELL_X32 FILLER_37_2847 ();
 FILLCELL_X32 FILLER_37_2879 ();
 FILLCELL_X32 FILLER_37_2911 ();
 FILLCELL_X32 FILLER_37_2943 ();
 FILLCELL_X32 FILLER_37_2975 ();
 FILLCELL_X32 FILLER_37_3007 ();
 FILLCELL_X32 FILLER_37_3039 ();
 FILLCELL_X32 FILLER_37_3071 ();
 FILLCELL_X32 FILLER_37_3103 ();
 FILLCELL_X32 FILLER_37_3135 ();
 FILLCELL_X32 FILLER_37_3167 ();
 FILLCELL_X32 FILLER_37_3199 ();
 FILLCELL_X32 FILLER_37_3231 ();
 FILLCELL_X32 FILLER_37_3263 ();
 FILLCELL_X32 FILLER_37_3295 ();
 FILLCELL_X32 FILLER_37_3327 ();
 FILLCELL_X32 FILLER_37_3359 ();
 FILLCELL_X32 FILLER_37_3391 ();
 FILLCELL_X32 FILLER_37_3423 ();
 FILLCELL_X32 FILLER_37_3455 ();
 FILLCELL_X32 FILLER_37_3487 ();
 FILLCELL_X32 FILLER_37_3519 ();
 FILLCELL_X32 FILLER_37_3551 ();
 FILLCELL_X32 FILLER_37_3583 ();
 FILLCELL_X32 FILLER_37_3615 ();
 FILLCELL_X32 FILLER_37_3647 ();
 FILLCELL_X32 FILLER_37_3679 ();
 FILLCELL_X16 FILLER_37_3711 ();
 FILLCELL_X8 FILLER_37_3727 ();
 FILLCELL_X2 FILLER_37_3735 ();
 FILLCELL_X1 FILLER_37_3737 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X32 FILLER_38_289 ();
 FILLCELL_X32 FILLER_38_321 ();
 FILLCELL_X32 FILLER_38_353 ();
 FILLCELL_X32 FILLER_38_385 ();
 FILLCELL_X32 FILLER_38_417 ();
 FILLCELL_X32 FILLER_38_449 ();
 FILLCELL_X32 FILLER_38_481 ();
 FILLCELL_X32 FILLER_38_513 ();
 FILLCELL_X32 FILLER_38_545 ();
 FILLCELL_X32 FILLER_38_577 ();
 FILLCELL_X16 FILLER_38_609 ();
 FILLCELL_X4 FILLER_38_625 ();
 FILLCELL_X2 FILLER_38_629 ();
 FILLCELL_X32 FILLER_38_632 ();
 FILLCELL_X32 FILLER_38_664 ();
 FILLCELL_X32 FILLER_38_696 ();
 FILLCELL_X32 FILLER_38_728 ();
 FILLCELL_X32 FILLER_38_760 ();
 FILLCELL_X32 FILLER_38_792 ();
 FILLCELL_X32 FILLER_38_824 ();
 FILLCELL_X32 FILLER_38_856 ();
 FILLCELL_X32 FILLER_38_888 ();
 FILLCELL_X32 FILLER_38_920 ();
 FILLCELL_X32 FILLER_38_952 ();
 FILLCELL_X32 FILLER_38_984 ();
 FILLCELL_X32 FILLER_38_1016 ();
 FILLCELL_X32 FILLER_38_1048 ();
 FILLCELL_X32 FILLER_38_1080 ();
 FILLCELL_X32 FILLER_38_1112 ();
 FILLCELL_X32 FILLER_38_1144 ();
 FILLCELL_X32 FILLER_38_1176 ();
 FILLCELL_X32 FILLER_38_1208 ();
 FILLCELL_X32 FILLER_38_1240 ();
 FILLCELL_X32 FILLER_38_1272 ();
 FILLCELL_X32 FILLER_38_1304 ();
 FILLCELL_X32 FILLER_38_1336 ();
 FILLCELL_X32 FILLER_38_1368 ();
 FILLCELL_X32 FILLER_38_1400 ();
 FILLCELL_X32 FILLER_38_1432 ();
 FILLCELL_X32 FILLER_38_1464 ();
 FILLCELL_X32 FILLER_38_1496 ();
 FILLCELL_X32 FILLER_38_1528 ();
 FILLCELL_X32 FILLER_38_1560 ();
 FILLCELL_X32 FILLER_38_1592 ();
 FILLCELL_X32 FILLER_38_1624 ();
 FILLCELL_X32 FILLER_38_1656 ();
 FILLCELL_X32 FILLER_38_1688 ();
 FILLCELL_X32 FILLER_38_1720 ();
 FILLCELL_X32 FILLER_38_1752 ();
 FILLCELL_X32 FILLER_38_1784 ();
 FILLCELL_X32 FILLER_38_1816 ();
 FILLCELL_X32 FILLER_38_1848 ();
 FILLCELL_X8 FILLER_38_1880 ();
 FILLCELL_X4 FILLER_38_1888 ();
 FILLCELL_X2 FILLER_38_1892 ();
 FILLCELL_X32 FILLER_38_1895 ();
 FILLCELL_X32 FILLER_38_1927 ();
 FILLCELL_X32 FILLER_38_1959 ();
 FILLCELL_X32 FILLER_38_1991 ();
 FILLCELL_X32 FILLER_38_2023 ();
 FILLCELL_X32 FILLER_38_2055 ();
 FILLCELL_X32 FILLER_38_2087 ();
 FILLCELL_X32 FILLER_38_2119 ();
 FILLCELL_X32 FILLER_38_2151 ();
 FILLCELL_X32 FILLER_38_2183 ();
 FILLCELL_X32 FILLER_38_2215 ();
 FILLCELL_X32 FILLER_38_2247 ();
 FILLCELL_X32 FILLER_38_2279 ();
 FILLCELL_X32 FILLER_38_2311 ();
 FILLCELL_X32 FILLER_38_2343 ();
 FILLCELL_X32 FILLER_38_2375 ();
 FILLCELL_X32 FILLER_38_2407 ();
 FILLCELL_X32 FILLER_38_2439 ();
 FILLCELL_X32 FILLER_38_2471 ();
 FILLCELL_X32 FILLER_38_2503 ();
 FILLCELL_X32 FILLER_38_2535 ();
 FILLCELL_X32 FILLER_38_2567 ();
 FILLCELL_X32 FILLER_38_2599 ();
 FILLCELL_X32 FILLER_38_2631 ();
 FILLCELL_X32 FILLER_38_2663 ();
 FILLCELL_X32 FILLER_38_2695 ();
 FILLCELL_X32 FILLER_38_2727 ();
 FILLCELL_X32 FILLER_38_2759 ();
 FILLCELL_X32 FILLER_38_2791 ();
 FILLCELL_X32 FILLER_38_2823 ();
 FILLCELL_X32 FILLER_38_2855 ();
 FILLCELL_X32 FILLER_38_2887 ();
 FILLCELL_X32 FILLER_38_2919 ();
 FILLCELL_X32 FILLER_38_2951 ();
 FILLCELL_X32 FILLER_38_2983 ();
 FILLCELL_X32 FILLER_38_3015 ();
 FILLCELL_X32 FILLER_38_3047 ();
 FILLCELL_X32 FILLER_38_3079 ();
 FILLCELL_X32 FILLER_38_3111 ();
 FILLCELL_X8 FILLER_38_3143 ();
 FILLCELL_X4 FILLER_38_3151 ();
 FILLCELL_X2 FILLER_38_3155 ();
 FILLCELL_X32 FILLER_38_3158 ();
 FILLCELL_X32 FILLER_38_3190 ();
 FILLCELL_X32 FILLER_38_3222 ();
 FILLCELL_X32 FILLER_38_3254 ();
 FILLCELL_X32 FILLER_38_3286 ();
 FILLCELL_X32 FILLER_38_3318 ();
 FILLCELL_X32 FILLER_38_3350 ();
 FILLCELL_X32 FILLER_38_3382 ();
 FILLCELL_X32 FILLER_38_3414 ();
 FILLCELL_X32 FILLER_38_3446 ();
 FILLCELL_X32 FILLER_38_3478 ();
 FILLCELL_X32 FILLER_38_3510 ();
 FILLCELL_X32 FILLER_38_3542 ();
 FILLCELL_X32 FILLER_38_3574 ();
 FILLCELL_X32 FILLER_38_3606 ();
 FILLCELL_X32 FILLER_38_3638 ();
 FILLCELL_X32 FILLER_38_3670 ();
 FILLCELL_X32 FILLER_38_3702 ();
 FILLCELL_X4 FILLER_38_3734 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X32 FILLER_39_289 ();
 FILLCELL_X32 FILLER_39_321 ();
 FILLCELL_X32 FILLER_39_353 ();
 FILLCELL_X32 FILLER_39_385 ();
 FILLCELL_X32 FILLER_39_417 ();
 FILLCELL_X32 FILLER_39_449 ();
 FILLCELL_X32 FILLER_39_481 ();
 FILLCELL_X32 FILLER_39_513 ();
 FILLCELL_X32 FILLER_39_545 ();
 FILLCELL_X32 FILLER_39_577 ();
 FILLCELL_X32 FILLER_39_609 ();
 FILLCELL_X32 FILLER_39_641 ();
 FILLCELL_X32 FILLER_39_673 ();
 FILLCELL_X32 FILLER_39_705 ();
 FILLCELL_X32 FILLER_39_737 ();
 FILLCELL_X32 FILLER_39_769 ();
 FILLCELL_X32 FILLER_39_801 ();
 FILLCELL_X32 FILLER_39_833 ();
 FILLCELL_X32 FILLER_39_865 ();
 FILLCELL_X32 FILLER_39_897 ();
 FILLCELL_X32 FILLER_39_929 ();
 FILLCELL_X32 FILLER_39_961 ();
 FILLCELL_X32 FILLER_39_993 ();
 FILLCELL_X32 FILLER_39_1025 ();
 FILLCELL_X32 FILLER_39_1057 ();
 FILLCELL_X32 FILLER_39_1089 ();
 FILLCELL_X32 FILLER_39_1121 ();
 FILLCELL_X32 FILLER_39_1153 ();
 FILLCELL_X32 FILLER_39_1185 ();
 FILLCELL_X32 FILLER_39_1217 ();
 FILLCELL_X8 FILLER_39_1249 ();
 FILLCELL_X4 FILLER_39_1257 ();
 FILLCELL_X2 FILLER_39_1261 ();
 FILLCELL_X32 FILLER_39_1264 ();
 FILLCELL_X32 FILLER_39_1296 ();
 FILLCELL_X32 FILLER_39_1328 ();
 FILLCELL_X32 FILLER_39_1360 ();
 FILLCELL_X32 FILLER_39_1392 ();
 FILLCELL_X32 FILLER_39_1424 ();
 FILLCELL_X32 FILLER_39_1456 ();
 FILLCELL_X32 FILLER_39_1488 ();
 FILLCELL_X32 FILLER_39_1520 ();
 FILLCELL_X32 FILLER_39_1552 ();
 FILLCELL_X32 FILLER_39_1584 ();
 FILLCELL_X32 FILLER_39_1616 ();
 FILLCELL_X32 FILLER_39_1648 ();
 FILLCELL_X32 FILLER_39_1680 ();
 FILLCELL_X32 FILLER_39_1712 ();
 FILLCELL_X32 FILLER_39_1744 ();
 FILLCELL_X32 FILLER_39_1776 ();
 FILLCELL_X32 FILLER_39_1808 ();
 FILLCELL_X32 FILLER_39_1840 ();
 FILLCELL_X32 FILLER_39_1872 ();
 FILLCELL_X32 FILLER_39_1904 ();
 FILLCELL_X32 FILLER_39_1936 ();
 FILLCELL_X32 FILLER_39_1968 ();
 FILLCELL_X32 FILLER_39_2000 ();
 FILLCELL_X32 FILLER_39_2032 ();
 FILLCELL_X32 FILLER_39_2064 ();
 FILLCELL_X32 FILLER_39_2096 ();
 FILLCELL_X32 FILLER_39_2128 ();
 FILLCELL_X32 FILLER_39_2160 ();
 FILLCELL_X32 FILLER_39_2192 ();
 FILLCELL_X32 FILLER_39_2224 ();
 FILLCELL_X32 FILLER_39_2256 ();
 FILLCELL_X32 FILLER_39_2288 ();
 FILLCELL_X32 FILLER_39_2320 ();
 FILLCELL_X32 FILLER_39_2352 ();
 FILLCELL_X32 FILLER_39_2384 ();
 FILLCELL_X32 FILLER_39_2416 ();
 FILLCELL_X32 FILLER_39_2448 ();
 FILLCELL_X32 FILLER_39_2480 ();
 FILLCELL_X8 FILLER_39_2512 ();
 FILLCELL_X4 FILLER_39_2520 ();
 FILLCELL_X2 FILLER_39_2524 ();
 FILLCELL_X32 FILLER_39_2527 ();
 FILLCELL_X32 FILLER_39_2559 ();
 FILLCELL_X32 FILLER_39_2591 ();
 FILLCELL_X32 FILLER_39_2623 ();
 FILLCELL_X32 FILLER_39_2655 ();
 FILLCELL_X32 FILLER_39_2687 ();
 FILLCELL_X32 FILLER_39_2719 ();
 FILLCELL_X32 FILLER_39_2751 ();
 FILLCELL_X32 FILLER_39_2783 ();
 FILLCELL_X32 FILLER_39_2815 ();
 FILLCELL_X32 FILLER_39_2847 ();
 FILLCELL_X32 FILLER_39_2879 ();
 FILLCELL_X32 FILLER_39_2911 ();
 FILLCELL_X32 FILLER_39_2943 ();
 FILLCELL_X32 FILLER_39_2975 ();
 FILLCELL_X32 FILLER_39_3007 ();
 FILLCELL_X32 FILLER_39_3039 ();
 FILLCELL_X32 FILLER_39_3071 ();
 FILLCELL_X32 FILLER_39_3103 ();
 FILLCELL_X32 FILLER_39_3135 ();
 FILLCELL_X32 FILLER_39_3167 ();
 FILLCELL_X32 FILLER_39_3199 ();
 FILLCELL_X32 FILLER_39_3231 ();
 FILLCELL_X32 FILLER_39_3263 ();
 FILLCELL_X32 FILLER_39_3295 ();
 FILLCELL_X32 FILLER_39_3327 ();
 FILLCELL_X32 FILLER_39_3359 ();
 FILLCELL_X32 FILLER_39_3391 ();
 FILLCELL_X32 FILLER_39_3423 ();
 FILLCELL_X32 FILLER_39_3455 ();
 FILLCELL_X32 FILLER_39_3487 ();
 FILLCELL_X32 FILLER_39_3519 ();
 FILLCELL_X32 FILLER_39_3551 ();
 FILLCELL_X32 FILLER_39_3583 ();
 FILLCELL_X32 FILLER_39_3615 ();
 FILLCELL_X32 FILLER_39_3647 ();
 FILLCELL_X32 FILLER_39_3679 ();
 FILLCELL_X16 FILLER_39_3711 ();
 FILLCELL_X8 FILLER_39_3727 ();
 FILLCELL_X2 FILLER_39_3735 ();
 FILLCELL_X1 FILLER_39_3737 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X32 FILLER_40_289 ();
 FILLCELL_X32 FILLER_40_321 ();
 FILLCELL_X32 FILLER_40_353 ();
 FILLCELL_X32 FILLER_40_385 ();
 FILLCELL_X32 FILLER_40_417 ();
 FILLCELL_X32 FILLER_40_449 ();
 FILLCELL_X32 FILLER_40_481 ();
 FILLCELL_X32 FILLER_40_513 ();
 FILLCELL_X32 FILLER_40_545 ();
 FILLCELL_X32 FILLER_40_577 ();
 FILLCELL_X16 FILLER_40_609 ();
 FILLCELL_X4 FILLER_40_625 ();
 FILLCELL_X2 FILLER_40_629 ();
 FILLCELL_X32 FILLER_40_632 ();
 FILLCELL_X32 FILLER_40_664 ();
 FILLCELL_X32 FILLER_40_696 ();
 FILLCELL_X32 FILLER_40_728 ();
 FILLCELL_X32 FILLER_40_760 ();
 FILLCELL_X32 FILLER_40_792 ();
 FILLCELL_X32 FILLER_40_824 ();
 FILLCELL_X32 FILLER_40_856 ();
 FILLCELL_X32 FILLER_40_888 ();
 FILLCELL_X32 FILLER_40_920 ();
 FILLCELL_X32 FILLER_40_952 ();
 FILLCELL_X32 FILLER_40_984 ();
 FILLCELL_X32 FILLER_40_1016 ();
 FILLCELL_X32 FILLER_40_1048 ();
 FILLCELL_X32 FILLER_40_1080 ();
 FILLCELL_X32 FILLER_40_1112 ();
 FILLCELL_X32 FILLER_40_1144 ();
 FILLCELL_X32 FILLER_40_1176 ();
 FILLCELL_X32 FILLER_40_1208 ();
 FILLCELL_X32 FILLER_40_1240 ();
 FILLCELL_X32 FILLER_40_1272 ();
 FILLCELL_X32 FILLER_40_1304 ();
 FILLCELL_X32 FILLER_40_1336 ();
 FILLCELL_X32 FILLER_40_1368 ();
 FILLCELL_X32 FILLER_40_1400 ();
 FILLCELL_X32 FILLER_40_1432 ();
 FILLCELL_X32 FILLER_40_1464 ();
 FILLCELL_X32 FILLER_40_1496 ();
 FILLCELL_X32 FILLER_40_1528 ();
 FILLCELL_X32 FILLER_40_1560 ();
 FILLCELL_X32 FILLER_40_1592 ();
 FILLCELL_X32 FILLER_40_1624 ();
 FILLCELL_X32 FILLER_40_1656 ();
 FILLCELL_X32 FILLER_40_1688 ();
 FILLCELL_X32 FILLER_40_1720 ();
 FILLCELL_X32 FILLER_40_1752 ();
 FILLCELL_X32 FILLER_40_1784 ();
 FILLCELL_X32 FILLER_40_1816 ();
 FILLCELL_X32 FILLER_40_1848 ();
 FILLCELL_X8 FILLER_40_1880 ();
 FILLCELL_X4 FILLER_40_1888 ();
 FILLCELL_X2 FILLER_40_1892 ();
 FILLCELL_X32 FILLER_40_1895 ();
 FILLCELL_X32 FILLER_40_1927 ();
 FILLCELL_X32 FILLER_40_1959 ();
 FILLCELL_X32 FILLER_40_1991 ();
 FILLCELL_X32 FILLER_40_2023 ();
 FILLCELL_X32 FILLER_40_2055 ();
 FILLCELL_X32 FILLER_40_2087 ();
 FILLCELL_X32 FILLER_40_2119 ();
 FILLCELL_X32 FILLER_40_2151 ();
 FILLCELL_X32 FILLER_40_2183 ();
 FILLCELL_X32 FILLER_40_2215 ();
 FILLCELL_X32 FILLER_40_2247 ();
 FILLCELL_X32 FILLER_40_2279 ();
 FILLCELL_X32 FILLER_40_2311 ();
 FILLCELL_X32 FILLER_40_2343 ();
 FILLCELL_X32 FILLER_40_2375 ();
 FILLCELL_X32 FILLER_40_2407 ();
 FILLCELL_X32 FILLER_40_2439 ();
 FILLCELL_X32 FILLER_40_2471 ();
 FILLCELL_X32 FILLER_40_2503 ();
 FILLCELL_X32 FILLER_40_2535 ();
 FILLCELL_X32 FILLER_40_2567 ();
 FILLCELL_X32 FILLER_40_2599 ();
 FILLCELL_X32 FILLER_40_2631 ();
 FILLCELL_X32 FILLER_40_2663 ();
 FILLCELL_X32 FILLER_40_2695 ();
 FILLCELL_X32 FILLER_40_2727 ();
 FILLCELL_X32 FILLER_40_2759 ();
 FILLCELL_X32 FILLER_40_2791 ();
 FILLCELL_X32 FILLER_40_2823 ();
 FILLCELL_X32 FILLER_40_2855 ();
 FILLCELL_X32 FILLER_40_2887 ();
 FILLCELL_X32 FILLER_40_2919 ();
 FILLCELL_X32 FILLER_40_2951 ();
 FILLCELL_X32 FILLER_40_2983 ();
 FILLCELL_X32 FILLER_40_3015 ();
 FILLCELL_X32 FILLER_40_3047 ();
 FILLCELL_X32 FILLER_40_3079 ();
 FILLCELL_X32 FILLER_40_3111 ();
 FILLCELL_X8 FILLER_40_3143 ();
 FILLCELL_X4 FILLER_40_3151 ();
 FILLCELL_X2 FILLER_40_3155 ();
 FILLCELL_X32 FILLER_40_3158 ();
 FILLCELL_X32 FILLER_40_3190 ();
 FILLCELL_X32 FILLER_40_3222 ();
 FILLCELL_X32 FILLER_40_3254 ();
 FILLCELL_X32 FILLER_40_3286 ();
 FILLCELL_X32 FILLER_40_3318 ();
 FILLCELL_X32 FILLER_40_3350 ();
 FILLCELL_X32 FILLER_40_3382 ();
 FILLCELL_X32 FILLER_40_3414 ();
 FILLCELL_X32 FILLER_40_3446 ();
 FILLCELL_X32 FILLER_40_3478 ();
 FILLCELL_X32 FILLER_40_3510 ();
 FILLCELL_X32 FILLER_40_3542 ();
 FILLCELL_X32 FILLER_40_3574 ();
 FILLCELL_X32 FILLER_40_3606 ();
 FILLCELL_X32 FILLER_40_3638 ();
 FILLCELL_X32 FILLER_40_3670 ();
 FILLCELL_X32 FILLER_40_3702 ();
 FILLCELL_X4 FILLER_40_3734 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X32 FILLER_41_321 ();
 FILLCELL_X32 FILLER_41_353 ();
 FILLCELL_X32 FILLER_41_385 ();
 FILLCELL_X32 FILLER_41_417 ();
 FILLCELL_X32 FILLER_41_449 ();
 FILLCELL_X32 FILLER_41_481 ();
 FILLCELL_X32 FILLER_41_513 ();
 FILLCELL_X32 FILLER_41_545 ();
 FILLCELL_X32 FILLER_41_577 ();
 FILLCELL_X32 FILLER_41_609 ();
 FILLCELL_X32 FILLER_41_641 ();
 FILLCELL_X32 FILLER_41_673 ();
 FILLCELL_X32 FILLER_41_705 ();
 FILLCELL_X32 FILLER_41_737 ();
 FILLCELL_X32 FILLER_41_769 ();
 FILLCELL_X32 FILLER_41_801 ();
 FILLCELL_X32 FILLER_41_833 ();
 FILLCELL_X32 FILLER_41_865 ();
 FILLCELL_X32 FILLER_41_897 ();
 FILLCELL_X32 FILLER_41_929 ();
 FILLCELL_X32 FILLER_41_961 ();
 FILLCELL_X32 FILLER_41_993 ();
 FILLCELL_X32 FILLER_41_1025 ();
 FILLCELL_X32 FILLER_41_1057 ();
 FILLCELL_X32 FILLER_41_1089 ();
 FILLCELL_X32 FILLER_41_1121 ();
 FILLCELL_X32 FILLER_41_1153 ();
 FILLCELL_X32 FILLER_41_1185 ();
 FILLCELL_X32 FILLER_41_1217 ();
 FILLCELL_X8 FILLER_41_1249 ();
 FILLCELL_X4 FILLER_41_1257 ();
 FILLCELL_X2 FILLER_41_1261 ();
 FILLCELL_X32 FILLER_41_1264 ();
 FILLCELL_X32 FILLER_41_1296 ();
 FILLCELL_X32 FILLER_41_1328 ();
 FILLCELL_X32 FILLER_41_1360 ();
 FILLCELL_X32 FILLER_41_1392 ();
 FILLCELL_X32 FILLER_41_1424 ();
 FILLCELL_X32 FILLER_41_1456 ();
 FILLCELL_X32 FILLER_41_1488 ();
 FILLCELL_X32 FILLER_41_1520 ();
 FILLCELL_X32 FILLER_41_1552 ();
 FILLCELL_X32 FILLER_41_1584 ();
 FILLCELL_X32 FILLER_41_1616 ();
 FILLCELL_X32 FILLER_41_1648 ();
 FILLCELL_X32 FILLER_41_1680 ();
 FILLCELL_X32 FILLER_41_1712 ();
 FILLCELL_X32 FILLER_41_1744 ();
 FILLCELL_X32 FILLER_41_1776 ();
 FILLCELL_X32 FILLER_41_1808 ();
 FILLCELL_X32 FILLER_41_1840 ();
 FILLCELL_X32 FILLER_41_1872 ();
 FILLCELL_X32 FILLER_41_1904 ();
 FILLCELL_X32 FILLER_41_1936 ();
 FILLCELL_X32 FILLER_41_1968 ();
 FILLCELL_X32 FILLER_41_2000 ();
 FILLCELL_X32 FILLER_41_2032 ();
 FILLCELL_X32 FILLER_41_2064 ();
 FILLCELL_X32 FILLER_41_2096 ();
 FILLCELL_X32 FILLER_41_2128 ();
 FILLCELL_X32 FILLER_41_2160 ();
 FILLCELL_X32 FILLER_41_2192 ();
 FILLCELL_X32 FILLER_41_2224 ();
 FILLCELL_X32 FILLER_41_2256 ();
 FILLCELL_X32 FILLER_41_2288 ();
 FILLCELL_X32 FILLER_41_2320 ();
 FILLCELL_X32 FILLER_41_2352 ();
 FILLCELL_X32 FILLER_41_2384 ();
 FILLCELL_X32 FILLER_41_2416 ();
 FILLCELL_X32 FILLER_41_2448 ();
 FILLCELL_X32 FILLER_41_2480 ();
 FILLCELL_X8 FILLER_41_2512 ();
 FILLCELL_X4 FILLER_41_2520 ();
 FILLCELL_X2 FILLER_41_2524 ();
 FILLCELL_X32 FILLER_41_2527 ();
 FILLCELL_X32 FILLER_41_2559 ();
 FILLCELL_X32 FILLER_41_2591 ();
 FILLCELL_X32 FILLER_41_2623 ();
 FILLCELL_X32 FILLER_41_2655 ();
 FILLCELL_X32 FILLER_41_2687 ();
 FILLCELL_X32 FILLER_41_2719 ();
 FILLCELL_X32 FILLER_41_2751 ();
 FILLCELL_X32 FILLER_41_2783 ();
 FILLCELL_X32 FILLER_41_2815 ();
 FILLCELL_X32 FILLER_41_2847 ();
 FILLCELL_X32 FILLER_41_2879 ();
 FILLCELL_X32 FILLER_41_2911 ();
 FILLCELL_X32 FILLER_41_2943 ();
 FILLCELL_X32 FILLER_41_2975 ();
 FILLCELL_X32 FILLER_41_3007 ();
 FILLCELL_X32 FILLER_41_3039 ();
 FILLCELL_X32 FILLER_41_3071 ();
 FILLCELL_X32 FILLER_41_3103 ();
 FILLCELL_X32 FILLER_41_3135 ();
 FILLCELL_X32 FILLER_41_3167 ();
 FILLCELL_X32 FILLER_41_3199 ();
 FILLCELL_X32 FILLER_41_3231 ();
 FILLCELL_X32 FILLER_41_3263 ();
 FILLCELL_X32 FILLER_41_3295 ();
 FILLCELL_X32 FILLER_41_3327 ();
 FILLCELL_X32 FILLER_41_3359 ();
 FILLCELL_X32 FILLER_41_3391 ();
 FILLCELL_X32 FILLER_41_3423 ();
 FILLCELL_X32 FILLER_41_3455 ();
 FILLCELL_X32 FILLER_41_3487 ();
 FILLCELL_X32 FILLER_41_3519 ();
 FILLCELL_X32 FILLER_41_3551 ();
 FILLCELL_X32 FILLER_41_3583 ();
 FILLCELL_X32 FILLER_41_3615 ();
 FILLCELL_X32 FILLER_41_3647 ();
 FILLCELL_X32 FILLER_41_3679 ();
 FILLCELL_X16 FILLER_41_3711 ();
 FILLCELL_X8 FILLER_41_3727 ();
 FILLCELL_X2 FILLER_41_3735 ();
 FILLCELL_X1 FILLER_41_3737 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X32 FILLER_42_321 ();
 FILLCELL_X32 FILLER_42_353 ();
 FILLCELL_X32 FILLER_42_385 ();
 FILLCELL_X32 FILLER_42_417 ();
 FILLCELL_X32 FILLER_42_449 ();
 FILLCELL_X32 FILLER_42_481 ();
 FILLCELL_X32 FILLER_42_513 ();
 FILLCELL_X32 FILLER_42_545 ();
 FILLCELL_X32 FILLER_42_577 ();
 FILLCELL_X16 FILLER_42_609 ();
 FILLCELL_X4 FILLER_42_625 ();
 FILLCELL_X2 FILLER_42_629 ();
 FILLCELL_X32 FILLER_42_632 ();
 FILLCELL_X32 FILLER_42_664 ();
 FILLCELL_X32 FILLER_42_696 ();
 FILLCELL_X32 FILLER_42_728 ();
 FILLCELL_X32 FILLER_42_760 ();
 FILLCELL_X32 FILLER_42_792 ();
 FILLCELL_X32 FILLER_42_824 ();
 FILLCELL_X32 FILLER_42_856 ();
 FILLCELL_X32 FILLER_42_888 ();
 FILLCELL_X32 FILLER_42_920 ();
 FILLCELL_X32 FILLER_42_952 ();
 FILLCELL_X32 FILLER_42_984 ();
 FILLCELL_X32 FILLER_42_1016 ();
 FILLCELL_X32 FILLER_42_1048 ();
 FILLCELL_X32 FILLER_42_1080 ();
 FILLCELL_X32 FILLER_42_1112 ();
 FILLCELL_X32 FILLER_42_1144 ();
 FILLCELL_X32 FILLER_42_1176 ();
 FILLCELL_X32 FILLER_42_1208 ();
 FILLCELL_X32 FILLER_42_1240 ();
 FILLCELL_X32 FILLER_42_1272 ();
 FILLCELL_X32 FILLER_42_1304 ();
 FILLCELL_X32 FILLER_42_1336 ();
 FILLCELL_X32 FILLER_42_1368 ();
 FILLCELL_X32 FILLER_42_1400 ();
 FILLCELL_X32 FILLER_42_1432 ();
 FILLCELL_X32 FILLER_42_1464 ();
 FILLCELL_X32 FILLER_42_1496 ();
 FILLCELL_X32 FILLER_42_1528 ();
 FILLCELL_X32 FILLER_42_1560 ();
 FILLCELL_X32 FILLER_42_1592 ();
 FILLCELL_X32 FILLER_42_1624 ();
 FILLCELL_X32 FILLER_42_1656 ();
 FILLCELL_X32 FILLER_42_1688 ();
 FILLCELL_X32 FILLER_42_1720 ();
 FILLCELL_X32 FILLER_42_1752 ();
 FILLCELL_X32 FILLER_42_1784 ();
 FILLCELL_X32 FILLER_42_1816 ();
 FILLCELL_X32 FILLER_42_1848 ();
 FILLCELL_X8 FILLER_42_1880 ();
 FILLCELL_X4 FILLER_42_1888 ();
 FILLCELL_X2 FILLER_42_1892 ();
 FILLCELL_X32 FILLER_42_1895 ();
 FILLCELL_X32 FILLER_42_1927 ();
 FILLCELL_X32 FILLER_42_1959 ();
 FILLCELL_X32 FILLER_42_1991 ();
 FILLCELL_X32 FILLER_42_2023 ();
 FILLCELL_X32 FILLER_42_2055 ();
 FILLCELL_X32 FILLER_42_2087 ();
 FILLCELL_X32 FILLER_42_2119 ();
 FILLCELL_X32 FILLER_42_2151 ();
 FILLCELL_X32 FILLER_42_2183 ();
 FILLCELL_X32 FILLER_42_2215 ();
 FILLCELL_X32 FILLER_42_2247 ();
 FILLCELL_X32 FILLER_42_2279 ();
 FILLCELL_X32 FILLER_42_2311 ();
 FILLCELL_X32 FILLER_42_2343 ();
 FILLCELL_X32 FILLER_42_2375 ();
 FILLCELL_X32 FILLER_42_2407 ();
 FILLCELL_X32 FILLER_42_2439 ();
 FILLCELL_X32 FILLER_42_2471 ();
 FILLCELL_X32 FILLER_42_2503 ();
 FILLCELL_X32 FILLER_42_2535 ();
 FILLCELL_X32 FILLER_42_2567 ();
 FILLCELL_X32 FILLER_42_2599 ();
 FILLCELL_X32 FILLER_42_2631 ();
 FILLCELL_X32 FILLER_42_2663 ();
 FILLCELL_X32 FILLER_42_2695 ();
 FILLCELL_X32 FILLER_42_2727 ();
 FILLCELL_X32 FILLER_42_2759 ();
 FILLCELL_X32 FILLER_42_2791 ();
 FILLCELL_X32 FILLER_42_2823 ();
 FILLCELL_X32 FILLER_42_2855 ();
 FILLCELL_X32 FILLER_42_2887 ();
 FILLCELL_X32 FILLER_42_2919 ();
 FILLCELL_X32 FILLER_42_2951 ();
 FILLCELL_X32 FILLER_42_2983 ();
 FILLCELL_X32 FILLER_42_3015 ();
 FILLCELL_X32 FILLER_42_3047 ();
 FILLCELL_X32 FILLER_42_3079 ();
 FILLCELL_X32 FILLER_42_3111 ();
 FILLCELL_X8 FILLER_42_3143 ();
 FILLCELL_X4 FILLER_42_3151 ();
 FILLCELL_X2 FILLER_42_3155 ();
 FILLCELL_X32 FILLER_42_3158 ();
 FILLCELL_X32 FILLER_42_3190 ();
 FILLCELL_X32 FILLER_42_3222 ();
 FILLCELL_X32 FILLER_42_3254 ();
 FILLCELL_X32 FILLER_42_3286 ();
 FILLCELL_X32 FILLER_42_3318 ();
 FILLCELL_X32 FILLER_42_3350 ();
 FILLCELL_X32 FILLER_42_3382 ();
 FILLCELL_X32 FILLER_42_3414 ();
 FILLCELL_X32 FILLER_42_3446 ();
 FILLCELL_X32 FILLER_42_3478 ();
 FILLCELL_X32 FILLER_42_3510 ();
 FILLCELL_X32 FILLER_42_3542 ();
 FILLCELL_X32 FILLER_42_3574 ();
 FILLCELL_X32 FILLER_42_3606 ();
 FILLCELL_X32 FILLER_42_3638 ();
 FILLCELL_X32 FILLER_42_3670 ();
 FILLCELL_X32 FILLER_42_3702 ();
 FILLCELL_X4 FILLER_42_3734 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X32 FILLER_43_193 ();
 FILLCELL_X32 FILLER_43_225 ();
 FILLCELL_X32 FILLER_43_257 ();
 FILLCELL_X32 FILLER_43_289 ();
 FILLCELL_X32 FILLER_43_321 ();
 FILLCELL_X32 FILLER_43_353 ();
 FILLCELL_X32 FILLER_43_385 ();
 FILLCELL_X32 FILLER_43_417 ();
 FILLCELL_X32 FILLER_43_449 ();
 FILLCELL_X32 FILLER_43_481 ();
 FILLCELL_X32 FILLER_43_513 ();
 FILLCELL_X32 FILLER_43_545 ();
 FILLCELL_X32 FILLER_43_577 ();
 FILLCELL_X32 FILLER_43_609 ();
 FILLCELL_X32 FILLER_43_641 ();
 FILLCELL_X32 FILLER_43_673 ();
 FILLCELL_X32 FILLER_43_705 ();
 FILLCELL_X32 FILLER_43_737 ();
 FILLCELL_X32 FILLER_43_769 ();
 FILLCELL_X32 FILLER_43_801 ();
 FILLCELL_X32 FILLER_43_833 ();
 FILLCELL_X32 FILLER_43_865 ();
 FILLCELL_X32 FILLER_43_897 ();
 FILLCELL_X32 FILLER_43_929 ();
 FILLCELL_X32 FILLER_43_961 ();
 FILLCELL_X32 FILLER_43_993 ();
 FILLCELL_X32 FILLER_43_1025 ();
 FILLCELL_X32 FILLER_43_1057 ();
 FILLCELL_X32 FILLER_43_1089 ();
 FILLCELL_X32 FILLER_43_1121 ();
 FILLCELL_X32 FILLER_43_1153 ();
 FILLCELL_X32 FILLER_43_1185 ();
 FILLCELL_X32 FILLER_43_1217 ();
 FILLCELL_X8 FILLER_43_1249 ();
 FILLCELL_X4 FILLER_43_1257 ();
 FILLCELL_X2 FILLER_43_1261 ();
 FILLCELL_X32 FILLER_43_1264 ();
 FILLCELL_X32 FILLER_43_1296 ();
 FILLCELL_X32 FILLER_43_1328 ();
 FILLCELL_X32 FILLER_43_1360 ();
 FILLCELL_X32 FILLER_43_1392 ();
 FILLCELL_X32 FILLER_43_1424 ();
 FILLCELL_X32 FILLER_43_1456 ();
 FILLCELL_X32 FILLER_43_1488 ();
 FILLCELL_X32 FILLER_43_1520 ();
 FILLCELL_X32 FILLER_43_1552 ();
 FILLCELL_X32 FILLER_43_1584 ();
 FILLCELL_X32 FILLER_43_1616 ();
 FILLCELL_X32 FILLER_43_1648 ();
 FILLCELL_X32 FILLER_43_1680 ();
 FILLCELL_X32 FILLER_43_1712 ();
 FILLCELL_X32 FILLER_43_1744 ();
 FILLCELL_X32 FILLER_43_1776 ();
 FILLCELL_X32 FILLER_43_1808 ();
 FILLCELL_X32 FILLER_43_1840 ();
 FILLCELL_X32 FILLER_43_1872 ();
 FILLCELL_X32 FILLER_43_1904 ();
 FILLCELL_X32 FILLER_43_1936 ();
 FILLCELL_X32 FILLER_43_1968 ();
 FILLCELL_X32 FILLER_43_2000 ();
 FILLCELL_X32 FILLER_43_2032 ();
 FILLCELL_X32 FILLER_43_2064 ();
 FILLCELL_X32 FILLER_43_2096 ();
 FILLCELL_X32 FILLER_43_2128 ();
 FILLCELL_X32 FILLER_43_2160 ();
 FILLCELL_X32 FILLER_43_2192 ();
 FILLCELL_X32 FILLER_43_2224 ();
 FILLCELL_X32 FILLER_43_2256 ();
 FILLCELL_X32 FILLER_43_2288 ();
 FILLCELL_X32 FILLER_43_2320 ();
 FILLCELL_X32 FILLER_43_2352 ();
 FILLCELL_X32 FILLER_43_2384 ();
 FILLCELL_X32 FILLER_43_2416 ();
 FILLCELL_X32 FILLER_43_2448 ();
 FILLCELL_X32 FILLER_43_2480 ();
 FILLCELL_X8 FILLER_43_2512 ();
 FILLCELL_X4 FILLER_43_2520 ();
 FILLCELL_X2 FILLER_43_2524 ();
 FILLCELL_X32 FILLER_43_2527 ();
 FILLCELL_X32 FILLER_43_2559 ();
 FILLCELL_X32 FILLER_43_2591 ();
 FILLCELL_X32 FILLER_43_2623 ();
 FILLCELL_X32 FILLER_43_2655 ();
 FILLCELL_X32 FILLER_43_2687 ();
 FILLCELL_X32 FILLER_43_2719 ();
 FILLCELL_X32 FILLER_43_2751 ();
 FILLCELL_X32 FILLER_43_2783 ();
 FILLCELL_X32 FILLER_43_2815 ();
 FILLCELL_X32 FILLER_43_2847 ();
 FILLCELL_X32 FILLER_43_2879 ();
 FILLCELL_X32 FILLER_43_2911 ();
 FILLCELL_X32 FILLER_43_2943 ();
 FILLCELL_X32 FILLER_43_2975 ();
 FILLCELL_X32 FILLER_43_3007 ();
 FILLCELL_X32 FILLER_43_3039 ();
 FILLCELL_X32 FILLER_43_3071 ();
 FILLCELL_X32 FILLER_43_3103 ();
 FILLCELL_X32 FILLER_43_3135 ();
 FILLCELL_X32 FILLER_43_3167 ();
 FILLCELL_X32 FILLER_43_3199 ();
 FILLCELL_X32 FILLER_43_3231 ();
 FILLCELL_X32 FILLER_43_3263 ();
 FILLCELL_X32 FILLER_43_3295 ();
 FILLCELL_X32 FILLER_43_3327 ();
 FILLCELL_X32 FILLER_43_3359 ();
 FILLCELL_X32 FILLER_43_3391 ();
 FILLCELL_X32 FILLER_43_3423 ();
 FILLCELL_X32 FILLER_43_3455 ();
 FILLCELL_X32 FILLER_43_3487 ();
 FILLCELL_X32 FILLER_43_3519 ();
 FILLCELL_X32 FILLER_43_3551 ();
 FILLCELL_X32 FILLER_43_3583 ();
 FILLCELL_X32 FILLER_43_3615 ();
 FILLCELL_X32 FILLER_43_3647 ();
 FILLCELL_X32 FILLER_43_3679 ();
 FILLCELL_X16 FILLER_43_3711 ();
 FILLCELL_X8 FILLER_43_3727 ();
 FILLCELL_X2 FILLER_43_3735 ();
 FILLCELL_X1 FILLER_43_3737 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X32 FILLER_44_193 ();
 FILLCELL_X32 FILLER_44_225 ();
 FILLCELL_X32 FILLER_44_257 ();
 FILLCELL_X32 FILLER_44_289 ();
 FILLCELL_X32 FILLER_44_321 ();
 FILLCELL_X32 FILLER_44_353 ();
 FILLCELL_X32 FILLER_44_385 ();
 FILLCELL_X32 FILLER_44_417 ();
 FILLCELL_X32 FILLER_44_449 ();
 FILLCELL_X32 FILLER_44_481 ();
 FILLCELL_X32 FILLER_44_513 ();
 FILLCELL_X32 FILLER_44_545 ();
 FILLCELL_X32 FILLER_44_577 ();
 FILLCELL_X16 FILLER_44_609 ();
 FILLCELL_X4 FILLER_44_625 ();
 FILLCELL_X2 FILLER_44_629 ();
 FILLCELL_X32 FILLER_44_632 ();
 FILLCELL_X32 FILLER_44_664 ();
 FILLCELL_X32 FILLER_44_696 ();
 FILLCELL_X32 FILLER_44_728 ();
 FILLCELL_X32 FILLER_44_760 ();
 FILLCELL_X32 FILLER_44_792 ();
 FILLCELL_X32 FILLER_44_824 ();
 FILLCELL_X32 FILLER_44_856 ();
 FILLCELL_X32 FILLER_44_888 ();
 FILLCELL_X32 FILLER_44_920 ();
 FILLCELL_X32 FILLER_44_952 ();
 FILLCELL_X32 FILLER_44_984 ();
 FILLCELL_X32 FILLER_44_1016 ();
 FILLCELL_X32 FILLER_44_1048 ();
 FILLCELL_X32 FILLER_44_1080 ();
 FILLCELL_X32 FILLER_44_1112 ();
 FILLCELL_X32 FILLER_44_1144 ();
 FILLCELL_X32 FILLER_44_1176 ();
 FILLCELL_X32 FILLER_44_1208 ();
 FILLCELL_X32 FILLER_44_1240 ();
 FILLCELL_X32 FILLER_44_1272 ();
 FILLCELL_X32 FILLER_44_1304 ();
 FILLCELL_X32 FILLER_44_1336 ();
 FILLCELL_X32 FILLER_44_1368 ();
 FILLCELL_X32 FILLER_44_1400 ();
 FILLCELL_X32 FILLER_44_1432 ();
 FILLCELL_X32 FILLER_44_1464 ();
 FILLCELL_X32 FILLER_44_1496 ();
 FILLCELL_X32 FILLER_44_1528 ();
 FILLCELL_X32 FILLER_44_1560 ();
 FILLCELL_X32 FILLER_44_1592 ();
 FILLCELL_X32 FILLER_44_1624 ();
 FILLCELL_X32 FILLER_44_1656 ();
 FILLCELL_X32 FILLER_44_1688 ();
 FILLCELL_X32 FILLER_44_1720 ();
 FILLCELL_X32 FILLER_44_1752 ();
 FILLCELL_X32 FILLER_44_1784 ();
 FILLCELL_X32 FILLER_44_1816 ();
 FILLCELL_X32 FILLER_44_1848 ();
 FILLCELL_X8 FILLER_44_1880 ();
 FILLCELL_X4 FILLER_44_1888 ();
 FILLCELL_X2 FILLER_44_1892 ();
 FILLCELL_X32 FILLER_44_1895 ();
 FILLCELL_X32 FILLER_44_1927 ();
 FILLCELL_X32 FILLER_44_1959 ();
 FILLCELL_X32 FILLER_44_1991 ();
 FILLCELL_X32 FILLER_44_2023 ();
 FILLCELL_X32 FILLER_44_2055 ();
 FILLCELL_X32 FILLER_44_2087 ();
 FILLCELL_X32 FILLER_44_2119 ();
 FILLCELL_X32 FILLER_44_2151 ();
 FILLCELL_X32 FILLER_44_2183 ();
 FILLCELL_X32 FILLER_44_2215 ();
 FILLCELL_X32 FILLER_44_2247 ();
 FILLCELL_X32 FILLER_44_2279 ();
 FILLCELL_X32 FILLER_44_2311 ();
 FILLCELL_X32 FILLER_44_2343 ();
 FILLCELL_X32 FILLER_44_2375 ();
 FILLCELL_X32 FILLER_44_2407 ();
 FILLCELL_X32 FILLER_44_2439 ();
 FILLCELL_X32 FILLER_44_2471 ();
 FILLCELL_X32 FILLER_44_2503 ();
 FILLCELL_X32 FILLER_44_2535 ();
 FILLCELL_X32 FILLER_44_2567 ();
 FILLCELL_X32 FILLER_44_2599 ();
 FILLCELL_X32 FILLER_44_2631 ();
 FILLCELL_X32 FILLER_44_2663 ();
 FILLCELL_X32 FILLER_44_2695 ();
 FILLCELL_X32 FILLER_44_2727 ();
 FILLCELL_X32 FILLER_44_2759 ();
 FILLCELL_X32 FILLER_44_2791 ();
 FILLCELL_X32 FILLER_44_2823 ();
 FILLCELL_X32 FILLER_44_2855 ();
 FILLCELL_X32 FILLER_44_2887 ();
 FILLCELL_X32 FILLER_44_2919 ();
 FILLCELL_X32 FILLER_44_2951 ();
 FILLCELL_X32 FILLER_44_2983 ();
 FILLCELL_X32 FILLER_44_3015 ();
 FILLCELL_X32 FILLER_44_3047 ();
 FILLCELL_X32 FILLER_44_3079 ();
 FILLCELL_X32 FILLER_44_3111 ();
 FILLCELL_X8 FILLER_44_3143 ();
 FILLCELL_X4 FILLER_44_3151 ();
 FILLCELL_X2 FILLER_44_3155 ();
 FILLCELL_X32 FILLER_44_3158 ();
 FILLCELL_X32 FILLER_44_3190 ();
 FILLCELL_X32 FILLER_44_3222 ();
 FILLCELL_X32 FILLER_44_3254 ();
 FILLCELL_X32 FILLER_44_3286 ();
 FILLCELL_X32 FILLER_44_3318 ();
 FILLCELL_X32 FILLER_44_3350 ();
 FILLCELL_X32 FILLER_44_3382 ();
 FILLCELL_X32 FILLER_44_3414 ();
 FILLCELL_X32 FILLER_44_3446 ();
 FILLCELL_X32 FILLER_44_3478 ();
 FILLCELL_X32 FILLER_44_3510 ();
 FILLCELL_X32 FILLER_44_3542 ();
 FILLCELL_X32 FILLER_44_3574 ();
 FILLCELL_X32 FILLER_44_3606 ();
 FILLCELL_X32 FILLER_44_3638 ();
 FILLCELL_X32 FILLER_44_3670 ();
 FILLCELL_X32 FILLER_44_3702 ();
 FILLCELL_X4 FILLER_44_3734 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X32 FILLER_45_161 ();
 FILLCELL_X32 FILLER_45_193 ();
 FILLCELL_X32 FILLER_45_225 ();
 FILLCELL_X32 FILLER_45_257 ();
 FILLCELL_X32 FILLER_45_289 ();
 FILLCELL_X32 FILLER_45_321 ();
 FILLCELL_X32 FILLER_45_353 ();
 FILLCELL_X32 FILLER_45_385 ();
 FILLCELL_X32 FILLER_45_417 ();
 FILLCELL_X32 FILLER_45_449 ();
 FILLCELL_X32 FILLER_45_481 ();
 FILLCELL_X32 FILLER_45_513 ();
 FILLCELL_X32 FILLER_45_545 ();
 FILLCELL_X32 FILLER_45_577 ();
 FILLCELL_X32 FILLER_45_609 ();
 FILLCELL_X32 FILLER_45_641 ();
 FILLCELL_X32 FILLER_45_673 ();
 FILLCELL_X32 FILLER_45_705 ();
 FILLCELL_X32 FILLER_45_737 ();
 FILLCELL_X32 FILLER_45_769 ();
 FILLCELL_X32 FILLER_45_801 ();
 FILLCELL_X32 FILLER_45_833 ();
 FILLCELL_X32 FILLER_45_865 ();
 FILLCELL_X32 FILLER_45_897 ();
 FILLCELL_X32 FILLER_45_929 ();
 FILLCELL_X32 FILLER_45_961 ();
 FILLCELL_X32 FILLER_45_993 ();
 FILLCELL_X32 FILLER_45_1025 ();
 FILLCELL_X32 FILLER_45_1057 ();
 FILLCELL_X32 FILLER_45_1089 ();
 FILLCELL_X32 FILLER_45_1121 ();
 FILLCELL_X32 FILLER_45_1153 ();
 FILLCELL_X32 FILLER_45_1185 ();
 FILLCELL_X32 FILLER_45_1217 ();
 FILLCELL_X8 FILLER_45_1249 ();
 FILLCELL_X4 FILLER_45_1257 ();
 FILLCELL_X2 FILLER_45_1261 ();
 FILLCELL_X32 FILLER_45_1264 ();
 FILLCELL_X32 FILLER_45_1296 ();
 FILLCELL_X32 FILLER_45_1328 ();
 FILLCELL_X32 FILLER_45_1360 ();
 FILLCELL_X32 FILLER_45_1392 ();
 FILLCELL_X32 FILLER_45_1424 ();
 FILLCELL_X32 FILLER_45_1456 ();
 FILLCELL_X32 FILLER_45_1488 ();
 FILLCELL_X32 FILLER_45_1520 ();
 FILLCELL_X32 FILLER_45_1552 ();
 FILLCELL_X32 FILLER_45_1584 ();
 FILLCELL_X32 FILLER_45_1616 ();
 FILLCELL_X32 FILLER_45_1648 ();
 FILLCELL_X32 FILLER_45_1680 ();
 FILLCELL_X32 FILLER_45_1712 ();
 FILLCELL_X32 FILLER_45_1744 ();
 FILLCELL_X32 FILLER_45_1776 ();
 FILLCELL_X32 FILLER_45_1808 ();
 FILLCELL_X32 FILLER_45_1840 ();
 FILLCELL_X32 FILLER_45_1872 ();
 FILLCELL_X32 FILLER_45_1904 ();
 FILLCELL_X32 FILLER_45_1936 ();
 FILLCELL_X32 FILLER_45_1968 ();
 FILLCELL_X32 FILLER_45_2000 ();
 FILLCELL_X32 FILLER_45_2032 ();
 FILLCELL_X32 FILLER_45_2064 ();
 FILLCELL_X32 FILLER_45_2096 ();
 FILLCELL_X32 FILLER_45_2128 ();
 FILLCELL_X32 FILLER_45_2160 ();
 FILLCELL_X32 FILLER_45_2192 ();
 FILLCELL_X32 FILLER_45_2224 ();
 FILLCELL_X32 FILLER_45_2256 ();
 FILLCELL_X32 FILLER_45_2288 ();
 FILLCELL_X32 FILLER_45_2320 ();
 FILLCELL_X32 FILLER_45_2352 ();
 FILLCELL_X32 FILLER_45_2384 ();
 FILLCELL_X32 FILLER_45_2416 ();
 FILLCELL_X32 FILLER_45_2448 ();
 FILLCELL_X32 FILLER_45_2480 ();
 FILLCELL_X8 FILLER_45_2512 ();
 FILLCELL_X4 FILLER_45_2520 ();
 FILLCELL_X2 FILLER_45_2524 ();
 FILLCELL_X32 FILLER_45_2527 ();
 FILLCELL_X32 FILLER_45_2559 ();
 FILLCELL_X32 FILLER_45_2591 ();
 FILLCELL_X32 FILLER_45_2623 ();
 FILLCELL_X32 FILLER_45_2655 ();
 FILLCELL_X32 FILLER_45_2687 ();
 FILLCELL_X32 FILLER_45_2719 ();
 FILLCELL_X32 FILLER_45_2751 ();
 FILLCELL_X32 FILLER_45_2783 ();
 FILLCELL_X32 FILLER_45_2815 ();
 FILLCELL_X32 FILLER_45_2847 ();
 FILLCELL_X32 FILLER_45_2879 ();
 FILLCELL_X32 FILLER_45_2911 ();
 FILLCELL_X32 FILLER_45_2943 ();
 FILLCELL_X32 FILLER_45_2975 ();
 FILLCELL_X32 FILLER_45_3007 ();
 FILLCELL_X32 FILLER_45_3039 ();
 FILLCELL_X32 FILLER_45_3071 ();
 FILLCELL_X32 FILLER_45_3103 ();
 FILLCELL_X32 FILLER_45_3135 ();
 FILLCELL_X32 FILLER_45_3167 ();
 FILLCELL_X32 FILLER_45_3199 ();
 FILLCELL_X32 FILLER_45_3231 ();
 FILLCELL_X32 FILLER_45_3263 ();
 FILLCELL_X32 FILLER_45_3295 ();
 FILLCELL_X32 FILLER_45_3327 ();
 FILLCELL_X32 FILLER_45_3359 ();
 FILLCELL_X32 FILLER_45_3391 ();
 FILLCELL_X32 FILLER_45_3423 ();
 FILLCELL_X32 FILLER_45_3455 ();
 FILLCELL_X32 FILLER_45_3487 ();
 FILLCELL_X32 FILLER_45_3519 ();
 FILLCELL_X32 FILLER_45_3551 ();
 FILLCELL_X32 FILLER_45_3583 ();
 FILLCELL_X32 FILLER_45_3615 ();
 FILLCELL_X32 FILLER_45_3647 ();
 FILLCELL_X32 FILLER_45_3679 ();
 FILLCELL_X16 FILLER_45_3711 ();
 FILLCELL_X8 FILLER_45_3727 ();
 FILLCELL_X2 FILLER_45_3735 ();
 FILLCELL_X1 FILLER_45_3737 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X32 FILLER_46_161 ();
 FILLCELL_X32 FILLER_46_193 ();
 FILLCELL_X32 FILLER_46_225 ();
 FILLCELL_X32 FILLER_46_257 ();
 FILLCELL_X32 FILLER_46_289 ();
 FILLCELL_X32 FILLER_46_321 ();
 FILLCELL_X32 FILLER_46_353 ();
 FILLCELL_X32 FILLER_46_385 ();
 FILLCELL_X32 FILLER_46_417 ();
 FILLCELL_X32 FILLER_46_449 ();
 FILLCELL_X32 FILLER_46_481 ();
 FILLCELL_X32 FILLER_46_513 ();
 FILLCELL_X32 FILLER_46_545 ();
 FILLCELL_X32 FILLER_46_577 ();
 FILLCELL_X16 FILLER_46_609 ();
 FILLCELL_X4 FILLER_46_625 ();
 FILLCELL_X2 FILLER_46_629 ();
 FILLCELL_X32 FILLER_46_632 ();
 FILLCELL_X32 FILLER_46_664 ();
 FILLCELL_X32 FILLER_46_696 ();
 FILLCELL_X32 FILLER_46_728 ();
 FILLCELL_X32 FILLER_46_760 ();
 FILLCELL_X32 FILLER_46_792 ();
 FILLCELL_X32 FILLER_46_824 ();
 FILLCELL_X32 FILLER_46_856 ();
 FILLCELL_X32 FILLER_46_888 ();
 FILLCELL_X32 FILLER_46_920 ();
 FILLCELL_X32 FILLER_46_952 ();
 FILLCELL_X32 FILLER_46_984 ();
 FILLCELL_X32 FILLER_46_1016 ();
 FILLCELL_X32 FILLER_46_1048 ();
 FILLCELL_X32 FILLER_46_1080 ();
 FILLCELL_X32 FILLER_46_1112 ();
 FILLCELL_X32 FILLER_46_1144 ();
 FILLCELL_X32 FILLER_46_1176 ();
 FILLCELL_X32 FILLER_46_1208 ();
 FILLCELL_X32 FILLER_46_1240 ();
 FILLCELL_X32 FILLER_46_1272 ();
 FILLCELL_X32 FILLER_46_1304 ();
 FILLCELL_X32 FILLER_46_1336 ();
 FILLCELL_X32 FILLER_46_1368 ();
 FILLCELL_X32 FILLER_46_1400 ();
 FILLCELL_X32 FILLER_46_1432 ();
 FILLCELL_X32 FILLER_46_1464 ();
 FILLCELL_X32 FILLER_46_1496 ();
 FILLCELL_X32 FILLER_46_1528 ();
 FILLCELL_X32 FILLER_46_1560 ();
 FILLCELL_X32 FILLER_46_1592 ();
 FILLCELL_X32 FILLER_46_1624 ();
 FILLCELL_X32 FILLER_46_1656 ();
 FILLCELL_X32 FILLER_46_1688 ();
 FILLCELL_X32 FILLER_46_1720 ();
 FILLCELL_X32 FILLER_46_1752 ();
 FILLCELL_X32 FILLER_46_1784 ();
 FILLCELL_X32 FILLER_46_1816 ();
 FILLCELL_X32 FILLER_46_1848 ();
 FILLCELL_X8 FILLER_46_1880 ();
 FILLCELL_X4 FILLER_46_1888 ();
 FILLCELL_X2 FILLER_46_1892 ();
 FILLCELL_X32 FILLER_46_1895 ();
 FILLCELL_X32 FILLER_46_1927 ();
 FILLCELL_X32 FILLER_46_1959 ();
 FILLCELL_X32 FILLER_46_1991 ();
 FILLCELL_X32 FILLER_46_2023 ();
 FILLCELL_X32 FILLER_46_2055 ();
 FILLCELL_X32 FILLER_46_2087 ();
 FILLCELL_X32 FILLER_46_2119 ();
 FILLCELL_X32 FILLER_46_2151 ();
 FILLCELL_X32 FILLER_46_2183 ();
 FILLCELL_X32 FILLER_46_2215 ();
 FILLCELL_X32 FILLER_46_2247 ();
 FILLCELL_X32 FILLER_46_2279 ();
 FILLCELL_X32 FILLER_46_2311 ();
 FILLCELL_X32 FILLER_46_2343 ();
 FILLCELL_X32 FILLER_46_2375 ();
 FILLCELL_X32 FILLER_46_2407 ();
 FILLCELL_X32 FILLER_46_2439 ();
 FILLCELL_X32 FILLER_46_2471 ();
 FILLCELL_X32 FILLER_46_2503 ();
 FILLCELL_X32 FILLER_46_2535 ();
 FILLCELL_X32 FILLER_46_2567 ();
 FILLCELL_X32 FILLER_46_2599 ();
 FILLCELL_X32 FILLER_46_2631 ();
 FILLCELL_X32 FILLER_46_2663 ();
 FILLCELL_X32 FILLER_46_2695 ();
 FILLCELL_X32 FILLER_46_2727 ();
 FILLCELL_X32 FILLER_46_2759 ();
 FILLCELL_X32 FILLER_46_2791 ();
 FILLCELL_X32 FILLER_46_2823 ();
 FILLCELL_X32 FILLER_46_2855 ();
 FILLCELL_X32 FILLER_46_2887 ();
 FILLCELL_X32 FILLER_46_2919 ();
 FILLCELL_X32 FILLER_46_2951 ();
 FILLCELL_X32 FILLER_46_2983 ();
 FILLCELL_X32 FILLER_46_3015 ();
 FILLCELL_X32 FILLER_46_3047 ();
 FILLCELL_X32 FILLER_46_3079 ();
 FILLCELL_X32 FILLER_46_3111 ();
 FILLCELL_X8 FILLER_46_3143 ();
 FILLCELL_X4 FILLER_46_3151 ();
 FILLCELL_X2 FILLER_46_3155 ();
 FILLCELL_X32 FILLER_46_3158 ();
 FILLCELL_X32 FILLER_46_3190 ();
 FILLCELL_X32 FILLER_46_3222 ();
 FILLCELL_X32 FILLER_46_3254 ();
 FILLCELL_X32 FILLER_46_3286 ();
 FILLCELL_X32 FILLER_46_3318 ();
 FILLCELL_X32 FILLER_46_3350 ();
 FILLCELL_X32 FILLER_46_3382 ();
 FILLCELL_X32 FILLER_46_3414 ();
 FILLCELL_X32 FILLER_46_3446 ();
 FILLCELL_X32 FILLER_46_3478 ();
 FILLCELL_X32 FILLER_46_3510 ();
 FILLCELL_X32 FILLER_46_3542 ();
 FILLCELL_X32 FILLER_46_3574 ();
 FILLCELL_X32 FILLER_46_3606 ();
 FILLCELL_X32 FILLER_46_3638 ();
 FILLCELL_X32 FILLER_46_3670 ();
 FILLCELL_X32 FILLER_46_3702 ();
 FILLCELL_X4 FILLER_46_3734 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X32 FILLER_47_129 ();
 FILLCELL_X32 FILLER_47_161 ();
 FILLCELL_X32 FILLER_47_193 ();
 FILLCELL_X32 FILLER_47_225 ();
 FILLCELL_X32 FILLER_47_257 ();
 FILLCELL_X32 FILLER_47_289 ();
 FILLCELL_X32 FILLER_47_321 ();
 FILLCELL_X32 FILLER_47_353 ();
 FILLCELL_X32 FILLER_47_385 ();
 FILLCELL_X32 FILLER_47_417 ();
 FILLCELL_X32 FILLER_47_449 ();
 FILLCELL_X32 FILLER_47_481 ();
 FILLCELL_X32 FILLER_47_513 ();
 FILLCELL_X32 FILLER_47_545 ();
 FILLCELL_X32 FILLER_47_577 ();
 FILLCELL_X32 FILLER_47_609 ();
 FILLCELL_X32 FILLER_47_641 ();
 FILLCELL_X32 FILLER_47_673 ();
 FILLCELL_X32 FILLER_47_705 ();
 FILLCELL_X32 FILLER_47_737 ();
 FILLCELL_X32 FILLER_47_769 ();
 FILLCELL_X32 FILLER_47_801 ();
 FILLCELL_X32 FILLER_47_833 ();
 FILLCELL_X32 FILLER_47_865 ();
 FILLCELL_X32 FILLER_47_897 ();
 FILLCELL_X32 FILLER_47_929 ();
 FILLCELL_X32 FILLER_47_961 ();
 FILLCELL_X32 FILLER_47_993 ();
 FILLCELL_X32 FILLER_47_1025 ();
 FILLCELL_X32 FILLER_47_1057 ();
 FILLCELL_X32 FILLER_47_1089 ();
 FILLCELL_X32 FILLER_47_1121 ();
 FILLCELL_X32 FILLER_47_1153 ();
 FILLCELL_X32 FILLER_47_1185 ();
 FILLCELL_X32 FILLER_47_1217 ();
 FILLCELL_X8 FILLER_47_1249 ();
 FILLCELL_X4 FILLER_47_1257 ();
 FILLCELL_X2 FILLER_47_1261 ();
 FILLCELL_X32 FILLER_47_1264 ();
 FILLCELL_X32 FILLER_47_1296 ();
 FILLCELL_X32 FILLER_47_1328 ();
 FILLCELL_X32 FILLER_47_1360 ();
 FILLCELL_X32 FILLER_47_1392 ();
 FILLCELL_X32 FILLER_47_1424 ();
 FILLCELL_X32 FILLER_47_1456 ();
 FILLCELL_X32 FILLER_47_1488 ();
 FILLCELL_X32 FILLER_47_1520 ();
 FILLCELL_X32 FILLER_47_1552 ();
 FILLCELL_X32 FILLER_47_1584 ();
 FILLCELL_X32 FILLER_47_1616 ();
 FILLCELL_X32 FILLER_47_1648 ();
 FILLCELL_X32 FILLER_47_1680 ();
 FILLCELL_X32 FILLER_47_1712 ();
 FILLCELL_X32 FILLER_47_1744 ();
 FILLCELL_X32 FILLER_47_1776 ();
 FILLCELL_X32 FILLER_47_1808 ();
 FILLCELL_X32 FILLER_47_1840 ();
 FILLCELL_X32 FILLER_47_1872 ();
 FILLCELL_X32 FILLER_47_1904 ();
 FILLCELL_X32 FILLER_47_1936 ();
 FILLCELL_X32 FILLER_47_1968 ();
 FILLCELL_X32 FILLER_47_2000 ();
 FILLCELL_X32 FILLER_47_2032 ();
 FILLCELL_X32 FILLER_47_2064 ();
 FILLCELL_X32 FILLER_47_2096 ();
 FILLCELL_X32 FILLER_47_2128 ();
 FILLCELL_X32 FILLER_47_2160 ();
 FILLCELL_X32 FILLER_47_2192 ();
 FILLCELL_X32 FILLER_47_2224 ();
 FILLCELL_X32 FILLER_47_2256 ();
 FILLCELL_X32 FILLER_47_2288 ();
 FILLCELL_X32 FILLER_47_2320 ();
 FILLCELL_X32 FILLER_47_2352 ();
 FILLCELL_X32 FILLER_47_2384 ();
 FILLCELL_X32 FILLER_47_2416 ();
 FILLCELL_X32 FILLER_47_2448 ();
 FILLCELL_X32 FILLER_47_2480 ();
 FILLCELL_X8 FILLER_47_2512 ();
 FILLCELL_X4 FILLER_47_2520 ();
 FILLCELL_X2 FILLER_47_2524 ();
 FILLCELL_X32 FILLER_47_2527 ();
 FILLCELL_X32 FILLER_47_2559 ();
 FILLCELL_X32 FILLER_47_2591 ();
 FILLCELL_X32 FILLER_47_2623 ();
 FILLCELL_X32 FILLER_47_2655 ();
 FILLCELL_X32 FILLER_47_2687 ();
 FILLCELL_X32 FILLER_47_2719 ();
 FILLCELL_X32 FILLER_47_2751 ();
 FILLCELL_X32 FILLER_47_2783 ();
 FILLCELL_X32 FILLER_47_2815 ();
 FILLCELL_X32 FILLER_47_2847 ();
 FILLCELL_X32 FILLER_47_2879 ();
 FILLCELL_X32 FILLER_47_2911 ();
 FILLCELL_X32 FILLER_47_2943 ();
 FILLCELL_X32 FILLER_47_2975 ();
 FILLCELL_X32 FILLER_47_3007 ();
 FILLCELL_X32 FILLER_47_3039 ();
 FILLCELL_X32 FILLER_47_3071 ();
 FILLCELL_X32 FILLER_47_3103 ();
 FILLCELL_X32 FILLER_47_3135 ();
 FILLCELL_X32 FILLER_47_3167 ();
 FILLCELL_X32 FILLER_47_3199 ();
 FILLCELL_X32 FILLER_47_3231 ();
 FILLCELL_X32 FILLER_47_3263 ();
 FILLCELL_X32 FILLER_47_3295 ();
 FILLCELL_X32 FILLER_47_3327 ();
 FILLCELL_X32 FILLER_47_3359 ();
 FILLCELL_X32 FILLER_47_3391 ();
 FILLCELL_X32 FILLER_47_3423 ();
 FILLCELL_X32 FILLER_47_3455 ();
 FILLCELL_X32 FILLER_47_3487 ();
 FILLCELL_X32 FILLER_47_3519 ();
 FILLCELL_X32 FILLER_47_3551 ();
 FILLCELL_X32 FILLER_47_3583 ();
 FILLCELL_X32 FILLER_47_3615 ();
 FILLCELL_X32 FILLER_47_3647 ();
 FILLCELL_X32 FILLER_47_3679 ();
 FILLCELL_X16 FILLER_47_3711 ();
 FILLCELL_X8 FILLER_47_3727 ();
 FILLCELL_X2 FILLER_47_3735 ();
 FILLCELL_X1 FILLER_47_3737 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X32 FILLER_48_65 ();
 FILLCELL_X32 FILLER_48_97 ();
 FILLCELL_X32 FILLER_48_129 ();
 FILLCELL_X32 FILLER_48_161 ();
 FILLCELL_X32 FILLER_48_193 ();
 FILLCELL_X32 FILLER_48_225 ();
 FILLCELL_X32 FILLER_48_257 ();
 FILLCELL_X32 FILLER_48_289 ();
 FILLCELL_X32 FILLER_48_321 ();
 FILLCELL_X32 FILLER_48_353 ();
 FILLCELL_X32 FILLER_48_385 ();
 FILLCELL_X32 FILLER_48_417 ();
 FILLCELL_X32 FILLER_48_449 ();
 FILLCELL_X32 FILLER_48_481 ();
 FILLCELL_X32 FILLER_48_513 ();
 FILLCELL_X32 FILLER_48_545 ();
 FILLCELL_X32 FILLER_48_577 ();
 FILLCELL_X16 FILLER_48_609 ();
 FILLCELL_X4 FILLER_48_625 ();
 FILLCELL_X2 FILLER_48_629 ();
 FILLCELL_X32 FILLER_48_632 ();
 FILLCELL_X32 FILLER_48_664 ();
 FILLCELL_X32 FILLER_48_696 ();
 FILLCELL_X32 FILLER_48_728 ();
 FILLCELL_X32 FILLER_48_760 ();
 FILLCELL_X32 FILLER_48_792 ();
 FILLCELL_X32 FILLER_48_824 ();
 FILLCELL_X32 FILLER_48_856 ();
 FILLCELL_X32 FILLER_48_888 ();
 FILLCELL_X32 FILLER_48_920 ();
 FILLCELL_X32 FILLER_48_952 ();
 FILLCELL_X32 FILLER_48_984 ();
 FILLCELL_X32 FILLER_48_1016 ();
 FILLCELL_X32 FILLER_48_1048 ();
 FILLCELL_X32 FILLER_48_1080 ();
 FILLCELL_X32 FILLER_48_1112 ();
 FILLCELL_X32 FILLER_48_1144 ();
 FILLCELL_X32 FILLER_48_1176 ();
 FILLCELL_X32 FILLER_48_1208 ();
 FILLCELL_X32 FILLER_48_1240 ();
 FILLCELL_X32 FILLER_48_1272 ();
 FILLCELL_X32 FILLER_48_1304 ();
 FILLCELL_X32 FILLER_48_1336 ();
 FILLCELL_X32 FILLER_48_1368 ();
 FILLCELL_X32 FILLER_48_1400 ();
 FILLCELL_X32 FILLER_48_1432 ();
 FILLCELL_X32 FILLER_48_1464 ();
 FILLCELL_X32 FILLER_48_1496 ();
 FILLCELL_X32 FILLER_48_1528 ();
 FILLCELL_X32 FILLER_48_1560 ();
 FILLCELL_X32 FILLER_48_1592 ();
 FILLCELL_X32 FILLER_48_1624 ();
 FILLCELL_X32 FILLER_48_1656 ();
 FILLCELL_X32 FILLER_48_1688 ();
 FILLCELL_X32 FILLER_48_1720 ();
 FILLCELL_X32 FILLER_48_1752 ();
 FILLCELL_X32 FILLER_48_1784 ();
 FILLCELL_X32 FILLER_48_1816 ();
 FILLCELL_X32 FILLER_48_1848 ();
 FILLCELL_X8 FILLER_48_1880 ();
 FILLCELL_X4 FILLER_48_1888 ();
 FILLCELL_X2 FILLER_48_1892 ();
 FILLCELL_X32 FILLER_48_1895 ();
 FILLCELL_X32 FILLER_48_1927 ();
 FILLCELL_X32 FILLER_48_1959 ();
 FILLCELL_X32 FILLER_48_1991 ();
 FILLCELL_X32 FILLER_48_2023 ();
 FILLCELL_X32 FILLER_48_2055 ();
 FILLCELL_X32 FILLER_48_2087 ();
 FILLCELL_X32 FILLER_48_2119 ();
 FILLCELL_X32 FILLER_48_2151 ();
 FILLCELL_X32 FILLER_48_2183 ();
 FILLCELL_X32 FILLER_48_2215 ();
 FILLCELL_X32 FILLER_48_2247 ();
 FILLCELL_X32 FILLER_48_2279 ();
 FILLCELL_X32 FILLER_48_2311 ();
 FILLCELL_X32 FILLER_48_2343 ();
 FILLCELL_X32 FILLER_48_2375 ();
 FILLCELL_X32 FILLER_48_2407 ();
 FILLCELL_X32 FILLER_48_2439 ();
 FILLCELL_X32 FILLER_48_2471 ();
 FILLCELL_X32 FILLER_48_2503 ();
 FILLCELL_X32 FILLER_48_2535 ();
 FILLCELL_X32 FILLER_48_2567 ();
 FILLCELL_X32 FILLER_48_2599 ();
 FILLCELL_X32 FILLER_48_2631 ();
 FILLCELL_X32 FILLER_48_2663 ();
 FILLCELL_X32 FILLER_48_2695 ();
 FILLCELL_X32 FILLER_48_2727 ();
 FILLCELL_X32 FILLER_48_2759 ();
 FILLCELL_X32 FILLER_48_2791 ();
 FILLCELL_X32 FILLER_48_2823 ();
 FILLCELL_X32 FILLER_48_2855 ();
 FILLCELL_X32 FILLER_48_2887 ();
 FILLCELL_X32 FILLER_48_2919 ();
 FILLCELL_X32 FILLER_48_2951 ();
 FILLCELL_X32 FILLER_48_2983 ();
 FILLCELL_X32 FILLER_48_3015 ();
 FILLCELL_X32 FILLER_48_3047 ();
 FILLCELL_X32 FILLER_48_3079 ();
 FILLCELL_X32 FILLER_48_3111 ();
 FILLCELL_X8 FILLER_48_3143 ();
 FILLCELL_X4 FILLER_48_3151 ();
 FILLCELL_X2 FILLER_48_3155 ();
 FILLCELL_X32 FILLER_48_3158 ();
 FILLCELL_X32 FILLER_48_3190 ();
 FILLCELL_X32 FILLER_48_3222 ();
 FILLCELL_X32 FILLER_48_3254 ();
 FILLCELL_X32 FILLER_48_3286 ();
 FILLCELL_X32 FILLER_48_3318 ();
 FILLCELL_X32 FILLER_48_3350 ();
 FILLCELL_X32 FILLER_48_3382 ();
 FILLCELL_X32 FILLER_48_3414 ();
 FILLCELL_X32 FILLER_48_3446 ();
 FILLCELL_X32 FILLER_48_3478 ();
 FILLCELL_X32 FILLER_48_3510 ();
 FILLCELL_X32 FILLER_48_3542 ();
 FILLCELL_X32 FILLER_48_3574 ();
 FILLCELL_X32 FILLER_48_3606 ();
 FILLCELL_X32 FILLER_48_3638 ();
 FILLCELL_X32 FILLER_48_3670 ();
 FILLCELL_X32 FILLER_48_3702 ();
 FILLCELL_X4 FILLER_48_3734 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X32 FILLER_49_97 ();
 FILLCELL_X32 FILLER_49_129 ();
 FILLCELL_X32 FILLER_49_161 ();
 FILLCELL_X32 FILLER_49_193 ();
 FILLCELL_X32 FILLER_49_225 ();
 FILLCELL_X32 FILLER_49_257 ();
 FILLCELL_X32 FILLER_49_289 ();
 FILLCELL_X32 FILLER_49_321 ();
 FILLCELL_X32 FILLER_49_353 ();
 FILLCELL_X32 FILLER_49_385 ();
 FILLCELL_X32 FILLER_49_417 ();
 FILLCELL_X32 FILLER_49_449 ();
 FILLCELL_X32 FILLER_49_481 ();
 FILLCELL_X32 FILLER_49_513 ();
 FILLCELL_X32 FILLER_49_545 ();
 FILLCELL_X32 FILLER_49_577 ();
 FILLCELL_X32 FILLER_49_609 ();
 FILLCELL_X32 FILLER_49_641 ();
 FILLCELL_X32 FILLER_49_673 ();
 FILLCELL_X32 FILLER_49_705 ();
 FILLCELL_X32 FILLER_49_737 ();
 FILLCELL_X32 FILLER_49_769 ();
 FILLCELL_X32 FILLER_49_801 ();
 FILLCELL_X32 FILLER_49_833 ();
 FILLCELL_X32 FILLER_49_865 ();
 FILLCELL_X32 FILLER_49_897 ();
 FILLCELL_X32 FILLER_49_929 ();
 FILLCELL_X32 FILLER_49_961 ();
 FILLCELL_X32 FILLER_49_993 ();
 FILLCELL_X32 FILLER_49_1025 ();
 FILLCELL_X32 FILLER_49_1057 ();
 FILLCELL_X32 FILLER_49_1089 ();
 FILLCELL_X32 FILLER_49_1121 ();
 FILLCELL_X32 FILLER_49_1153 ();
 FILLCELL_X32 FILLER_49_1185 ();
 FILLCELL_X32 FILLER_49_1217 ();
 FILLCELL_X8 FILLER_49_1249 ();
 FILLCELL_X4 FILLER_49_1257 ();
 FILLCELL_X2 FILLER_49_1261 ();
 FILLCELL_X32 FILLER_49_1264 ();
 FILLCELL_X32 FILLER_49_1296 ();
 FILLCELL_X32 FILLER_49_1328 ();
 FILLCELL_X32 FILLER_49_1360 ();
 FILLCELL_X32 FILLER_49_1392 ();
 FILLCELL_X32 FILLER_49_1424 ();
 FILLCELL_X32 FILLER_49_1456 ();
 FILLCELL_X32 FILLER_49_1488 ();
 FILLCELL_X32 FILLER_49_1520 ();
 FILLCELL_X32 FILLER_49_1552 ();
 FILLCELL_X32 FILLER_49_1584 ();
 FILLCELL_X32 FILLER_49_1616 ();
 FILLCELL_X32 FILLER_49_1648 ();
 FILLCELL_X32 FILLER_49_1680 ();
 FILLCELL_X32 FILLER_49_1712 ();
 FILLCELL_X32 FILLER_49_1744 ();
 FILLCELL_X32 FILLER_49_1776 ();
 FILLCELL_X32 FILLER_49_1808 ();
 FILLCELL_X32 FILLER_49_1840 ();
 FILLCELL_X32 FILLER_49_1872 ();
 FILLCELL_X32 FILLER_49_1904 ();
 FILLCELL_X32 FILLER_49_1936 ();
 FILLCELL_X32 FILLER_49_1968 ();
 FILLCELL_X32 FILLER_49_2000 ();
 FILLCELL_X32 FILLER_49_2032 ();
 FILLCELL_X32 FILLER_49_2064 ();
 FILLCELL_X32 FILLER_49_2096 ();
 FILLCELL_X32 FILLER_49_2128 ();
 FILLCELL_X32 FILLER_49_2160 ();
 FILLCELL_X32 FILLER_49_2192 ();
 FILLCELL_X32 FILLER_49_2224 ();
 FILLCELL_X32 FILLER_49_2256 ();
 FILLCELL_X32 FILLER_49_2288 ();
 FILLCELL_X32 FILLER_49_2320 ();
 FILLCELL_X32 FILLER_49_2352 ();
 FILLCELL_X32 FILLER_49_2384 ();
 FILLCELL_X32 FILLER_49_2416 ();
 FILLCELL_X32 FILLER_49_2448 ();
 FILLCELL_X32 FILLER_49_2480 ();
 FILLCELL_X8 FILLER_49_2512 ();
 FILLCELL_X4 FILLER_49_2520 ();
 FILLCELL_X2 FILLER_49_2524 ();
 FILLCELL_X32 FILLER_49_2527 ();
 FILLCELL_X32 FILLER_49_2559 ();
 FILLCELL_X32 FILLER_49_2591 ();
 FILLCELL_X32 FILLER_49_2623 ();
 FILLCELL_X32 FILLER_49_2655 ();
 FILLCELL_X32 FILLER_49_2687 ();
 FILLCELL_X32 FILLER_49_2719 ();
 FILLCELL_X32 FILLER_49_2751 ();
 FILLCELL_X32 FILLER_49_2783 ();
 FILLCELL_X32 FILLER_49_2815 ();
 FILLCELL_X32 FILLER_49_2847 ();
 FILLCELL_X32 FILLER_49_2879 ();
 FILLCELL_X32 FILLER_49_2911 ();
 FILLCELL_X32 FILLER_49_2943 ();
 FILLCELL_X32 FILLER_49_2975 ();
 FILLCELL_X32 FILLER_49_3007 ();
 FILLCELL_X32 FILLER_49_3039 ();
 FILLCELL_X32 FILLER_49_3071 ();
 FILLCELL_X32 FILLER_49_3103 ();
 FILLCELL_X32 FILLER_49_3135 ();
 FILLCELL_X32 FILLER_49_3167 ();
 FILLCELL_X32 FILLER_49_3199 ();
 FILLCELL_X32 FILLER_49_3231 ();
 FILLCELL_X32 FILLER_49_3263 ();
 FILLCELL_X32 FILLER_49_3295 ();
 FILLCELL_X32 FILLER_49_3327 ();
 FILLCELL_X32 FILLER_49_3359 ();
 FILLCELL_X32 FILLER_49_3391 ();
 FILLCELL_X32 FILLER_49_3423 ();
 FILLCELL_X32 FILLER_49_3455 ();
 FILLCELL_X32 FILLER_49_3487 ();
 FILLCELL_X32 FILLER_49_3519 ();
 FILLCELL_X32 FILLER_49_3551 ();
 FILLCELL_X32 FILLER_49_3583 ();
 FILLCELL_X32 FILLER_49_3615 ();
 FILLCELL_X32 FILLER_49_3647 ();
 FILLCELL_X32 FILLER_49_3679 ();
 FILLCELL_X16 FILLER_49_3711 ();
 FILLCELL_X8 FILLER_49_3727 ();
 FILLCELL_X2 FILLER_49_3735 ();
 FILLCELL_X1 FILLER_49_3737 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X32 FILLER_50_65 ();
 FILLCELL_X32 FILLER_50_97 ();
 FILLCELL_X32 FILLER_50_129 ();
 FILLCELL_X32 FILLER_50_161 ();
 FILLCELL_X32 FILLER_50_193 ();
 FILLCELL_X32 FILLER_50_225 ();
 FILLCELL_X32 FILLER_50_257 ();
 FILLCELL_X32 FILLER_50_289 ();
 FILLCELL_X32 FILLER_50_321 ();
 FILLCELL_X32 FILLER_50_353 ();
 FILLCELL_X32 FILLER_50_385 ();
 FILLCELL_X32 FILLER_50_417 ();
 FILLCELL_X32 FILLER_50_449 ();
 FILLCELL_X32 FILLER_50_481 ();
 FILLCELL_X32 FILLER_50_513 ();
 FILLCELL_X32 FILLER_50_545 ();
 FILLCELL_X32 FILLER_50_577 ();
 FILLCELL_X16 FILLER_50_609 ();
 FILLCELL_X4 FILLER_50_625 ();
 FILLCELL_X2 FILLER_50_629 ();
 FILLCELL_X32 FILLER_50_632 ();
 FILLCELL_X32 FILLER_50_664 ();
 FILLCELL_X32 FILLER_50_696 ();
 FILLCELL_X32 FILLER_50_728 ();
 FILLCELL_X32 FILLER_50_760 ();
 FILLCELL_X32 FILLER_50_792 ();
 FILLCELL_X32 FILLER_50_824 ();
 FILLCELL_X32 FILLER_50_856 ();
 FILLCELL_X32 FILLER_50_888 ();
 FILLCELL_X32 FILLER_50_920 ();
 FILLCELL_X32 FILLER_50_952 ();
 FILLCELL_X32 FILLER_50_984 ();
 FILLCELL_X32 FILLER_50_1016 ();
 FILLCELL_X32 FILLER_50_1048 ();
 FILLCELL_X32 FILLER_50_1080 ();
 FILLCELL_X32 FILLER_50_1112 ();
 FILLCELL_X32 FILLER_50_1144 ();
 FILLCELL_X32 FILLER_50_1176 ();
 FILLCELL_X32 FILLER_50_1208 ();
 FILLCELL_X32 FILLER_50_1240 ();
 FILLCELL_X32 FILLER_50_1272 ();
 FILLCELL_X32 FILLER_50_1304 ();
 FILLCELL_X32 FILLER_50_1336 ();
 FILLCELL_X32 FILLER_50_1368 ();
 FILLCELL_X32 FILLER_50_1400 ();
 FILLCELL_X32 FILLER_50_1432 ();
 FILLCELL_X32 FILLER_50_1464 ();
 FILLCELL_X32 FILLER_50_1496 ();
 FILLCELL_X32 FILLER_50_1528 ();
 FILLCELL_X32 FILLER_50_1560 ();
 FILLCELL_X32 FILLER_50_1592 ();
 FILLCELL_X32 FILLER_50_1624 ();
 FILLCELL_X32 FILLER_50_1656 ();
 FILLCELL_X32 FILLER_50_1688 ();
 FILLCELL_X32 FILLER_50_1720 ();
 FILLCELL_X32 FILLER_50_1752 ();
 FILLCELL_X32 FILLER_50_1784 ();
 FILLCELL_X32 FILLER_50_1816 ();
 FILLCELL_X32 FILLER_50_1848 ();
 FILLCELL_X8 FILLER_50_1880 ();
 FILLCELL_X4 FILLER_50_1888 ();
 FILLCELL_X2 FILLER_50_1892 ();
 FILLCELL_X32 FILLER_50_1895 ();
 FILLCELL_X32 FILLER_50_1927 ();
 FILLCELL_X32 FILLER_50_1959 ();
 FILLCELL_X32 FILLER_50_1991 ();
 FILLCELL_X32 FILLER_50_2023 ();
 FILLCELL_X32 FILLER_50_2055 ();
 FILLCELL_X32 FILLER_50_2087 ();
 FILLCELL_X32 FILLER_50_2119 ();
 FILLCELL_X32 FILLER_50_2151 ();
 FILLCELL_X32 FILLER_50_2183 ();
 FILLCELL_X32 FILLER_50_2215 ();
 FILLCELL_X32 FILLER_50_2247 ();
 FILLCELL_X32 FILLER_50_2279 ();
 FILLCELL_X32 FILLER_50_2311 ();
 FILLCELL_X32 FILLER_50_2343 ();
 FILLCELL_X32 FILLER_50_2375 ();
 FILLCELL_X32 FILLER_50_2407 ();
 FILLCELL_X32 FILLER_50_2439 ();
 FILLCELL_X32 FILLER_50_2471 ();
 FILLCELL_X32 FILLER_50_2503 ();
 FILLCELL_X32 FILLER_50_2535 ();
 FILLCELL_X32 FILLER_50_2567 ();
 FILLCELL_X32 FILLER_50_2599 ();
 FILLCELL_X32 FILLER_50_2631 ();
 FILLCELL_X32 FILLER_50_2663 ();
 FILLCELL_X32 FILLER_50_2695 ();
 FILLCELL_X32 FILLER_50_2727 ();
 FILLCELL_X32 FILLER_50_2759 ();
 FILLCELL_X32 FILLER_50_2791 ();
 FILLCELL_X32 FILLER_50_2823 ();
 FILLCELL_X32 FILLER_50_2855 ();
 FILLCELL_X32 FILLER_50_2887 ();
 FILLCELL_X32 FILLER_50_2919 ();
 FILLCELL_X32 FILLER_50_2951 ();
 FILLCELL_X32 FILLER_50_2983 ();
 FILLCELL_X32 FILLER_50_3015 ();
 FILLCELL_X32 FILLER_50_3047 ();
 FILLCELL_X32 FILLER_50_3079 ();
 FILLCELL_X32 FILLER_50_3111 ();
 FILLCELL_X8 FILLER_50_3143 ();
 FILLCELL_X4 FILLER_50_3151 ();
 FILLCELL_X2 FILLER_50_3155 ();
 FILLCELL_X32 FILLER_50_3158 ();
 FILLCELL_X32 FILLER_50_3190 ();
 FILLCELL_X32 FILLER_50_3222 ();
 FILLCELL_X32 FILLER_50_3254 ();
 FILLCELL_X32 FILLER_50_3286 ();
 FILLCELL_X32 FILLER_50_3318 ();
 FILLCELL_X32 FILLER_50_3350 ();
 FILLCELL_X32 FILLER_50_3382 ();
 FILLCELL_X32 FILLER_50_3414 ();
 FILLCELL_X32 FILLER_50_3446 ();
 FILLCELL_X32 FILLER_50_3478 ();
 FILLCELL_X32 FILLER_50_3510 ();
 FILLCELL_X32 FILLER_50_3542 ();
 FILLCELL_X32 FILLER_50_3574 ();
 FILLCELL_X32 FILLER_50_3606 ();
 FILLCELL_X32 FILLER_50_3638 ();
 FILLCELL_X32 FILLER_50_3670 ();
 FILLCELL_X32 FILLER_50_3702 ();
 FILLCELL_X4 FILLER_50_3734 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X32 FILLER_51_65 ();
 FILLCELL_X32 FILLER_51_97 ();
 FILLCELL_X32 FILLER_51_129 ();
 FILLCELL_X32 FILLER_51_161 ();
 FILLCELL_X32 FILLER_51_193 ();
 FILLCELL_X32 FILLER_51_225 ();
 FILLCELL_X32 FILLER_51_257 ();
 FILLCELL_X32 FILLER_51_289 ();
 FILLCELL_X32 FILLER_51_321 ();
 FILLCELL_X32 FILLER_51_353 ();
 FILLCELL_X32 FILLER_51_385 ();
 FILLCELL_X32 FILLER_51_417 ();
 FILLCELL_X32 FILLER_51_449 ();
 FILLCELL_X32 FILLER_51_481 ();
 FILLCELL_X32 FILLER_51_513 ();
 FILLCELL_X32 FILLER_51_545 ();
 FILLCELL_X32 FILLER_51_577 ();
 FILLCELL_X32 FILLER_51_609 ();
 FILLCELL_X32 FILLER_51_641 ();
 FILLCELL_X32 FILLER_51_673 ();
 FILLCELL_X32 FILLER_51_705 ();
 FILLCELL_X32 FILLER_51_737 ();
 FILLCELL_X32 FILLER_51_769 ();
 FILLCELL_X32 FILLER_51_801 ();
 FILLCELL_X32 FILLER_51_833 ();
 FILLCELL_X32 FILLER_51_865 ();
 FILLCELL_X32 FILLER_51_897 ();
 FILLCELL_X32 FILLER_51_929 ();
 FILLCELL_X32 FILLER_51_961 ();
 FILLCELL_X32 FILLER_51_993 ();
 FILLCELL_X32 FILLER_51_1025 ();
 FILLCELL_X32 FILLER_51_1057 ();
 FILLCELL_X32 FILLER_51_1089 ();
 FILLCELL_X32 FILLER_51_1121 ();
 FILLCELL_X32 FILLER_51_1153 ();
 FILLCELL_X32 FILLER_51_1185 ();
 FILLCELL_X32 FILLER_51_1217 ();
 FILLCELL_X8 FILLER_51_1249 ();
 FILLCELL_X4 FILLER_51_1257 ();
 FILLCELL_X2 FILLER_51_1261 ();
 FILLCELL_X32 FILLER_51_1264 ();
 FILLCELL_X32 FILLER_51_1296 ();
 FILLCELL_X32 FILLER_51_1328 ();
 FILLCELL_X32 FILLER_51_1360 ();
 FILLCELL_X32 FILLER_51_1392 ();
 FILLCELL_X32 FILLER_51_1424 ();
 FILLCELL_X32 FILLER_51_1456 ();
 FILLCELL_X32 FILLER_51_1488 ();
 FILLCELL_X32 FILLER_51_1520 ();
 FILLCELL_X32 FILLER_51_1552 ();
 FILLCELL_X32 FILLER_51_1584 ();
 FILLCELL_X32 FILLER_51_1616 ();
 FILLCELL_X32 FILLER_51_1648 ();
 FILLCELL_X32 FILLER_51_1680 ();
 FILLCELL_X32 FILLER_51_1712 ();
 FILLCELL_X32 FILLER_51_1744 ();
 FILLCELL_X32 FILLER_51_1776 ();
 FILLCELL_X32 FILLER_51_1808 ();
 FILLCELL_X32 FILLER_51_1840 ();
 FILLCELL_X32 FILLER_51_1872 ();
 FILLCELL_X32 FILLER_51_1904 ();
 FILLCELL_X32 FILLER_51_1936 ();
 FILLCELL_X32 FILLER_51_1968 ();
 FILLCELL_X32 FILLER_51_2000 ();
 FILLCELL_X32 FILLER_51_2032 ();
 FILLCELL_X32 FILLER_51_2064 ();
 FILLCELL_X32 FILLER_51_2096 ();
 FILLCELL_X32 FILLER_51_2128 ();
 FILLCELL_X32 FILLER_51_2160 ();
 FILLCELL_X32 FILLER_51_2192 ();
 FILLCELL_X32 FILLER_51_2224 ();
 FILLCELL_X32 FILLER_51_2256 ();
 FILLCELL_X32 FILLER_51_2288 ();
 FILLCELL_X32 FILLER_51_2320 ();
 FILLCELL_X32 FILLER_51_2352 ();
 FILLCELL_X32 FILLER_51_2384 ();
 FILLCELL_X32 FILLER_51_2416 ();
 FILLCELL_X32 FILLER_51_2448 ();
 FILLCELL_X32 FILLER_51_2480 ();
 FILLCELL_X8 FILLER_51_2512 ();
 FILLCELL_X4 FILLER_51_2520 ();
 FILLCELL_X2 FILLER_51_2524 ();
 FILLCELL_X32 FILLER_51_2527 ();
 FILLCELL_X32 FILLER_51_2559 ();
 FILLCELL_X32 FILLER_51_2591 ();
 FILLCELL_X32 FILLER_51_2623 ();
 FILLCELL_X32 FILLER_51_2655 ();
 FILLCELL_X32 FILLER_51_2687 ();
 FILLCELL_X32 FILLER_51_2719 ();
 FILLCELL_X32 FILLER_51_2751 ();
 FILLCELL_X32 FILLER_51_2783 ();
 FILLCELL_X32 FILLER_51_2815 ();
 FILLCELL_X32 FILLER_51_2847 ();
 FILLCELL_X32 FILLER_51_2879 ();
 FILLCELL_X32 FILLER_51_2911 ();
 FILLCELL_X32 FILLER_51_2943 ();
 FILLCELL_X32 FILLER_51_2975 ();
 FILLCELL_X32 FILLER_51_3007 ();
 FILLCELL_X32 FILLER_51_3039 ();
 FILLCELL_X32 FILLER_51_3071 ();
 FILLCELL_X32 FILLER_51_3103 ();
 FILLCELL_X32 FILLER_51_3135 ();
 FILLCELL_X32 FILLER_51_3167 ();
 FILLCELL_X32 FILLER_51_3199 ();
 FILLCELL_X32 FILLER_51_3231 ();
 FILLCELL_X32 FILLER_51_3263 ();
 FILLCELL_X32 FILLER_51_3295 ();
 FILLCELL_X32 FILLER_51_3327 ();
 FILLCELL_X32 FILLER_51_3359 ();
 FILLCELL_X32 FILLER_51_3391 ();
 FILLCELL_X32 FILLER_51_3423 ();
 FILLCELL_X32 FILLER_51_3455 ();
 FILLCELL_X32 FILLER_51_3487 ();
 FILLCELL_X32 FILLER_51_3519 ();
 FILLCELL_X32 FILLER_51_3551 ();
 FILLCELL_X32 FILLER_51_3583 ();
 FILLCELL_X32 FILLER_51_3615 ();
 FILLCELL_X32 FILLER_51_3647 ();
 FILLCELL_X32 FILLER_51_3679 ();
 FILLCELL_X16 FILLER_51_3711 ();
 FILLCELL_X8 FILLER_51_3727 ();
 FILLCELL_X2 FILLER_51_3735 ();
 FILLCELL_X1 FILLER_51_3737 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X32 FILLER_52_65 ();
 FILLCELL_X32 FILLER_52_97 ();
 FILLCELL_X32 FILLER_52_129 ();
 FILLCELL_X32 FILLER_52_161 ();
 FILLCELL_X32 FILLER_52_193 ();
 FILLCELL_X32 FILLER_52_225 ();
 FILLCELL_X32 FILLER_52_257 ();
 FILLCELL_X32 FILLER_52_289 ();
 FILLCELL_X32 FILLER_52_321 ();
 FILLCELL_X32 FILLER_52_353 ();
 FILLCELL_X32 FILLER_52_385 ();
 FILLCELL_X32 FILLER_52_417 ();
 FILLCELL_X32 FILLER_52_449 ();
 FILLCELL_X32 FILLER_52_481 ();
 FILLCELL_X32 FILLER_52_513 ();
 FILLCELL_X32 FILLER_52_545 ();
 FILLCELL_X32 FILLER_52_577 ();
 FILLCELL_X16 FILLER_52_609 ();
 FILLCELL_X4 FILLER_52_625 ();
 FILLCELL_X2 FILLER_52_629 ();
 FILLCELL_X32 FILLER_52_632 ();
 FILLCELL_X32 FILLER_52_664 ();
 FILLCELL_X32 FILLER_52_696 ();
 FILLCELL_X32 FILLER_52_728 ();
 FILLCELL_X32 FILLER_52_760 ();
 FILLCELL_X32 FILLER_52_792 ();
 FILLCELL_X32 FILLER_52_824 ();
 FILLCELL_X32 FILLER_52_856 ();
 FILLCELL_X32 FILLER_52_888 ();
 FILLCELL_X32 FILLER_52_920 ();
 FILLCELL_X32 FILLER_52_952 ();
 FILLCELL_X32 FILLER_52_984 ();
 FILLCELL_X32 FILLER_52_1016 ();
 FILLCELL_X32 FILLER_52_1048 ();
 FILLCELL_X32 FILLER_52_1080 ();
 FILLCELL_X32 FILLER_52_1112 ();
 FILLCELL_X32 FILLER_52_1144 ();
 FILLCELL_X32 FILLER_52_1176 ();
 FILLCELL_X32 FILLER_52_1208 ();
 FILLCELL_X32 FILLER_52_1240 ();
 FILLCELL_X32 FILLER_52_1272 ();
 FILLCELL_X32 FILLER_52_1304 ();
 FILLCELL_X32 FILLER_52_1336 ();
 FILLCELL_X32 FILLER_52_1368 ();
 FILLCELL_X32 FILLER_52_1400 ();
 FILLCELL_X32 FILLER_52_1432 ();
 FILLCELL_X32 FILLER_52_1464 ();
 FILLCELL_X32 FILLER_52_1496 ();
 FILLCELL_X32 FILLER_52_1528 ();
 FILLCELL_X32 FILLER_52_1560 ();
 FILLCELL_X32 FILLER_52_1592 ();
 FILLCELL_X32 FILLER_52_1624 ();
 FILLCELL_X32 FILLER_52_1656 ();
 FILLCELL_X32 FILLER_52_1688 ();
 FILLCELL_X32 FILLER_52_1720 ();
 FILLCELL_X32 FILLER_52_1752 ();
 FILLCELL_X32 FILLER_52_1784 ();
 FILLCELL_X32 FILLER_52_1816 ();
 FILLCELL_X32 FILLER_52_1848 ();
 FILLCELL_X8 FILLER_52_1880 ();
 FILLCELL_X4 FILLER_52_1888 ();
 FILLCELL_X2 FILLER_52_1892 ();
 FILLCELL_X32 FILLER_52_1895 ();
 FILLCELL_X32 FILLER_52_1927 ();
 FILLCELL_X32 FILLER_52_1959 ();
 FILLCELL_X32 FILLER_52_1991 ();
 FILLCELL_X32 FILLER_52_2023 ();
 FILLCELL_X32 FILLER_52_2055 ();
 FILLCELL_X32 FILLER_52_2087 ();
 FILLCELL_X32 FILLER_52_2119 ();
 FILLCELL_X32 FILLER_52_2151 ();
 FILLCELL_X32 FILLER_52_2183 ();
 FILLCELL_X32 FILLER_52_2215 ();
 FILLCELL_X32 FILLER_52_2247 ();
 FILLCELL_X32 FILLER_52_2279 ();
 FILLCELL_X32 FILLER_52_2311 ();
 FILLCELL_X32 FILLER_52_2343 ();
 FILLCELL_X32 FILLER_52_2375 ();
 FILLCELL_X32 FILLER_52_2407 ();
 FILLCELL_X32 FILLER_52_2439 ();
 FILLCELL_X32 FILLER_52_2471 ();
 FILLCELL_X32 FILLER_52_2503 ();
 FILLCELL_X32 FILLER_52_2535 ();
 FILLCELL_X32 FILLER_52_2567 ();
 FILLCELL_X32 FILLER_52_2599 ();
 FILLCELL_X32 FILLER_52_2631 ();
 FILLCELL_X32 FILLER_52_2663 ();
 FILLCELL_X32 FILLER_52_2695 ();
 FILLCELL_X32 FILLER_52_2727 ();
 FILLCELL_X32 FILLER_52_2759 ();
 FILLCELL_X32 FILLER_52_2791 ();
 FILLCELL_X32 FILLER_52_2823 ();
 FILLCELL_X32 FILLER_52_2855 ();
 FILLCELL_X32 FILLER_52_2887 ();
 FILLCELL_X32 FILLER_52_2919 ();
 FILLCELL_X32 FILLER_52_2951 ();
 FILLCELL_X32 FILLER_52_2983 ();
 FILLCELL_X32 FILLER_52_3015 ();
 FILLCELL_X32 FILLER_52_3047 ();
 FILLCELL_X32 FILLER_52_3079 ();
 FILLCELL_X32 FILLER_52_3111 ();
 FILLCELL_X8 FILLER_52_3143 ();
 FILLCELL_X4 FILLER_52_3151 ();
 FILLCELL_X2 FILLER_52_3155 ();
 FILLCELL_X32 FILLER_52_3158 ();
 FILLCELL_X32 FILLER_52_3190 ();
 FILLCELL_X32 FILLER_52_3222 ();
 FILLCELL_X32 FILLER_52_3254 ();
 FILLCELL_X32 FILLER_52_3286 ();
 FILLCELL_X32 FILLER_52_3318 ();
 FILLCELL_X32 FILLER_52_3350 ();
 FILLCELL_X32 FILLER_52_3382 ();
 FILLCELL_X32 FILLER_52_3414 ();
 FILLCELL_X32 FILLER_52_3446 ();
 FILLCELL_X32 FILLER_52_3478 ();
 FILLCELL_X32 FILLER_52_3510 ();
 FILLCELL_X32 FILLER_52_3542 ();
 FILLCELL_X32 FILLER_52_3574 ();
 FILLCELL_X32 FILLER_52_3606 ();
 FILLCELL_X32 FILLER_52_3638 ();
 FILLCELL_X32 FILLER_52_3670 ();
 FILLCELL_X32 FILLER_52_3702 ();
 FILLCELL_X4 FILLER_52_3734 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X32 FILLER_53_97 ();
 FILLCELL_X32 FILLER_53_129 ();
 FILLCELL_X32 FILLER_53_161 ();
 FILLCELL_X32 FILLER_53_193 ();
 FILLCELL_X32 FILLER_53_225 ();
 FILLCELL_X32 FILLER_53_257 ();
 FILLCELL_X32 FILLER_53_289 ();
 FILLCELL_X32 FILLER_53_321 ();
 FILLCELL_X32 FILLER_53_353 ();
 FILLCELL_X32 FILLER_53_385 ();
 FILLCELL_X32 FILLER_53_417 ();
 FILLCELL_X32 FILLER_53_449 ();
 FILLCELL_X32 FILLER_53_481 ();
 FILLCELL_X32 FILLER_53_513 ();
 FILLCELL_X32 FILLER_53_545 ();
 FILLCELL_X32 FILLER_53_577 ();
 FILLCELL_X32 FILLER_53_609 ();
 FILLCELL_X32 FILLER_53_641 ();
 FILLCELL_X32 FILLER_53_673 ();
 FILLCELL_X32 FILLER_53_705 ();
 FILLCELL_X32 FILLER_53_737 ();
 FILLCELL_X32 FILLER_53_769 ();
 FILLCELL_X32 FILLER_53_801 ();
 FILLCELL_X32 FILLER_53_833 ();
 FILLCELL_X32 FILLER_53_865 ();
 FILLCELL_X32 FILLER_53_897 ();
 FILLCELL_X32 FILLER_53_929 ();
 FILLCELL_X32 FILLER_53_961 ();
 FILLCELL_X32 FILLER_53_993 ();
 FILLCELL_X32 FILLER_53_1025 ();
 FILLCELL_X32 FILLER_53_1057 ();
 FILLCELL_X32 FILLER_53_1089 ();
 FILLCELL_X32 FILLER_53_1121 ();
 FILLCELL_X32 FILLER_53_1153 ();
 FILLCELL_X32 FILLER_53_1185 ();
 FILLCELL_X32 FILLER_53_1217 ();
 FILLCELL_X8 FILLER_53_1249 ();
 FILLCELL_X4 FILLER_53_1257 ();
 FILLCELL_X2 FILLER_53_1261 ();
 FILLCELL_X32 FILLER_53_1264 ();
 FILLCELL_X32 FILLER_53_1296 ();
 FILLCELL_X32 FILLER_53_1328 ();
 FILLCELL_X32 FILLER_53_1360 ();
 FILLCELL_X32 FILLER_53_1392 ();
 FILLCELL_X32 FILLER_53_1424 ();
 FILLCELL_X32 FILLER_53_1456 ();
 FILLCELL_X32 FILLER_53_1488 ();
 FILLCELL_X32 FILLER_53_1520 ();
 FILLCELL_X32 FILLER_53_1552 ();
 FILLCELL_X32 FILLER_53_1584 ();
 FILLCELL_X32 FILLER_53_1616 ();
 FILLCELL_X32 FILLER_53_1648 ();
 FILLCELL_X32 FILLER_53_1680 ();
 FILLCELL_X32 FILLER_53_1712 ();
 FILLCELL_X32 FILLER_53_1744 ();
 FILLCELL_X32 FILLER_53_1776 ();
 FILLCELL_X32 FILLER_53_1808 ();
 FILLCELL_X32 FILLER_53_1840 ();
 FILLCELL_X32 FILLER_53_1872 ();
 FILLCELL_X32 FILLER_53_1904 ();
 FILLCELL_X32 FILLER_53_1936 ();
 FILLCELL_X32 FILLER_53_1968 ();
 FILLCELL_X32 FILLER_53_2000 ();
 FILLCELL_X32 FILLER_53_2032 ();
 FILLCELL_X32 FILLER_53_2064 ();
 FILLCELL_X32 FILLER_53_2096 ();
 FILLCELL_X32 FILLER_53_2128 ();
 FILLCELL_X32 FILLER_53_2160 ();
 FILLCELL_X32 FILLER_53_2192 ();
 FILLCELL_X32 FILLER_53_2224 ();
 FILLCELL_X32 FILLER_53_2256 ();
 FILLCELL_X32 FILLER_53_2288 ();
 FILLCELL_X32 FILLER_53_2320 ();
 FILLCELL_X32 FILLER_53_2352 ();
 FILLCELL_X32 FILLER_53_2384 ();
 FILLCELL_X32 FILLER_53_2416 ();
 FILLCELL_X32 FILLER_53_2448 ();
 FILLCELL_X32 FILLER_53_2480 ();
 FILLCELL_X8 FILLER_53_2512 ();
 FILLCELL_X4 FILLER_53_2520 ();
 FILLCELL_X2 FILLER_53_2524 ();
 FILLCELL_X32 FILLER_53_2527 ();
 FILLCELL_X32 FILLER_53_2559 ();
 FILLCELL_X32 FILLER_53_2591 ();
 FILLCELL_X32 FILLER_53_2623 ();
 FILLCELL_X32 FILLER_53_2655 ();
 FILLCELL_X32 FILLER_53_2687 ();
 FILLCELL_X32 FILLER_53_2719 ();
 FILLCELL_X32 FILLER_53_2751 ();
 FILLCELL_X32 FILLER_53_2783 ();
 FILLCELL_X32 FILLER_53_2815 ();
 FILLCELL_X32 FILLER_53_2847 ();
 FILLCELL_X32 FILLER_53_2879 ();
 FILLCELL_X32 FILLER_53_2911 ();
 FILLCELL_X32 FILLER_53_2943 ();
 FILLCELL_X32 FILLER_53_2975 ();
 FILLCELL_X32 FILLER_53_3007 ();
 FILLCELL_X32 FILLER_53_3039 ();
 FILLCELL_X32 FILLER_53_3071 ();
 FILLCELL_X32 FILLER_53_3103 ();
 FILLCELL_X32 FILLER_53_3135 ();
 FILLCELL_X32 FILLER_53_3167 ();
 FILLCELL_X32 FILLER_53_3199 ();
 FILLCELL_X32 FILLER_53_3231 ();
 FILLCELL_X32 FILLER_53_3263 ();
 FILLCELL_X32 FILLER_53_3295 ();
 FILLCELL_X32 FILLER_53_3327 ();
 FILLCELL_X32 FILLER_53_3359 ();
 FILLCELL_X32 FILLER_53_3391 ();
 FILLCELL_X32 FILLER_53_3423 ();
 FILLCELL_X32 FILLER_53_3455 ();
 FILLCELL_X32 FILLER_53_3487 ();
 FILLCELL_X32 FILLER_53_3519 ();
 FILLCELL_X32 FILLER_53_3551 ();
 FILLCELL_X32 FILLER_53_3583 ();
 FILLCELL_X32 FILLER_53_3615 ();
 FILLCELL_X32 FILLER_53_3647 ();
 FILLCELL_X32 FILLER_53_3679 ();
 FILLCELL_X16 FILLER_53_3711 ();
 FILLCELL_X8 FILLER_53_3727 ();
 FILLCELL_X2 FILLER_53_3735 ();
 FILLCELL_X1 FILLER_53_3737 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X32 FILLER_54_33 ();
 FILLCELL_X32 FILLER_54_65 ();
 FILLCELL_X32 FILLER_54_97 ();
 FILLCELL_X32 FILLER_54_129 ();
 FILLCELL_X32 FILLER_54_161 ();
 FILLCELL_X32 FILLER_54_193 ();
 FILLCELL_X32 FILLER_54_225 ();
 FILLCELL_X32 FILLER_54_257 ();
 FILLCELL_X32 FILLER_54_289 ();
 FILLCELL_X32 FILLER_54_321 ();
 FILLCELL_X32 FILLER_54_353 ();
 FILLCELL_X32 FILLER_54_385 ();
 FILLCELL_X32 FILLER_54_417 ();
 FILLCELL_X32 FILLER_54_449 ();
 FILLCELL_X32 FILLER_54_481 ();
 FILLCELL_X32 FILLER_54_513 ();
 FILLCELL_X32 FILLER_54_545 ();
 FILLCELL_X32 FILLER_54_577 ();
 FILLCELL_X16 FILLER_54_609 ();
 FILLCELL_X4 FILLER_54_625 ();
 FILLCELL_X2 FILLER_54_629 ();
 FILLCELL_X32 FILLER_54_632 ();
 FILLCELL_X32 FILLER_54_664 ();
 FILLCELL_X32 FILLER_54_696 ();
 FILLCELL_X32 FILLER_54_728 ();
 FILLCELL_X32 FILLER_54_760 ();
 FILLCELL_X32 FILLER_54_792 ();
 FILLCELL_X32 FILLER_54_824 ();
 FILLCELL_X32 FILLER_54_856 ();
 FILLCELL_X32 FILLER_54_888 ();
 FILLCELL_X32 FILLER_54_920 ();
 FILLCELL_X32 FILLER_54_952 ();
 FILLCELL_X32 FILLER_54_984 ();
 FILLCELL_X32 FILLER_54_1016 ();
 FILLCELL_X32 FILLER_54_1048 ();
 FILLCELL_X32 FILLER_54_1080 ();
 FILLCELL_X32 FILLER_54_1112 ();
 FILLCELL_X32 FILLER_54_1144 ();
 FILLCELL_X32 FILLER_54_1176 ();
 FILLCELL_X32 FILLER_54_1208 ();
 FILLCELL_X32 FILLER_54_1240 ();
 FILLCELL_X32 FILLER_54_1272 ();
 FILLCELL_X32 FILLER_54_1304 ();
 FILLCELL_X32 FILLER_54_1336 ();
 FILLCELL_X32 FILLER_54_1368 ();
 FILLCELL_X32 FILLER_54_1400 ();
 FILLCELL_X32 FILLER_54_1432 ();
 FILLCELL_X32 FILLER_54_1464 ();
 FILLCELL_X32 FILLER_54_1496 ();
 FILLCELL_X32 FILLER_54_1528 ();
 FILLCELL_X32 FILLER_54_1560 ();
 FILLCELL_X32 FILLER_54_1592 ();
 FILLCELL_X32 FILLER_54_1624 ();
 FILLCELL_X32 FILLER_54_1656 ();
 FILLCELL_X32 FILLER_54_1688 ();
 FILLCELL_X32 FILLER_54_1720 ();
 FILLCELL_X32 FILLER_54_1752 ();
 FILLCELL_X32 FILLER_54_1784 ();
 FILLCELL_X32 FILLER_54_1816 ();
 FILLCELL_X32 FILLER_54_1848 ();
 FILLCELL_X8 FILLER_54_1880 ();
 FILLCELL_X4 FILLER_54_1888 ();
 FILLCELL_X2 FILLER_54_1892 ();
 FILLCELL_X32 FILLER_54_1895 ();
 FILLCELL_X32 FILLER_54_1927 ();
 FILLCELL_X32 FILLER_54_1959 ();
 FILLCELL_X32 FILLER_54_1991 ();
 FILLCELL_X32 FILLER_54_2023 ();
 FILLCELL_X32 FILLER_54_2055 ();
 FILLCELL_X32 FILLER_54_2087 ();
 FILLCELL_X32 FILLER_54_2119 ();
 FILLCELL_X32 FILLER_54_2151 ();
 FILLCELL_X32 FILLER_54_2183 ();
 FILLCELL_X32 FILLER_54_2215 ();
 FILLCELL_X32 FILLER_54_2247 ();
 FILLCELL_X32 FILLER_54_2279 ();
 FILLCELL_X32 FILLER_54_2311 ();
 FILLCELL_X32 FILLER_54_2343 ();
 FILLCELL_X32 FILLER_54_2375 ();
 FILLCELL_X32 FILLER_54_2407 ();
 FILLCELL_X32 FILLER_54_2439 ();
 FILLCELL_X32 FILLER_54_2471 ();
 FILLCELL_X32 FILLER_54_2503 ();
 FILLCELL_X32 FILLER_54_2535 ();
 FILLCELL_X32 FILLER_54_2567 ();
 FILLCELL_X32 FILLER_54_2599 ();
 FILLCELL_X32 FILLER_54_2631 ();
 FILLCELL_X32 FILLER_54_2663 ();
 FILLCELL_X32 FILLER_54_2695 ();
 FILLCELL_X32 FILLER_54_2727 ();
 FILLCELL_X32 FILLER_54_2759 ();
 FILLCELL_X32 FILLER_54_2791 ();
 FILLCELL_X32 FILLER_54_2823 ();
 FILLCELL_X32 FILLER_54_2855 ();
 FILLCELL_X32 FILLER_54_2887 ();
 FILLCELL_X32 FILLER_54_2919 ();
 FILLCELL_X32 FILLER_54_2951 ();
 FILLCELL_X32 FILLER_54_2983 ();
 FILLCELL_X32 FILLER_54_3015 ();
 FILLCELL_X32 FILLER_54_3047 ();
 FILLCELL_X32 FILLER_54_3079 ();
 FILLCELL_X32 FILLER_54_3111 ();
 FILLCELL_X8 FILLER_54_3143 ();
 FILLCELL_X4 FILLER_54_3151 ();
 FILLCELL_X2 FILLER_54_3155 ();
 FILLCELL_X32 FILLER_54_3158 ();
 FILLCELL_X32 FILLER_54_3190 ();
 FILLCELL_X32 FILLER_54_3222 ();
 FILLCELL_X32 FILLER_54_3254 ();
 FILLCELL_X32 FILLER_54_3286 ();
 FILLCELL_X32 FILLER_54_3318 ();
 FILLCELL_X32 FILLER_54_3350 ();
 FILLCELL_X32 FILLER_54_3382 ();
 FILLCELL_X32 FILLER_54_3414 ();
 FILLCELL_X32 FILLER_54_3446 ();
 FILLCELL_X32 FILLER_54_3478 ();
 FILLCELL_X32 FILLER_54_3510 ();
 FILLCELL_X32 FILLER_54_3542 ();
 FILLCELL_X32 FILLER_54_3574 ();
 FILLCELL_X32 FILLER_54_3606 ();
 FILLCELL_X32 FILLER_54_3638 ();
 FILLCELL_X32 FILLER_54_3670 ();
 FILLCELL_X32 FILLER_54_3702 ();
 FILLCELL_X4 FILLER_54_3734 ();
 FILLCELL_X32 FILLER_55_1 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X32 FILLER_55_65 ();
 FILLCELL_X32 FILLER_55_97 ();
 FILLCELL_X32 FILLER_55_129 ();
 FILLCELL_X32 FILLER_55_161 ();
 FILLCELL_X32 FILLER_55_193 ();
 FILLCELL_X32 FILLER_55_225 ();
 FILLCELL_X32 FILLER_55_257 ();
 FILLCELL_X32 FILLER_55_289 ();
 FILLCELL_X32 FILLER_55_321 ();
 FILLCELL_X32 FILLER_55_353 ();
 FILLCELL_X32 FILLER_55_385 ();
 FILLCELL_X32 FILLER_55_417 ();
 FILLCELL_X32 FILLER_55_449 ();
 FILLCELL_X32 FILLER_55_481 ();
 FILLCELL_X32 FILLER_55_513 ();
 FILLCELL_X32 FILLER_55_545 ();
 FILLCELL_X32 FILLER_55_577 ();
 FILLCELL_X32 FILLER_55_609 ();
 FILLCELL_X32 FILLER_55_641 ();
 FILLCELL_X32 FILLER_55_673 ();
 FILLCELL_X32 FILLER_55_705 ();
 FILLCELL_X32 FILLER_55_737 ();
 FILLCELL_X32 FILLER_55_769 ();
 FILLCELL_X32 FILLER_55_801 ();
 FILLCELL_X32 FILLER_55_833 ();
 FILLCELL_X32 FILLER_55_865 ();
 FILLCELL_X32 FILLER_55_897 ();
 FILLCELL_X32 FILLER_55_929 ();
 FILLCELL_X32 FILLER_55_961 ();
 FILLCELL_X32 FILLER_55_993 ();
 FILLCELL_X32 FILLER_55_1025 ();
 FILLCELL_X32 FILLER_55_1057 ();
 FILLCELL_X32 FILLER_55_1089 ();
 FILLCELL_X32 FILLER_55_1121 ();
 FILLCELL_X32 FILLER_55_1153 ();
 FILLCELL_X32 FILLER_55_1185 ();
 FILLCELL_X32 FILLER_55_1217 ();
 FILLCELL_X8 FILLER_55_1249 ();
 FILLCELL_X4 FILLER_55_1257 ();
 FILLCELL_X2 FILLER_55_1261 ();
 FILLCELL_X32 FILLER_55_1264 ();
 FILLCELL_X32 FILLER_55_1296 ();
 FILLCELL_X32 FILLER_55_1328 ();
 FILLCELL_X32 FILLER_55_1360 ();
 FILLCELL_X32 FILLER_55_1392 ();
 FILLCELL_X32 FILLER_55_1424 ();
 FILLCELL_X32 FILLER_55_1456 ();
 FILLCELL_X32 FILLER_55_1488 ();
 FILLCELL_X32 FILLER_55_1520 ();
 FILLCELL_X32 FILLER_55_1552 ();
 FILLCELL_X32 FILLER_55_1584 ();
 FILLCELL_X32 FILLER_55_1616 ();
 FILLCELL_X32 FILLER_55_1648 ();
 FILLCELL_X32 FILLER_55_1680 ();
 FILLCELL_X32 FILLER_55_1712 ();
 FILLCELL_X32 FILLER_55_1744 ();
 FILLCELL_X32 FILLER_55_1776 ();
 FILLCELL_X32 FILLER_55_1808 ();
 FILLCELL_X32 FILLER_55_1840 ();
 FILLCELL_X32 FILLER_55_1872 ();
 FILLCELL_X32 FILLER_55_1904 ();
 FILLCELL_X32 FILLER_55_1936 ();
 FILLCELL_X32 FILLER_55_1968 ();
 FILLCELL_X32 FILLER_55_2000 ();
 FILLCELL_X32 FILLER_55_2032 ();
 FILLCELL_X32 FILLER_55_2064 ();
 FILLCELL_X32 FILLER_55_2096 ();
 FILLCELL_X32 FILLER_55_2128 ();
 FILLCELL_X32 FILLER_55_2160 ();
 FILLCELL_X32 FILLER_55_2192 ();
 FILLCELL_X32 FILLER_55_2224 ();
 FILLCELL_X32 FILLER_55_2256 ();
 FILLCELL_X32 FILLER_55_2288 ();
 FILLCELL_X32 FILLER_55_2320 ();
 FILLCELL_X32 FILLER_55_2352 ();
 FILLCELL_X32 FILLER_55_2384 ();
 FILLCELL_X32 FILLER_55_2416 ();
 FILLCELL_X32 FILLER_55_2448 ();
 FILLCELL_X32 FILLER_55_2480 ();
 FILLCELL_X8 FILLER_55_2512 ();
 FILLCELL_X4 FILLER_55_2520 ();
 FILLCELL_X2 FILLER_55_2524 ();
 FILLCELL_X32 FILLER_55_2527 ();
 FILLCELL_X32 FILLER_55_2559 ();
 FILLCELL_X32 FILLER_55_2591 ();
 FILLCELL_X32 FILLER_55_2623 ();
 FILLCELL_X32 FILLER_55_2655 ();
 FILLCELL_X32 FILLER_55_2687 ();
 FILLCELL_X32 FILLER_55_2719 ();
 FILLCELL_X32 FILLER_55_2751 ();
 FILLCELL_X32 FILLER_55_2783 ();
 FILLCELL_X32 FILLER_55_2815 ();
 FILLCELL_X32 FILLER_55_2847 ();
 FILLCELL_X32 FILLER_55_2879 ();
 FILLCELL_X32 FILLER_55_2911 ();
 FILLCELL_X32 FILLER_55_2943 ();
 FILLCELL_X32 FILLER_55_2975 ();
 FILLCELL_X32 FILLER_55_3007 ();
 FILLCELL_X32 FILLER_55_3039 ();
 FILLCELL_X32 FILLER_55_3071 ();
 FILLCELL_X32 FILLER_55_3103 ();
 FILLCELL_X32 FILLER_55_3135 ();
 FILLCELL_X32 FILLER_55_3167 ();
 FILLCELL_X32 FILLER_55_3199 ();
 FILLCELL_X32 FILLER_55_3231 ();
 FILLCELL_X32 FILLER_55_3263 ();
 FILLCELL_X32 FILLER_55_3295 ();
 FILLCELL_X32 FILLER_55_3327 ();
 FILLCELL_X32 FILLER_55_3359 ();
 FILLCELL_X32 FILLER_55_3391 ();
 FILLCELL_X32 FILLER_55_3423 ();
 FILLCELL_X32 FILLER_55_3455 ();
 FILLCELL_X32 FILLER_55_3487 ();
 FILLCELL_X32 FILLER_55_3519 ();
 FILLCELL_X32 FILLER_55_3551 ();
 FILLCELL_X32 FILLER_55_3583 ();
 FILLCELL_X32 FILLER_55_3615 ();
 FILLCELL_X32 FILLER_55_3647 ();
 FILLCELL_X32 FILLER_55_3679 ();
 FILLCELL_X16 FILLER_55_3711 ();
 FILLCELL_X8 FILLER_55_3727 ();
 FILLCELL_X2 FILLER_55_3735 ();
 FILLCELL_X1 FILLER_55_3737 ();
 FILLCELL_X32 FILLER_56_1 ();
 FILLCELL_X32 FILLER_56_33 ();
 FILLCELL_X32 FILLER_56_65 ();
 FILLCELL_X32 FILLER_56_97 ();
 FILLCELL_X32 FILLER_56_129 ();
 FILLCELL_X32 FILLER_56_161 ();
 FILLCELL_X32 FILLER_56_193 ();
 FILLCELL_X32 FILLER_56_225 ();
 FILLCELL_X32 FILLER_56_257 ();
 FILLCELL_X32 FILLER_56_289 ();
 FILLCELL_X32 FILLER_56_321 ();
 FILLCELL_X32 FILLER_56_353 ();
 FILLCELL_X32 FILLER_56_385 ();
 FILLCELL_X32 FILLER_56_417 ();
 FILLCELL_X32 FILLER_56_449 ();
 FILLCELL_X32 FILLER_56_481 ();
 FILLCELL_X32 FILLER_56_513 ();
 FILLCELL_X32 FILLER_56_545 ();
 FILLCELL_X32 FILLER_56_577 ();
 FILLCELL_X16 FILLER_56_609 ();
 FILLCELL_X4 FILLER_56_625 ();
 FILLCELL_X2 FILLER_56_629 ();
 FILLCELL_X32 FILLER_56_632 ();
 FILLCELL_X32 FILLER_56_664 ();
 FILLCELL_X32 FILLER_56_696 ();
 FILLCELL_X32 FILLER_56_728 ();
 FILLCELL_X32 FILLER_56_760 ();
 FILLCELL_X32 FILLER_56_792 ();
 FILLCELL_X32 FILLER_56_824 ();
 FILLCELL_X32 FILLER_56_856 ();
 FILLCELL_X32 FILLER_56_888 ();
 FILLCELL_X32 FILLER_56_920 ();
 FILLCELL_X32 FILLER_56_952 ();
 FILLCELL_X32 FILLER_56_984 ();
 FILLCELL_X32 FILLER_56_1016 ();
 FILLCELL_X32 FILLER_56_1048 ();
 FILLCELL_X32 FILLER_56_1080 ();
 FILLCELL_X32 FILLER_56_1112 ();
 FILLCELL_X32 FILLER_56_1144 ();
 FILLCELL_X32 FILLER_56_1176 ();
 FILLCELL_X32 FILLER_56_1208 ();
 FILLCELL_X32 FILLER_56_1240 ();
 FILLCELL_X32 FILLER_56_1272 ();
 FILLCELL_X32 FILLER_56_1304 ();
 FILLCELL_X32 FILLER_56_1336 ();
 FILLCELL_X32 FILLER_56_1368 ();
 FILLCELL_X32 FILLER_56_1400 ();
 FILLCELL_X32 FILLER_56_1432 ();
 FILLCELL_X32 FILLER_56_1464 ();
 FILLCELL_X32 FILLER_56_1496 ();
 FILLCELL_X32 FILLER_56_1528 ();
 FILLCELL_X32 FILLER_56_1560 ();
 FILLCELL_X32 FILLER_56_1592 ();
 FILLCELL_X32 FILLER_56_1624 ();
 FILLCELL_X32 FILLER_56_1656 ();
 FILLCELL_X32 FILLER_56_1688 ();
 FILLCELL_X32 FILLER_56_1720 ();
 FILLCELL_X32 FILLER_56_1752 ();
 FILLCELL_X32 FILLER_56_1784 ();
 FILLCELL_X32 FILLER_56_1816 ();
 FILLCELL_X32 FILLER_56_1848 ();
 FILLCELL_X8 FILLER_56_1880 ();
 FILLCELL_X4 FILLER_56_1888 ();
 FILLCELL_X2 FILLER_56_1892 ();
 FILLCELL_X32 FILLER_56_1895 ();
 FILLCELL_X32 FILLER_56_1927 ();
 FILLCELL_X32 FILLER_56_1959 ();
 FILLCELL_X32 FILLER_56_1991 ();
 FILLCELL_X32 FILLER_56_2023 ();
 FILLCELL_X32 FILLER_56_2055 ();
 FILLCELL_X32 FILLER_56_2087 ();
 FILLCELL_X32 FILLER_56_2119 ();
 FILLCELL_X32 FILLER_56_2151 ();
 FILLCELL_X32 FILLER_56_2183 ();
 FILLCELL_X32 FILLER_56_2215 ();
 FILLCELL_X32 FILLER_56_2247 ();
 FILLCELL_X32 FILLER_56_2279 ();
 FILLCELL_X32 FILLER_56_2311 ();
 FILLCELL_X32 FILLER_56_2343 ();
 FILLCELL_X32 FILLER_56_2375 ();
 FILLCELL_X32 FILLER_56_2407 ();
 FILLCELL_X32 FILLER_56_2439 ();
 FILLCELL_X32 FILLER_56_2471 ();
 FILLCELL_X32 FILLER_56_2503 ();
 FILLCELL_X32 FILLER_56_2535 ();
 FILLCELL_X32 FILLER_56_2567 ();
 FILLCELL_X32 FILLER_56_2599 ();
 FILLCELL_X32 FILLER_56_2631 ();
 FILLCELL_X32 FILLER_56_2663 ();
 FILLCELL_X32 FILLER_56_2695 ();
 FILLCELL_X32 FILLER_56_2727 ();
 FILLCELL_X32 FILLER_56_2759 ();
 FILLCELL_X32 FILLER_56_2791 ();
 FILLCELL_X32 FILLER_56_2823 ();
 FILLCELL_X32 FILLER_56_2855 ();
 FILLCELL_X32 FILLER_56_2887 ();
 FILLCELL_X32 FILLER_56_2919 ();
 FILLCELL_X32 FILLER_56_2951 ();
 FILLCELL_X32 FILLER_56_2983 ();
 FILLCELL_X32 FILLER_56_3015 ();
 FILLCELL_X32 FILLER_56_3047 ();
 FILLCELL_X32 FILLER_56_3079 ();
 FILLCELL_X32 FILLER_56_3111 ();
 FILLCELL_X8 FILLER_56_3143 ();
 FILLCELL_X4 FILLER_56_3151 ();
 FILLCELL_X2 FILLER_56_3155 ();
 FILLCELL_X32 FILLER_56_3158 ();
 FILLCELL_X32 FILLER_56_3190 ();
 FILLCELL_X32 FILLER_56_3222 ();
 FILLCELL_X32 FILLER_56_3254 ();
 FILLCELL_X32 FILLER_56_3286 ();
 FILLCELL_X32 FILLER_56_3318 ();
 FILLCELL_X32 FILLER_56_3350 ();
 FILLCELL_X32 FILLER_56_3382 ();
 FILLCELL_X32 FILLER_56_3414 ();
 FILLCELL_X32 FILLER_56_3446 ();
 FILLCELL_X32 FILLER_56_3478 ();
 FILLCELL_X32 FILLER_56_3510 ();
 FILLCELL_X32 FILLER_56_3542 ();
 FILLCELL_X32 FILLER_56_3574 ();
 FILLCELL_X32 FILLER_56_3606 ();
 FILLCELL_X32 FILLER_56_3638 ();
 FILLCELL_X32 FILLER_56_3670 ();
 FILLCELL_X32 FILLER_56_3702 ();
 FILLCELL_X4 FILLER_56_3734 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X32 FILLER_57_33 ();
 FILLCELL_X32 FILLER_57_65 ();
 FILLCELL_X32 FILLER_57_97 ();
 FILLCELL_X32 FILLER_57_129 ();
 FILLCELL_X32 FILLER_57_161 ();
 FILLCELL_X32 FILLER_57_193 ();
 FILLCELL_X32 FILLER_57_225 ();
 FILLCELL_X32 FILLER_57_257 ();
 FILLCELL_X32 FILLER_57_289 ();
 FILLCELL_X32 FILLER_57_321 ();
 FILLCELL_X32 FILLER_57_353 ();
 FILLCELL_X32 FILLER_57_385 ();
 FILLCELL_X32 FILLER_57_417 ();
 FILLCELL_X32 FILLER_57_449 ();
 FILLCELL_X32 FILLER_57_481 ();
 FILLCELL_X32 FILLER_57_513 ();
 FILLCELL_X32 FILLER_57_545 ();
 FILLCELL_X32 FILLER_57_577 ();
 FILLCELL_X32 FILLER_57_609 ();
 FILLCELL_X32 FILLER_57_641 ();
 FILLCELL_X32 FILLER_57_673 ();
 FILLCELL_X32 FILLER_57_705 ();
 FILLCELL_X32 FILLER_57_737 ();
 FILLCELL_X32 FILLER_57_769 ();
 FILLCELL_X32 FILLER_57_801 ();
 FILLCELL_X32 FILLER_57_833 ();
 FILLCELL_X32 FILLER_57_865 ();
 FILLCELL_X32 FILLER_57_897 ();
 FILLCELL_X32 FILLER_57_929 ();
 FILLCELL_X32 FILLER_57_961 ();
 FILLCELL_X32 FILLER_57_993 ();
 FILLCELL_X32 FILLER_57_1025 ();
 FILLCELL_X32 FILLER_57_1057 ();
 FILLCELL_X32 FILLER_57_1089 ();
 FILLCELL_X32 FILLER_57_1121 ();
 FILLCELL_X32 FILLER_57_1153 ();
 FILLCELL_X32 FILLER_57_1185 ();
 FILLCELL_X32 FILLER_57_1217 ();
 FILLCELL_X8 FILLER_57_1249 ();
 FILLCELL_X4 FILLER_57_1257 ();
 FILLCELL_X2 FILLER_57_1261 ();
 FILLCELL_X32 FILLER_57_1264 ();
 FILLCELL_X32 FILLER_57_1296 ();
 FILLCELL_X32 FILLER_57_1328 ();
 FILLCELL_X32 FILLER_57_1360 ();
 FILLCELL_X32 FILLER_57_1392 ();
 FILLCELL_X32 FILLER_57_1424 ();
 FILLCELL_X32 FILLER_57_1456 ();
 FILLCELL_X32 FILLER_57_1488 ();
 FILLCELL_X32 FILLER_57_1520 ();
 FILLCELL_X32 FILLER_57_1552 ();
 FILLCELL_X32 FILLER_57_1584 ();
 FILLCELL_X32 FILLER_57_1616 ();
 FILLCELL_X32 FILLER_57_1648 ();
 FILLCELL_X32 FILLER_57_1680 ();
 FILLCELL_X32 FILLER_57_1712 ();
 FILLCELL_X32 FILLER_57_1744 ();
 FILLCELL_X32 FILLER_57_1776 ();
 FILLCELL_X32 FILLER_57_1808 ();
 FILLCELL_X32 FILLER_57_1840 ();
 FILLCELL_X32 FILLER_57_1872 ();
 FILLCELL_X32 FILLER_57_1904 ();
 FILLCELL_X32 FILLER_57_1936 ();
 FILLCELL_X32 FILLER_57_1968 ();
 FILLCELL_X32 FILLER_57_2000 ();
 FILLCELL_X32 FILLER_57_2032 ();
 FILLCELL_X32 FILLER_57_2064 ();
 FILLCELL_X32 FILLER_57_2096 ();
 FILLCELL_X32 FILLER_57_2128 ();
 FILLCELL_X32 FILLER_57_2160 ();
 FILLCELL_X32 FILLER_57_2192 ();
 FILLCELL_X32 FILLER_57_2224 ();
 FILLCELL_X32 FILLER_57_2256 ();
 FILLCELL_X32 FILLER_57_2288 ();
 FILLCELL_X32 FILLER_57_2320 ();
 FILLCELL_X32 FILLER_57_2352 ();
 FILLCELL_X32 FILLER_57_2384 ();
 FILLCELL_X32 FILLER_57_2416 ();
 FILLCELL_X32 FILLER_57_2448 ();
 FILLCELL_X32 FILLER_57_2480 ();
 FILLCELL_X8 FILLER_57_2512 ();
 FILLCELL_X4 FILLER_57_2520 ();
 FILLCELL_X2 FILLER_57_2524 ();
 FILLCELL_X32 FILLER_57_2527 ();
 FILLCELL_X32 FILLER_57_2559 ();
 FILLCELL_X32 FILLER_57_2591 ();
 FILLCELL_X32 FILLER_57_2623 ();
 FILLCELL_X32 FILLER_57_2655 ();
 FILLCELL_X32 FILLER_57_2687 ();
 FILLCELL_X32 FILLER_57_2719 ();
 FILLCELL_X32 FILLER_57_2751 ();
 FILLCELL_X32 FILLER_57_2783 ();
 FILLCELL_X32 FILLER_57_2815 ();
 FILLCELL_X32 FILLER_57_2847 ();
 FILLCELL_X32 FILLER_57_2879 ();
 FILLCELL_X32 FILLER_57_2911 ();
 FILLCELL_X32 FILLER_57_2943 ();
 FILLCELL_X32 FILLER_57_2975 ();
 FILLCELL_X32 FILLER_57_3007 ();
 FILLCELL_X32 FILLER_57_3039 ();
 FILLCELL_X32 FILLER_57_3071 ();
 FILLCELL_X32 FILLER_57_3103 ();
 FILLCELL_X32 FILLER_57_3135 ();
 FILLCELL_X32 FILLER_57_3167 ();
 FILLCELL_X32 FILLER_57_3199 ();
 FILLCELL_X32 FILLER_57_3231 ();
 FILLCELL_X32 FILLER_57_3263 ();
 FILLCELL_X32 FILLER_57_3295 ();
 FILLCELL_X32 FILLER_57_3327 ();
 FILLCELL_X32 FILLER_57_3359 ();
 FILLCELL_X32 FILLER_57_3391 ();
 FILLCELL_X32 FILLER_57_3423 ();
 FILLCELL_X32 FILLER_57_3455 ();
 FILLCELL_X32 FILLER_57_3487 ();
 FILLCELL_X32 FILLER_57_3519 ();
 FILLCELL_X32 FILLER_57_3551 ();
 FILLCELL_X32 FILLER_57_3583 ();
 FILLCELL_X32 FILLER_57_3615 ();
 FILLCELL_X32 FILLER_57_3647 ();
 FILLCELL_X32 FILLER_57_3679 ();
 FILLCELL_X16 FILLER_57_3711 ();
 FILLCELL_X8 FILLER_57_3727 ();
 FILLCELL_X2 FILLER_57_3735 ();
 FILLCELL_X1 FILLER_57_3737 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X32 FILLER_58_33 ();
 FILLCELL_X32 FILLER_58_65 ();
 FILLCELL_X32 FILLER_58_97 ();
 FILLCELL_X32 FILLER_58_129 ();
 FILLCELL_X32 FILLER_58_161 ();
 FILLCELL_X32 FILLER_58_193 ();
 FILLCELL_X32 FILLER_58_225 ();
 FILLCELL_X32 FILLER_58_257 ();
 FILLCELL_X32 FILLER_58_289 ();
 FILLCELL_X32 FILLER_58_321 ();
 FILLCELL_X32 FILLER_58_353 ();
 FILLCELL_X32 FILLER_58_385 ();
 FILLCELL_X32 FILLER_58_417 ();
 FILLCELL_X32 FILLER_58_449 ();
 FILLCELL_X32 FILLER_58_481 ();
 FILLCELL_X32 FILLER_58_513 ();
 FILLCELL_X32 FILLER_58_545 ();
 FILLCELL_X32 FILLER_58_577 ();
 FILLCELL_X16 FILLER_58_609 ();
 FILLCELL_X4 FILLER_58_625 ();
 FILLCELL_X2 FILLER_58_629 ();
 FILLCELL_X32 FILLER_58_632 ();
 FILLCELL_X32 FILLER_58_664 ();
 FILLCELL_X32 FILLER_58_696 ();
 FILLCELL_X32 FILLER_58_728 ();
 FILLCELL_X32 FILLER_58_760 ();
 FILLCELL_X32 FILLER_58_792 ();
 FILLCELL_X32 FILLER_58_824 ();
 FILLCELL_X32 FILLER_58_856 ();
 FILLCELL_X32 FILLER_58_888 ();
 FILLCELL_X32 FILLER_58_920 ();
 FILLCELL_X32 FILLER_58_952 ();
 FILLCELL_X32 FILLER_58_984 ();
 FILLCELL_X32 FILLER_58_1016 ();
 FILLCELL_X32 FILLER_58_1048 ();
 FILLCELL_X32 FILLER_58_1080 ();
 FILLCELL_X32 FILLER_58_1112 ();
 FILLCELL_X32 FILLER_58_1144 ();
 FILLCELL_X32 FILLER_58_1176 ();
 FILLCELL_X32 FILLER_58_1208 ();
 FILLCELL_X32 FILLER_58_1240 ();
 FILLCELL_X32 FILLER_58_1272 ();
 FILLCELL_X32 FILLER_58_1304 ();
 FILLCELL_X32 FILLER_58_1336 ();
 FILLCELL_X32 FILLER_58_1368 ();
 FILLCELL_X32 FILLER_58_1400 ();
 FILLCELL_X32 FILLER_58_1432 ();
 FILLCELL_X32 FILLER_58_1464 ();
 FILLCELL_X32 FILLER_58_1496 ();
 FILLCELL_X32 FILLER_58_1528 ();
 FILLCELL_X32 FILLER_58_1560 ();
 FILLCELL_X32 FILLER_58_1592 ();
 FILLCELL_X32 FILLER_58_1624 ();
 FILLCELL_X32 FILLER_58_1656 ();
 FILLCELL_X32 FILLER_58_1688 ();
 FILLCELL_X32 FILLER_58_1720 ();
 FILLCELL_X32 FILLER_58_1752 ();
 FILLCELL_X32 FILLER_58_1784 ();
 FILLCELL_X32 FILLER_58_1816 ();
 FILLCELL_X32 FILLER_58_1848 ();
 FILLCELL_X8 FILLER_58_1880 ();
 FILLCELL_X4 FILLER_58_1888 ();
 FILLCELL_X2 FILLER_58_1892 ();
 FILLCELL_X32 FILLER_58_1895 ();
 FILLCELL_X32 FILLER_58_1927 ();
 FILLCELL_X32 FILLER_58_1959 ();
 FILLCELL_X32 FILLER_58_1991 ();
 FILLCELL_X32 FILLER_58_2023 ();
 FILLCELL_X32 FILLER_58_2055 ();
 FILLCELL_X32 FILLER_58_2087 ();
 FILLCELL_X32 FILLER_58_2119 ();
 FILLCELL_X32 FILLER_58_2151 ();
 FILLCELL_X32 FILLER_58_2183 ();
 FILLCELL_X32 FILLER_58_2215 ();
 FILLCELL_X32 FILLER_58_2247 ();
 FILLCELL_X32 FILLER_58_2279 ();
 FILLCELL_X32 FILLER_58_2311 ();
 FILLCELL_X32 FILLER_58_2343 ();
 FILLCELL_X32 FILLER_58_2375 ();
 FILLCELL_X32 FILLER_58_2407 ();
 FILLCELL_X32 FILLER_58_2439 ();
 FILLCELL_X32 FILLER_58_2471 ();
 FILLCELL_X32 FILLER_58_2503 ();
 FILLCELL_X32 FILLER_58_2535 ();
 FILLCELL_X32 FILLER_58_2567 ();
 FILLCELL_X32 FILLER_58_2599 ();
 FILLCELL_X32 FILLER_58_2631 ();
 FILLCELL_X32 FILLER_58_2663 ();
 FILLCELL_X32 FILLER_58_2695 ();
 FILLCELL_X32 FILLER_58_2727 ();
 FILLCELL_X32 FILLER_58_2759 ();
 FILLCELL_X32 FILLER_58_2791 ();
 FILLCELL_X32 FILLER_58_2823 ();
 FILLCELL_X32 FILLER_58_2855 ();
 FILLCELL_X32 FILLER_58_2887 ();
 FILLCELL_X32 FILLER_58_2919 ();
 FILLCELL_X32 FILLER_58_2951 ();
 FILLCELL_X32 FILLER_58_2983 ();
 FILLCELL_X32 FILLER_58_3015 ();
 FILLCELL_X32 FILLER_58_3047 ();
 FILLCELL_X32 FILLER_58_3079 ();
 FILLCELL_X32 FILLER_58_3111 ();
 FILLCELL_X8 FILLER_58_3143 ();
 FILLCELL_X4 FILLER_58_3151 ();
 FILLCELL_X2 FILLER_58_3155 ();
 FILLCELL_X32 FILLER_58_3158 ();
 FILLCELL_X32 FILLER_58_3190 ();
 FILLCELL_X32 FILLER_58_3222 ();
 FILLCELL_X32 FILLER_58_3254 ();
 FILLCELL_X32 FILLER_58_3286 ();
 FILLCELL_X32 FILLER_58_3318 ();
 FILLCELL_X32 FILLER_58_3350 ();
 FILLCELL_X32 FILLER_58_3382 ();
 FILLCELL_X32 FILLER_58_3414 ();
 FILLCELL_X32 FILLER_58_3446 ();
 FILLCELL_X32 FILLER_58_3478 ();
 FILLCELL_X32 FILLER_58_3510 ();
 FILLCELL_X32 FILLER_58_3542 ();
 FILLCELL_X32 FILLER_58_3574 ();
 FILLCELL_X32 FILLER_58_3606 ();
 FILLCELL_X32 FILLER_58_3638 ();
 FILLCELL_X32 FILLER_58_3670 ();
 FILLCELL_X32 FILLER_58_3702 ();
 FILLCELL_X4 FILLER_58_3734 ();
 FILLCELL_X32 FILLER_59_1 ();
 FILLCELL_X32 FILLER_59_33 ();
 FILLCELL_X32 FILLER_59_65 ();
 FILLCELL_X32 FILLER_59_97 ();
 FILLCELL_X32 FILLER_59_129 ();
 FILLCELL_X32 FILLER_59_161 ();
 FILLCELL_X32 FILLER_59_193 ();
 FILLCELL_X32 FILLER_59_225 ();
 FILLCELL_X32 FILLER_59_257 ();
 FILLCELL_X32 FILLER_59_289 ();
 FILLCELL_X32 FILLER_59_321 ();
 FILLCELL_X32 FILLER_59_353 ();
 FILLCELL_X32 FILLER_59_385 ();
 FILLCELL_X32 FILLER_59_417 ();
 FILLCELL_X32 FILLER_59_449 ();
 FILLCELL_X32 FILLER_59_481 ();
 FILLCELL_X32 FILLER_59_513 ();
 FILLCELL_X32 FILLER_59_545 ();
 FILLCELL_X32 FILLER_59_577 ();
 FILLCELL_X32 FILLER_59_609 ();
 FILLCELL_X32 FILLER_59_641 ();
 FILLCELL_X32 FILLER_59_673 ();
 FILLCELL_X32 FILLER_59_705 ();
 FILLCELL_X32 FILLER_59_737 ();
 FILLCELL_X32 FILLER_59_769 ();
 FILLCELL_X32 FILLER_59_801 ();
 FILLCELL_X32 FILLER_59_833 ();
 FILLCELL_X32 FILLER_59_865 ();
 FILLCELL_X32 FILLER_59_897 ();
 FILLCELL_X32 FILLER_59_929 ();
 FILLCELL_X32 FILLER_59_961 ();
 FILLCELL_X32 FILLER_59_993 ();
 FILLCELL_X32 FILLER_59_1025 ();
 FILLCELL_X32 FILLER_59_1057 ();
 FILLCELL_X32 FILLER_59_1089 ();
 FILLCELL_X32 FILLER_59_1121 ();
 FILLCELL_X32 FILLER_59_1153 ();
 FILLCELL_X32 FILLER_59_1185 ();
 FILLCELL_X32 FILLER_59_1217 ();
 FILLCELL_X8 FILLER_59_1249 ();
 FILLCELL_X4 FILLER_59_1257 ();
 FILLCELL_X2 FILLER_59_1261 ();
 FILLCELL_X32 FILLER_59_1264 ();
 FILLCELL_X32 FILLER_59_1296 ();
 FILLCELL_X32 FILLER_59_1328 ();
 FILLCELL_X32 FILLER_59_1360 ();
 FILLCELL_X32 FILLER_59_1392 ();
 FILLCELL_X32 FILLER_59_1424 ();
 FILLCELL_X32 FILLER_59_1456 ();
 FILLCELL_X32 FILLER_59_1488 ();
 FILLCELL_X32 FILLER_59_1520 ();
 FILLCELL_X32 FILLER_59_1552 ();
 FILLCELL_X32 FILLER_59_1584 ();
 FILLCELL_X32 FILLER_59_1616 ();
 FILLCELL_X32 FILLER_59_1648 ();
 FILLCELL_X32 FILLER_59_1680 ();
 FILLCELL_X32 FILLER_59_1712 ();
 FILLCELL_X32 FILLER_59_1744 ();
 FILLCELL_X32 FILLER_59_1776 ();
 FILLCELL_X32 FILLER_59_1808 ();
 FILLCELL_X32 FILLER_59_1840 ();
 FILLCELL_X32 FILLER_59_1872 ();
 FILLCELL_X32 FILLER_59_1904 ();
 FILLCELL_X32 FILLER_59_1936 ();
 FILLCELL_X32 FILLER_59_1968 ();
 FILLCELL_X32 FILLER_59_2000 ();
 FILLCELL_X32 FILLER_59_2032 ();
 FILLCELL_X32 FILLER_59_2064 ();
 FILLCELL_X32 FILLER_59_2096 ();
 FILLCELL_X32 FILLER_59_2128 ();
 FILLCELL_X32 FILLER_59_2160 ();
 FILLCELL_X32 FILLER_59_2192 ();
 FILLCELL_X32 FILLER_59_2224 ();
 FILLCELL_X32 FILLER_59_2256 ();
 FILLCELL_X32 FILLER_59_2288 ();
 FILLCELL_X32 FILLER_59_2320 ();
 FILLCELL_X32 FILLER_59_2352 ();
 FILLCELL_X32 FILLER_59_2384 ();
 FILLCELL_X32 FILLER_59_2416 ();
 FILLCELL_X32 FILLER_59_2448 ();
 FILLCELL_X32 FILLER_59_2480 ();
 FILLCELL_X8 FILLER_59_2512 ();
 FILLCELL_X4 FILLER_59_2520 ();
 FILLCELL_X2 FILLER_59_2524 ();
 FILLCELL_X32 FILLER_59_2527 ();
 FILLCELL_X32 FILLER_59_2559 ();
 FILLCELL_X32 FILLER_59_2591 ();
 FILLCELL_X32 FILLER_59_2623 ();
 FILLCELL_X32 FILLER_59_2655 ();
 FILLCELL_X32 FILLER_59_2687 ();
 FILLCELL_X32 FILLER_59_2719 ();
 FILLCELL_X32 FILLER_59_2751 ();
 FILLCELL_X32 FILLER_59_2783 ();
 FILLCELL_X32 FILLER_59_2815 ();
 FILLCELL_X32 FILLER_59_2847 ();
 FILLCELL_X32 FILLER_59_2879 ();
 FILLCELL_X32 FILLER_59_2911 ();
 FILLCELL_X32 FILLER_59_2943 ();
 FILLCELL_X32 FILLER_59_2975 ();
 FILLCELL_X32 FILLER_59_3007 ();
 FILLCELL_X32 FILLER_59_3039 ();
 FILLCELL_X32 FILLER_59_3071 ();
 FILLCELL_X32 FILLER_59_3103 ();
 FILLCELL_X32 FILLER_59_3135 ();
 FILLCELL_X32 FILLER_59_3167 ();
 FILLCELL_X32 FILLER_59_3199 ();
 FILLCELL_X32 FILLER_59_3231 ();
 FILLCELL_X32 FILLER_59_3263 ();
 FILLCELL_X32 FILLER_59_3295 ();
 FILLCELL_X32 FILLER_59_3327 ();
 FILLCELL_X32 FILLER_59_3359 ();
 FILLCELL_X32 FILLER_59_3391 ();
 FILLCELL_X32 FILLER_59_3423 ();
 FILLCELL_X32 FILLER_59_3455 ();
 FILLCELL_X32 FILLER_59_3487 ();
 FILLCELL_X32 FILLER_59_3519 ();
 FILLCELL_X32 FILLER_59_3551 ();
 FILLCELL_X32 FILLER_59_3583 ();
 FILLCELL_X32 FILLER_59_3615 ();
 FILLCELL_X32 FILLER_59_3647 ();
 FILLCELL_X32 FILLER_59_3679 ();
 FILLCELL_X16 FILLER_59_3711 ();
 FILLCELL_X8 FILLER_59_3727 ();
 FILLCELL_X2 FILLER_59_3735 ();
 FILLCELL_X1 FILLER_59_3737 ();
 FILLCELL_X32 FILLER_60_1 ();
 FILLCELL_X32 FILLER_60_33 ();
 FILLCELL_X32 FILLER_60_65 ();
 FILLCELL_X32 FILLER_60_97 ();
 FILLCELL_X32 FILLER_60_129 ();
 FILLCELL_X32 FILLER_60_161 ();
 FILLCELL_X32 FILLER_60_193 ();
 FILLCELL_X32 FILLER_60_225 ();
 FILLCELL_X32 FILLER_60_257 ();
 FILLCELL_X32 FILLER_60_289 ();
 FILLCELL_X32 FILLER_60_321 ();
 FILLCELL_X32 FILLER_60_353 ();
 FILLCELL_X32 FILLER_60_385 ();
 FILLCELL_X32 FILLER_60_417 ();
 FILLCELL_X32 FILLER_60_449 ();
 FILLCELL_X32 FILLER_60_481 ();
 FILLCELL_X32 FILLER_60_513 ();
 FILLCELL_X32 FILLER_60_545 ();
 FILLCELL_X32 FILLER_60_577 ();
 FILLCELL_X16 FILLER_60_609 ();
 FILLCELL_X4 FILLER_60_625 ();
 FILLCELL_X2 FILLER_60_629 ();
 FILLCELL_X32 FILLER_60_632 ();
 FILLCELL_X32 FILLER_60_664 ();
 FILLCELL_X32 FILLER_60_696 ();
 FILLCELL_X32 FILLER_60_728 ();
 FILLCELL_X32 FILLER_60_760 ();
 FILLCELL_X32 FILLER_60_792 ();
 FILLCELL_X32 FILLER_60_824 ();
 FILLCELL_X32 FILLER_60_856 ();
 FILLCELL_X32 FILLER_60_888 ();
 FILLCELL_X32 FILLER_60_920 ();
 FILLCELL_X32 FILLER_60_952 ();
 FILLCELL_X32 FILLER_60_984 ();
 FILLCELL_X32 FILLER_60_1016 ();
 FILLCELL_X32 FILLER_60_1048 ();
 FILLCELL_X32 FILLER_60_1080 ();
 FILLCELL_X32 FILLER_60_1112 ();
 FILLCELL_X32 FILLER_60_1144 ();
 FILLCELL_X32 FILLER_60_1176 ();
 FILLCELL_X32 FILLER_60_1208 ();
 FILLCELL_X32 FILLER_60_1240 ();
 FILLCELL_X32 FILLER_60_1272 ();
 FILLCELL_X32 FILLER_60_1304 ();
 FILLCELL_X32 FILLER_60_1336 ();
 FILLCELL_X32 FILLER_60_1368 ();
 FILLCELL_X32 FILLER_60_1400 ();
 FILLCELL_X32 FILLER_60_1432 ();
 FILLCELL_X32 FILLER_60_1464 ();
 FILLCELL_X32 FILLER_60_1496 ();
 FILLCELL_X32 FILLER_60_1528 ();
 FILLCELL_X32 FILLER_60_1560 ();
 FILLCELL_X32 FILLER_60_1592 ();
 FILLCELL_X32 FILLER_60_1624 ();
 FILLCELL_X32 FILLER_60_1656 ();
 FILLCELL_X32 FILLER_60_1688 ();
 FILLCELL_X32 FILLER_60_1720 ();
 FILLCELL_X32 FILLER_60_1752 ();
 FILLCELL_X32 FILLER_60_1784 ();
 FILLCELL_X32 FILLER_60_1816 ();
 FILLCELL_X32 FILLER_60_1848 ();
 FILLCELL_X8 FILLER_60_1880 ();
 FILLCELL_X4 FILLER_60_1888 ();
 FILLCELL_X2 FILLER_60_1892 ();
 FILLCELL_X32 FILLER_60_1895 ();
 FILLCELL_X32 FILLER_60_1927 ();
 FILLCELL_X32 FILLER_60_1959 ();
 FILLCELL_X32 FILLER_60_1991 ();
 FILLCELL_X32 FILLER_60_2023 ();
 FILLCELL_X32 FILLER_60_2055 ();
 FILLCELL_X32 FILLER_60_2087 ();
 FILLCELL_X32 FILLER_60_2119 ();
 FILLCELL_X32 FILLER_60_2151 ();
 FILLCELL_X32 FILLER_60_2183 ();
 FILLCELL_X32 FILLER_60_2215 ();
 FILLCELL_X32 FILLER_60_2247 ();
 FILLCELL_X32 FILLER_60_2279 ();
 FILLCELL_X32 FILLER_60_2311 ();
 FILLCELL_X32 FILLER_60_2343 ();
 FILLCELL_X32 FILLER_60_2375 ();
 FILLCELL_X32 FILLER_60_2407 ();
 FILLCELL_X32 FILLER_60_2439 ();
 FILLCELL_X32 FILLER_60_2471 ();
 FILLCELL_X32 FILLER_60_2503 ();
 FILLCELL_X32 FILLER_60_2535 ();
 FILLCELL_X32 FILLER_60_2567 ();
 FILLCELL_X32 FILLER_60_2599 ();
 FILLCELL_X32 FILLER_60_2631 ();
 FILLCELL_X32 FILLER_60_2663 ();
 FILLCELL_X32 FILLER_60_2695 ();
 FILLCELL_X32 FILLER_60_2727 ();
 FILLCELL_X32 FILLER_60_2759 ();
 FILLCELL_X32 FILLER_60_2791 ();
 FILLCELL_X32 FILLER_60_2823 ();
 FILLCELL_X32 FILLER_60_2855 ();
 FILLCELL_X32 FILLER_60_2887 ();
 FILLCELL_X32 FILLER_60_2919 ();
 FILLCELL_X32 FILLER_60_2951 ();
 FILLCELL_X32 FILLER_60_2983 ();
 FILLCELL_X32 FILLER_60_3015 ();
 FILLCELL_X32 FILLER_60_3047 ();
 FILLCELL_X32 FILLER_60_3079 ();
 FILLCELL_X32 FILLER_60_3111 ();
 FILLCELL_X8 FILLER_60_3143 ();
 FILLCELL_X4 FILLER_60_3151 ();
 FILLCELL_X2 FILLER_60_3155 ();
 FILLCELL_X32 FILLER_60_3158 ();
 FILLCELL_X32 FILLER_60_3190 ();
 FILLCELL_X32 FILLER_60_3222 ();
 FILLCELL_X32 FILLER_60_3254 ();
 FILLCELL_X32 FILLER_60_3286 ();
 FILLCELL_X32 FILLER_60_3318 ();
 FILLCELL_X32 FILLER_60_3350 ();
 FILLCELL_X32 FILLER_60_3382 ();
 FILLCELL_X32 FILLER_60_3414 ();
 FILLCELL_X32 FILLER_60_3446 ();
 FILLCELL_X32 FILLER_60_3478 ();
 FILLCELL_X32 FILLER_60_3510 ();
 FILLCELL_X32 FILLER_60_3542 ();
 FILLCELL_X32 FILLER_60_3574 ();
 FILLCELL_X32 FILLER_60_3606 ();
 FILLCELL_X32 FILLER_60_3638 ();
 FILLCELL_X32 FILLER_60_3670 ();
 FILLCELL_X32 FILLER_60_3702 ();
 FILLCELL_X4 FILLER_60_3734 ();
 FILLCELL_X32 FILLER_61_1 ();
 FILLCELL_X32 FILLER_61_33 ();
 FILLCELL_X32 FILLER_61_65 ();
 FILLCELL_X32 FILLER_61_97 ();
 FILLCELL_X32 FILLER_61_129 ();
 FILLCELL_X32 FILLER_61_161 ();
 FILLCELL_X32 FILLER_61_193 ();
 FILLCELL_X32 FILLER_61_225 ();
 FILLCELL_X32 FILLER_61_257 ();
 FILLCELL_X32 FILLER_61_289 ();
 FILLCELL_X32 FILLER_61_321 ();
 FILLCELL_X32 FILLER_61_353 ();
 FILLCELL_X32 FILLER_61_385 ();
 FILLCELL_X32 FILLER_61_417 ();
 FILLCELL_X32 FILLER_61_449 ();
 FILLCELL_X32 FILLER_61_481 ();
 FILLCELL_X32 FILLER_61_513 ();
 FILLCELL_X32 FILLER_61_545 ();
 FILLCELL_X32 FILLER_61_577 ();
 FILLCELL_X32 FILLER_61_609 ();
 FILLCELL_X32 FILLER_61_641 ();
 FILLCELL_X32 FILLER_61_673 ();
 FILLCELL_X32 FILLER_61_705 ();
 FILLCELL_X32 FILLER_61_737 ();
 FILLCELL_X32 FILLER_61_769 ();
 FILLCELL_X32 FILLER_61_801 ();
 FILLCELL_X32 FILLER_61_833 ();
 FILLCELL_X32 FILLER_61_865 ();
 FILLCELL_X32 FILLER_61_897 ();
 FILLCELL_X32 FILLER_61_929 ();
 FILLCELL_X32 FILLER_61_961 ();
 FILLCELL_X32 FILLER_61_993 ();
 FILLCELL_X32 FILLER_61_1025 ();
 FILLCELL_X32 FILLER_61_1057 ();
 FILLCELL_X32 FILLER_61_1089 ();
 FILLCELL_X32 FILLER_61_1121 ();
 FILLCELL_X32 FILLER_61_1153 ();
 FILLCELL_X32 FILLER_61_1185 ();
 FILLCELL_X32 FILLER_61_1217 ();
 FILLCELL_X8 FILLER_61_1249 ();
 FILLCELL_X4 FILLER_61_1257 ();
 FILLCELL_X2 FILLER_61_1261 ();
 FILLCELL_X32 FILLER_61_1264 ();
 FILLCELL_X32 FILLER_61_1296 ();
 FILLCELL_X32 FILLER_61_1328 ();
 FILLCELL_X32 FILLER_61_1360 ();
 FILLCELL_X32 FILLER_61_1392 ();
 FILLCELL_X32 FILLER_61_1424 ();
 FILLCELL_X32 FILLER_61_1456 ();
 FILLCELL_X32 FILLER_61_1488 ();
 FILLCELL_X32 FILLER_61_1520 ();
 FILLCELL_X32 FILLER_61_1552 ();
 FILLCELL_X32 FILLER_61_1584 ();
 FILLCELL_X32 FILLER_61_1616 ();
 FILLCELL_X32 FILLER_61_1648 ();
 FILLCELL_X32 FILLER_61_1680 ();
 FILLCELL_X32 FILLER_61_1712 ();
 FILLCELL_X32 FILLER_61_1744 ();
 FILLCELL_X32 FILLER_61_1776 ();
 FILLCELL_X32 FILLER_61_1808 ();
 FILLCELL_X32 FILLER_61_1840 ();
 FILLCELL_X32 FILLER_61_1872 ();
 FILLCELL_X32 FILLER_61_1904 ();
 FILLCELL_X32 FILLER_61_1936 ();
 FILLCELL_X32 FILLER_61_1968 ();
 FILLCELL_X32 FILLER_61_2000 ();
 FILLCELL_X32 FILLER_61_2032 ();
 FILLCELL_X32 FILLER_61_2064 ();
 FILLCELL_X32 FILLER_61_2096 ();
 FILLCELL_X32 FILLER_61_2128 ();
 FILLCELL_X32 FILLER_61_2160 ();
 FILLCELL_X32 FILLER_61_2192 ();
 FILLCELL_X32 FILLER_61_2224 ();
 FILLCELL_X32 FILLER_61_2256 ();
 FILLCELL_X32 FILLER_61_2288 ();
 FILLCELL_X32 FILLER_61_2320 ();
 FILLCELL_X32 FILLER_61_2352 ();
 FILLCELL_X32 FILLER_61_2384 ();
 FILLCELL_X32 FILLER_61_2416 ();
 FILLCELL_X32 FILLER_61_2448 ();
 FILLCELL_X32 FILLER_61_2480 ();
 FILLCELL_X8 FILLER_61_2512 ();
 FILLCELL_X4 FILLER_61_2520 ();
 FILLCELL_X2 FILLER_61_2524 ();
 FILLCELL_X32 FILLER_61_2527 ();
 FILLCELL_X32 FILLER_61_2559 ();
 FILLCELL_X32 FILLER_61_2591 ();
 FILLCELL_X32 FILLER_61_2623 ();
 FILLCELL_X32 FILLER_61_2655 ();
 FILLCELL_X32 FILLER_61_2687 ();
 FILLCELL_X32 FILLER_61_2719 ();
 FILLCELL_X32 FILLER_61_2751 ();
 FILLCELL_X32 FILLER_61_2783 ();
 FILLCELL_X32 FILLER_61_2815 ();
 FILLCELL_X32 FILLER_61_2847 ();
 FILLCELL_X32 FILLER_61_2879 ();
 FILLCELL_X32 FILLER_61_2911 ();
 FILLCELL_X32 FILLER_61_2943 ();
 FILLCELL_X32 FILLER_61_2975 ();
 FILLCELL_X32 FILLER_61_3007 ();
 FILLCELL_X32 FILLER_61_3039 ();
 FILLCELL_X32 FILLER_61_3071 ();
 FILLCELL_X32 FILLER_61_3103 ();
 FILLCELL_X32 FILLER_61_3135 ();
 FILLCELL_X32 FILLER_61_3167 ();
 FILLCELL_X32 FILLER_61_3199 ();
 FILLCELL_X32 FILLER_61_3231 ();
 FILLCELL_X32 FILLER_61_3263 ();
 FILLCELL_X32 FILLER_61_3295 ();
 FILLCELL_X32 FILLER_61_3327 ();
 FILLCELL_X32 FILLER_61_3359 ();
 FILLCELL_X32 FILLER_61_3391 ();
 FILLCELL_X32 FILLER_61_3423 ();
 FILLCELL_X32 FILLER_61_3455 ();
 FILLCELL_X32 FILLER_61_3487 ();
 FILLCELL_X32 FILLER_61_3519 ();
 FILLCELL_X32 FILLER_61_3551 ();
 FILLCELL_X32 FILLER_61_3583 ();
 FILLCELL_X32 FILLER_61_3615 ();
 FILLCELL_X32 FILLER_61_3647 ();
 FILLCELL_X32 FILLER_61_3679 ();
 FILLCELL_X16 FILLER_61_3711 ();
 FILLCELL_X8 FILLER_61_3727 ();
 FILLCELL_X2 FILLER_61_3735 ();
 FILLCELL_X1 FILLER_61_3737 ();
 FILLCELL_X32 FILLER_62_1 ();
 FILLCELL_X32 FILLER_62_33 ();
 FILLCELL_X32 FILLER_62_65 ();
 FILLCELL_X32 FILLER_62_97 ();
 FILLCELL_X32 FILLER_62_129 ();
 FILLCELL_X32 FILLER_62_161 ();
 FILLCELL_X32 FILLER_62_193 ();
 FILLCELL_X32 FILLER_62_225 ();
 FILLCELL_X32 FILLER_62_257 ();
 FILLCELL_X32 FILLER_62_289 ();
 FILLCELL_X32 FILLER_62_321 ();
 FILLCELL_X32 FILLER_62_353 ();
 FILLCELL_X32 FILLER_62_385 ();
 FILLCELL_X32 FILLER_62_417 ();
 FILLCELL_X32 FILLER_62_449 ();
 FILLCELL_X32 FILLER_62_481 ();
 FILLCELL_X32 FILLER_62_513 ();
 FILLCELL_X32 FILLER_62_545 ();
 FILLCELL_X32 FILLER_62_577 ();
 FILLCELL_X16 FILLER_62_609 ();
 FILLCELL_X4 FILLER_62_625 ();
 FILLCELL_X2 FILLER_62_629 ();
 FILLCELL_X32 FILLER_62_632 ();
 FILLCELL_X32 FILLER_62_664 ();
 FILLCELL_X32 FILLER_62_696 ();
 FILLCELL_X32 FILLER_62_728 ();
 FILLCELL_X32 FILLER_62_760 ();
 FILLCELL_X32 FILLER_62_792 ();
 FILLCELL_X32 FILLER_62_824 ();
 FILLCELL_X32 FILLER_62_856 ();
 FILLCELL_X32 FILLER_62_888 ();
 FILLCELL_X32 FILLER_62_920 ();
 FILLCELL_X32 FILLER_62_952 ();
 FILLCELL_X32 FILLER_62_984 ();
 FILLCELL_X32 FILLER_62_1016 ();
 FILLCELL_X32 FILLER_62_1048 ();
 FILLCELL_X32 FILLER_62_1080 ();
 FILLCELL_X32 FILLER_62_1112 ();
 FILLCELL_X32 FILLER_62_1144 ();
 FILLCELL_X32 FILLER_62_1176 ();
 FILLCELL_X32 FILLER_62_1208 ();
 FILLCELL_X32 FILLER_62_1240 ();
 FILLCELL_X32 FILLER_62_1272 ();
 FILLCELL_X32 FILLER_62_1304 ();
 FILLCELL_X32 FILLER_62_1336 ();
 FILLCELL_X32 FILLER_62_1368 ();
 FILLCELL_X32 FILLER_62_1400 ();
 FILLCELL_X32 FILLER_62_1432 ();
 FILLCELL_X32 FILLER_62_1464 ();
 FILLCELL_X32 FILLER_62_1496 ();
 FILLCELL_X32 FILLER_62_1528 ();
 FILLCELL_X32 FILLER_62_1560 ();
 FILLCELL_X32 FILLER_62_1592 ();
 FILLCELL_X32 FILLER_62_1624 ();
 FILLCELL_X32 FILLER_62_1656 ();
 FILLCELL_X32 FILLER_62_1688 ();
 FILLCELL_X32 FILLER_62_1720 ();
 FILLCELL_X32 FILLER_62_1752 ();
 FILLCELL_X32 FILLER_62_1784 ();
 FILLCELL_X32 FILLER_62_1816 ();
 FILLCELL_X32 FILLER_62_1848 ();
 FILLCELL_X8 FILLER_62_1880 ();
 FILLCELL_X4 FILLER_62_1888 ();
 FILLCELL_X2 FILLER_62_1892 ();
 FILLCELL_X32 FILLER_62_1895 ();
 FILLCELL_X32 FILLER_62_1927 ();
 FILLCELL_X32 FILLER_62_1959 ();
 FILLCELL_X32 FILLER_62_1991 ();
 FILLCELL_X32 FILLER_62_2023 ();
 FILLCELL_X32 FILLER_62_2055 ();
 FILLCELL_X32 FILLER_62_2087 ();
 FILLCELL_X32 FILLER_62_2119 ();
 FILLCELL_X32 FILLER_62_2151 ();
 FILLCELL_X32 FILLER_62_2183 ();
 FILLCELL_X32 FILLER_62_2215 ();
 FILLCELL_X32 FILLER_62_2247 ();
 FILLCELL_X32 FILLER_62_2279 ();
 FILLCELL_X32 FILLER_62_2311 ();
 FILLCELL_X32 FILLER_62_2343 ();
 FILLCELL_X32 FILLER_62_2375 ();
 FILLCELL_X32 FILLER_62_2407 ();
 FILLCELL_X32 FILLER_62_2439 ();
 FILLCELL_X32 FILLER_62_2471 ();
 FILLCELL_X32 FILLER_62_2503 ();
 FILLCELL_X32 FILLER_62_2535 ();
 FILLCELL_X32 FILLER_62_2567 ();
 FILLCELL_X32 FILLER_62_2599 ();
 FILLCELL_X32 FILLER_62_2631 ();
 FILLCELL_X32 FILLER_62_2663 ();
 FILLCELL_X32 FILLER_62_2695 ();
 FILLCELL_X32 FILLER_62_2727 ();
 FILLCELL_X32 FILLER_62_2759 ();
 FILLCELL_X32 FILLER_62_2791 ();
 FILLCELL_X32 FILLER_62_2823 ();
 FILLCELL_X32 FILLER_62_2855 ();
 FILLCELL_X32 FILLER_62_2887 ();
 FILLCELL_X32 FILLER_62_2919 ();
 FILLCELL_X32 FILLER_62_2951 ();
 FILLCELL_X32 FILLER_62_2983 ();
 FILLCELL_X32 FILLER_62_3015 ();
 FILLCELL_X32 FILLER_62_3047 ();
 FILLCELL_X32 FILLER_62_3079 ();
 FILLCELL_X32 FILLER_62_3111 ();
 FILLCELL_X8 FILLER_62_3143 ();
 FILLCELL_X4 FILLER_62_3151 ();
 FILLCELL_X2 FILLER_62_3155 ();
 FILLCELL_X32 FILLER_62_3158 ();
 FILLCELL_X32 FILLER_62_3190 ();
 FILLCELL_X32 FILLER_62_3222 ();
 FILLCELL_X32 FILLER_62_3254 ();
 FILLCELL_X32 FILLER_62_3286 ();
 FILLCELL_X32 FILLER_62_3318 ();
 FILLCELL_X32 FILLER_62_3350 ();
 FILLCELL_X32 FILLER_62_3382 ();
 FILLCELL_X32 FILLER_62_3414 ();
 FILLCELL_X32 FILLER_62_3446 ();
 FILLCELL_X32 FILLER_62_3478 ();
 FILLCELL_X32 FILLER_62_3510 ();
 FILLCELL_X32 FILLER_62_3542 ();
 FILLCELL_X32 FILLER_62_3574 ();
 FILLCELL_X32 FILLER_62_3606 ();
 FILLCELL_X32 FILLER_62_3638 ();
 FILLCELL_X32 FILLER_62_3670 ();
 FILLCELL_X32 FILLER_62_3702 ();
 FILLCELL_X4 FILLER_62_3734 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X32 FILLER_63_33 ();
 FILLCELL_X32 FILLER_63_65 ();
 FILLCELL_X32 FILLER_63_97 ();
 FILLCELL_X32 FILLER_63_129 ();
 FILLCELL_X32 FILLER_63_161 ();
 FILLCELL_X32 FILLER_63_193 ();
 FILLCELL_X32 FILLER_63_225 ();
 FILLCELL_X32 FILLER_63_257 ();
 FILLCELL_X32 FILLER_63_289 ();
 FILLCELL_X32 FILLER_63_321 ();
 FILLCELL_X32 FILLER_63_353 ();
 FILLCELL_X32 FILLER_63_385 ();
 FILLCELL_X32 FILLER_63_417 ();
 FILLCELL_X32 FILLER_63_449 ();
 FILLCELL_X32 FILLER_63_481 ();
 FILLCELL_X32 FILLER_63_513 ();
 FILLCELL_X32 FILLER_63_545 ();
 FILLCELL_X32 FILLER_63_577 ();
 FILLCELL_X32 FILLER_63_609 ();
 FILLCELL_X32 FILLER_63_641 ();
 FILLCELL_X32 FILLER_63_673 ();
 FILLCELL_X32 FILLER_63_705 ();
 FILLCELL_X32 FILLER_63_737 ();
 FILLCELL_X32 FILLER_63_769 ();
 FILLCELL_X32 FILLER_63_801 ();
 FILLCELL_X32 FILLER_63_833 ();
 FILLCELL_X32 FILLER_63_865 ();
 FILLCELL_X32 FILLER_63_897 ();
 FILLCELL_X32 FILLER_63_929 ();
 FILLCELL_X32 FILLER_63_961 ();
 FILLCELL_X32 FILLER_63_993 ();
 FILLCELL_X32 FILLER_63_1025 ();
 FILLCELL_X32 FILLER_63_1057 ();
 FILLCELL_X32 FILLER_63_1089 ();
 FILLCELL_X32 FILLER_63_1121 ();
 FILLCELL_X32 FILLER_63_1153 ();
 FILLCELL_X32 FILLER_63_1185 ();
 FILLCELL_X32 FILLER_63_1217 ();
 FILLCELL_X8 FILLER_63_1249 ();
 FILLCELL_X4 FILLER_63_1257 ();
 FILLCELL_X2 FILLER_63_1261 ();
 FILLCELL_X32 FILLER_63_1264 ();
 FILLCELL_X32 FILLER_63_1296 ();
 FILLCELL_X32 FILLER_63_1328 ();
 FILLCELL_X32 FILLER_63_1360 ();
 FILLCELL_X32 FILLER_63_1392 ();
 FILLCELL_X32 FILLER_63_1424 ();
 FILLCELL_X32 FILLER_63_1456 ();
 FILLCELL_X32 FILLER_63_1488 ();
 FILLCELL_X32 FILLER_63_1520 ();
 FILLCELL_X32 FILLER_63_1552 ();
 FILLCELL_X32 FILLER_63_1584 ();
 FILLCELL_X32 FILLER_63_1616 ();
 FILLCELL_X32 FILLER_63_1648 ();
 FILLCELL_X32 FILLER_63_1680 ();
 FILLCELL_X32 FILLER_63_1712 ();
 FILLCELL_X32 FILLER_63_1744 ();
 FILLCELL_X32 FILLER_63_1776 ();
 FILLCELL_X32 FILLER_63_1808 ();
 FILLCELL_X32 FILLER_63_1840 ();
 FILLCELL_X32 FILLER_63_1872 ();
 FILLCELL_X32 FILLER_63_1904 ();
 FILLCELL_X32 FILLER_63_1936 ();
 FILLCELL_X32 FILLER_63_1968 ();
 FILLCELL_X32 FILLER_63_2000 ();
 FILLCELL_X32 FILLER_63_2032 ();
 FILLCELL_X32 FILLER_63_2064 ();
 FILLCELL_X32 FILLER_63_2096 ();
 FILLCELL_X32 FILLER_63_2128 ();
 FILLCELL_X32 FILLER_63_2160 ();
 FILLCELL_X32 FILLER_63_2192 ();
 FILLCELL_X32 FILLER_63_2224 ();
 FILLCELL_X32 FILLER_63_2256 ();
 FILLCELL_X32 FILLER_63_2288 ();
 FILLCELL_X32 FILLER_63_2320 ();
 FILLCELL_X32 FILLER_63_2352 ();
 FILLCELL_X32 FILLER_63_2384 ();
 FILLCELL_X32 FILLER_63_2416 ();
 FILLCELL_X32 FILLER_63_2448 ();
 FILLCELL_X32 FILLER_63_2480 ();
 FILLCELL_X8 FILLER_63_2512 ();
 FILLCELL_X4 FILLER_63_2520 ();
 FILLCELL_X2 FILLER_63_2524 ();
 FILLCELL_X32 FILLER_63_2527 ();
 FILLCELL_X32 FILLER_63_2559 ();
 FILLCELL_X32 FILLER_63_2591 ();
 FILLCELL_X32 FILLER_63_2623 ();
 FILLCELL_X32 FILLER_63_2655 ();
 FILLCELL_X32 FILLER_63_2687 ();
 FILLCELL_X32 FILLER_63_2719 ();
 FILLCELL_X32 FILLER_63_2751 ();
 FILLCELL_X32 FILLER_63_2783 ();
 FILLCELL_X32 FILLER_63_2815 ();
 FILLCELL_X32 FILLER_63_2847 ();
 FILLCELL_X32 FILLER_63_2879 ();
 FILLCELL_X32 FILLER_63_2911 ();
 FILLCELL_X32 FILLER_63_2943 ();
 FILLCELL_X32 FILLER_63_2975 ();
 FILLCELL_X32 FILLER_63_3007 ();
 FILLCELL_X32 FILLER_63_3039 ();
 FILLCELL_X32 FILLER_63_3071 ();
 FILLCELL_X32 FILLER_63_3103 ();
 FILLCELL_X32 FILLER_63_3135 ();
 FILLCELL_X32 FILLER_63_3167 ();
 FILLCELL_X32 FILLER_63_3199 ();
 FILLCELL_X32 FILLER_63_3231 ();
 FILLCELL_X32 FILLER_63_3263 ();
 FILLCELL_X32 FILLER_63_3295 ();
 FILLCELL_X32 FILLER_63_3327 ();
 FILLCELL_X32 FILLER_63_3359 ();
 FILLCELL_X32 FILLER_63_3391 ();
 FILLCELL_X32 FILLER_63_3423 ();
 FILLCELL_X32 FILLER_63_3455 ();
 FILLCELL_X32 FILLER_63_3487 ();
 FILLCELL_X32 FILLER_63_3519 ();
 FILLCELL_X32 FILLER_63_3551 ();
 FILLCELL_X32 FILLER_63_3583 ();
 FILLCELL_X32 FILLER_63_3615 ();
 FILLCELL_X32 FILLER_63_3647 ();
 FILLCELL_X32 FILLER_63_3679 ();
 FILLCELL_X16 FILLER_63_3711 ();
 FILLCELL_X8 FILLER_63_3727 ();
 FILLCELL_X2 FILLER_63_3735 ();
 FILLCELL_X1 FILLER_63_3737 ();
 FILLCELL_X32 FILLER_64_1 ();
 FILLCELL_X32 FILLER_64_33 ();
 FILLCELL_X32 FILLER_64_65 ();
 FILLCELL_X32 FILLER_64_97 ();
 FILLCELL_X32 FILLER_64_129 ();
 FILLCELL_X32 FILLER_64_161 ();
 FILLCELL_X32 FILLER_64_193 ();
 FILLCELL_X32 FILLER_64_225 ();
 FILLCELL_X32 FILLER_64_257 ();
 FILLCELL_X32 FILLER_64_289 ();
 FILLCELL_X32 FILLER_64_321 ();
 FILLCELL_X32 FILLER_64_353 ();
 FILLCELL_X32 FILLER_64_385 ();
 FILLCELL_X32 FILLER_64_417 ();
 FILLCELL_X32 FILLER_64_449 ();
 FILLCELL_X32 FILLER_64_481 ();
 FILLCELL_X32 FILLER_64_513 ();
 FILLCELL_X32 FILLER_64_545 ();
 FILLCELL_X32 FILLER_64_577 ();
 FILLCELL_X16 FILLER_64_609 ();
 FILLCELL_X4 FILLER_64_625 ();
 FILLCELL_X2 FILLER_64_629 ();
 FILLCELL_X32 FILLER_64_632 ();
 FILLCELL_X32 FILLER_64_664 ();
 FILLCELL_X32 FILLER_64_696 ();
 FILLCELL_X32 FILLER_64_728 ();
 FILLCELL_X32 FILLER_64_760 ();
 FILLCELL_X32 FILLER_64_792 ();
 FILLCELL_X32 FILLER_64_824 ();
 FILLCELL_X32 FILLER_64_856 ();
 FILLCELL_X32 FILLER_64_888 ();
 FILLCELL_X32 FILLER_64_920 ();
 FILLCELL_X32 FILLER_64_952 ();
 FILLCELL_X32 FILLER_64_984 ();
 FILLCELL_X32 FILLER_64_1016 ();
 FILLCELL_X32 FILLER_64_1048 ();
 FILLCELL_X32 FILLER_64_1080 ();
 FILLCELL_X32 FILLER_64_1112 ();
 FILLCELL_X32 FILLER_64_1144 ();
 FILLCELL_X32 FILLER_64_1176 ();
 FILLCELL_X32 FILLER_64_1208 ();
 FILLCELL_X32 FILLER_64_1240 ();
 FILLCELL_X32 FILLER_64_1272 ();
 FILLCELL_X32 FILLER_64_1304 ();
 FILLCELL_X32 FILLER_64_1336 ();
 FILLCELL_X32 FILLER_64_1368 ();
 FILLCELL_X32 FILLER_64_1400 ();
 FILLCELL_X32 FILLER_64_1432 ();
 FILLCELL_X32 FILLER_64_1464 ();
 FILLCELL_X32 FILLER_64_1496 ();
 FILLCELL_X32 FILLER_64_1528 ();
 FILLCELL_X32 FILLER_64_1560 ();
 FILLCELL_X32 FILLER_64_1592 ();
 FILLCELL_X32 FILLER_64_1624 ();
 FILLCELL_X32 FILLER_64_1656 ();
 FILLCELL_X32 FILLER_64_1688 ();
 FILLCELL_X32 FILLER_64_1720 ();
 FILLCELL_X32 FILLER_64_1752 ();
 FILLCELL_X32 FILLER_64_1784 ();
 FILLCELL_X32 FILLER_64_1816 ();
 FILLCELL_X32 FILLER_64_1848 ();
 FILLCELL_X8 FILLER_64_1880 ();
 FILLCELL_X4 FILLER_64_1888 ();
 FILLCELL_X2 FILLER_64_1892 ();
 FILLCELL_X32 FILLER_64_1895 ();
 FILLCELL_X32 FILLER_64_1927 ();
 FILLCELL_X32 FILLER_64_1959 ();
 FILLCELL_X32 FILLER_64_1991 ();
 FILLCELL_X32 FILLER_64_2023 ();
 FILLCELL_X32 FILLER_64_2055 ();
 FILLCELL_X32 FILLER_64_2087 ();
 FILLCELL_X32 FILLER_64_2119 ();
 FILLCELL_X32 FILLER_64_2151 ();
 FILLCELL_X32 FILLER_64_2183 ();
 FILLCELL_X32 FILLER_64_2215 ();
 FILLCELL_X32 FILLER_64_2247 ();
 FILLCELL_X32 FILLER_64_2279 ();
 FILLCELL_X32 FILLER_64_2311 ();
 FILLCELL_X32 FILLER_64_2343 ();
 FILLCELL_X32 FILLER_64_2375 ();
 FILLCELL_X32 FILLER_64_2407 ();
 FILLCELL_X32 FILLER_64_2439 ();
 FILLCELL_X32 FILLER_64_2471 ();
 FILLCELL_X32 FILLER_64_2503 ();
 FILLCELL_X32 FILLER_64_2535 ();
 FILLCELL_X32 FILLER_64_2567 ();
 FILLCELL_X32 FILLER_64_2599 ();
 FILLCELL_X32 FILLER_64_2631 ();
 FILLCELL_X32 FILLER_64_2663 ();
 FILLCELL_X32 FILLER_64_2695 ();
 FILLCELL_X32 FILLER_64_2727 ();
 FILLCELL_X32 FILLER_64_2759 ();
 FILLCELL_X32 FILLER_64_2791 ();
 FILLCELL_X32 FILLER_64_2823 ();
 FILLCELL_X32 FILLER_64_2855 ();
 FILLCELL_X32 FILLER_64_2887 ();
 FILLCELL_X32 FILLER_64_2919 ();
 FILLCELL_X32 FILLER_64_2951 ();
 FILLCELL_X32 FILLER_64_2983 ();
 FILLCELL_X32 FILLER_64_3015 ();
 FILLCELL_X32 FILLER_64_3047 ();
 FILLCELL_X32 FILLER_64_3079 ();
 FILLCELL_X32 FILLER_64_3111 ();
 FILLCELL_X8 FILLER_64_3143 ();
 FILLCELL_X4 FILLER_64_3151 ();
 FILLCELL_X2 FILLER_64_3155 ();
 FILLCELL_X32 FILLER_64_3158 ();
 FILLCELL_X32 FILLER_64_3190 ();
 FILLCELL_X32 FILLER_64_3222 ();
 FILLCELL_X32 FILLER_64_3254 ();
 FILLCELL_X32 FILLER_64_3286 ();
 FILLCELL_X32 FILLER_64_3318 ();
 FILLCELL_X32 FILLER_64_3350 ();
 FILLCELL_X32 FILLER_64_3382 ();
 FILLCELL_X32 FILLER_64_3414 ();
 FILLCELL_X32 FILLER_64_3446 ();
 FILLCELL_X32 FILLER_64_3478 ();
 FILLCELL_X32 FILLER_64_3510 ();
 FILLCELL_X32 FILLER_64_3542 ();
 FILLCELL_X32 FILLER_64_3574 ();
 FILLCELL_X32 FILLER_64_3606 ();
 FILLCELL_X32 FILLER_64_3638 ();
 FILLCELL_X32 FILLER_64_3670 ();
 FILLCELL_X32 FILLER_64_3702 ();
 FILLCELL_X4 FILLER_64_3734 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X32 FILLER_65_33 ();
 FILLCELL_X32 FILLER_65_65 ();
 FILLCELL_X32 FILLER_65_97 ();
 FILLCELL_X32 FILLER_65_129 ();
 FILLCELL_X32 FILLER_65_161 ();
 FILLCELL_X32 FILLER_65_193 ();
 FILLCELL_X32 FILLER_65_225 ();
 FILLCELL_X32 FILLER_65_257 ();
 FILLCELL_X32 FILLER_65_289 ();
 FILLCELL_X32 FILLER_65_321 ();
 FILLCELL_X32 FILLER_65_353 ();
 FILLCELL_X32 FILLER_65_385 ();
 FILLCELL_X32 FILLER_65_417 ();
 FILLCELL_X32 FILLER_65_449 ();
 FILLCELL_X32 FILLER_65_481 ();
 FILLCELL_X32 FILLER_65_513 ();
 FILLCELL_X32 FILLER_65_545 ();
 FILLCELL_X32 FILLER_65_577 ();
 FILLCELL_X32 FILLER_65_609 ();
 FILLCELL_X32 FILLER_65_641 ();
 FILLCELL_X32 FILLER_65_673 ();
 FILLCELL_X32 FILLER_65_705 ();
 FILLCELL_X32 FILLER_65_737 ();
 FILLCELL_X32 FILLER_65_769 ();
 FILLCELL_X32 FILLER_65_801 ();
 FILLCELL_X32 FILLER_65_833 ();
 FILLCELL_X32 FILLER_65_865 ();
 FILLCELL_X32 FILLER_65_897 ();
 FILLCELL_X32 FILLER_65_929 ();
 FILLCELL_X32 FILLER_65_961 ();
 FILLCELL_X32 FILLER_65_993 ();
 FILLCELL_X32 FILLER_65_1025 ();
 FILLCELL_X32 FILLER_65_1057 ();
 FILLCELL_X32 FILLER_65_1089 ();
 FILLCELL_X32 FILLER_65_1121 ();
 FILLCELL_X32 FILLER_65_1153 ();
 FILLCELL_X32 FILLER_65_1185 ();
 FILLCELL_X32 FILLER_65_1217 ();
 FILLCELL_X8 FILLER_65_1249 ();
 FILLCELL_X4 FILLER_65_1257 ();
 FILLCELL_X2 FILLER_65_1261 ();
 FILLCELL_X32 FILLER_65_1264 ();
 FILLCELL_X32 FILLER_65_1296 ();
 FILLCELL_X32 FILLER_65_1328 ();
 FILLCELL_X32 FILLER_65_1360 ();
 FILLCELL_X32 FILLER_65_1392 ();
 FILLCELL_X32 FILLER_65_1424 ();
 FILLCELL_X32 FILLER_65_1456 ();
 FILLCELL_X32 FILLER_65_1488 ();
 FILLCELL_X32 FILLER_65_1520 ();
 FILLCELL_X32 FILLER_65_1552 ();
 FILLCELL_X32 FILLER_65_1584 ();
 FILLCELL_X32 FILLER_65_1616 ();
 FILLCELL_X32 FILLER_65_1648 ();
 FILLCELL_X32 FILLER_65_1680 ();
 FILLCELL_X32 FILLER_65_1712 ();
 FILLCELL_X32 FILLER_65_1744 ();
 FILLCELL_X32 FILLER_65_1776 ();
 FILLCELL_X32 FILLER_65_1808 ();
 FILLCELL_X32 FILLER_65_1840 ();
 FILLCELL_X32 FILLER_65_1872 ();
 FILLCELL_X32 FILLER_65_1904 ();
 FILLCELL_X32 FILLER_65_1936 ();
 FILLCELL_X32 FILLER_65_1968 ();
 FILLCELL_X32 FILLER_65_2000 ();
 FILLCELL_X32 FILLER_65_2032 ();
 FILLCELL_X32 FILLER_65_2064 ();
 FILLCELL_X32 FILLER_65_2096 ();
 FILLCELL_X32 FILLER_65_2128 ();
 FILLCELL_X32 FILLER_65_2160 ();
 FILLCELL_X32 FILLER_65_2192 ();
 FILLCELL_X32 FILLER_65_2224 ();
 FILLCELL_X32 FILLER_65_2256 ();
 FILLCELL_X32 FILLER_65_2288 ();
 FILLCELL_X32 FILLER_65_2320 ();
 FILLCELL_X32 FILLER_65_2352 ();
 FILLCELL_X32 FILLER_65_2384 ();
 FILLCELL_X32 FILLER_65_2416 ();
 FILLCELL_X32 FILLER_65_2448 ();
 FILLCELL_X32 FILLER_65_2480 ();
 FILLCELL_X8 FILLER_65_2512 ();
 FILLCELL_X4 FILLER_65_2520 ();
 FILLCELL_X2 FILLER_65_2524 ();
 FILLCELL_X32 FILLER_65_2527 ();
 FILLCELL_X32 FILLER_65_2559 ();
 FILLCELL_X32 FILLER_65_2591 ();
 FILLCELL_X32 FILLER_65_2623 ();
 FILLCELL_X32 FILLER_65_2655 ();
 FILLCELL_X32 FILLER_65_2687 ();
 FILLCELL_X32 FILLER_65_2719 ();
 FILLCELL_X32 FILLER_65_2751 ();
 FILLCELL_X32 FILLER_65_2783 ();
 FILLCELL_X32 FILLER_65_2815 ();
 FILLCELL_X32 FILLER_65_2847 ();
 FILLCELL_X32 FILLER_65_2879 ();
 FILLCELL_X32 FILLER_65_2911 ();
 FILLCELL_X32 FILLER_65_2943 ();
 FILLCELL_X32 FILLER_65_2975 ();
 FILLCELL_X32 FILLER_65_3007 ();
 FILLCELL_X32 FILLER_65_3039 ();
 FILLCELL_X32 FILLER_65_3071 ();
 FILLCELL_X32 FILLER_65_3103 ();
 FILLCELL_X32 FILLER_65_3135 ();
 FILLCELL_X32 FILLER_65_3167 ();
 FILLCELL_X32 FILLER_65_3199 ();
 FILLCELL_X32 FILLER_65_3231 ();
 FILLCELL_X32 FILLER_65_3263 ();
 FILLCELL_X32 FILLER_65_3295 ();
 FILLCELL_X32 FILLER_65_3327 ();
 FILLCELL_X32 FILLER_65_3359 ();
 FILLCELL_X32 FILLER_65_3391 ();
 FILLCELL_X32 FILLER_65_3423 ();
 FILLCELL_X32 FILLER_65_3455 ();
 FILLCELL_X32 FILLER_65_3487 ();
 FILLCELL_X32 FILLER_65_3519 ();
 FILLCELL_X32 FILLER_65_3551 ();
 FILLCELL_X32 FILLER_65_3583 ();
 FILLCELL_X32 FILLER_65_3615 ();
 FILLCELL_X32 FILLER_65_3647 ();
 FILLCELL_X32 FILLER_65_3679 ();
 FILLCELL_X16 FILLER_65_3711 ();
 FILLCELL_X8 FILLER_65_3727 ();
 FILLCELL_X2 FILLER_65_3735 ();
 FILLCELL_X1 FILLER_65_3737 ();
 FILLCELL_X32 FILLER_66_1 ();
 FILLCELL_X32 FILLER_66_33 ();
 FILLCELL_X32 FILLER_66_65 ();
 FILLCELL_X32 FILLER_66_97 ();
 FILLCELL_X32 FILLER_66_129 ();
 FILLCELL_X32 FILLER_66_161 ();
 FILLCELL_X32 FILLER_66_193 ();
 FILLCELL_X32 FILLER_66_225 ();
 FILLCELL_X32 FILLER_66_257 ();
 FILLCELL_X32 FILLER_66_289 ();
 FILLCELL_X32 FILLER_66_321 ();
 FILLCELL_X32 FILLER_66_353 ();
 FILLCELL_X32 FILLER_66_385 ();
 FILLCELL_X32 FILLER_66_417 ();
 FILLCELL_X32 FILLER_66_449 ();
 FILLCELL_X32 FILLER_66_481 ();
 FILLCELL_X32 FILLER_66_513 ();
 FILLCELL_X32 FILLER_66_545 ();
 FILLCELL_X32 FILLER_66_577 ();
 FILLCELL_X16 FILLER_66_609 ();
 FILLCELL_X4 FILLER_66_625 ();
 FILLCELL_X2 FILLER_66_629 ();
 FILLCELL_X32 FILLER_66_632 ();
 FILLCELL_X32 FILLER_66_664 ();
 FILLCELL_X32 FILLER_66_696 ();
 FILLCELL_X32 FILLER_66_728 ();
 FILLCELL_X32 FILLER_66_760 ();
 FILLCELL_X32 FILLER_66_792 ();
 FILLCELL_X32 FILLER_66_824 ();
 FILLCELL_X32 FILLER_66_856 ();
 FILLCELL_X32 FILLER_66_888 ();
 FILLCELL_X32 FILLER_66_920 ();
 FILLCELL_X32 FILLER_66_952 ();
 FILLCELL_X32 FILLER_66_984 ();
 FILLCELL_X32 FILLER_66_1016 ();
 FILLCELL_X32 FILLER_66_1048 ();
 FILLCELL_X32 FILLER_66_1080 ();
 FILLCELL_X32 FILLER_66_1112 ();
 FILLCELL_X32 FILLER_66_1144 ();
 FILLCELL_X32 FILLER_66_1176 ();
 FILLCELL_X32 FILLER_66_1208 ();
 FILLCELL_X32 FILLER_66_1240 ();
 FILLCELL_X32 FILLER_66_1272 ();
 FILLCELL_X32 FILLER_66_1304 ();
 FILLCELL_X32 FILLER_66_1336 ();
 FILLCELL_X32 FILLER_66_1368 ();
 FILLCELL_X32 FILLER_66_1400 ();
 FILLCELL_X32 FILLER_66_1432 ();
 FILLCELL_X32 FILLER_66_1464 ();
 FILLCELL_X32 FILLER_66_1496 ();
 FILLCELL_X32 FILLER_66_1528 ();
 FILLCELL_X32 FILLER_66_1560 ();
 FILLCELL_X32 FILLER_66_1592 ();
 FILLCELL_X32 FILLER_66_1624 ();
 FILLCELL_X32 FILLER_66_1656 ();
 FILLCELL_X32 FILLER_66_1688 ();
 FILLCELL_X32 FILLER_66_1720 ();
 FILLCELL_X32 FILLER_66_1752 ();
 FILLCELL_X32 FILLER_66_1784 ();
 FILLCELL_X32 FILLER_66_1816 ();
 FILLCELL_X32 FILLER_66_1848 ();
 FILLCELL_X8 FILLER_66_1880 ();
 FILLCELL_X4 FILLER_66_1888 ();
 FILLCELL_X2 FILLER_66_1892 ();
 FILLCELL_X32 FILLER_66_1895 ();
 FILLCELL_X32 FILLER_66_1927 ();
 FILLCELL_X32 FILLER_66_1959 ();
 FILLCELL_X32 FILLER_66_1991 ();
 FILLCELL_X32 FILLER_66_2023 ();
 FILLCELL_X32 FILLER_66_2055 ();
 FILLCELL_X32 FILLER_66_2087 ();
 FILLCELL_X32 FILLER_66_2119 ();
 FILLCELL_X32 FILLER_66_2151 ();
 FILLCELL_X32 FILLER_66_2183 ();
 FILLCELL_X32 FILLER_66_2215 ();
 FILLCELL_X32 FILLER_66_2247 ();
 FILLCELL_X32 FILLER_66_2279 ();
 FILLCELL_X32 FILLER_66_2311 ();
 FILLCELL_X32 FILLER_66_2343 ();
 FILLCELL_X32 FILLER_66_2375 ();
 FILLCELL_X32 FILLER_66_2407 ();
 FILLCELL_X32 FILLER_66_2439 ();
 FILLCELL_X32 FILLER_66_2471 ();
 FILLCELL_X32 FILLER_66_2503 ();
 FILLCELL_X32 FILLER_66_2535 ();
 FILLCELL_X32 FILLER_66_2567 ();
 FILLCELL_X32 FILLER_66_2599 ();
 FILLCELL_X32 FILLER_66_2631 ();
 FILLCELL_X32 FILLER_66_2663 ();
 FILLCELL_X32 FILLER_66_2695 ();
 FILLCELL_X32 FILLER_66_2727 ();
 FILLCELL_X32 FILLER_66_2759 ();
 FILLCELL_X32 FILLER_66_2791 ();
 FILLCELL_X32 FILLER_66_2823 ();
 FILLCELL_X32 FILLER_66_2855 ();
 FILLCELL_X32 FILLER_66_2887 ();
 FILLCELL_X32 FILLER_66_2919 ();
 FILLCELL_X32 FILLER_66_2951 ();
 FILLCELL_X32 FILLER_66_2983 ();
 FILLCELL_X32 FILLER_66_3015 ();
 FILLCELL_X32 FILLER_66_3047 ();
 FILLCELL_X32 FILLER_66_3079 ();
 FILLCELL_X32 FILLER_66_3111 ();
 FILLCELL_X8 FILLER_66_3143 ();
 FILLCELL_X4 FILLER_66_3151 ();
 FILLCELL_X2 FILLER_66_3155 ();
 FILLCELL_X32 FILLER_66_3158 ();
 FILLCELL_X32 FILLER_66_3190 ();
 FILLCELL_X32 FILLER_66_3222 ();
 FILLCELL_X32 FILLER_66_3254 ();
 FILLCELL_X32 FILLER_66_3286 ();
 FILLCELL_X32 FILLER_66_3318 ();
 FILLCELL_X32 FILLER_66_3350 ();
 FILLCELL_X32 FILLER_66_3382 ();
 FILLCELL_X32 FILLER_66_3414 ();
 FILLCELL_X32 FILLER_66_3446 ();
 FILLCELL_X32 FILLER_66_3478 ();
 FILLCELL_X32 FILLER_66_3510 ();
 FILLCELL_X32 FILLER_66_3542 ();
 FILLCELL_X32 FILLER_66_3574 ();
 FILLCELL_X32 FILLER_66_3606 ();
 FILLCELL_X32 FILLER_66_3638 ();
 FILLCELL_X32 FILLER_66_3670 ();
 FILLCELL_X32 FILLER_66_3702 ();
 FILLCELL_X4 FILLER_66_3734 ();
 FILLCELL_X32 FILLER_67_1 ();
 FILLCELL_X32 FILLER_67_33 ();
 FILLCELL_X32 FILLER_67_65 ();
 FILLCELL_X32 FILLER_67_97 ();
 FILLCELL_X32 FILLER_67_129 ();
 FILLCELL_X32 FILLER_67_161 ();
 FILLCELL_X32 FILLER_67_193 ();
 FILLCELL_X32 FILLER_67_225 ();
 FILLCELL_X32 FILLER_67_257 ();
 FILLCELL_X32 FILLER_67_289 ();
 FILLCELL_X32 FILLER_67_321 ();
 FILLCELL_X32 FILLER_67_353 ();
 FILLCELL_X32 FILLER_67_385 ();
 FILLCELL_X32 FILLER_67_417 ();
 FILLCELL_X32 FILLER_67_449 ();
 FILLCELL_X32 FILLER_67_481 ();
 FILLCELL_X32 FILLER_67_513 ();
 FILLCELL_X32 FILLER_67_545 ();
 FILLCELL_X32 FILLER_67_577 ();
 FILLCELL_X32 FILLER_67_609 ();
 FILLCELL_X32 FILLER_67_641 ();
 FILLCELL_X32 FILLER_67_673 ();
 FILLCELL_X32 FILLER_67_705 ();
 FILLCELL_X32 FILLER_67_737 ();
 FILLCELL_X32 FILLER_67_769 ();
 FILLCELL_X32 FILLER_67_801 ();
 FILLCELL_X32 FILLER_67_833 ();
 FILLCELL_X32 FILLER_67_865 ();
 FILLCELL_X32 FILLER_67_897 ();
 FILLCELL_X32 FILLER_67_929 ();
 FILLCELL_X32 FILLER_67_961 ();
 FILLCELL_X32 FILLER_67_993 ();
 FILLCELL_X32 FILLER_67_1025 ();
 FILLCELL_X32 FILLER_67_1057 ();
 FILLCELL_X32 FILLER_67_1089 ();
 FILLCELL_X32 FILLER_67_1121 ();
 FILLCELL_X32 FILLER_67_1153 ();
 FILLCELL_X32 FILLER_67_1185 ();
 FILLCELL_X32 FILLER_67_1217 ();
 FILLCELL_X8 FILLER_67_1249 ();
 FILLCELL_X4 FILLER_67_1257 ();
 FILLCELL_X2 FILLER_67_1261 ();
 FILLCELL_X32 FILLER_67_1264 ();
 FILLCELL_X32 FILLER_67_1296 ();
 FILLCELL_X32 FILLER_67_1328 ();
 FILLCELL_X32 FILLER_67_1360 ();
 FILLCELL_X32 FILLER_67_1392 ();
 FILLCELL_X32 FILLER_67_1424 ();
 FILLCELL_X32 FILLER_67_1456 ();
 FILLCELL_X32 FILLER_67_1488 ();
 FILLCELL_X32 FILLER_67_1520 ();
 FILLCELL_X32 FILLER_67_1552 ();
 FILLCELL_X32 FILLER_67_1584 ();
 FILLCELL_X32 FILLER_67_1616 ();
 FILLCELL_X32 FILLER_67_1648 ();
 FILLCELL_X32 FILLER_67_1680 ();
 FILLCELL_X32 FILLER_67_1712 ();
 FILLCELL_X32 FILLER_67_1744 ();
 FILLCELL_X32 FILLER_67_1776 ();
 FILLCELL_X32 FILLER_67_1808 ();
 FILLCELL_X32 FILLER_67_1840 ();
 FILLCELL_X32 FILLER_67_1872 ();
 FILLCELL_X32 FILLER_67_1904 ();
 FILLCELL_X32 FILLER_67_1936 ();
 FILLCELL_X32 FILLER_67_1968 ();
 FILLCELL_X32 FILLER_67_2000 ();
 FILLCELL_X32 FILLER_67_2032 ();
 FILLCELL_X32 FILLER_67_2064 ();
 FILLCELL_X32 FILLER_67_2096 ();
 FILLCELL_X32 FILLER_67_2128 ();
 FILLCELL_X32 FILLER_67_2160 ();
 FILLCELL_X32 FILLER_67_2192 ();
 FILLCELL_X32 FILLER_67_2224 ();
 FILLCELL_X32 FILLER_67_2256 ();
 FILLCELL_X32 FILLER_67_2288 ();
 FILLCELL_X32 FILLER_67_2320 ();
 FILLCELL_X32 FILLER_67_2352 ();
 FILLCELL_X32 FILLER_67_2384 ();
 FILLCELL_X32 FILLER_67_2416 ();
 FILLCELL_X32 FILLER_67_2448 ();
 FILLCELL_X32 FILLER_67_2480 ();
 FILLCELL_X8 FILLER_67_2512 ();
 FILLCELL_X4 FILLER_67_2520 ();
 FILLCELL_X2 FILLER_67_2524 ();
 FILLCELL_X32 FILLER_67_2527 ();
 FILLCELL_X32 FILLER_67_2559 ();
 FILLCELL_X32 FILLER_67_2591 ();
 FILLCELL_X32 FILLER_67_2623 ();
 FILLCELL_X32 FILLER_67_2655 ();
 FILLCELL_X32 FILLER_67_2687 ();
 FILLCELL_X32 FILLER_67_2719 ();
 FILLCELL_X32 FILLER_67_2751 ();
 FILLCELL_X32 FILLER_67_2783 ();
 FILLCELL_X32 FILLER_67_2815 ();
 FILLCELL_X32 FILLER_67_2847 ();
 FILLCELL_X32 FILLER_67_2879 ();
 FILLCELL_X32 FILLER_67_2911 ();
 FILLCELL_X32 FILLER_67_2943 ();
 FILLCELL_X32 FILLER_67_2975 ();
 FILLCELL_X32 FILLER_67_3007 ();
 FILLCELL_X32 FILLER_67_3039 ();
 FILLCELL_X32 FILLER_67_3071 ();
 FILLCELL_X32 FILLER_67_3103 ();
 FILLCELL_X32 FILLER_67_3135 ();
 FILLCELL_X32 FILLER_67_3167 ();
 FILLCELL_X32 FILLER_67_3199 ();
 FILLCELL_X32 FILLER_67_3231 ();
 FILLCELL_X32 FILLER_67_3263 ();
 FILLCELL_X32 FILLER_67_3295 ();
 FILLCELL_X32 FILLER_67_3327 ();
 FILLCELL_X32 FILLER_67_3359 ();
 FILLCELL_X32 FILLER_67_3391 ();
 FILLCELL_X32 FILLER_67_3423 ();
 FILLCELL_X32 FILLER_67_3455 ();
 FILLCELL_X32 FILLER_67_3487 ();
 FILLCELL_X32 FILLER_67_3519 ();
 FILLCELL_X32 FILLER_67_3551 ();
 FILLCELL_X32 FILLER_67_3583 ();
 FILLCELL_X32 FILLER_67_3615 ();
 FILLCELL_X32 FILLER_67_3647 ();
 FILLCELL_X32 FILLER_67_3679 ();
 FILLCELL_X16 FILLER_67_3711 ();
 FILLCELL_X8 FILLER_67_3727 ();
 FILLCELL_X2 FILLER_67_3735 ();
 FILLCELL_X1 FILLER_67_3737 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X32 FILLER_68_33 ();
 FILLCELL_X32 FILLER_68_65 ();
 FILLCELL_X32 FILLER_68_97 ();
 FILLCELL_X32 FILLER_68_129 ();
 FILLCELL_X32 FILLER_68_161 ();
 FILLCELL_X32 FILLER_68_193 ();
 FILLCELL_X32 FILLER_68_225 ();
 FILLCELL_X32 FILLER_68_257 ();
 FILLCELL_X32 FILLER_68_289 ();
 FILLCELL_X32 FILLER_68_321 ();
 FILLCELL_X32 FILLER_68_353 ();
 FILLCELL_X32 FILLER_68_385 ();
 FILLCELL_X32 FILLER_68_417 ();
 FILLCELL_X32 FILLER_68_449 ();
 FILLCELL_X32 FILLER_68_481 ();
 FILLCELL_X32 FILLER_68_513 ();
 FILLCELL_X32 FILLER_68_545 ();
 FILLCELL_X32 FILLER_68_577 ();
 FILLCELL_X16 FILLER_68_609 ();
 FILLCELL_X4 FILLER_68_625 ();
 FILLCELL_X2 FILLER_68_629 ();
 FILLCELL_X32 FILLER_68_632 ();
 FILLCELL_X32 FILLER_68_664 ();
 FILLCELL_X32 FILLER_68_696 ();
 FILLCELL_X32 FILLER_68_728 ();
 FILLCELL_X32 FILLER_68_760 ();
 FILLCELL_X32 FILLER_68_792 ();
 FILLCELL_X32 FILLER_68_824 ();
 FILLCELL_X32 FILLER_68_856 ();
 FILLCELL_X32 FILLER_68_888 ();
 FILLCELL_X32 FILLER_68_920 ();
 FILLCELL_X32 FILLER_68_952 ();
 FILLCELL_X32 FILLER_68_984 ();
 FILLCELL_X32 FILLER_68_1016 ();
 FILLCELL_X32 FILLER_68_1048 ();
 FILLCELL_X32 FILLER_68_1080 ();
 FILLCELL_X32 FILLER_68_1112 ();
 FILLCELL_X32 FILLER_68_1144 ();
 FILLCELL_X32 FILLER_68_1176 ();
 FILLCELL_X32 FILLER_68_1208 ();
 FILLCELL_X32 FILLER_68_1240 ();
 FILLCELL_X32 FILLER_68_1272 ();
 FILLCELL_X32 FILLER_68_1304 ();
 FILLCELL_X32 FILLER_68_1336 ();
 FILLCELL_X32 FILLER_68_1368 ();
 FILLCELL_X32 FILLER_68_1400 ();
 FILLCELL_X32 FILLER_68_1432 ();
 FILLCELL_X32 FILLER_68_1464 ();
 FILLCELL_X32 FILLER_68_1496 ();
 FILLCELL_X32 FILLER_68_1528 ();
 FILLCELL_X32 FILLER_68_1560 ();
 FILLCELL_X32 FILLER_68_1592 ();
 FILLCELL_X32 FILLER_68_1624 ();
 FILLCELL_X32 FILLER_68_1656 ();
 FILLCELL_X32 FILLER_68_1688 ();
 FILLCELL_X32 FILLER_68_1720 ();
 FILLCELL_X32 FILLER_68_1752 ();
 FILLCELL_X32 FILLER_68_1784 ();
 FILLCELL_X32 FILLER_68_1816 ();
 FILLCELL_X32 FILLER_68_1848 ();
 FILLCELL_X8 FILLER_68_1880 ();
 FILLCELL_X4 FILLER_68_1888 ();
 FILLCELL_X2 FILLER_68_1892 ();
 FILLCELL_X32 FILLER_68_1895 ();
 FILLCELL_X32 FILLER_68_1927 ();
 FILLCELL_X32 FILLER_68_1959 ();
 FILLCELL_X32 FILLER_68_1991 ();
 FILLCELL_X32 FILLER_68_2023 ();
 FILLCELL_X32 FILLER_68_2055 ();
 FILLCELL_X32 FILLER_68_2087 ();
 FILLCELL_X32 FILLER_68_2119 ();
 FILLCELL_X32 FILLER_68_2151 ();
 FILLCELL_X32 FILLER_68_2183 ();
 FILLCELL_X32 FILLER_68_2215 ();
 FILLCELL_X32 FILLER_68_2247 ();
 FILLCELL_X32 FILLER_68_2279 ();
 FILLCELL_X32 FILLER_68_2311 ();
 FILLCELL_X32 FILLER_68_2343 ();
 FILLCELL_X32 FILLER_68_2375 ();
 FILLCELL_X32 FILLER_68_2407 ();
 FILLCELL_X32 FILLER_68_2439 ();
 FILLCELL_X32 FILLER_68_2471 ();
 FILLCELL_X32 FILLER_68_2503 ();
 FILLCELL_X32 FILLER_68_2535 ();
 FILLCELL_X32 FILLER_68_2567 ();
 FILLCELL_X32 FILLER_68_2599 ();
 FILLCELL_X32 FILLER_68_2631 ();
 FILLCELL_X32 FILLER_68_2663 ();
 FILLCELL_X32 FILLER_68_2695 ();
 FILLCELL_X32 FILLER_68_2727 ();
 FILLCELL_X32 FILLER_68_2759 ();
 FILLCELL_X32 FILLER_68_2791 ();
 FILLCELL_X32 FILLER_68_2823 ();
 FILLCELL_X32 FILLER_68_2855 ();
 FILLCELL_X32 FILLER_68_2887 ();
 FILLCELL_X32 FILLER_68_2919 ();
 FILLCELL_X32 FILLER_68_2951 ();
 FILLCELL_X32 FILLER_68_2983 ();
 FILLCELL_X32 FILLER_68_3015 ();
 FILLCELL_X32 FILLER_68_3047 ();
 FILLCELL_X32 FILLER_68_3079 ();
 FILLCELL_X32 FILLER_68_3111 ();
 FILLCELL_X8 FILLER_68_3143 ();
 FILLCELL_X4 FILLER_68_3151 ();
 FILLCELL_X2 FILLER_68_3155 ();
 FILLCELL_X32 FILLER_68_3158 ();
 FILLCELL_X32 FILLER_68_3190 ();
 FILLCELL_X32 FILLER_68_3222 ();
 FILLCELL_X32 FILLER_68_3254 ();
 FILLCELL_X32 FILLER_68_3286 ();
 FILLCELL_X32 FILLER_68_3318 ();
 FILLCELL_X32 FILLER_68_3350 ();
 FILLCELL_X32 FILLER_68_3382 ();
 FILLCELL_X32 FILLER_68_3414 ();
 FILLCELL_X32 FILLER_68_3446 ();
 FILLCELL_X32 FILLER_68_3478 ();
 FILLCELL_X32 FILLER_68_3510 ();
 FILLCELL_X32 FILLER_68_3542 ();
 FILLCELL_X32 FILLER_68_3574 ();
 FILLCELL_X32 FILLER_68_3606 ();
 FILLCELL_X32 FILLER_68_3638 ();
 FILLCELL_X32 FILLER_68_3670 ();
 FILLCELL_X32 FILLER_68_3702 ();
 FILLCELL_X4 FILLER_68_3734 ();
 FILLCELL_X32 FILLER_69_1 ();
 FILLCELL_X32 FILLER_69_33 ();
 FILLCELL_X32 FILLER_69_65 ();
 FILLCELL_X32 FILLER_69_97 ();
 FILLCELL_X32 FILLER_69_129 ();
 FILLCELL_X32 FILLER_69_161 ();
 FILLCELL_X32 FILLER_69_193 ();
 FILLCELL_X32 FILLER_69_225 ();
 FILLCELL_X32 FILLER_69_257 ();
 FILLCELL_X32 FILLER_69_289 ();
 FILLCELL_X32 FILLER_69_321 ();
 FILLCELL_X32 FILLER_69_353 ();
 FILLCELL_X32 FILLER_69_385 ();
 FILLCELL_X32 FILLER_69_417 ();
 FILLCELL_X32 FILLER_69_449 ();
 FILLCELL_X32 FILLER_69_481 ();
 FILLCELL_X32 FILLER_69_513 ();
 FILLCELL_X32 FILLER_69_545 ();
 FILLCELL_X32 FILLER_69_577 ();
 FILLCELL_X32 FILLER_69_609 ();
 FILLCELL_X32 FILLER_69_641 ();
 FILLCELL_X32 FILLER_69_673 ();
 FILLCELL_X32 FILLER_69_705 ();
 FILLCELL_X32 FILLER_69_737 ();
 FILLCELL_X32 FILLER_69_769 ();
 FILLCELL_X32 FILLER_69_801 ();
 FILLCELL_X32 FILLER_69_833 ();
 FILLCELL_X32 FILLER_69_865 ();
 FILLCELL_X32 FILLER_69_897 ();
 FILLCELL_X32 FILLER_69_929 ();
 FILLCELL_X32 FILLER_69_961 ();
 FILLCELL_X32 FILLER_69_993 ();
 FILLCELL_X32 FILLER_69_1025 ();
 FILLCELL_X32 FILLER_69_1057 ();
 FILLCELL_X32 FILLER_69_1089 ();
 FILLCELL_X32 FILLER_69_1121 ();
 FILLCELL_X32 FILLER_69_1153 ();
 FILLCELL_X32 FILLER_69_1185 ();
 FILLCELL_X32 FILLER_69_1217 ();
 FILLCELL_X8 FILLER_69_1249 ();
 FILLCELL_X4 FILLER_69_1257 ();
 FILLCELL_X2 FILLER_69_1261 ();
 FILLCELL_X32 FILLER_69_1264 ();
 FILLCELL_X32 FILLER_69_1296 ();
 FILLCELL_X32 FILLER_69_1328 ();
 FILLCELL_X32 FILLER_69_1360 ();
 FILLCELL_X32 FILLER_69_1392 ();
 FILLCELL_X32 FILLER_69_1424 ();
 FILLCELL_X32 FILLER_69_1456 ();
 FILLCELL_X32 FILLER_69_1488 ();
 FILLCELL_X32 FILLER_69_1520 ();
 FILLCELL_X32 FILLER_69_1552 ();
 FILLCELL_X32 FILLER_69_1584 ();
 FILLCELL_X32 FILLER_69_1616 ();
 FILLCELL_X32 FILLER_69_1648 ();
 FILLCELL_X32 FILLER_69_1680 ();
 FILLCELL_X32 FILLER_69_1712 ();
 FILLCELL_X32 FILLER_69_1744 ();
 FILLCELL_X32 FILLER_69_1776 ();
 FILLCELL_X32 FILLER_69_1808 ();
 FILLCELL_X32 FILLER_69_1840 ();
 FILLCELL_X32 FILLER_69_1872 ();
 FILLCELL_X32 FILLER_69_1904 ();
 FILLCELL_X32 FILLER_69_1936 ();
 FILLCELL_X32 FILLER_69_1968 ();
 FILLCELL_X32 FILLER_69_2000 ();
 FILLCELL_X32 FILLER_69_2032 ();
 FILLCELL_X32 FILLER_69_2064 ();
 FILLCELL_X32 FILLER_69_2096 ();
 FILLCELL_X32 FILLER_69_2128 ();
 FILLCELL_X32 FILLER_69_2160 ();
 FILLCELL_X32 FILLER_69_2192 ();
 FILLCELL_X32 FILLER_69_2224 ();
 FILLCELL_X32 FILLER_69_2256 ();
 FILLCELL_X32 FILLER_69_2288 ();
 FILLCELL_X32 FILLER_69_2320 ();
 FILLCELL_X32 FILLER_69_2352 ();
 FILLCELL_X32 FILLER_69_2384 ();
 FILLCELL_X32 FILLER_69_2416 ();
 FILLCELL_X32 FILLER_69_2448 ();
 FILLCELL_X32 FILLER_69_2480 ();
 FILLCELL_X8 FILLER_69_2512 ();
 FILLCELL_X4 FILLER_69_2520 ();
 FILLCELL_X2 FILLER_69_2524 ();
 FILLCELL_X32 FILLER_69_2527 ();
 FILLCELL_X32 FILLER_69_2559 ();
 FILLCELL_X32 FILLER_69_2591 ();
 FILLCELL_X32 FILLER_69_2623 ();
 FILLCELL_X32 FILLER_69_2655 ();
 FILLCELL_X32 FILLER_69_2687 ();
 FILLCELL_X32 FILLER_69_2719 ();
 FILLCELL_X32 FILLER_69_2751 ();
 FILLCELL_X32 FILLER_69_2783 ();
 FILLCELL_X32 FILLER_69_2815 ();
 FILLCELL_X32 FILLER_69_2847 ();
 FILLCELL_X32 FILLER_69_2879 ();
 FILLCELL_X32 FILLER_69_2911 ();
 FILLCELL_X32 FILLER_69_2943 ();
 FILLCELL_X32 FILLER_69_2975 ();
 FILLCELL_X32 FILLER_69_3007 ();
 FILLCELL_X32 FILLER_69_3039 ();
 FILLCELL_X32 FILLER_69_3071 ();
 FILLCELL_X32 FILLER_69_3103 ();
 FILLCELL_X32 FILLER_69_3135 ();
 FILLCELL_X32 FILLER_69_3167 ();
 FILLCELL_X32 FILLER_69_3199 ();
 FILLCELL_X32 FILLER_69_3231 ();
 FILLCELL_X32 FILLER_69_3263 ();
 FILLCELL_X32 FILLER_69_3295 ();
 FILLCELL_X32 FILLER_69_3327 ();
 FILLCELL_X32 FILLER_69_3359 ();
 FILLCELL_X32 FILLER_69_3391 ();
 FILLCELL_X32 FILLER_69_3423 ();
 FILLCELL_X32 FILLER_69_3455 ();
 FILLCELL_X32 FILLER_69_3487 ();
 FILLCELL_X32 FILLER_69_3519 ();
 FILLCELL_X32 FILLER_69_3551 ();
 FILLCELL_X32 FILLER_69_3583 ();
 FILLCELL_X32 FILLER_69_3615 ();
 FILLCELL_X32 FILLER_69_3647 ();
 FILLCELL_X32 FILLER_69_3679 ();
 FILLCELL_X16 FILLER_69_3711 ();
 FILLCELL_X8 FILLER_69_3727 ();
 FILLCELL_X2 FILLER_69_3735 ();
 FILLCELL_X1 FILLER_69_3737 ();
 FILLCELL_X32 FILLER_70_1 ();
 FILLCELL_X32 FILLER_70_33 ();
 FILLCELL_X32 FILLER_70_65 ();
 FILLCELL_X32 FILLER_70_97 ();
 FILLCELL_X32 FILLER_70_129 ();
 FILLCELL_X32 FILLER_70_161 ();
 FILLCELL_X32 FILLER_70_193 ();
 FILLCELL_X32 FILLER_70_225 ();
 FILLCELL_X32 FILLER_70_257 ();
 FILLCELL_X32 FILLER_70_289 ();
 FILLCELL_X32 FILLER_70_321 ();
 FILLCELL_X32 FILLER_70_353 ();
 FILLCELL_X32 FILLER_70_385 ();
 FILLCELL_X32 FILLER_70_417 ();
 FILLCELL_X32 FILLER_70_449 ();
 FILLCELL_X32 FILLER_70_481 ();
 FILLCELL_X32 FILLER_70_513 ();
 FILLCELL_X32 FILLER_70_545 ();
 FILLCELL_X32 FILLER_70_577 ();
 FILLCELL_X16 FILLER_70_609 ();
 FILLCELL_X4 FILLER_70_625 ();
 FILLCELL_X2 FILLER_70_629 ();
 FILLCELL_X32 FILLER_70_632 ();
 FILLCELL_X32 FILLER_70_664 ();
 FILLCELL_X32 FILLER_70_696 ();
 FILLCELL_X32 FILLER_70_728 ();
 FILLCELL_X32 FILLER_70_760 ();
 FILLCELL_X32 FILLER_70_792 ();
 FILLCELL_X32 FILLER_70_824 ();
 FILLCELL_X32 FILLER_70_856 ();
 FILLCELL_X32 FILLER_70_888 ();
 FILLCELL_X32 FILLER_70_920 ();
 FILLCELL_X32 FILLER_70_952 ();
 FILLCELL_X32 FILLER_70_984 ();
 FILLCELL_X32 FILLER_70_1016 ();
 FILLCELL_X32 FILLER_70_1048 ();
 FILLCELL_X32 FILLER_70_1080 ();
 FILLCELL_X32 FILLER_70_1112 ();
 FILLCELL_X32 FILLER_70_1144 ();
 FILLCELL_X32 FILLER_70_1176 ();
 FILLCELL_X32 FILLER_70_1208 ();
 FILLCELL_X32 FILLER_70_1240 ();
 FILLCELL_X32 FILLER_70_1272 ();
 FILLCELL_X32 FILLER_70_1304 ();
 FILLCELL_X32 FILLER_70_1336 ();
 FILLCELL_X32 FILLER_70_1368 ();
 FILLCELL_X32 FILLER_70_1400 ();
 FILLCELL_X32 FILLER_70_1432 ();
 FILLCELL_X32 FILLER_70_1464 ();
 FILLCELL_X32 FILLER_70_1496 ();
 FILLCELL_X32 FILLER_70_1528 ();
 FILLCELL_X32 FILLER_70_1560 ();
 FILLCELL_X32 FILLER_70_1592 ();
 FILLCELL_X32 FILLER_70_1624 ();
 FILLCELL_X32 FILLER_70_1656 ();
 FILLCELL_X32 FILLER_70_1688 ();
 FILLCELL_X32 FILLER_70_1720 ();
 FILLCELL_X32 FILLER_70_1752 ();
 FILLCELL_X32 FILLER_70_1784 ();
 FILLCELL_X32 FILLER_70_1816 ();
 FILLCELL_X32 FILLER_70_1848 ();
 FILLCELL_X8 FILLER_70_1880 ();
 FILLCELL_X4 FILLER_70_1888 ();
 FILLCELL_X2 FILLER_70_1892 ();
 FILLCELL_X32 FILLER_70_1895 ();
 FILLCELL_X32 FILLER_70_1927 ();
 FILLCELL_X32 FILLER_70_1959 ();
 FILLCELL_X32 FILLER_70_1991 ();
 FILLCELL_X32 FILLER_70_2023 ();
 FILLCELL_X32 FILLER_70_2055 ();
 FILLCELL_X32 FILLER_70_2087 ();
 FILLCELL_X32 FILLER_70_2119 ();
 FILLCELL_X32 FILLER_70_2151 ();
 FILLCELL_X32 FILLER_70_2183 ();
 FILLCELL_X32 FILLER_70_2215 ();
 FILLCELL_X32 FILLER_70_2247 ();
 FILLCELL_X32 FILLER_70_2279 ();
 FILLCELL_X32 FILLER_70_2311 ();
 FILLCELL_X32 FILLER_70_2343 ();
 FILLCELL_X32 FILLER_70_2375 ();
 FILLCELL_X32 FILLER_70_2407 ();
 FILLCELL_X32 FILLER_70_2439 ();
 FILLCELL_X32 FILLER_70_2471 ();
 FILLCELL_X32 FILLER_70_2503 ();
 FILLCELL_X32 FILLER_70_2535 ();
 FILLCELL_X32 FILLER_70_2567 ();
 FILLCELL_X32 FILLER_70_2599 ();
 FILLCELL_X32 FILLER_70_2631 ();
 FILLCELL_X32 FILLER_70_2663 ();
 FILLCELL_X32 FILLER_70_2695 ();
 FILLCELL_X32 FILLER_70_2727 ();
 FILLCELL_X32 FILLER_70_2759 ();
 FILLCELL_X32 FILLER_70_2791 ();
 FILLCELL_X32 FILLER_70_2823 ();
 FILLCELL_X32 FILLER_70_2855 ();
 FILLCELL_X32 FILLER_70_2887 ();
 FILLCELL_X32 FILLER_70_2919 ();
 FILLCELL_X32 FILLER_70_2951 ();
 FILLCELL_X32 FILLER_70_2983 ();
 FILLCELL_X32 FILLER_70_3015 ();
 FILLCELL_X32 FILLER_70_3047 ();
 FILLCELL_X32 FILLER_70_3079 ();
 FILLCELL_X32 FILLER_70_3111 ();
 FILLCELL_X8 FILLER_70_3143 ();
 FILLCELL_X4 FILLER_70_3151 ();
 FILLCELL_X2 FILLER_70_3155 ();
 FILLCELL_X32 FILLER_70_3158 ();
 FILLCELL_X32 FILLER_70_3190 ();
 FILLCELL_X32 FILLER_70_3222 ();
 FILLCELL_X32 FILLER_70_3254 ();
 FILLCELL_X32 FILLER_70_3286 ();
 FILLCELL_X32 FILLER_70_3318 ();
 FILLCELL_X32 FILLER_70_3350 ();
 FILLCELL_X32 FILLER_70_3382 ();
 FILLCELL_X32 FILLER_70_3414 ();
 FILLCELL_X32 FILLER_70_3446 ();
 FILLCELL_X32 FILLER_70_3478 ();
 FILLCELL_X32 FILLER_70_3510 ();
 FILLCELL_X32 FILLER_70_3542 ();
 FILLCELL_X32 FILLER_70_3574 ();
 FILLCELL_X32 FILLER_70_3606 ();
 FILLCELL_X32 FILLER_70_3638 ();
 FILLCELL_X32 FILLER_70_3670 ();
 FILLCELL_X32 FILLER_70_3702 ();
 FILLCELL_X4 FILLER_70_3734 ();
 FILLCELL_X32 FILLER_71_1 ();
 FILLCELL_X32 FILLER_71_33 ();
 FILLCELL_X32 FILLER_71_65 ();
 FILLCELL_X32 FILLER_71_97 ();
 FILLCELL_X32 FILLER_71_129 ();
 FILLCELL_X32 FILLER_71_161 ();
 FILLCELL_X32 FILLER_71_193 ();
 FILLCELL_X32 FILLER_71_225 ();
 FILLCELL_X32 FILLER_71_257 ();
 FILLCELL_X32 FILLER_71_289 ();
 FILLCELL_X32 FILLER_71_321 ();
 FILLCELL_X32 FILLER_71_353 ();
 FILLCELL_X32 FILLER_71_385 ();
 FILLCELL_X32 FILLER_71_417 ();
 FILLCELL_X32 FILLER_71_449 ();
 FILLCELL_X32 FILLER_71_481 ();
 FILLCELL_X32 FILLER_71_513 ();
 FILLCELL_X32 FILLER_71_545 ();
 FILLCELL_X32 FILLER_71_577 ();
 FILLCELL_X32 FILLER_71_609 ();
 FILLCELL_X32 FILLER_71_641 ();
 FILLCELL_X32 FILLER_71_673 ();
 FILLCELL_X32 FILLER_71_705 ();
 FILLCELL_X32 FILLER_71_737 ();
 FILLCELL_X32 FILLER_71_769 ();
 FILLCELL_X32 FILLER_71_801 ();
 FILLCELL_X32 FILLER_71_833 ();
 FILLCELL_X32 FILLER_71_865 ();
 FILLCELL_X32 FILLER_71_897 ();
 FILLCELL_X32 FILLER_71_929 ();
 FILLCELL_X32 FILLER_71_961 ();
 FILLCELL_X32 FILLER_71_993 ();
 FILLCELL_X32 FILLER_71_1025 ();
 FILLCELL_X32 FILLER_71_1057 ();
 FILLCELL_X32 FILLER_71_1089 ();
 FILLCELL_X32 FILLER_71_1121 ();
 FILLCELL_X32 FILLER_71_1153 ();
 FILLCELL_X32 FILLER_71_1185 ();
 FILLCELL_X32 FILLER_71_1217 ();
 FILLCELL_X8 FILLER_71_1249 ();
 FILLCELL_X4 FILLER_71_1257 ();
 FILLCELL_X2 FILLER_71_1261 ();
 FILLCELL_X32 FILLER_71_1264 ();
 FILLCELL_X32 FILLER_71_1296 ();
 FILLCELL_X32 FILLER_71_1328 ();
 FILLCELL_X32 FILLER_71_1360 ();
 FILLCELL_X32 FILLER_71_1392 ();
 FILLCELL_X32 FILLER_71_1424 ();
 FILLCELL_X32 FILLER_71_1456 ();
 FILLCELL_X32 FILLER_71_1488 ();
 FILLCELL_X32 FILLER_71_1520 ();
 FILLCELL_X32 FILLER_71_1552 ();
 FILLCELL_X32 FILLER_71_1584 ();
 FILLCELL_X32 FILLER_71_1616 ();
 FILLCELL_X32 FILLER_71_1648 ();
 FILLCELL_X32 FILLER_71_1680 ();
 FILLCELL_X32 FILLER_71_1712 ();
 FILLCELL_X32 FILLER_71_1744 ();
 FILLCELL_X32 FILLER_71_1776 ();
 FILLCELL_X32 FILLER_71_1808 ();
 FILLCELL_X32 FILLER_71_1840 ();
 FILLCELL_X32 FILLER_71_1872 ();
 FILLCELL_X32 FILLER_71_1904 ();
 FILLCELL_X32 FILLER_71_1936 ();
 FILLCELL_X32 FILLER_71_1968 ();
 FILLCELL_X32 FILLER_71_2000 ();
 FILLCELL_X32 FILLER_71_2032 ();
 FILLCELL_X32 FILLER_71_2064 ();
 FILLCELL_X32 FILLER_71_2096 ();
 FILLCELL_X32 FILLER_71_2128 ();
 FILLCELL_X32 FILLER_71_2160 ();
 FILLCELL_X32 FILLER_71_2192 ();
 FILLCELL_X32 FILLER_71_2224 ();
 FILLCELL_X32 FILLER_71_2256 ();
 FILLCELL_X32 FILLER_71_2288 ();
 FILLCELL_X32 FILLER_71_2320 ();
 FILLCELL_X32 FILLER_71_2352 ();
 FILLCELL_X32 FILLER_71_2384 ();
 FILLCELL_X32 FILLER_71_2416 ();
 FILLCELL_X32 FILLER_71_2448 ();
 FILLCELL_X32 FILLER_71_2480 ();
 FILLCELL_X8 FILLER_71_2512 ();
 FILLCELL_X4 FILLER_71_2520 ();
 FILLCELL_X2 FILLER_71_2524 ();
 FILLCELL_X32 FILLER_71_2527 ();
 FILLCELL_X32 FILLER_71_2559 ();
 FILLCELL_X32 FILLER_71_2591 ();
 FILLCELL_X32 FILLER_71_2623 ();
 FILLCELL_X32 FILLER_71_2655 ();
 FILLCELL_X32 FILLER_71_2687 ();
 FILLCELL_X32 FILLER_71_2719 ();
 FILLCELL_X32 FILLER_71_2751 ();
 FILLCELL_X32 FILLER_71_2783 ();
 FILLCELL_X32 FILLER_71_2815 ();
 FILLCELL_X32 FILLER_71_2847 ();
 FILLCELL_X32 FILLER_71_2879 ();
 FILLCELL_X32 FILLER_71_2911 ();
 FILLCELL_X32 FILLER_71_2943 ();
 FILLCELL_X32 FILLER_71_2975 ();
 FILLCELL_X32 FILLER_71_3007 ();
 FILLCELL_X32 FILLER_71_3039 ();
 FILLCELL_X32 FILLER_71_3071 ();
 FILLCELL_X32 FILLER_71_3103 ();
 FILLCELL_X32 FILLER_71_3135 ();
 FILLCELL_X32 FILLER_71_3167 ();
 FILLCELL_X32 FILLER_71_3199 ();
 FILLCELL_X32 FILLER_71_3231 ();
 FILLCELL_X32 FILLER_71_3263 ();
 FILLCELL_X32 FILLER_71_3295 ();
 FILLCELL_X32 FILLER_71_3327 ();
 FILLCELL_X32 FILLER_71_3359 ();
 FILLCELL_X32 FILLER_71_3391 ();
 FILLCELL_X32 FILLER_71_3423 ();
 FILLCELL_X32 FILLER_71_3455 ();
 FILLCELL_X32 FILLER_71_3487 ();
 FILLCELL_X32 FILLER_71_3519 ();
 FILLCELL_X32 FILLER_71_3551 ();
 FILLCELL_X32 FILLER_71_3583 ();
 FILLCELL_X32 FILLER_71_3615 ();
 FILLCELL_X32 FILLER_71_3647 ();
 FILLCELL_X32 FILLER_71_3679 ();
 FILLCELL_X16 FILLER_71_3711 ();
 FILLCELL_X8 FILLER_71_3727 ();
 FILLCELL_X2 FILLER_71_3735 ();
 FILLCELL_X1 FILLER_71_3737 ();
 FILLCELL_X32 FILLER_72_1 ();
 FILLCELL_X32 FILLER_72_33 ();
 FILLCELL_X32 FILLER_72_65 ();
 FILLCELL_X32 FILLER_72_97 ();
 FILLCELL_X32 FILLER_72_129 ();
 FILLCELL_X32 FILLER_72_161 ();
 FILLCELL_X32 FILLER_72_193 ();
 FILLCELL_X32 FILLER_72_225 ();
 FILLCELL_X32 FILLER_72_257 ();
 FILLCELL_X32 FILLER_72_289 ();
 FILLCELL_X32 FILLER_72_321 ();
 FILLCELL_X32 FILLER_72_353 ();
 FILLCELL_X32 FILLER_72_385 ();
 FILLCELL_X32 FILLER_72_417 ();
 FILLCELL_X32 FILLER_72_449 ();
 FILLCELL_X32 FILLER_72_481 ();
 FILLCELL_X32 FILLER_72_513 ();
 FILLCELL_X32 FILLER_72_545 ();
 FILLCELL_X32 FILLER_72_577 ();
 FILLCELL_X16 FILLER_72_609 ();
 FILLCELL_X4 FILLER_72_625 ();
 FILLCELL_X2 FILLER_72_629 ();
 FILLCELL_X32 FILLER_72_632 ();
 FILLCELL_X32 FILLER_72_664 ();
 FILLCELL_X32 FILLER_72_696 ();
 FILLCELL_X32 FILLER_72_728 ();
 FILLCELL_X32 FILLER_72_760 ();
 FILLCELL_X32 FILLER_72_792 ();
 FILLCELL_X32 FILLER_72_824 ();
 FILLCELL_X32 FILLER_72_856 ();
 FILLCELL_X32 FILLER_72_888 ();
 FILLCELL_X32 FILLER_72_920 ();
 FILLCELL_X32 FILLER_72_952 ();
 FILLCELL_X32 FILLER_72_984 ();
 FILLCELL_X32 FILLER_72_1016 ();
 FILLCELL_X32 FILLER_72_1048 ();
 FILLCELL_X32 FILLER_72_1080 ();
 FILLCELL_X32 FILLER_72_1112 ();
 FILLCELL_X32 FILLER_72_1144 ();
 FILLCELL_X32 FILLER_72_1176 ();
 FILLCELL_X32 FILLER_72_1208 ();
 FILLCELL_X32 FILLER_72_1240 ();
 FILLCELL_X32 FILLER_72_1272 ();
 FILLCELL_X32 FILLER_72_1304 ();
 FILLCELL_X32 FILLER_72_1336 ();
 FILLCELL_X32 FILLER_72_1368 ();
 FILLCELL_X32 FILLER_72_1400 ();
 FILLCELL_X32 FILLER_72_1432 ();
 FILLCELL_X32 FILLER_72_1464 ();
 FILLCELL_X32 FILLER_72_1496 ();
 FILLCELL_X32 FILLER_72_1528 ();
 FILLCELL_X32 FILLER_72_1560 ();
 FILLCELL_X32 FILLER_72_1592 ();
 FILLCELL_X32 FILLER_72_1624 ();
 FILLCELL_X32 FILLER_72_1656 ();
 FILLCELL_X32 FILLER_72_1688 ();
 FILLCELL_X32 FILLER_72_1720 ();
 FILLCELL_X32 FILLER_72_1752 ();
 FILLCELL_X32 FILLER_72_1784 ();
 FILLCELL_X32 FILLER_72_1816 ();
 FILLCELL_X32 FILLER_72_1848 ();
 FILLCELL_X8 FILLER_72_1880 ();
 FILLCELL_X4 FILLER_72_1888 ();
 FILLCELL_X2 FILLER_72_1892 ();
 FILLCELL_X32 FILLER_72_1895 ();
 FILLCELL_X32 FILLER_72_1927 ();
 FILLCELL_X32 FILLER_72_1959 ();
 FILLCELL_X32 FILLER_72_1991 ();
 FILLCELL_X32 FILLER_72_2023 ();
 FILLCELL_X32 FILLER_72_2055 ();
 FILLCELL_X32 FILLER_72_2087 ();
 FILLCELL_X32 FILLER_72_2119 ();
 FILLCELL_X32 FILLER_72_2151 ();
 FILLCELL_X32 FILLER_72_2183 ();
 FILLCELL_X32 FILLER_72_2215 ();
 FILLCELL_X32 FILLER_72_2247 ();
 FILLCELL_X32 FILLER_72_2279 ();
 FILLCELL_X32 FILLER_72_2311 ();
 FILLCELL_X32 FILLER_72_2343 ();
 FILLCELL_X32 FILLER_72_2375 ();
 FILLCELL_X32 FILLER_72_2407 ();
 FILLCELL_X32 FILLER_72_2439 ();
 FILLCELL_X32 FILLER_72_2471 ();
 FILLCELL_X32 FILLER_72_2503 ();
 FILLCELL_X32 FILLER_72_2535 ();
 FILLCELL_X32 FILLER_72_2567 ();
 FILLCELL_X32 FILLER_72_2599 ();
 FILLCELL_X32 FILLER_72_2631 ();
 FILLCELL_X32 FILLER_72_2663 ();
 FILLCELL_X32 FILLER_72_2695 ();
 FILLCELL_X32 FILLER_72_2727 ();
 FILLCELL_X32 FILLER_72_2759 ();
 FILLCELL_X32 FILLER_72_2791 ();
 FILLCELL_X32 FILLER_72_2823 ();
 FILLCELL_X32 FILLER_72_2855 ();
 FILLCELL_X32 FILLER_72_2887 ();
 FILLCELL_X32 FILLER_72_2919 ();
 FILLCELL_X32 FILLER_72_2951 ();
 FILLCELL_X32 FILLER_72_2983 ();
 FILLCELL_X32 FILLER_72_3015 ();
 FILLCELL_X32 FILLER_72_3047 ();
 FILLCELL_X32 FILLER_72_3079 ();
 FILLCELL_X32 FILLER_72_3111 ();
 FILLCELL_X8 FILLER_72_3143 ();
 FILLCELL_X4 FILLER_72_3151 ();
 FILLCELL_X2 FILLER_72_3155 ();
 FILLCELL_X32 FILLER_72_3158 ();
 FILLCELL_X32 FILLER_72_3190 ();
 FILLCELL_X32 FILLER_72_3222 ();
 FILLCELL_X32 FILLER_72_3254 ();
 FILLCELL_X32 FILLER_72_3286 ();
 FILLCELL_X32 FILLER_72_3318 ();
 FILLCELL_X32 FILLER_72_3350 ();
 FILLCELL_X32 FILLER_72_3382 ();
 FILLCELL_X32 FILLER_72_3414 ();
 FILLCELL_X32 FILLER_72_3446 ();
 FILLCELL_X32 FILLER_72_3478 ();
 FILLCELL_X32 FILLER_72_3510 ();
 FILLCELL_X32 FILLER_72_3542 ();
 FILLCELL_X32 FILLER_72_3574 ();
 FILLCELL_X32 FILLER_72_3606 ();
 FILLCELL_X32 FILLER_72_3638 ();
 FILLCELL_X32 FILLER_72_3670 ();
 FILLCELL_X32 FILLER_72_3702 ();
 FILLCELL_X4 FILLER_72_3734 ();
 FILLCELL_X32 FILLER_73_1 ();
 FILLCELL_X32 FILLER_73_33 ();
 FILLCELL_X32 FILLER_73_65 ();
 FILLCELL_X32 FILLER_73_97 ();
 FILLCELL_X32 FILLER_73_129 ();
 FILLCELL_X32 FILLER_73_161 ();
 FILLCELL_X32 FILLER_73_193 ();
 FILLCELL_X32 FILLER_73_225 ();
 FILLCELL_X32 FILLER_73_257 ();
 FILLCELL_X32 FILLER_73_289 ();
 FILLCELL_X32 FILLER_73_321 ();
 FILLCELL_X32 FILLER_73_353 ();
 FILLCELL_X32 FILLER_73_385 ();
 FILLCELL_X32 FILLER_73_417 ();
 FILLCELL_X32 FILLER_73_449 ();
 FILLCELL_X32 FILLER_73_481 ();
 FILLCELL_X32 FILLER_73_513 ();
 FILLCELL_X32 FILLER_73_545 ();
 FILLCELL_X32 FILLER_73_577 ();
 FILLCELL_X32 FILLER_73_609 ();
 FILLCELL_X32 FILLER_73_641 ();
 FILLCELL_X32 FILLER_73_673 ();
 FILLCELL_X32 FILLER_73_705 ();
 FILLCELL_X32 FILLER_73_737 ();
 FILLCELL_X32 FILLER_73_769 ();
 FILLCELL_X32 FILLER_73_801 ();
 FILLCELL_X32 FILLER_73_833 ();
 FILLCELL_X32 FILLER_73_865 ();
 FILLCELL_X32 FILLER_73_897 ();
 FILLCELL_X32 FILLER_73_929 ();
 FILLCELL_X32 FILLER_73_961 ();
 FILLCELL_X32 FILLER_73_993 ();
 FILLCELL_X32 FILLER_73_1025 ();
 FILLCELL_X32 FILLER_73_1057 ();
 FILLCELL_X32 FILLER_73_1089 ();
 FILLCELL_X32 FILLER_73_1121 ();
 FILLCELL_X32 FILLER_73_1153 ();
 FILLCELL_X32 FILLER_73_1185 ();
 FILLCELL_X32 FILLER_73_1217 ();
 FILLCELL_X8 FILLER_73_1249 ();
 FILLCELL_X4 FILLER_73_1257 ();
 FILLCELL_X2 FILLER_73_1261 ();
 FILLCELL_X32 FILLER_73_1264 ();
 FILLCELL_X32 FILLER_73_1296 ();
 FILLCELL_X32 FILLER_73_1328 ();
 FILLCELL_X32 FILLER_73_1360 ();
 FILLCELL_X32 FILLER_73_1392 ();
 FILLCELL_X32 FILLER_73_1424 ();
 FILLCELL_X32 FILLER_73_1456 ();
 FILLCELL_X32 FILLER_73_1488 ();
 FILLCELL_X32 FILLER_73_1520 ();
 FILLCELL_X32 FILLER_73_1552 ();
 FILLCELL_X32 FILLER_73_1584 ();
 FILLCELL_X32 FILLER_73_1616 ();
 FILLCELL_X32 FILLER_73_1648 ();
 FILLCELL_X32 FILLER_73_1680 ();
 FILLCELL_X32 FILLER_73_1712 ();
 FILLCELL_X32 FILLER_73_1744 ();
 FILLCELL_X32 FILLER_73_1776 ();
 FILLCELL_X32 FILLER_73_1808 ();
 FILLCELL_X32 FILLER_73_1840 ();
 FILLCELL_X32 FILLER_73_1872 ();
 FILLCELL_X32 FILLER_73_1904 ();
 FILLCELL_X32 FILLER_73_1936 ();
 FILLCELL_X32 FILLER_73_1968 ();
 FILLCELL_X32 FILLER_73_2000 ();
 FILLCELL_X32 FILLER_73_2032 ();
 FILLCELL_X32 FILLER_73_2064 ();
 FILLCELL_X32 FILLER_73_2096 ();
 FILLCELL_X32 FILLER_73_2128 ();
 FILLCELL_X32 FILLER_73_2160 ();
 FILLCELL_X32 FILLER_73_2192 ();
 FILLCELL_X32 FILLER_73_2224 ();
 FILLCELL_X32 FILLER_73_2256 ();
 FILLCELL_X32 FILLER_73_2288 ();
 FILLCELL_X32 FILLER_73_2320 ();
 FILLCELL_X32 FILLER_73_2352 ();
 FILLCELL_X32 FILLER_73_2384 ();
 FILLCELL_X32 FILLER_73_2416 ();
 FILLCELL_X32 FILLER_73_2448 ();
 FILLCELL_X32 FILLER_73_2480 ();
 FILLCELL_X8 FILLER_73_2512 ();
 FILLCELL_X4 FILLER_73_2520 ();
 FILLCELL_X2 FILLER_73_2524 ();
 FILLCELL_X32 FILLER_73_2527 ();
 FILLCELL_X32 FILLER_73_2559 ();
 FILLCELL_X32 FILLER_73_2591 ();
 FILLCELL_X32 FILLER_73_2623 ();
 FILLCELL_X32 FILLER_73_2655 ();
 FILLCELL_X32 FILLER_73_2687 ();
 FILLCELL_X32 FILLER_73_2719 ();
 FILLCELL_X32 FILLER_73_2751 ();
 FILLCELL_X32 FILLER_73_2783 ();
 FILLCELL_X32 FILLER_73_2815 ();
 FILLCELL_X32 FILLER_73_2847 ();
 FILLCELL_X32 FILLER_73_2879 ();
 FILLCELL_X32 FILLER_73_2911 ();
 FILLCELL_X32 FILLER_73_2943 ();
 FILLCELL_X32 FILLER_73_2975 ();
 FILLCELL_X32 FILLER_73_3007 ();
 FILLCELL_X32 FILLER_73_3039 ();
 FILLCELL_X32 FILLER_73_3071 ();
 FILLCELL_X32 FILLER_73_3103 ();
 FILLCELL_X32 FILLER_73_3135 ();
 FILLCELL_X32 FILLER_73_3167 ();
 FILLCELL_X32 FILLER_73_3199 ();
 FILLCELL_X32 FILLER_73_3231 ();
 FILLCELL_X32 FILLER_73_3263 ();
 FILLCELL_X32 FILLER_73_3295 ();
 FILLCELL_X32 FILLER_73_3327 ();
 FILLCELL_X32 FILLER_73_3359 ();
 FILLCELL_X32 FILLER_73_3391 ();
 FILLCELL_X32 FILLER_73_3423 ();
 FILLCELL_X32 FILLER_73_3455 ();
 FILLCELL_X32 FILLER_73_3487 ();
 FILLCELL_X32 FILLER_73_3519 ();
 FILLCELL_X32 FILLER_73_3551 ();
 FILLCELL_X32 FILLER_73_3583 ();
 FILLCELL_X32 FILLER_73_3615 ();
 FILLCELL_X32 FILLER_73_3647 ();
 FILLCELL_X32 FILLER_73_3679 ();
 FILLCELL_X16 FILLER_73_3711 ();
 FILLCELL_X8 FILLER_73_3727 ();
 FILLCELL_X2 FILLER_73_3735 ();
 FILLCELL_X1 FILLER_73_3737 ();
 FILLCELL_X32 FILLER_74_1 ();
 FILLCELL_X32 FILLER_74_33 ();
 FILLCELL_X32 FILLER_74_65 ();
 FILLCELL_X32 FILLER_74_97 ();
 FILLCELL_X32 FILLER_74_129 ();
 FILLCELL_X32 FILLER_74_161 ();
 FILLCELL_X32 FILLER_74_193 ();
 FILLCELL_X32 FILLER_74_225 ();
 FILLCELL_X32 FILLER_74_257 ();
 FILLCELL_X32 FILLER_74_289 ();
 FILLCELL_X32 FILLER_74_321 ();
 FILLCELL_X32 FILLER_74_353 ();
 FILLCELL_X32 FILLER_74_385 ();
 FILLCELL_X32 FILLER_74_417 ();
 FILLCELL_X32 FILLER_74_449 ();
 FILLCELL_X32 FILLER_74_481 ();
 FILLCELL_X32 FILLER_74_513 ();
 FILLCELL_X32 FILLER_74_545 ();
 FILLCELL_X32 FILLER_74_577 ();
 FILLCELL_X16 FILLER_74_609 ();
 FILLCELL_X4 FILLER_74_625 ();
 FILLCELL_X2 FILLER_74_629 ();
 FILLCELL_X32 FILLER_74_632 ();
 FILLCELL_X32 FILLER_74_664 ();
 FILLCELL_X32 FILLER_74_696 ();
 FILLCELL_X32 FILLER_74_728 ();
 FILLCELL_X32 FILLER_74_760 ();
 FILLCELL_X32 FILLER_74_792 ();
 FILLCELL_X32 FILLER_74_824 ();
 FILLCELL_X32 FILLER_74_856 ();
 FILLCELL_X32 FILLER_74_888 ();
 FILLCELL_X32 FILLER_74_920 ();
 FILLCELL_X32 FILLER_74_952 ();
 FILLCELL_X32 FILLER_74_984 ();
 FILLCELL_X32 FILLER_74_1016 ();
 FILLCELL_X32 FILLER_74_1048 ();
 FILLCELL_X32 FILLER_74_1080 ();
 FILLCELL_X32 FILLER_74_1112 ();
 FILLCELL_X32 FILLER_74_1144 ();
 FILLCELL_X32 FILLER_74_1176 ();
 FILLCELL_X32 FILLER_74_1208 ();
 FILLCELL_X32 FILLER_74_1240 ();
 FILLCELL_X32 FILLER_74_1272 ();
 FILLCELL_X32 FILLER_74_1304 ();
 FILLCELL_X32 FILLER_74_1336 ();
 FILLCELL_X32 FILLER_74_1368 ();
 FILLCELL_X32 FILLER_74_1400 ();
 FILLCELL_X32 FILLER_74_1432 ();
 FILLCELL_X32 FILLER_74_1464 ();
 FILLCELL_X32 FILLER_74_1496 ();
 FILLCELL_X32 FILLER_74_1528 ();
 FILLCELL_X32 FILLER_74_1560 ();
 FILLCELL_X32 FILLER_74_1592 ();
 FILLCELL_X32 FILLER_74_1624 ();
 FILLCELL_X32 FILLER_74_1656 ();
 FILLCELL_X32 FILLER_74_1688 ();
 FILLCELL_X32 FILLER_74_1720 ();
 FILLCELL_X32 FILLER_74_1752 ();
 FILLCELL_X32 FILLER_74_1784 ();
 FILLCELL_X32 FILLER_74_1816 ();
 FILLCELL_X32 FILLER_74_1848 ();
 FILLCELL_X8 FILLER_74_1880 ();
 FILLCELL_X4 FILLER_74_1888 ();
 FILLCELL_X2 FILLER_74_1892 ();
 FILLCELL_X32 FILLER_74_1895 ();
 FILLCELL_X32 FILLER_74_1927 ();
 FILLCELL_X32 FILLER_74_1959 ();
 FILLCELL_X32 FILLER_74_1991 ();
 FILLCELL_X32 FILLER_74_2023 ();
 FILLCELL_X32 FILLER_74_2055 ();
 FILLCELL_X32 FILLER_74_2087 ();
 FILLCELL_X32 FILLER_74_2119 ();
 FILLCELL_X32 FILLER_74_2151 ();
 FILLCELL_X32 FILLER_74_2183 ();
 FILLCELL_X32 FILLER_74_2215 ();
 FILLCELL_X32 FILLER_74_2247 ();
 FILLCELL_X32 FILLER_74_2279 ();
 FILLCELL_X32 FILLER_74_2311 ();
 FILLCELL_X32 FILLER_74_2343 ();
 FILLCELL_X32 FILLER_74_2375 ();
 FILLCELL_X32 FILLER_74_2407 ();
 FILLCELL_X32 FILLER_74_2439 ();
 FILLCELL_X32 FILLER_74_2471 ();
 FILLCELL_X32 FILLER_74_2503 ();
 FILLCELL_X32 FILLER_74_2535 ();
 FILLCELL_X32 FILLER_74_2567 ();
 FILLCELL_X32 FILLER_74_2599 ();
 FILLCELL_X32 FILLER_74_2631 ();
 FILLCELL_X32 FILLER_74_2663 ();
 FILLCELL_X32 FILLER_74_2695 ();
 FILLCELL_X32 FILLER_74_2727 ();
 FILLCELL_X32 FILLER_74_2759 ();
 FILLCELL_X32 FILLER_74_2791 ();
 FILLCELL_X32 FILLER_74_2823 ();
 FILLCELL_X32 FILLER_74_2855 ();
 FILLCELL_X32 FILLER_74_2887 ();
 FILLCELL_X32 FILLER_74_2919 ();
 FILLCELL_X32 FILLER_74_2951 ();
 FILLCELL_X32 FILLER_74_2983 ();
 FILLCELL_X32 FILLER_74_3015 ();
 FILLCELL_X32 FILLER_74_3047 ();
 FILLCELL_X32 FILLER_74_3079 ();
 FILLCELL_X32 FILLER_74_3111 ();
 FILLCELL_X8 FILLER_74_3143 ();
 FILLCELL_X4 FILLER_74_3151 ();
 FILLCELL_X2 FILLER_74_3155 ();
 FILLCELL_X32 FILLER_74_3158 ();
 FILLCELL_X32 FILLER_74_3190 ();
 FILLCELL_X32 FILLER_74_3222 ();
 FILLCELL_X32 FILLER_74_3254 ();
 FILLCELL_X32 FILLER_74_3286 ();
 FILLCELL_X32 FILLER_74_3318 ();
 FILLCELL_X32 FILLER_74_3350 ();
 FILLCELL_X32 FILLER_74_3382 ();
 FILLCELL_X32 FILLER_74_3414 ();
 FILLCELL_X32 FILLER_74_3446 ();
 FILLCELL_X32 FILLER_74_3478 ();
 FILLCELL_X32 FILLER_74_3510 ();
 FILLCELL_X32 FILLER_74_3542 ();
 FILLCELL_X32 FILLER_74_3574 ();
 FILLCELL_X32 FILLER_74_3606 ();
 FILLCELL_X32 FILLER_74_3638 ();
 FILLCELL_X32 FILLER_74_3670 ();
 FILLCELL_X32 FILLER_74_3702 ();
 FILLCELL_X4 FILLER_74_3734 ();
 FILLCELL_X32 FILLER_75_1 ();
 FILLCELL_X32 FILLER_75_33 ();
 FILLCELL_X32 FILLER_75_65 ();
 FILLCELL_X32 FILLER_75_97 ();
 FILLCELL_X32 FILLER_75_129 ();
 FILLCELL_X32 FILLER_75_161 ();
 FILLCELL_X32 FILLER_75_193 ();
 FILLCELL_X32 FILLER_75_225 ();
 FILLCELL_X32 FILLER_75_257 ();
 FILLCELL_X32 FILLER_75_289 ();
 FILLCELL_X32 FILLER_75_321 ();
 FILLCELL_X32 FILLER_75_353 ();
 FILLCELL_X32 FILLER_75_385 ();
 FILLCELL_X32 FILLER_75_417 ();
 FILLCELL_X32 FILLER_75_449 ();
 FILLCELL_X32 FILLER_75_481 ();
 FILLCELL_X32 FILLER_75_513 ();
 FILLCELL_X32 FILLER_75_545 ();
 FILLCELL_X32 FILLER_75_577 ();
 FILLCELL_X32 FILLER_75_609 ();
 FILLCELL_X32 FILLER_75_641 ();
 FILLCELL_X32 FILLER_75_673 ();
 FILLCELL_X32 FILLER_75_705 ();
 FILLCELL_X32 FILLER_75_737 ();
 FILLCELL_X32 FILLER_75_769 ();
 FILLCELL_X32 FILLER_75_801 ();
 FILLCELL_X32 FILLER_75_833 ();
 FILLCELL_X32 FILLER_75_865 ();
 FILLCELL_X32 FILLER_75_897 ();
 FILLCELL_X32 FILLER_75_929 ();
 FILLCELL_X32 FILLER_75_961 ();
 FILLCELL_X32 FILLER_75_993 ();
 FILLCELL_X32 FILLER_75_1025 ();
 FILLCELL_X32 FILLER_75_1057 ();
 FILLCELL_X32 FILLER_75_1089 ();
 FILLCELL_X32 FILLER_75_1121 ();
 FILLCELL_X32 FILLER_75_1153 ();
 FILLCELL_X32 FILLER_75_1185 ();
 FILLCELL_X32 FILLER_75_1217 ();
 FILLCELL_X8 FILLER_75_1249 ();
 FILLCELL_X4 FILLER_75_1257 ();
 FILLCELL_X2 FILLER_75_1261 ();
 FILLCELL_X32 FILLER_75_1264 ();
 FILLCELL_X32 FILLER_75_1296 ();
 FILLCELL_X32 FILLER_75_1328 ();
 FILLCELL_X32 FILLER_75_1360 ();
 FILLCELL_X32 FILLER_75_1392 ();
 FILLCELL_X32 FILLER_75_1424 ();
 FILLCELL_X32 FILLER_75_1456 ();
 FILLCELL_X32 FILLER_75_1488 ();
 FILLCELL_X32 FILLER_75_1520 ();
 FILLCELL_X32 FILLER_75_1552 ();
 FILLCELL_X32 FILLER_75_1584 ();
 FILLCELL_X32 FILLER_75_1616 ();
 FILLCELL_X32 FILLER_75_1648 ();
 FILLCELL_X32 FILLER_75_1680 ();
 FILLCELL_X32 FILLER_75_1712 ();
 FILLCELL_X32 FILLER_75_1744 ();
 FILLCELL_X32 FILLER_75_1776 ();
 FILLCELL_X32 FILLER_75_1808 ();
 FILLCELL_X32 FILLER_75_1840 ();
 FILLCELL_X32 FILLER_75_1872 ();
 FILLCELL_X32 FILLER_75_1904 ();
 FILLCELL_X32 FILLER_75_1936 ();
 FILLCELL_X32 FILLER_75_1968 ();
 FILLCELL_X32 FILLER_75_2000 ();
 FILLCELL_X32 FILLER_75_2032 ();
 FILLCELL_X32 FILLER_75_2064 ();
 FILLCELL_X32 FILLER_75_2096 ();
 FILLCELL_X32 FILLER_75_2128 ();
 FILLCELL_X32 FILLER_75_2160 ();
 FILLCELL_X32 FILLER_75_2192 ();
 FILLCELL_X32 FILLER_75_2224 ();
 FILLCELL_X32 FILLER_75_2256 ();
 FILLCELL_X32 FILLER_75_2288 ();
 FILLCELL_X32 FILLER_75_2320 ();
 FILLCELL_X32 FILLER_75_2352 ();
 FILLCELL_X32 FILLER_75_2384 ();
 FILLCELL_X32 FILLER_75_2416 ();
 FILLCELL_X32 FILLER_75_2448 ();
 FILLCELL_X32 FILLER_75_2480 ();
 FILLCELL_X8 FILLER_75_2512 ();
 FILLCELL_X4 FILLER_75_2520 ();
 FILLCELL_X2 FILLER_75_2524 ();
 FILLCELL_X32 FILLER_75_2527 ();
 FILLCELL_X32 FILLER_75_2559 ();
 FILLCELL_X32 FILLER_75_2591 ();
 FILLCELL_X32 FILLER_75_2623 ();
 FILLCELL_X32 FILLER_75_2655 ();
 FILLCELL_X32 FILLER_75_2687 ();
 FILLCELL_X32 FILLER_75_2719 ();
 FILLCELL_X32 FILLER_75_2751 ();
 FILLCELL_X32 FILLER_75_2783 ();
 FILLCELL_X32 FILLER_75_2815 ();
 FILLCELL_X32 FILLER_75_2847 ();
 FILLCELL_X32 FILLER_75_2879 ();
 FILLCELL_X32 FILLER_75_2911 ();
 FILLCELL_X32 FILLER_75_2943 ();
 FILLCELL_X32 FILLER_75_2975 ();
 FILLCELL_X32 FILLER_75_3007 ();
 FILLCELL_X32 FILLER_75_3039 ();
 FILLCELL_X32 FILLER_75_3071 ();
 FILLCELL_X32 FILLER_75_3103 ();
 FILLCELL_X32 FILLER_75_3135 ();
 FILLCELL_X32 FILLER_75_3167 ();
 FILLCELL_X32 FILLER_75_3199 ();
 FILLCELL_X32 FILLER_75_3231 ();
 FILLCELL_X32 FILLER_75_3263 ();
 FILLCELL_X32 FILLER_75_3295 ();
 FILLCELL_X32 FILLER_75_3327 ();
 FILLCELL_X32 FILLER_75_3359 ();
 FILLCELL_X32 FILLER_75_3391 ();
 FILLCELL_X32 FILLER_75_3423 ();
 FILLCELL_X32 FILLER_75_3455 ();
 FILLCELL_X32 FILLER_75_3487 ();
 FILLCELL_X32 FILLER_75_3519 ();
 FILLCELL_X32 FILLER_75_3551 ();
 FILLCELL_X32 FILLER_75_3583 ();
 FILLCELL_X32 FILLER_75_3615 ();
 FILLCELL_X32 FILLER_75_3647 ();
 FILLCELL_X32 FILLER_75_3679 ();
 FILLCELL_X16 FILLER_75_3711 ();
 FILLCELL_X8 FILLER_75_3727 ();
 FILLCELL_X2 FILLER_75_3735 ();
 FILLCELL_X1 FILLER_75_3737 ();
 FILLCELL_X32 FILLER_76_1 ();
 FILLCELL_X32 FILLER_76_33 ();
 FILLCELL_X32 FILLER_76_65 ();
 FILLCELL_X32 FILLER_76_97 ();
 FILLCELL_X32 FILLER_76_129 ();
 FILLCELL_X32 FILLER_76_161 ();
 FILLCELL_X32 FILLER_76_193 ();
 FILLCELL_X32 FILLER_76_225 ();
 FILLCELL_X32 FILLER_76_257 ();
 FILLCELL_X32 FILLER_76_289 ();
 FILLCELL_X32 FILLER_76_321 ();
 FILLCELL_X32 FILLER_76_353 ();
 FILLCELL_X32 FILLER_76_385 ();
 FILLCELL_X32 FILLER_76_417 ();
 FILLCELL_X32 FILLER_76_449 ();
 FILLCELL_X32 FILLER_76_481 ();
 FILLCELL_X32 FILLER_76_513 ();
 FILLCELL_X32 FILLER_76_545 ();
 FILLCELL_X32 FILLER_76_577 ();
 FILLCELL_X16 FILLER_76_609 ();
 FILLCELL_X4 FILLER_76_625 ();
 FILLCELL_X2 FILLER_76_629 ();
 FILLCELL_X32 FILLER_76_632 ();
 FILLCELL_X32 FILLER_76_664 ();
 FILLCELL_X32 FILLER_76_696 ();
 FILLCELL_X32 FILLER_76_728 ();
 FILLCELL_X32 FILLER_76_760 ();
 FILLCELL_X32 FILLER_76_792 ();
 FILLCELL_X32 FILLER_76_824 ();
 FILLCELL_X32 FILLER_76_856 ();
 FILLCELL_X32 FILLER_76_888 ();
 FILLCELL_X32 FILLER_76_920 ();
 FILLCELL_X32 FILLER_76_952 ();
 FILLCELL_X32 FILLER_76_984 ();
 FILLCELL_X32 FILLER_76_1016 ();
 FILLCELL_X32 FILLER_76_1048 ();
 FILLCELL_X32 FILLER_76_1080 ();
 FILLCELL_X32 FILLER_76_1112 ();
 FILLCELL_X32 FILLER_76_1144 ();
 FILLCELL_X32 FILLER_76_1176 ();
 FILLCELL_X32 FILLER_76_1208 ();
 FILLCELL_X32 FILLER_76_1240 ();
 FILLCELL_X32 FILLER_76_1272 ();
 FILLCELL_X32 FILLER_76_1304 ();
 FILLCELL_X32 FILLER_76_1336 ();
 FILLCELL_X32 FILLER_76_1368 ();
 FILLCELL_X32 FILLER_76_1400 ();
 FILLCELL_X32 FILLER_76_1432 ();
 FILLCELL_X32 FILLER_76_1464 ();
 FILLCELL_X32 FILLER_76_1496 ();
 FILLCELL_X32 FILLER_76_1528 ();
 FILLCELL_X32 FILLER_76_1560 ();
 FILLCELL_X32 FILLER_76_1592 ();
 FILLCELL_X32 FILLER_76_1624 ();
 FILLCELL_X32 FILLER_76_1656 ();
 FILLCELL_X32 FILLER_76_1688 ();
 FILLCELL_X32 FILLER_76_1720 ();
 FILLCELL_X32 FILLER_76_1752 ();
 FILLCELL_X32 FILLER_76_1784 ();
 FILLCELL_X32 FILLER_76_1816 ();
 FILLCELL_X32 FILLER_76_1848 ();
 FILLCELL_X8 FILLER_76_1880 ();
 FILLCELL_X4 FILLER_76_1888 ();
 FILLCELL_X2 FILLER_76_1892 ();
 FILLCELL_X32 FILLER_76_1895 ();
 FILLCELL_X32 FILLER_76_1927 ();
 FILLCELL_X32 FILLER_76_1959 ();
 FILLCELL_X32 FILLER_76_1991 ();
 FILLCELL_X32 FILLER_76_2023 ();
 FILLCELL_X32 FILLER_76_2055 ();
 FILLCELL_X32 FILLER_76_2087 ();
 FILLCELL_X32 FILLER_76_2119 ();
 FILLCELL_X32 FILLER_76_2151 ();
 FILLCELL_X32 FILLER_76_2183 ();
 FILLCELL_X32 FILLER_76_2215 ();
 FILLCELL_X32 FILLER_76_2247 ();
 FILLCELL_X32 FILLER_76_2279 ();
 FILLCELL_X32 FILLER_76_2311 ();
 FILLCELL_X32 FILLER_76_2343 ();
 FILLCELL_X32 FILLER_76_2375 ();
 FILLCELL_X32 FILLER_76_2407 ();
 FILLCELL_X32 FILLER_76_2439 ();
 FILLCELL_X32 FILLER_76_2471 ();
 FILLCELL_X32 FILLER_76_2503 ();
 FILLCELL_X32 FILLER_76_2535 ();
 FILLCELL_X32 FILLER_76_2567 ();
 FILLCELL_X32 FILLER_76_2599 ();
 FILLCELL_X32 FILLER_76_2631 ();
 FILLCELL_X32 FILLER_76_2663 ();
 FILLCELL_X32 FILLER_76_2695 ();
 FILLCELL_X32 FILLER_76_2727 ();
 FILLCELL_X32 FILLER_76_2759 ();
 FILLCELL_X32 FILLER_76_2791 ();
 FILLCELL_X32 FILLER_76_2823 ();
 FILLCELL_X32 FILLER_76_2855 ();
 FILLCELL_X32 FILLER_76_2887 ();
 FILLCELL_X32 FILLER_76_2919 ();
 FILLCELL_X32 FILLER_76_2951 ();
 FILLCELL_X32 FILLER_76_2983 ();
 FILLCELL_X32 FILLER_76_3015 ();
 FILLCELL_X32 FILLER_76_3047 ();
 FILLCELL_X32 FILLER_76_3079 ();
 FILLCELL_X32 FILLER_76_3111 ();
 FILLCELL_X8 FILLER_76_3143 ();
 FILLCELL_X4 FILLER_76_3151 ();
 FILLCELL_X2 FILLER_76_3155 ();
 FILLCELL_X32 FILLER_76_3158 ();
 FILLCELL_X32 FILLER_76_3190 ();
 FILLCELL_X32 FILLER_76_3222 ();
 FILLCELL_X32 FILLER_76_3254 ();
 FILLCELL_X32 FILLER_76_3286 ();
 FILLCELL_X32 FILLER_76_3318 ();
 FILLCELL_X32 FILLER_76_3350 ();
 FILLCELL_X32 FILLER_76_3382 ();
 FILLCELL_X32 FILLER_76_3414 ();
 FILLCELL_X32 FILLER_76_3446 ();
 FILLCELL_X32 FILLER_76_3478 ();
 FILLCELL_X32 FILLER_76_3510 ();
 FILLCELL_X32 FILLER_76_3542 ();
 FILLCELL_X32 FILLER_76_3574 ();
 FILLCELL_X32 FILLER_76_3606 ();
 FILLCELL_X32 FILLER_76_3638 ();
 FILLCELL_X32 FILLER_76_3670 ();
 FILLCELL_X32 FILLER_76_3702 ();
 FILLCELL_X4 FILLER_76_3734 ();
 FILLCELL_X32 FILLER_77_1 ();
 FILLCELL_X32 FILLER_77_33 ();
 FILLCELL_X32 FILLER_77_65 ();
 FILLCELL_X32 FILLER_77_97 ();
 FILLCELL_X32 FILLER_77_129 ();
 FILLCELL_X32 FILLER_77_161 ();
 FILLCELL_X32 FILLER_77_193 ();
 FILLCELL_X32 FILLER_77_225 ();
 FILLCELL_X32 FILLER_77_257 ();
 FILLCELL_X32 FILLER_77_289 ();
 FILLCELL_X32 FILLER_77_321 ();
 FILLCELL_X32 FILLER_77_353 ();
 FILLCELL_X32 FILLER_77_385 ();
 FILLCELL_X32 FILLER_77_417 ();
 FILLCELL_X32 FILLER_77_449 ();
 FILLCELL_X32 FILLER_77_481 ();
 FILLCELL_X32 FILLER_77_513 ();
 FILLCELL_X32 FILLER_77_545 ();
 FILLCELL_X32 FILLER_77_577 ();
 FILLCELL_X32 FILLER_77_609 ();
 FILLCELL_X32 FILLER_77_641 ();
 FILLCELL_X32 FILLER_77_673 ();
 FILLCELL_X32 FILLER_77_705 ();
 FILLCELL_X32 FILLER_77_737 ();
 FILLCELL_X32 FILLER_77_769 ();
 FILLCELL_X32 FILLER_77_801 ();
 FILLCELL_X32 FILLER_77_833 ();
 FILLCELL_X32 FILLER_77_865 ();
 FILLCELL_X32 FILLER_77_897 ();
 FILLCELL_X32 FILLER_77_929 ();
 FILLCELL_X32 FILLER_77_961 ();
 FILLCELL_X32 FILLER_77_993 ();
 FILLCELL_X32 FILLER_77_1025 ();
 FILLCELL_X32 FILLER_77_1057 ();
 FILLCELL_X32 FILLER_77_1089 ();
 FILLCELL_X32 FILLER_77_1121 ();
 FILLCELL_X32 FILLER_77_1153 ();
 FILLCELL_X32 FILLER_77_1185 ();
 FILLCELL_X32 FILLER_77_1217 ();
 FILLCELL_X8 FILLER_77_1249 ();
 FILLCELL_X4 FILLER_77_1257 ();
 FILLCELL_X2 FILLER_77_1261 ();
 FILLCELL_X32 FILLER_77_1264 ();
 FILLCELL_X32 FILLER_77_1296 ();
 FILLCELL_X32 FILLER_77_1328 ();
 FILLCELL_X32 FILLER_77_1360 ();
 FILLCELL_X32 FILLER_77_1392 ();
 FILLCELL_X32 FILLER_77_1424 ();
 FILLCELL_X32 FILLER_77_1456 ();
 FILLCELL_X32 FILLER_77_1488 ();
 FILLCELL_X32 FILLER_77_1520 ();
 FILLCELL_X32 FILLER_77_1552 ();
 FILLCELL_X32 FILLER_77_1584 ();
 FILLCELL_X32 FILLER_77_1616 ();
 FILLCELL_X32 FILLER_77_1648 ();
 FILLCELL_X32 FILLER_77_1680 ();
 FILLCELL_X32 FILLER_77_1712 ();
 FILLCELL_X32 FILLER_77_1744 ();
 FILLCELL_X32 FILLER_77_1776 ();
 FILLCELL_X32 FILLER_77_1808 ();
 FILLCELL_X32 FILLER_77_1840 ();
 FILLCELL_X32 FILLER_77_1872 ();
 FILLCELL_X32 FILLER_77_1904 ();
 FILLCELL_X32 FILLER_77_1936 ();
 FILLCELL_X32 FILLER_77_1968 ();
 FILLCELL_X32 FILLER_77_2000 ();
 FILLCELL_X32 FILLER_77_2032 ();
 FILLCELL_X32 FILLER_77_2064 ();
 FILLCELL_X32 FILLER_77_2096 ();
 FILLCELL_X32 FILLER_77_2128 ();
 FILLCELL_X32 FILLER_77_2160 ();
 FILLCELL_X32 FILLER_77_2192 ();
 FILLCELL_X32 FILLER_77_2224 ();
 FILLCELL_X32 FILLER_77_2256 ();
 FILLCELL_X32 FILLER_77_2288 ();
 FILLCELL_X32 FILLER_77_2320 ();
 FILLCELL_X32 FILLER_77_2352 ();
 FILLCELL_X32 FILLER_77_2384 ();
 FILLCELL_X32 FILLER_77_2416 ();
 FILLCELL_X32 FILLER_77_2448 ();
 FILLCELL_X32 FILLER_77_2480 ();
 FILLCELL_X8 FILLER_77_2512 ();
 FILLCELL_X4 FILLER_77_2520 ();
 FILLCELL_X2 FILLER_77_2524 ();
 FILLCELL_X32 FILLER_77_2527 ();
 FILLCELL_X32 FILLER_77_2559 ();
 FILLCELL_X32 FILLER_77_2591 ();
 FILLCELL_X32 FILLER_77_2623 ();
 FILLCELL_X32 FILLER_77_2655 ();
 FILLCELL_X32 FILLER_77_2687 ();
 FILLCELL_X32 FILLER_77_2719 ();
 FILLCELL_X32 FILLER_77_2751 ();
 FILLCELL_X32 FILLER_77_2783 ();
 FILLCELL_X32 FILLER_77_2815 ();
 FILLCELL_X32 FILLER_77_2847 ();
 FILLCELL_X32 FILLER_77_2879 ();
 FILLCELL_X32 FILLER_77_2911 ();
 FILLCELL_X32 FILLER_77_2943 ();
 FILLCELL_X32 FILLER_77_2975 ();
 FILLCELL_X32 FILLER_77_3007 ();
 FILLCELL_X32 FILLER_77_3039 ();
 FILLCELL_X32 FILLER_77_3071 ();
 FILLCELL_X32 FILLER_77_3103 ();
 FILLCELL_X32 FILLER_77_3135 ();
 FILLCELL_X32 FILLER_77_3167 ();
 FILLCELL_X32 FILLER_77_3199 ();
 FILLCELL_X32 FILLER_77_3231 ();
 FILLCELL_X32 FILLER_77_3263 ();
 FILLCELL_X32 FILLER_77_3295 ();
 FILLCELL_X32 FILLER_77_3327 ();
 FILLCELL_X32 FILLER_77_3359 ();
 FILLCELL_X32 FILLER_77_3391 ();
 FILLCELL_X32 FILLER_77_3423 ();
 FILLCELL_X32 FILLER_77_3455 ();
 FILLCELL_X32 FILLER_77_3487 ();
 FILLCELL_X32 FILLER_77_3519 ();
 FILLCELL_X32 FILLER_77_3551 ();
 FILLCELL_X32 FILLER_77_3583 ();
 FILLCELL_X32 FILLER_77_3615 ();
 FILLCELL_X32 FILLER_77_3647 ();
 FILLCELL_X32 FILLER_77_3679 ();
 FILLCELL_X16 FILLER_77_3711 ();
 FILLCELL_X8 FILLER_77_3727 ();
 FILLCELL_X2 FILLER_77_3735 ();
 FILLCELL_X1 FILLER_77_3737 ();
 FILLCELL_X32 FILLER_78_1 ();
 FILLCELL_X32 FILLER_78_33 ();
 FILLCELL_X32 FILLER_78_65 ();
 FILLCELL_X32 FILLER_78_97 ();
 FILLCELL_X32 FILLER_78_129 ();
 FILLCELL_X32 FILLER_78_161 ();
 FILLCELL_X32 FILLER_78_193 ();
 FILLCELL_X32 FILLER_78_225 ();
 FILLCELL_X32 FILLER_78_257 ();
 FILLCELL_X32 FILLER_78_289 ();
 FILLCELL_X32 FILLER_78_321 ();
 FILLCELL_X32 FILLER_78_353 ();
 FILLCELL_X32 FILLER_78_385 ();
 FILLCELL_X32 FILLER_78_417 ();
 FILLCELL_X32 FILLER_78_449 ();
 FILLCELL_X32 FILLER_78_481 ();
 FILLCELL_X32 FILLER_78_513 ();
 FILLCELL_X32 FILLER_78_545 ();
 FILLCELL_X32 FILLER_78_577 ();
 FILLCELL_X16 FILLER_78_609 ();
 FILLCELL_X4 FILLER_78_625 ();
 FILLCELL_X2 FILLER_78_629 ();
 FILLCELL_X32 FILLER_78_632 ();
 FILLCELL_X32 FILLER_78_664 ();
 FILLCELL_X32 FILLER_78_696 ();
 FILLCELL_X32 FILLER_78_728 ();
 FILLCELL_X32 FILLER_78_760 ();
 FILLCELL_X32 FILLER_78_792 ();
 FILLCELL_X32 FILLER_78_824 ();
 FILLCELL_X32 FILLER_78_856 ();
 FILLCELL_X32 FILLER_78_888 ();
 FILLCELL_X32 FILLER_78_920 ();
 FILLCELL_X32 FILLER_78_952 ();
 FILLCELL_X32 FILLER_78_984 ();
 FILLCELL_X32 FILLER_78_1016 ();
 FILLCELL_X32 FILLER_78_1048 ();
 FILLCELL_X32 FILLER_78_1080 ();
 FILLCELL_X32 FILLER_78_1112 ();
 FILLCELL_X32 FILLER_78_1144 ();
 FILLCELL_X32 FILLER_78_1176 ();
 FILLCELL_X32 FILLER_78_1208 ();
 FILLCELL_X32 FILLER_78_1240 ();
 FILLCELL_X32 FILLER_78_1272 ();
 FILLCELL_X32 FILLER_78_1304 ();
 FILLCELL_X32 FILLER_78_1336 ();
 FILLCELL_X32 FILLER_78_1368 ();
 FILLCELL_X32 FILLER_78_1400 ();
 FILLCELL_X32 FILLER_78_1432 ();
 FILLCELL_X32 FILLER_78_1464 ();
 FILLCELL_X32 FILLER_78_1496 ();
 FILLCELL_X32 FILLER_78_1528 ();
 FILLCELL_X32 FILLER_78_1560 ();
 FILLCELL_X32 FILLER_78_1592 ();
 FILLCELL_X32 FILLER_78_1624 ();
 FILLCELL_X32 FILLER_78_1656 ();
 FILLCELL_X32 FILLER_78_1688 ();
 FILLCELL_X32 FILLER_78_1720 ();
 FILLCELL_X32 FILLER_78_1752 ();
 FILLCELL_X32 FILLER_78_1784 ();
 FILLCELL_X32 FILLER_78_1816 ();
 FILLCELL_X32 FILLER_78_1848 ();
 FILLCELL_X8 FILLER_78_1880 ();
 FILLCELL_X4 FILLER_78_1888 ();
 FILLCELL_X2 FILLER_78_1892 ();
 FILLCELL_X32 FILLER_78_1895 ();
 FILLCELL_X32 FILLER_78_1927 ();
 FILLCELL_X32 FILLER_78_1959 ();
 FILLCELL_X32 FILLER_78_1991 ();
 FILLCELL_X32 FILLER_78_2023 ();
 FILLCELL_X32 FILLER_78_2055 ();
 FILLCELL_X32 FILLER_78_2087 ();
 FILLCELL_X32 FILLER_78_2119 ();
 FILLCELL_X32 FILLER_78_2151 ();
 FILLCELL_X32 FILLER_78_2183 ();
 FILLCELL_X32 FILLER_78_2215 ();
 FILLCELL_X32 FILLER_78_2247 ();
 FILLCELL_X32 FILLER_78_2279 ();
 FILLCELL_X32 FILLER_78_2311 ();
 FILLCELL_X32 FILLER_78_2343 ();
 FILLCELL_X32 FILLER_78_2375 ();
 FILLCELL_X32 FILLER_78_2407 ();
 FILLCELL_X32 FILLER_78_2439 ();
 FILLCELL_X32 FILLER_78_2471 ();
 FILLCELL_X32 FILLER_78_2503 ();
 FILLCELL_X32 FILLER_78_2535 ();
 FILLCELL_X32 FILLER_78_2567 ();
 FILLCELL_X32 FILLER_78_2599 ();
 FILLCELL_X32 FILLER_78_2631 ();
 FILLCELL_X32 FILLER_78_2663 ();
 FILLCELL_X32 FILLER_78_2695 ();
 FILLCELL_X32 FILLER_78_2727 ();
 FILLCELL_X32 FILLER_78_2759 ();
 FILLCELL_X32 FILLER_78_2791 ();
 FILLCELL_X32 FILLER_78_2823 ();
 FILLCELL_X32 FILLER_78_2855 ();
 FILLCELL_X32 FILLER_78_2887 ();
 FILLCELL_X32 FILLER_78_2919 ();
 FILLCELL_X32 FILLER_78_2951 ();
 FILLCELL_X32 FILLER_78_2983 ();
 FILLCELL_X32 FILLER_78_3015 ();
 FILLCELL_X32 FILLER_78_3047 ();
 FILLCELL_X32 FILLER_78_3079 ();
 FILLCELL_X32 FILLER_78_3111 ();
 FILLCELL_X8 FILLER_78_3143 ();
 FILLCELL_X4 FILLER_78_3151 ();
 FILLCELL_X2 FILLER_78_3155 ();
 FILLCELL_X32 FILLER_78_3158 ();
 FILLCELL_X32 FILLER_78_3190 ();
 FILLCELL_X32 FILLER_78_3222 ();
 FILLCELL_X32 FILLER_78_3254 ();
 FILLCELL_X32 FILLER_78_3286 ();
 FILLCELL_X32 FILLER_78_3318 ();
 FILLCELL_X32 FILLER_78_3350 ();
 FILLCELL_X32 FILLER_78_3382 ();
 FILLCELL_X32 FILLER_78_3414 ();
 FILLCELL_X32 FILLER_78_3446 ();
 FILLCELL_X32 FILLER_78_3478 ();
 FILLCELL_X32 FILLER_78_3510 ();
 FILLCELL_X32 FILLER_78_3542 ();
 FILLCELL_X32 FILLER_78_3574 ();
 FILLCELL_X32 FILLER_78_3606 ();
 FILLCELL_X32 FILLER_78_3638 ();
 FILLCELL_X32 FILLER_78_3670 ();
 FILLCELL_X32 FILLER_78_3702 ();
 FILLCELL_X4 FILLER_78_3734 ();
 FILLCELL_X32 FILLER_79_1 ();
 FILLCELL_X32 FILLER_79_33 ();
 FILLCELL_X32 FILLER_79_65 ();
 FILLCELL_X32 FILLER_79_97 ();
 FILLCELL_X32 FILLER_79_129 ();
 FILLCELL_X32 FILLER_79_161 ();
 FILLCELL_X32 FILLER_79_193 ();
 FILLCELL_X32 FILLER_79_225 ();
 FILLCELL_X32 FILLER_79_257 ();
 FILLCELL_X32 FILLER_79_289 ();
 FILLCELL_X32 FILLER_79_321 ();
 FILLCELL_X32 FILLER_79_353 ();
 FILLCELL_X32 FILLER_79_385 ();
 FILLCELL_X32 FILLER_79_417 ();
 FILLCELL_X32 FILLER_79_449 ();
 FILLCELL_X32 FILLER_79_481 ();
 FILLCELL_X32 FILLER_79_513 ();
 FILLCELL_X32 FILLER_79_545 ();
 FILLCELL_X32 FILLER_79_577 ();
 FILLCELL_X32 FILLER_79_609 ();
 FILLCELL_X32 FILLER_79_641 ();
 FILLCELL_X32 FILLER_79_673 ();
 FILLCELL_X32 FILLER_79_705 ();
 FILLCELL_X32 FILLER_79_737 ();
 FILLCELL_X32 FILLER_79_769 ();
 FILLCELL_X32 FILLER_79_801 ();
 FILLCELL_X32 FILLER_79_833 ();
 FILLCELL_X32 FILLER_79_865 ();
 FILLCELL_X32 FILLER_79_897 ();
 FILLCELL_X32 FILLER_79_929 ();
 FILLCELL_X32 FILLER_79_961 ();
 FILLCELL_X32 FILLER_79_993 ();
 FILLCELL_X32 FILLER_79_1025 ();
 FILLCELL_X32 FILLER_79_1057 ();
 FILLCELL_X32 FILLER_79_1089 ();
 FILLCELL_X32 FILLER_79_1121 ();
 FILLCELL_X32 FILLER_79_1153 ();
 FILLCELL_X32 FILLER_79_1185 ();
 FILLCELL_X32 FILLER_79_1217 ();
 FILLCELL_X8 FILLER_79_1249 ();
 FILLCELL_X4 FILLER_79_1257 ();
 FILLCELL_X2 FILLER_79_1261 ();
 FILLCELL_X32 FILLER_79_1264 ();
 FILLCELL_X32 FILLER_79_1296 ();
 FILLCELL_X32 FILLER_79_1328 ();
 FILLCELL_X32 FILLER_79_1360 ();
 FILLCELL_X32 FILLER_79_1392 ();
 FILLCELL_X32 FILLER_79_1424 ();
 FILLCELL_X32 FILLER_79_1456 ();
 FILLCELL_X32 FILLER_79_1488 ();
 FILLCELL_X32 FILLER_79_1520 ();
 FILLCELL_X32 FILLER_79_1552 ();
 FILLCELL_X32 FILLER_79_1584 ();
 FILLCELL_X32 FILLER_79_1616 ();
 FILLCELL_X32 FILLER_79_1648 ();
 FILLCELL_X32 FILLER_79_1680 ();
 FILLCELL_X32 FILLER_79_1712 ();
 FILLCELL_X32 FILLER_79_1744 ();
 FILLCELL_X32 FILLER_79_1776 ();
 FILLCELL_X32 FILLER_79_1808 ();
 FILLCELL_X32 FILLER_79_1840 ();
 FILLCELL_X32 FILLER_79_1872 ();
 FILLCELL_X32 FILLER_79_1904 ();
 FILLCELL_X32 FILLER_79_1936 ();
 FILLCELL_X32 FILLER_79_1968 ();
 FILLCELL_X32 FILLER_79_2000 ();
 FILLCELL_X32 FILLER_79_2032 ();
 FILLCELL_X32 FILLER_79_2064 ();
 FILLCELL_X32 FILLER_79_2096 ();
 FILLCELL_X32 FILLER_79_2128 ();
 FILLCELL_X32 FILLER_79_2160 ();
 FILLCELL_X32 FILLER_79_2192 ();
 FILLCELL_X32 FILLER_79_2224 ();
 FILLCELL_X32 FILLER_79_2256 ();
 FILLCELL_X32 FILLER_79_2288 ();
 FILLCELL_X32 FILLER_79_2320 ();
 FILLCELL_X32 FILLER_79_2352 ();
 FILLCELL_X32 FILLER_79_2384 ();
 FILLCELL_X32 FILLER_79_2416 ();
 FILLCELL_X32 FILLER_79_2448 ();
 FILLCELL_X32 FILLER_79_2480 ();
 FILLCELL_X8 FILLER_79_2512 ();
 FILLCELL_X4 FILLER_79_2520 ();
 FILLCELL_X2 FILLER_79_2524 ();
 FILLCELL_X32 FILLER_79_2527 ();
 FILLCELL_X32 FILLER_79_2559 ();
 FILLCELL_X32 FILLER_79_2591 ();
 FILLCELL_X32 FILLER_79_2623 ();
 FILLCELL_X32 FILLER_79_2655 ();
 FILLCELL_X32 FILLER_79_2687 ();
 FILLCELL_X32 FILLER_79_2719 ();
 FILLCELL_X32 FILLER_79_2751 ();
 FILLCELL_X32 FILLER_79_2783 ();
 FILLCELL_X32 FILLER_79_2815 ();
 FILLCELL_X32 FILLER_79_2847 ();
 FILLCELL_X32 FILLER_79_2879 ();
 FILLCELL_X32 FILLER_79_2911 ();
 FILLCELL_X32 FILLER_79_2943 ();
 FILLCELL_X32 FILLER_79_2975 ();
 FILLCELL_X32 FILLER_79_3007 ();
 FILLCELL_X32 FILLER_79_3039 ();
 FILLCELL_X32 FILLER_79_3071 ();
 FILLCELL_X32 FILLER_79_3103 ();
 FILLCELL_X32 FILLER_79_3135 ();
 FILLCELL_X32 FILLER_79_3167 ();
 FILLCELL_X32 FILLER_79_3199 ();
 FILLCELL_X32 FILLER_79_3231 ();
 FILLCELL_X32 FILLER_79_3263 ();
 FILLCELL_X32 FILLER_79_3295 ();
 FILLCELL_X32 FILLER_79_3327 ();
 FILLCELL_X32 FILLER_79_3359 ();
 FILLCELL_X32 FILLER_79_3391 ();
 FILLCELL_X32 FILLER_79_3423 ();
 FILLCELL_X32 FILLER_79_3455 ();
 FILLCELL_X32 FILLER_79_3487 ();
 FILLCELL_X32 FILLER_79_3519 ();
 FILLCELL_X32 FILLER_79_3551 ();
 FILLCELL_X32 FILLER_79_3583 ();
 FILLCELL_X32 FILLER_79_3615 ();
 FILLCELL_X32 FILLER_79_3647 ();
 FILLCELL_X32 FILLER_79_3679 ();
 FILLCELL_X16 FILLER_79_3711 ();
 FILLCELL_X8 FILLER_79_3727 ();
 FILLCELL_X2 FILLER_79_3735 ();
 FILLCELL_X1 FILLER_79_3737 ();
 FILLCELL_X32 FILLER_80_1 ();
 FILLCELL_X32 FILLER_80_33 ();
 FILLCELL_X32 FILLER_80_65 ();
 FILLCELL_X32 FILLER_80_97 ();
 FILLCELL_X32 FILLER_80_129 ();
 FILLCELL_X32 FILLER_80_161 ();
 FILLCELL_X32 FILLER_80_193 ();
 FILLCELL_X32 FILLER_80_225 ();
 FILLCELL_X32 FILLER_80_257 ();
 FILLCELL_X32 FILLER_80_289 ();
 FILLCELL_X32 FILLER_80_321 ();
 FILLCELL_X32 FILLER_80_353 ();
 FILLCELL_X32 FILLER_80_385 ();
 FILLCELL_X32 FILLER_80_417 ();
 FILLCELL_X32 FILLER_80_449 ();
 FILLCELL_X32 FILLER_80_481 ();
 FILLCELL_X32 FILLER_80_513 ();
 FILLCELL_X32 FILLER_80_545 ();
 FILLCELL_X32 FILLER_80_577 ();
 FILLCELL_X16 FILLER_80_609 ();
 FILLCELL_X4 FILLER_80_625 ();
 FILLCELL_X2 FILLER_80_629 ();
 FILLCELL_X32 FILLER_80_632 ();
 FILLCELL_X32 FILLER_80_664 ();
 FILLCELL_X32 FILLER_80_696 ();
 FILLCELL_X32 FILLER_80_728 ();
 FILLCELL_X32 FILLER_80_760 ();
 FILLCELL_X32 FILLER_80_792 ();
 FILLCELL_X32 FILLER_80_824 ();
 FILLCELL_X32 FILLER_80_856 ();
 FILLCELL_X32 FILLER_80_888 ();
 FILLCELL_X32 FILLER_80_920 ();
 FILLCELL_X32 FILLER_80_952 ();
 FILLCELL_X32 FILLER_80_984 ();
 FILLCELL_X32 FILLER_80_1016 ();
 FILLCELL_X32 FILLER_80_1048 ();
 FILLCELL_X32 FILLER_80_1080 ();
 FILLCELL_X32 FILLER_80_1112 ();
 FILLCELL_X32 FILLER_80_1144 ();
 FILLCELL_X32 FILLER_80_1176 ();
 FILLCELL_X32 FILLER_80_1208 ();
 FILLCELL_X32 FILLER_80_1240 ();
 FILLCELL_X32 FILLER_80_1272 ();
 FILLCELL_X32 FILLER_80_1304 ();
 FILLCELL_X32 FILLER_80_1336 ();
 FILLCELL_X32 FILLER_80_1368 ();
 FILLCELL_X32 FILLER_80_1400 ();
 FILLCELL_X32 FILLER_80_1432 ();
 FILLCELL_X32 FILLER_80_1464 ();
 FILLCELL_X32 FILLER_80_1496 ();
 FILLCELL_X32 FILLER_80_1528 ();
 FILLCELL_X32 FILLER_80_1560 ();
 FILLCELL_X32 FILLER_80_1592 ();
 FILLCELL_X32 FILLER_80_1624 ();
 FILLCELL_X32 FILLER_80_1656 ();
 FILLCELL_X32 FILLER_80_1688 ();
 FILLCELL_X32 FILLER_80_1720 ();
 FILLCELL_X32 FILLER_80_1752 ();
 FILLCELL_X32 FILLER_80_1784 ();
 FILLCELL_X32 FILLER_80_1816 ();
 FILLCELL_X32 FILLER_80_1848 ();
 FILLCELL_X8 FILLER_80_1880 ();
 FILLCELL_X4 FILLER_80_1888 ();
 FILLCELL_X2 FILLER_80_1892 ();
 FILLCELL_X32 FILLER_80_1895 ();
 FILLCELL_X32 FILLER_80_1927 ();
 FILLCELL_X32 FILLER_80_1959 ();
 FILLCELL_X32 FILLER_80_1991 ();
 FILLCELL_X32 FILLER_80_2023 ();
 FILLCELL_X32 FILLER_80_2055 ();
 FILLCELL_X32 FILLER_80_2087 ();
 FILLCELL_X32 FILLER_80_2119 ();
 FILLCELL_X32 FILLER_80_2151 ();
 FILLCELL_X32 FILLER_80_2183 ();
 FILLCELL_X32 FILLER_80_2215 ();
 FILLCELL_X32 FILLER_80_2247 ();
 FILLCELL_X32 FILLER_80_2279 ();
 FILLCELL_X32 FILLER_80_2311 ();
 FILLCELL_X32 FILLER_80_2343 ();
 FILLCELL_X32 FILLER_80_2375 ();
 FILLCELL_X32 FILLER_80_2407 ();
 FILLCELL_X32 FILLER_80_2439 ();
 FILLCELL_X32 FILLER_80_2471 ();
 FILLCELL_X32 FILLER_80_2503 ();
 FILLCELL_X32 FILLER_80_2535 ();
 FILLCELL_X32 FILLER_80_2567 ();
 FILLCELL_X32 FILLER_80_2599 ();
 FILLCELL_X32 FILLER_80_2631 ();
 FILLCELL_X32 FILLER_80_2663 ();
 FILLCELL_X32 FILLER_80_2695 ();
 FILLCELL_X32 FILLER_80_2727 ();
 FILLCELL_X32 FILLER_80_2759 ();
 FILLCELL_X32 FILLER_80_2791 ();
 FILLCELL_X32 FILLER_80_2823 ();
 FILLCELL_X32 FILLER_80_2855 ();
 FILLCELL_X32 FILLER_80_2887 ();
 FILLCELL_X32 FILLER_80_2919 ();
 FILLCELL_X32 FILLER_80_2951 ();
 FILLCELL_X32 FILLER_80_2983 ();
 FILLCELL_X32 FILLER_80_3015 ();
 FILLCELL_X32 FILLER_80_3047 ();
 FILLCELL_X32 FILLER_80_3079 ();
 FILLCELL_X32 FILLER_80_3111 ();
 FILLCELL_X8 FILLER_80_3143 ();
 FILLCELL_X4 FILLER_80_3151 ();
 FILLCELL_X2 FILLER_80_3155 ();
 FILLCELL_X32 FILLER_80_3158 ();
 FILLCELL_X32 FILLER_80_3190 ();
 FILLCELL_X32 FILLER_80_3222 ();
 FILLCELL_X32 FILLER_80_3254 ();
 FILLCELL_X32 FILLER_80_3286 ();
 FILLCELL_X32 FILLER_80_3318 ();
 FILLCELL_X32 FILLER_80_3350 ();
 FILLCELL_X32 FILLER_80_3382 ();
 FILLCELL_X32 FILLER_80_3414 ();
 FILLCELL_X32 FILLER_80_3446 ();
 FILLCELL_X32 FILLER_80_3478 ();
 FILLCELL_X32 FILLER_80_3510 ();
 FILLCELL_X32 FILLER_80_3542 ();
 FILLCELL_X32 FILLER_80_3574 ();
 FILLCELL_X32 FILLER_80_3606 ();
 FILLCELL_X32 FILLER_80_3638 ();
 FILLCELL_X32 FILLER_80_3670 ();
 FILLCELL_X32 FILLER_80_3702 ();
 FILLCELL_X4 FILLER_80_3734 ();
 FILLCELL_X32 FILLER_81_1 ();
 FILLCELL_X32 FILLER_81_33 ();
 FILLCELL_X32 FILLER_81_65 ();
 FILLCELL_X32 FILLER_81_97 ();
 FILLCELL_X32 FILLER_81_129 ();
 FILLCELL_X32 FILLER_81_161 ();
 FILLCELL_X32 FILLER_81_193 ();
 FILLCELL_X32 FILLER_81_225 ();
 FILLCELL_X32 FILLER_81_257 ();
 FILLCELL_X32 FILLER_81_289 ();
 FILLCELL_X32 FILLER_81_321 ();
 FILLCELL_X32 FILLER_81_353 ();
 FILLCELL_X32 FILLER_81_385 ();
 FILLCELL_X32 FILLER_81_417 ();
 FILLCELL_X32 FILLER_81_449 ();
 FILLCELL_X32 FILLER_81_481 ();
 FILLCELL_X32 FILLER_81_513 ();
 FILLCELL_X32 FILLER_81_545 ();
 FILLCELL_X32 FILLER_81_577 ();
 FILLCELL_X32 FILLER_81_609 ();
 FILLCELL_X32 FILLER_81_641 ();
 FILLCELL_X32 FILLER_81_673 ();
 FILLCELL_X32 FILLER_81_705 ();
 FILLCELL_X32 FILLER_81_737 ();
 FILLCELL_X32 FILLER_81_769 ();
 FILLCELL_X32 FILLER_81_801 ();
 FILLCELL_X32 FILLER_81_833 ();
 FILLCELL_X32 FILLER_81_865 ();
 FILLCELL_X32 FILLER_81_897 ();
 FILLCELL_X32 FILLER_81_929 ();
 FILLCELL_X32 FILLER_81_961 ();
 FILLCELL_X32 FILLER_81_993 ();
 FILLCELL_X32 FILLER_81_1025 ();
 FILLCELL_X32 FILLER_81_1057 ();
 FILLCELL_X32 FILLER_81_1089 ();
 FILLCELL_X32 FILLER_81_1121 ();
 FILLCELL_X32 FILLER_81_1153 ();
 FILLCELL_X32 FILLER_81_1185 ();
 FILLCELL_X32 FILLER_81_1217 ();
 FILLCELL_X8 FILLER_81_1249 ();
 FILLCELL_X4 FILLER_81_1257 ();
 FILLCELL_X2 FILLER_81_1261 ();
 FILLCELL_X32 FILLER_81_1264 ();
 FILLCELL_X32 FILLER_81_1296 ();
 FILLCELL_X32 FILLER_81_1328 ();
 FILLCELL_X32 FILLER_81_1360 ();
 FILLCELL_X32 FILLER_81_1392 ();
 FILLCELL_X32 FILLER_81_1424 ();
 FILLCELL_X32 FILLER_81_1456 ();
 FILLCELL_X32 FILLER_81_1488 ();
 FILLCELL_X32 FILLER_81_1520 ();
 FILLCELL_X32 FILLER_81_1552 ();
 FILLCELL_X32 FILLER_81_1584 ();
 FILLCELL_X32 FILLER_81_1616 ();
 FILLCELL_X32 FILLER_81_1648 ();
 FILLCELL_X32 FILLER_81_1680 ();
 FILLCELL_X32 FILLER_81_1712 ();
 FILLCELL_X32 FILLER_81_1744 ();
 FILLCELL_X32 FILLER_81_1776 ();
 FILLCELL_X32 FILLER_81_1808 ();
 FILLCELL_X32 FILLER_81_1840 ();
 FILLCELL_X32 FILLER_81_1872 ();
 FILLCELL_X32 FILLER_81_1904 ();
 FILLCELL_X32 FILLER_81_1936 ();
 FILLCELL_X32 FILLER_81_1968 ();
 FILLCELL_X32 FILLER_81_2000 ();
 FILLCELL_X32 FILLER_81_2032 ();
 FILLCELL_X32 FILLER_81_2064 ();
 FILLCELL_X32 FILLER_81_2096 ();
 FILLCELL_X32 FILLER_81_2128 ();
 FILLCELL_X32 FILLER_81_2160 ();
 FILLCELL_X32 FILLER_81_2192 ();
 FILLCELL_X32 FILLER_81_2224 ();
 FILLCELL_X32 FILLER_81_2256 ();
 FILLCELL_X32 FILLER_81_2288 ();
 FILLCELL_X32 FILLER_81_2320 ();
 FILLCELL_X32 FILLER_81_2352 ();
 FILLCELL_X32 FILLER_81_2384 ();
 FILLCELL_X32 FILLER_81_2416 ();
 FILLCELL_X32 FILLER_81_2448 ();
 FILLCELL_X32 FILLER_81_2480 ();
 FILLCELL_X8 FILLER_81_2512 ();
 FILLCELL_X4 FILLER_81_2520 ();
 FILLCELL_X2 FILLER_81_2524 ();
 FILLCELL_X32 FILLER_81_2527 ();
 FILLCELL_X32 FILLER_81_2559 ();
 FILLCELL_X32 FILLER_81_2591 ();
 FILLCELL_X32 FILLER_81_2623 ();
 FILLCELL_X32 FILLER_81_2655 ();
 FILLCELL_X32 FILLER_81_2687 ();
 FILLCELL_X32 FILLER_81_2719 ();
 FILLCELL_X32 FILLER_81_2751 ();
 FILLCELL_X32 FILLER_81_2783 ();
 FILLCELL_X32 FILLER_81_2815 ();
 FILLCELL_X32 FILLER_81_2847 ();
 FILLCELL_X32 FILLER_81_2879 ();
 FILLCELL_X32 FILLER_81_2911 ();
 FILLCELL_X32 FILLER_81_2943 ();
 FILLCELL_X32 FILLER_81_2975 ();
 FILLCELL_X32 FILLER_81_3007 ();
 FILLCELL_X32 FILLER_81_3039 ();
 FILLCELL_X32 FILLER_81_3071 ();
 FILLCELL_X32 FILLER_81_3103 ();
 FILLCELL_X32 FILLER_81_3135 ();
 FILLCELL_X32 FILLER_81_3167 ();
 FILLCELL_X32 FILLER_81_3199 ();
 FILLCELL_X32 FILLER_81_3231 ();
 FILLCELL_X32 FILLER_81_3263 ();
 FILLCELL_X32 FILLER_81_3295 ();
 FILLCELL_X32 FILLER_81_3327 ();
 FILLCELL_X32 FILLER_81_3359 ();
 FILLCELL_X32 FILLER_81_3391 ();
 FILLCELL_X32 FILLER_81_3423 ();
 FILLCELL_X32 FILLER_81_3455 ();
 FILLCELL_X32 FILLER_81_3487 ();
 FILLCELL_X32 FILLER_81_3519 ();
 FILLCELL_X32 FILLER_81_3551 ();
 FILLCELL_X32 FILLER_81_3583 ();
 FILLCELL_X32 FILLER_81_3615 ();
 FILLCELL_X32 FILLER_81_3647 ();
 FILLCELL_X32 FILLER_81_3679 ();
 FILLCELL_X16 FILLER_81_3711 ();
 FILLCELL_X8 FILLER_81_3727 ();
 FILLCELL_X2 FILLER_81_3735 ();
 FILLCELL_X1 FILLER_81_3737 ();
 FILLCELL_X32 FILLER_82_1 ();
 FILLCELL_X32 FILLER_82_33 ();
 FILLCELL_X32 FILLER_82_65 ();
 FILLCELL_X32 FILLER_82_97 ();
 FILLCELL_X32 FILLER_82_129 ();
 FILLCELL_X32 FILLER_82_161 ();
 FILLCELL_X32 FILLER_82_193 ();
 FILLCELL_X32 FILLER_82_225 ();
 FILLCELL_X32 FILLER_82_257 ();
 FILLCELL_X32 FILLER_82_289 ();
 FILLCELL_X32 FILLER_82_321 ();
 FILLCELL_X32 FILLER_82_353 ();
 FILLCELL_X32 FILLER_82_385 ();
 FILLCELL_X32 FILLER_82_417 ();
 FILLCELL_X32 FILLER_82_449 ();
 FILLCELL_X32 FILLER_82_481 ();
 FILLCELL_X32 FILLER_82_513 ();
 FILLCELL_X32 FILLER_82_545 ();
 FILLCELL_X32 FILLER_82_577 ();
 FILLCELL_X16 FILLER_82_609 ();
 FILLCELL_X4 FILLER_82_625 ();
 FILLCELL_X2 FILLER_82_629 ();
 FILLCELL_X32 FILLER_82_632 ();
 FILLCELL_X32 FILLER_82_664 ();
 FILLCELL_X32 FILLER_82_696 ();
 FILLCELL_X32 FILLER_82_728 ();
 FILLCELL_X32 FILLER_82_760 ();
 FILLCELL_X32 FILLER_82_792 ();
 FILLCELL_X32 FILLER_82_824 ();
 FILLCELL_X32 FILLER_82_856 ();
 FILLCELL_X32 FILLER_82_888 ();
 FILLCELL_X32 FILLER_82_920 ();
 FILLCELL_X32 FILLER_82_952 ();
 FILLCELL_X32 FILLER_82_984 ();
 FILLCELL_X32 FILLER_82_1016 ();
 FILLCELL_X32 FILLER_82_1048 ();
 FILLCELL_X32 FILLER_82_1080 ();
 FILLCELL_X32 FILLER_82_1112 ();
 FILLCELL_X32 FILLER_82_1144 ();
 FILLCELL_X32 FILLER_82_1176 ();
 FILLCELL_X32 FILLER_82_1208 ();
 FILLCELL_X32 FILLER_82_1240 ();
 FILLCELL_X32 FILLER_82_1272 ();
 FILLCELL_X32 FILLER_82_1304 ();
 FILLCELL_X32 FILLER_82_1336 ();
 FILLCELL_X32 FILLER_82_1368 ();
 FILLCELL_X32 FILLER_82_1400 ();
 FILLCELL_X32 FILLER_82_1432 ();
 FILLCELL_X32 FILLER_82_1464 ();
 FILLCELL_X32 FILLER_82_1496 ();
 FILLCELL_X32 FILLER_82_1528 ();
 FILLCELL_X32 FILLER_82_1560 ();
 FILLCELL_X32 FILLER_82_1592 ();
 FILLCELL_X32 FILLER_82_1624 ();
 FILLCELL_X32 FILLER_82_1656 ();
 FILLCELL_X32 FILLER_82_1688 ();
 FILLCELL_X32 FILLER_82_1720 ();
 FILLCELL_X32 FILLER_82_1752 ();
 FILLCELL_X32 FILLER_82_1784 ();
 FILLCELL_X32 FILLER_82_1816 ();
 FILLCELL_X32 FILLER_82_1848 ();
 FILLCELL_X8 FILLER_82_1880 ();
 FILLCELL_X4 FILLER_82_1888 ();
 FILLCELL_X2 FILLER_82_1892 ();
 FILLCELL_X32 FILLER_82_1895 ();
 FILLCELL_X32 FILLER_82_1927 ();
 FILLCELL_X32 FILLER_82_1959 ();
 FILLCELL_X32 FILLER_82_1991 ();
 FILLCELL_X32 FILLER_82_2023 ();
 FILLCELL_X32 FILLER_82_2055 ();
 FILLCELL_X32 FILLER_82_2087 ();
 FILLCELL_X32 FILLER_82_2119 ();
 FILLCELL_X32 FILLER_82_2151 ();
 FILLCELL_X32 FILLER_82_2183 ();
 FILLCELL_X32 FILLER_82_2215 ();
 FILLCELL_X32 FILLER_82_2247 ();
 FILLCELL_X32 FILLER_82_2279 ();
 FILLCELL_X32 FILLER_82_2311 ();
 FILLCELL_X32 FILLER_82_2343 ();
 FILLCELL_X32 FILLER_82_2375 ();
 FILLCELL_X32 FILLER_82_2407 ();
 FILLCELL_X32 FILLER_82_2439 ();
 FILLCELL_X32 FILLER_82_2471 ();
 FILLCELL_X32 FILLER_82_2503 ();
 FILLCELL_X32 FILLER_82_2535 ();
 FILLCELL_X32 FILLER_82_2567 ();
 FILLCELL_X32 FILLER_82_2599 ();
 FILLCELL_X32 FILLER_82_2631 ();
 FILLCELL_X32 FILLER_82_2663 ();
 FILLCELL_X32 FILLER_82_2695 ();
 FILLCELL_X32 FILLER_82_2727 ();
 FILLCELL_X32 FILLER_82_2759 ();
 FILLCELL_X32 FILLER_82_2791 ();
 FILLCELL_X32 FILLER_82_2823 ();
 FILLCELL_X32 FILLER_82_2855 ();
 FILLCELL_X32 FILLER_82_2887 ();
 FILLCELL_X32 FILLER_82_2919 ();
 FILLCELL_X32 FILLER_82_2951 ();
 FILLCELL_X32 FILLER_82_2983 ();
 FILLCELL_X32 FILLER_82_3015 ();
 FILLCELL_X32 FILLER_82_3047 ();
 FILLCELL_X32 FILLER_82_3079 ();
 FILLCELL_X32 FILLER_82_3111 ();
 FILLCELL_X8 FILLER_82_3143 ();
 FILLCELL_X4 FILLER_82_3151 ();
 FILLCELL_X2 FILLER_82_3155 ();
 FILLCELL_X32 FILLER_82_3158 ();
 FILLCELL_X32 FILLER_82_3190 ();
 FILLCELL_X32 FILLER_82_3222 ();
 FILLCELL_X32 FILLER_82_3254 ();
 FILLCELL_X32 FILLER_82_3286 ();
 FILLCELL_X32 FILLER_82_3318 ();
 FILLCELL_X32 FILLER_82_3350 ();
 FILLCELL_X32 FILLER_82_3382 ();
 FILLCELL_X32 FILLER_82_3414 ();
 FILLCELL_X32 FILLER_82_3446 ();
 FILLCELL_X32 FILLER_82_3478 ();
 FILLCELL_X32 FILLER_82_3510 ();
 FILLCELL_X32 FILLER_82_3542 ();
 FILLCELL_X32 FILLER_82_3574 ();
 FILLCELL_X32 FILLER_82_3606 ();
 FILLCELL_X32 FILLER_82_3638 ();
 FILLCELL_X32 FILLER_82_3670 ();
 FILLCELL_X32 FILLER_82_3702 ();
 FILLCELL_X4 FILLER_82_3734 ();
 FILLCELL_X32 FILLER_83_1 ();
 FILLCELL_X32 FILLER_83_33 ();
 FILLCELL_X32 FILLER_83_65 ();
 FILLCELL_X32 FILLER_83_97 ();
 FILLCELL_X32 FILLER_83_129 ();
 FILLCELL_X32 FILLER_83_161 ();
 FILLCELL_X32 FILLER_83_193 ();
 FILLCELL_X32 FILLER_83_225 ();
 FILLCELL_X32 FILLER_83_257 ();
 FILLCELL_X32 FILLER_83_289 ();
 FILLCELL_X32 FILLER_83_321 ();
 FILLCELL_X32 FILLER_83_353 ();
 FILLCELL_X32 FILLER_83_385 ();
 FILLCELL_X32 FILLER_83_417 ();
 FILLCELL_X32 FILLER_83_449 ();
 FILLCELL_X32 FILLER_83_481 ();
 FILLCELL_X32 FILLER_83_513 ();
 FILLCELL_X32 FILLER_83_545 ();
 FILLCELL_X32 FILLER_83_577 ();
 FILLCELL_X32 FILLER_83_609 ();
 FILLCELL_X32 FILLER_83_641 ();
 FILLCELL_X32 FILLER_83_673 ();
 FILLCELL_X32 FILLER_83_705 ();
 FILLCELL_X32 FILLER_83_737 ();
 FILLCELL_X32 FILLER_83_769 ();
 FILLCELL_X32 FILLER_83_801 ();
 FILLCELL_X32 FILLER_83_833 ();
 FILLCELL_X32 FILLER_83_865 ();
 FILLCELL_X32 FILLER_83_897 ();
 FILLCELL_X32 FILLER_83_929 ();
 FILLCELL_X32 FILLER_83_961 ();
 FILLCELL_X32 FILLER_83_993 ();
 FILLCELL_X32 FILLER_83_1025 ();
 FILLCELL_X32 FILLER_83_1057 ();
 FILLCELL_X32 FILLER_83_1089 ();
 FILLCELL_X32 FILLER_83_1121 ();
 FILLCELL_X32 FILLER_83_1153 ();
 FILLCELL_X32 FILLER_83_1185 ();
 FILLCELL_X32 FILLER_83_1217 ();
 FILLCELL_X8 FILLER_83_1249 ();
 FILLCELL_X4 FILLER_83_1257 ();
 FILLCELL_X2 FILLER_83_1261 ();
 FILLCELL_X32 FILLER_83_1264 ();
 FILLCELL_X32 FILLER_83_1296 ();
 FILLCELL_X32 FILLER_83_1328 ();
 FILLCELL_X32 FILLER_83_1360 ();
 FILLCELL_X32 FILLER_83_1392 ();
 FILLCELL_X32 FILLER_83_1424 ();
 FILLCELL_X32 FILLER_83_1456 ();
 FILLCELL_X32 FILLER_83_1488 ();
 FILLCELL_X32 FILLER_83_1520 ();
 FILLCELL_X32 FILLER_83_1552 ();
 FILLCELL_X32 FILLER_83_1584 ();
 FILLCELL_X32 FILLER_83_1616 ();
 FILLCELL_X32 FILLER_83_1648 ();
 FILLCELL_X32 FILLER_83_1680 ();
 FILLCELL_X32 FILLER_83_1712 ();
 FILLCELL_X32 FILLER_83_1744 ();
 FILLCELL_X32 FILLER_83_1776 ();
 FILLCELL_X32 FILLER_83_1808 ();
 FILLCELL_X32 FILLER_83_1840 ();
 FILLCELL_X32 FILLER_83_1872 ();
 FILLCELL_X32 FILLER_83_1904 ();
 FILLCELL_X32 FILLER_83_1936 ();
 FILLCELL_X32 FILLER_83_1968 ();
 FILLCELL_X32 FILLER_83_2000 ();
 FILLCELL_X32 FILLER_83_2032 ();
 FILLCELL_X32 FILLER_83_2064 ();
 FILLCELL_X32 FILLER_83_2096 ();
 FILLCELL_X32 FILLER_83_2128 ();
 FILLCELL_X32 FILLER_83_2160 ();
 FILLCELL_X32 FILLER_83_2192 ();
 FILLCELL_X32 FILLER_83_2224 ();
 FILLCELL_X32 FILLER_83_2256 ();
 FILLCELL_X32 FILLER_83_2288 ();
 FILLCELL_X32 FILLER_83_2320 ();
 FILLCELL_X32 FILLER_83_2352 ();
 FILLCELL_X32 FILLER_83_2384 ();
 FILLCELL_X32 FILLER_83_2416 ();
 FILLCELL_X32 FILLER_83_2448 ();
 FILLCELL_X32 FILLER_83_2480 ();
 FILLCELL_X8 FILLER_83_2512 ();
 FILLCELL_X4 FILLER_83_2520 ();
 FILLCELL_X2 FILLER_83_2524 ();
 FILLCELL_X32 FILLER_83_2527 ();
 FILLCELL_X32 FILLER_83_2559 ();
 FILLCELL_X32 FILLER_83_2591 ();
 FILLCELL_X32 FILLER_83_2623 ();
 FILLCELL_X32 FILLER_83_2655 ();
 FILLCELL_X32 FILLER_83_2687 ();
 FILLCELL_X32 FILLER_83_2719 ();
 FILLCELL_X32 FILLER_83_2751 ();
 FILLCELL_X32 FILLER_83_2783 ();
 FILLCELL_X32 FILLER_83_2815 ();
 FILLCELL_X32 FILLER_83_2847 ();
 FILLCELL_X32 FILLER_83_2879 ();
 FILLCELL_X32 FILLER_83_2911 ();
 FILLCELL_X32 FILLER_83_2943 ();
 FILLCELL_X32 FILLER_83_2975 ();
 FILLCELL_X32 FILLER_83_3007 ();
 FILLCELL_X32 FILLER_83_3039 ();
 FILLCELL_X32 FILLER_83_3071 ();
 FILLCELL_X32 FILLER_83_3103 ();
 FILLCELL_X32 FILLER_83_3135 ();
 FILLCELL_X32 FILLER_83_3167 ();
 FILLCELL_X32 FILLER_83_3199 ();
 FILLCELL_X32 FILLER_83_3231 ();
 FILLCELL_X32 FILLER_83_3263 ();
 FILLCELL_X32 FILLER_83_3295 ();
 FILLCELL_X32 FILLER_83_3327 ();
 FILLCELL_X32 FILLER_83_3359 ();
 FILLCELL_X32 FILLER_83_3391 ();
 FILLCELL_X32 FILLER_83_3423 ();
 FILLCELL_X32 FILLER_83_3455 ();
 FILLCELL_X32 FILLER_83_3487 ();
 FILLCELL_X32 FILLER_83_3519 ();
 FILLCELL_X32 FILLER_83_3551 ();
 FILLCELL_X32 FILLER_83_3583 ();
 FILLCELL_X32 FILLER_83_3615 ();
 FILLCELL_X32 FILLER_83_3647 ();
 FILLCELL_X32 FILLER_83_3679 ();
 FILLCELL_X16 FILLER_83_3711 ();
 FILLCELL_X8 FILLER_83_3727 ();
 FILLCELL_X2 FILLER_83_3735 ();
 FILLCELL_X1 FILLER_83_3737 ();
 FILLCELL_X32 FILLER_84_1 ();
 FILLCELL_X32 FILLER_84_33 ();
 FILLCELL_X32 FILLER_84_65 ();
 FILLCELL_X32 FILLER_84_97 ();
 FILLCELL_X32 FILLER_84_129 ();
 FILLCELL_X32 FILLER_84_161 ();
 FILLCELL_X32 FILLER_84_193 ();
 FILLCELL_X32 FILLER_84_225 ();
 FILLCELL_X32 FILLER_84_257 ();
 FILLCELL_X32 FILLER_84_289 ();
 FILLCELL_X32 FILLER_84_321 ();
 FILLCELL_X32 FILLER_84_353 ();
 FILLCELL_X32 FILLER_84_385 ();
 FILLCELL_X32 FILLER_84_417 ();
 FILLCELL_X32 FILLER_84_449 ();
 FILLCELL_X32 FILLER_84_481 ();
 FILLCELL_X32 FILLER_84_513 ();
 FILLCELL_X32 FILLER_84_545 ();
 FILLCELL_X32 FILLER_84_577 ();
 FILLCELL_X16 FILLER_84_609 ();
 FILLCELL_X4 FILLER_84_625 ();
 FILLCELL_X2 FILLER_84_629 ();
 FILLCELL_X32 FILLER_84_632 ();
 FILLCELL_X32 FILLER_84_664 ();
 FILLCELL_X32 FILLER_84_696 ();
 FILLCELL_X32 FILLER_84_728 ();
 FILLCELL_X32 FILLER_84_760 ();
 FILLCELL_X32 FILLER_84_792 ();
 FILLCELL_X32 FILLER_84_824 ();
 FILLCELL_X32 FILLER_84_856 ();
 FILLCELL_X32 FILLER_84_888 ();
 FILLCELL_X32 FILLER_84_920 ();
 FILLCELL_X32 FILLER_84_952 ();
 FILLCELL_X32 FILLER_84_984 ();
 FILLCELL_X32 FILLER_84_1016 ();
 FILLCELL_X32 FILLER_84_1048 ();
 FILLCELL_X32 FILLER_84_1080 ();
 FILLCELL_X32 FILLER_84_1112 ();
 FILLCELL_X32 FILLER_84_1144 ();
 FILLCELL_X32 FILLER_84_1176 ();
 FILLCELL_X32 FILLER_84_1208 ();
 FILLCELL_X32 FILLER_84_1240 ();
 FILLCELL_X32 FILLER_84_1272 ();
 FILLCELL_X32 FILLER_84_1304 ();
 FILLCELL_X32 FILLER_84_1336 ();
 FILLCELL_X32 FILLER_84_1368 ();
 FILLCELL_X32 FILLER_84_1400 ();
 FILLCELL_X32 FILLER_84_1432 ();
 FILLCELL_X32 FILLER_84_1464 ();
 FILLCELL_X32 FILLER_84_1496 ();
 FILLCELL_X32 FILLER_84_1528 ();
 FILLCELL_X32 FILLER_84_1560 ();
 FILLCELL_X32 FILLER_84_1592 ();
 FILLCELL_X32 FILLER_84_1624 ();
 FILLCELL_X32 FILLER_84_1656 ();
 FILLCELL_X32 FILLER_84_1688 ();
 FILLCELL_X32 FILLER_84_1720 ();
 FILLCELL_X32 FILLER_84_1752 ();
 FILLCELL_X32 FILLER_84_1784 ();
 FILLCELL_X32 FILLER_84_1816 ();
 FILLCELL_X32 FILLER_84_1848 ();
 FILLCELL_X8 FILLER_84_1880 ();
 FILLCELL_X4 FILLER_84_1888 ();
 FILLCELL_X2 FILLER_84_1892 ();
 FILLCELL_X32 FILLER_84_1895 ();
 FILLCELL_X32 FILLER_84_1927 ();
 FILLCELL_X32 FILLER_84_1959 ();
 FILLCELL_X32 FILLER_84_1991 ();
 FILLCELL_X32 FILLER_84_2023 ();
 FILLCELL_X32 FILLER_84_2055 ();
 FILLCELL_X32 FILLER_84_2087 ();
 FILLCELL_X32 FILLER_84_2119 ();
 FILLCELL_X32 FILLER_84_2151 ();
 FILLCELL_X32 FILLER_84_2183 ();
 FILLCELL_X32 FILLER_84_2215 ();
 FILLCELL_X32 FILLER_84_2247 ();
 FILLCELL_X32 FILLER_84_2279 ();
 FILLCELL_X32 FILLER_84_2311 ();
 FILLCELL_X32 FILLER_84_2343 ();
 FILLCELL_X32 FILLER_84_2375 ();
 FILLCELL_X32 FILLER_84_2407 ();
 FILLCELL_X32 FILLER_84_2439 ();
 FILLCELL_X32 FILLER_84_2471 ();
 FILLCELL_X32 FILLER_84_2503 ();
 FILLCELL_X32 FILLER_84_2535 ();
 FILLCELL_X32 FILLER_84_2567 ();
 FILLCELL_X32 FILLER_84_2599 ();
 FILLCELL_X32 FILLER_84_2631 ();
 FILLCELL_X32 FILLER_84_2663 ();
 FILLCELL_X32 FILLER_84_2695 ();
 FILLCELL_X32 FILLER_84_2727 ();
 FILLCELL_X32 FILLER_84_2759 ();
 FILLCELL_X32 FILLER_84_2791 ();
 FILLCELL_X32 FILLER_84_2823 ();
 FILLCELL_X32 FILLER_84_2855 ();
 FILLCELL_X32 FILLER_84_2887 ();
 FILLCELL_X32 FILLER_84_2919 ();
 FILLCELL_X32 FILLER_84_2951 ();
 FILLCELL_X32 FILLER_84_2983 ();
 FILLCELL_X32 FILLER_84_3015 ();
 FILLCELL_X32 FILLER_84_3047 ();
 FILLCELL_X32 FILLER_84_3079 ();
 FILLCELL_X32 FILLER_84_3111 ();
 FILLCELL_X8 FILLER_84_3143 ();
 FILLCELL_X4 FILLER_84_3151 ();
 FILLCELL_X2 FILLER_84_3155 ();
 FILLCELL_X32 FILLER_84_3158 ();
 FILLCELL_X32 FILLER_84_3190 ();
 FILLCELL_X32 FILLER_84_3222 ();
 FILLCELL_X32 FILLER_84_3254 ();
 FILLCELL_X32 FILLER_84_3286 ();
 FILLCELL_X32 FILLER_84_3318 ();
 FILLCELL_X32 FILLER_84_3350 ();
 FILLCELL_X32 FILLER_84_3382 ();
 FILLCELL_X32 FILLER_84_3414 ();
 FILLCELL_X32 FILLER_84_3446 ();
 FILLCELL_X32 FILLER_84_3478 ();
 FILLCELL_X32 FILLER_84_3510 ();
 FILLCELL_X32 FILLER_84_3542 ();
 FILLCELL_X32 FILLER_84_3574 ();
 FILLCELL_X32 FILLER_84_3606 ();
 FILLCELL_X32 FILLER_84_3638 ();
 FILLCELL_X32 FILLER_84_3670 ();
 FILLCELL_X32 FILLER_84_3702 ();
 FILLCELL_X4 FILLER_84_3734 ();
 FILLCELL_X32 FILLER_85_1 ();
 FILLCELL_X32 FILLER_85_33 ();
 FILLCELL_X32 FILLER_85_65 ();
 FILLCELL_X32 FILLER_85_97 ();
 FILLCELL_X32 FILLER_85_129 ();
 FILLCELL_X32 FILLER_85_161 ();
 FILLCELL_X32 FILLER_85_193 ();
 FILLCELL_X32 FILLER_85_225 ();
 FILLCELL_X32 FILLER_85_257 ();
 FILLCELL_X32 FILLER_85_289 ();
 FILLCELL_X32 FILLER_85_321 ();
 FILLCELL_X32 FILLER_85_353 ();
 FILLCELL_X32 FILLER_85_385 ();
 FILLCELL_X32 FILLER_85_417 ();
 FILLCELL_X32 FILLER_85_449 ();
 FILLCELL_X32 FILLER_85_481 ();
 FILLCELL_X32 FILLER_85_513 ();
 FILLCELL_X32 FILLER_85_545 ();
 FILLCELL_X32 FILLER_85_577 ();
 FILLCELL_X32 FILLER_85_609 ();
 FILLCELL_X32 FILLER_85_641 ();
 FILLCELL_X32 FILLER_85_673 ();
 FILLCELL_X32 FILLER_85_705 ();
 FILLCELL_X32 FILLER_85_737 ();
 FILLCELL_X32 FILLER_85_769 ();
 FILLCELL_X32 FILLER_85_801 ();
 FILLCELL_X32 FILLER_85_833 ();
 FILLCELL_X32 FILLER_85_865 ();
 FILLCELL_X32 FILLER_85_897 ();
 FILLCELL_X32 FILLER_85_929 ();
 FILLCELL_X32 FILLER_85_961 ();
 FILLCELL_X32 FILLER_85_993 ();
 FILLCELL_X32 FILLER_85_1025 ();
 FILLCELL_X32 FILLER_85_1057 ();
 FILLCELL_X32 FILLER_85_1089 ();
 FILLCELL_X32 FILLER_85_1121 ();
 FILLCELL_X32 FILLER_85_1153 ();
 FILLCELL_X32 FILLER_85_1185 ();
 FILLCELL_X32 FILLER_85_1217 ();
 FILLCELL_X8 FILLER_85_1249 ();
 FILLCELL_X4 FILLER_85_1257 ();
 FILLCELL_X2 FILLER_85_1261 ();
 FILLCELL_X32 FILLER_85_1264 ();
 FILLCELL_X32 FILLER_85_1296 ();
 FILLCELL_X32 FILLER_85_1328 ();
 FILLCELL_X32 FILLER_85_1360 ();
 FILLCELL_X32 FILLER_85_1392 ();
 FILLCELL_X32 FILLER_85_1424 ();
 FILLCELL_X32 FILLER_85_1456 ();
 FILLCELL_X32 FILLER_85_1488 ();
 FILLCELL_X32 FILLER_85_1520 ();
 FILLCELL_X32 FILLER_85_1552 ();
 FILLCELL_X32 FILLER_85_1584 ();
 FILLCELL_X32 FILLER_85_1616 ();
 FILLCELL_X32 FILLER_85_1648 ();
 FILLCELL_X32 FILLER_85_1680 ();
 FILLCELL_X32 FILLER_85_1712 ();
 FILLCELL_X32 FILLER_85_1744 ();
 FILLCELL_X32 FILLER_85_1776 ();
 FILLCELL_X32 FILLER_85_1808 ();
 FILLCELL_X32 FILLER_85_1840 ();
 FILLCELL_X32 FILLER_85_1872 ();
 FILLCELL_X32 FILLER_85_1904 ();
 FILLCELL_X32 FILLER_85_1936 ();
 FILLCELL_X32 FILLER_85_1968 ();
 FILLCELL_X32 FILLER_85_2000 ();
 FILLCELL_X32 FILLER_85_2032 ();
 FILLCELL_X32 FILLER_85_2064 ();
 FILLCELL_X32 FILLER_85_2096 ();
 FILLCELL_X32 FILLER_85_2128 ();
 FILLCELL_X32 FILLER_85_2160 ();
 FILLCELL_X32 FILLER_85_2192 ();
 FILLCELL_X32 FILLER_85_2224 ();
 FILLCELL_X32 FILLER_85_2256 ();
 FILLCELL_X32 FILLER_85_2288 ();
 FILLCELL_X32 FILLER_85_2320 ();
 FILLCELL_X32 FILLER_85_2352 ();
 FILLCELL_X32 FILLER_85_2384 ();
 FILLCELL_X32 FILLER_85_2416 ();
 FILLCELL_X32 FILLER_85_2448 ();
 FILLCELL_X32 FILLER_85_2480 ();
 FILLCELL_X8 FILLER_85_2512 ();
 FILLCELL_X4 FILLER_85_2520 ();
 FILLCELL_X2 FILLER_85_2524 ();
 FILLCELL_X32 FILLER_85_2527 ();
 FILLCELL_X32 FILLER_85_2559 ();
 FILLCELL_X32 FILLER_85_2591 ();
 FILLCELL_X32 FILLER_85_2623 ();
 FILLCELL_X32 FILLER_85_2655 ();
 FILLCELL_X32 FILLER_85_2687 ();
 FILLCELL_X32 FILLER_85_2719 ();
 FILLCELL_X32 FILLER_85_2751 ();
 FILLCELL_X32 FILLER_85_2783 ();
 FILLCELL_X32 FILLER_85_2815 ();
 FILLCELL_X32 FILLER_85_2847 ();
 FILLCELL_X32 FILLER_85_2879 ();
 FILLCELL_X32 FILLER_85_2911 ();
 FILLCELL_X32 FILLER_85_2943 ();
 FILLCELL_X32 FILLER_85_2975 ();
 FILLCELL_X32 FILLER_85_3007 ();
 FILLCELL_X32 FILLER_85_3039 ();
 FILLCELL_X32 FILLER_85_3071 ();
 FILLCELL_X32 FILLER_85_3103 ();
 FILLCELL_X32 FILLER_85_3135 ();
 FILLCELL_X32 FILLER_85_3167 ();
 FILLCELL_X32 FILLER_85_3199 ();
 FILLCELL_X32 FILLER_85_3231 ();
 FILLCELL_X32 FILLER_85_3263 ();
 FILLCELL_X32 FILLER_85_3295 ();
 FILLCELL_X32 FILLER_85_3327 ();
 FILLCELL_X32 FILLER_85_3359 ();
 FILLCELL_X32 FILLER_85_3391 ();
 FILLCELL_X32 FILLER_85_3423 ();
 FILLCELL_X32 FILLER_85_3455 ();
 FILLCELL_X32 FILLER_85_3487 ();
 FILLCELL_X32 FILLER_85_3519 ();
 FILLCELL_X32 FILLER_85_3551 ();
 FILLCELL_X32 FILLER_85_3583 ();
 FILLCELL_X32 FILLER_85_3615 ();
 FILLCELL_X32 FILLER_85_3647 ();
 FILLCELL_X32 FILLER_85_3679 ();
 FILLCELL_X16 FILLER_85_3711 ();
 FILLCELL_X8 FILLER_85_3727 ();
 FILLCELL_X2 FILLER_85_3735 ();
 FILLCELL_X1 FILLER_85_3737 ();
 FILLCELL_X32 FILLER_86_1 ();
 FILLCELL_X32 FILLER_86_33 ();
 FILLCELL_X32 FILLER_86_65 ();
 FILLCELL_X32 FILLER_86_97 ();
 FILLCELL_X32 FILLER_86_129 ();
 FILLCELL_X32 FILLER_86_161 ();
 FILLCELL_X32 FILLER_86_193 ();
 FILLCELL_X32 FILLER_86_225 ();
 FILLCELL_X32 FILLER_86_257 ();
 FILLCELL_X32 FILLER_86_289 ();
 FILLCELL_X32 FILLER_86_321 ();
 FILLCELL_X32 FILLER_86_353 ();
 FILLCELL_X32 FILLER_86_385 ();
 FILLCELL_X32 FILLER_86_417 ();
 FILLCELL_X32 FILLER_86_449 ();
 FILLCELL_X32 FILLER_86_481 ();
 FILLCELL_X32 FILLER_86_513 ();
 FILLCELL_X32 FILLER_86_545 ();
 FILLCELL_X32 FILLER_86_577 ();
 FILLCELL_X16 FILLER_86_609 ();
 FILLCELL_X4 FILLER_86_625 ();
 FILLCELL_X2 FILLER_86_629 ();
 FILLCELL_X32 FILLER_86_632 ();
 FILLCELL_X32 FILLER_86_664 ();
 FILLCELL_X32 FILLER_86_696 ();
 FILLCELL_X32 FILLER_86_728 ();
 FILLCELL_X32 FILLER_86_760 ();
 FILLCELL_X32 FILLER_86_792 ();
 FILLCELL_X32 FILLER_86_824 ();
 FILLCELL_X32 FILLER_86_856 ();
 FILLCELL_X32 FILLER_86_888 ();
 FILLCELL_X32 FILLER_86_920 ();
 FILLCELL_X32 FILLER_86_952 ();
 FILLCELL_X32 FILLER_86_984 ();
 FILLCELL_X32 FILLER_86_1016 ();
 FILLCELL_X32 FILLER_86_1048 ();
 FILLCELL_X32 FILLER_86_1080 ();
 FILLCELL_X32 FILLER_86_1112 ();
 FILLCELL_X32 FILLER_86_1144 ();
 FILLCELL_X32 FILLER_86_1176 ();
 FILLCELL_X32 FILLER_86_1208 ();
 FILLCELL_X32 FILLER_86_1240 ();
 FILLCELL_X32 FILLER_86_1272 ();
 FILLCELL_X32 FILLER_86_1304 ();
 FILLCELL_X32 FILLER_86_1336 ();
 FILLCELL_X32 FILLER_86_1368 ();
 FILLCELL_X32 FILLER_86_1400 ();
 FILLCELL_X32 FILLER_86_1432 ();
 FILLCELL_X32 FILLER_86_1464 ();
 FILLCELL_X32 FILLER_86_1496 ();
 FILLCELL_X32 FILLER_86_1528 ();
 FILLCELL_X32 FILLER_86_1560 ();
 FILLCELL_X32 FILLER_86_1592 ();
 FILLCELL_X32 FILLER_86_1624 ();
 FILLCELL_X32 FILLER_86_1656 ();
 FILLCELL_X32 FILLER_86_1688 ();
 FILLCELL_X32 FILLER_86_1720 ();
 FILLCELL_X32 FILLER_86_1752 ();
 FILLCELL_X32 FILLER_86_1784 ();
 FILLCELL_X32 FILLER_86_1816 ();
 FILLCELL_X32 FILLER_86_1848 ();
 FILLCELL_X8 FILLER_86_1880 ();
 FILLCELL_X4 FILLER_86_1888 ();
 FILLCELL_X2 FILLER_86_1892 ();
 FILLCELL_X32 FILLER_86_1895 ();
 FILLCELL_X32 FILLER_86_1927 ();
 FILLCELL_X32 FILLER_86_1959 ();
 FILLCELL_X32 FILLER_86_1991 ();
 FILLCELL_X32 FILLER_86_2023 ();
 FILLCELL_X32 FILLER_86_2055 ();
 FILLCELL_X32 FILLER_86_2087 ();
 FILLCELL_X32 FILLER_86_2119 ();
 FILLCELL_X32 FILLER_86_2151 ();
 FILLCELL_X32 FILLER_86_2183 ();
 FILLCELL_X32 FILLER_86_2215 ();
 FILLCELL_X32 FILLER_86_2247 ();
 FILLCELL_X32 FILLER_86_2279 ();
 FILLCELL_X32 FILLER_86_2311 ();
 FILLCELL_X32 FILLER_86_2343 ();
 FILLCELL_X32 FILLER_86_2375 ();
 FILLCELL_X32 FILLER_86_2407 ();
 FILLCELL_X32 FILLER_86_2439 ();
 FILLCELL_X32 FILLER_86_2471 ();
 FILLCELL_X32 FILLER_86_2503 ();
 FILLCELL_X32 FILLER_86_2535 ();
 FILLCELL_X32 FILLER_86_2567 ();
 FILLCELL_X32 FILLER_86_2599 ();
 FILLCELL_X32 FILLER_86_2631 ();
 FILLCELL_X32 FILLER_86_2663 ();
 FILLCELL_X32 FILLER_86_2695 ();
 FILLCELL_X32 FILLER_86_2727 ();
 FILLCELL_X32 FILLER_86_2759 ();
 FILLCELL_X32 FILLER_86_2791 ();
 FILLCELL_X32 FILLER_86_2823 ();
 FILLCELL_X32 FILLER_86_2855 ();
 FILLCELL_X32 FILLER_86_2887 ();
 FILLCELL_X32 FILLER_86_2919 ();
 FILLCELL_X32 FILLER_86_2951 ();
 FILLCELL_X32 FILLER_86_2983 ();
 FILLCELL_X32 FILLER_86_3015 ();
 FILLCELL_X32 FILLER_86_3047 ();
 FILLCELL_X32 FILLER_86_3079 ();
 FILLCELL_X32 FILLER_86_3111 ();
 FILLCELL_X8 FILLER_86_3143 ();
 FILLCELL_X4 FILLER_86_3151 ();
 FILLCELL_X2 FILLER_86_3155 ();
 FILLCELL_X32 FILLER_86_3158 ();
 FILLCELL_X32 FILLER_86_3190 ();
 FILLCELL_X32 FILLER_86_3222 ();
 FILLCELL_X32 FILLER_86_3254 ();
 FILLCELL_X32 FILLER_86_3286 ();
 FILLCELL_X32 FILLER_86_3318 ();
 FILLCELL_X32 FILLER_86_3350 ();
 FILLCELL_X32 FILLER_86_3382 ();
 FILLCELL_X32 FILLER_86_3414 ();
 FILLCELL_X32 FILLER_86_3446 ();
 FILLCELL_X32 FILLER_86_3478 ();
 FILLCELL_X32 FILLER_86_3510 ();
 FILLCELL_X32 FILLER_86_3542 ();
 FILLCELL_X32 FILLER_86_3574 ();
 FILLCELL_X32 FILLER_86_3606 ();
 FILLCELL_X32 FILLER_86_3638 ();
 FILLCELL_X32 FILLER_86_3670 ();
 FILLCELL_X32 FILLER_86_3702 ();
 FILLCELL_X4 FILLER_86_3734 ();
 FILLCELL_X32 FILLER_87_1 ();
 FILLCELL_X32 FILLER_87_33 ();
 FILLCELL_X32 FILLER_87_65 ();
 FILLCELL_X32 FILLER_87_97 ();
 FILLCELL_X32 FILLER_87_129 ();
 FILLCELL_X32 FILLER_87_161 ();
 FILLCELL_X32 FILLER_87_193 ();
 FILLCELL_X32 FILLER_87_225 ();
 FILLCELL_X32 FILLER_87_257 ();
 FILLCELL_X32 FILLER_87_289 ();
 FILLCELL_X32 FILLER_87_321 ();
 FILLCELL_X32 FILLER_87_353 ();
 FILLCELL_X32 FILLER_87_385 ();
 FILLCELL_X32 FILLER_87_417 ();
 FILLCELL_X32 FILLER_87_449 ();
 FILLCELL_X32 FILLER_87_481 ();
 FILLCELL_X32 FILLER_87_513 ();
 FILLCELL_X32 FILLER_87_545 ();
 FILLCELL_X32 FILLER_87_577 ();
 FILLCELL_X32 FILLER_87_609 ();
 FILLCELL_X32 FILLER_87_641 ();
 FILLCELL_X32 FILLER_87_673 ();
 FILLCELL_X32 FILLER_87_705 ();
 FILLCELL_X32 FILLER_87_737 ();
 FILLCELL_X32 FILLER_87_769 ();
 FILLCELL_X32 FILLER_87_801 ();
 FILLCELL_X32 FILLER_87_833 ();
 FILLCELL_X32 FILLER_87_865 ();
 FILLCELL_X32 FILLER_87_897 ();
 FILLCELL_X32 FILLER_87_929 ();
 FILLCELL_X32 FILLER_87_961 ();
 FILLCELL_X32 FILLER_87_993 ();
 FILLCELL_X32 FILLER_87_1025 ();
 FILLCELL_X32 FILLER_87_1057 ();
 FILLCELL_X32 FILLER_87_1089 ();
 FILLCELL_X32 FILLER_87_1121 ();
 FILLCELL_X32 FILLER_87_1153 ();
 FILLCELL_X32 FILLER_87_1185 ();
 FILLCELL_X32 FILLER_87_1217 ();
 FILLCELL_X8 FILLER_87_1249 ();
 FILLCELL_X4 FILLER_87_1257 ();
 FILLCELL_X2 FILLER_87_1261 ();
 FILLCELL_X32 FILLER_87_1264 ();
 FILLCELL_X32 FILLER_87_1296 ();
 FILLCELL_X32 FILLER_87_1328 ();
 FILLCELL_X32 FILLER_87_1360 ();
 FILLCELL_X32 FILLER_87_1392 ();
 FILLCELL_X32 FILLER_87_1424 ();
 FILLCELL_X32 FILLER_87_1456 ();
 FILLCELL_X32 FILLER_87_1488 ();
 FILLCELL_X32 FILLER_87_1520 ();
 FILLCELL_X32 FILLER_87_1552 ();
 FILLCELL_X32 FILLER_87_1584 ();
 FILLCELL_X32 FILLER_87_1616 ();
 FILLCELL_X32 FILLER_87_1648 ();
 FILLCELL_X32 FILLER_87_1680 ();
 FILLCELL_X32 FILLER_87_1712 ();
 FILLCELL_X32 FILLER_87_1744 ();
 FILLCELL_X32 FILLER_87_1776 ();
 FILLCELL_X32 FILLER_87_1808 ();
 FILLCELL_X32 FILLER_87_1840 ();
 FILLCELL_X32 FILLER_87_1872 ();
 FILLCELL_X32 FILLER_87_1904 ();
 FILLCELL_X32 FILLER_87_1936 ();
 FILLCELL_X32 FILLER_87_1968 ();
 FILLCELL_X32 FILLER_87_2000 ();
 FILLCELL_X32 FILLER_87_2032 ();
 FILLCELL_X32 FILLER_87_2064 ();
 FILLCELL_X32 FILLER_87_2096 ();
 FILLCELL_X32 FILLER_87_2128 ();
 FILLCELL_X32 FILLER_87_2160 ();
 FILLCELL_X32 FILLER_87_2192 ();
 FILLCELL_X32 FILLER_87_2224 ();
 FILLCELL_X32 FILLER_87_2256 ();
 FILLCELL_X32 FILLER_87_2288 ();
 FILLCELL_X32 FILLER_87_2320 ();
 FILLCELL_X32 FILLER_87_2352 ();
 FILLCELL_X32 FILLER_87_2384 ();
 FILLCELL_X32 FILLER_87_2416 ();
 FILLCELL_X32 FILLER_87_2448 ();
 FILLCELL_X32 FILLER_87_2480 ();
 FILLCELL_X8 FILLER_87_2512 ();
 FILLCELL_X4 FILLER_87_2520 ();
 FILLCELL_X2 FILLER_87_2524 ();
 FILLCELL_X32 FILLER_87_2527 ();
 FILLCELL_X32 FILLER_87_2559 ();
 FILLCELL_X32 FILLER_87_2591 ();
 FILLCELL_X32 FILLER_87_2623 ();
 FILLCELL_X32 FILLER_87_2655 ();
 FILLCELL_X32 FILLER_87_2687 ();
 FILLCELL_X32 FILLER_87_2719 ();
 FILLCELL_X32 FILLER_87_2751 ();
 FILLCELL_X32 FILLER_87_2783 ();
 FILLCELL_X32 FILLER_87_2815 ();
 FILLCELL_X32 FILLER_87_2847 ();
 FILLCELL_X32 FILLER_87_2879 ();
 FILLCELL_X32 FILLER_87_2911 ();
 FILLCELL_X32 FILLER_87_2943 ();
 FILLCELL_X32 FILLER_87_2975 ();
 FILLCELL_X32 FILLER_87_3007 ();
 FILLCELL_X32 FILLER_87_3039 ();
 FILLCELL_X32 FILLER_87_3071 ();
 FILLCELL_X32 FILLER_87_3103 ();
 FILLCELL_X32 FILLER_87_3135 ();
 FILLCELL_X32 FILLER_87_3167 ();
 FILLCELL_X32 FILLER_87_3199 ();
 FILLCELL_X32 FILLER_87_3231 ();
 FILLCELL_X32 FILLER_87_3263 ();
 FILLCELL_X32 FILLER_87_3295 ();
 FILLCELL_X32 FILLER_87_3327 ();
 FILLCELL_X32 FILLER_87_3359 ();
 FILLCELL_X32 FILLER_87_3391 ();
 FILLCELL_X32 FILLER_87_3423 ();
 FILLCELL_X32 FILLER_87_3455 ();
 FILLCELL_X32 FILLER_87_3487 ();
 FILLCELL_X32 FILLER_87_3519 ();
 FILLCELL_X32 FILLER_87_3551 ();
 FILLCELL_X32 FILLER_87_3583 ();
 FILLCELL_X32 FILLER_87_3615 ();
 FILLCELL_X32 FILLER_87_3647 ();
 FILLCELL_X32 FILLER_87_3679 ();
 FILLCELL_X16 FILLER_87_3711 ();
 FILLCELL_X8 FILLER_87_3727 ();
 FILLCELL_X2 FILLER_87_3735 ();
 FILLCELL_X1 FILLER_87_3737 ();
 FILLCELL_X32 FILLER_88_1 ();
 FILLCELL_X32 FILLER_88_33 ();
 FILLCELL_X32 FILLER_88_65 ();
 FILLCELL_X32 FILLER_88_97 ();
 FILLCELL_X32 FILLER_88_129 ();
 FILLCELL_X32 FILLER_88_161 ();
 FILLCELL_X32 FILLER_88_193 ();
 FILLCELL_X32 FILLER_88_225 ();
 FILLCELL_X32 FILLER_88_257 ();
 FILLCELL_X32 FILLER_88_289 ();
 FILLCELL_X32 FILLER_88_321 ();
 FILLCELL_X32 FILLER_88_353 ();
 FILLCELL_X32 FILLER_88_385 ();
 FILLCELL_X32 FILLER_88_417 ();
 FILLCELL_X32 FILLER_88_449 ();
 FILLCELL_X32 FILLER_88_481 ();
 FILLCELL_X32 FILLER_88_513 ();
 FILLCELL_X32 FILLER_88_545 ();
 FILLCELL_X32 FILLER_88_577 ();
 FILLCELL_X16 FILLER_88_609 ();
 FILLCELL_X4 FILLER_88_625 ();
 FILLCELL_X2 FILLER_88_629 ();
 FILLCELL_X32 FILLER_88_632 ();
 FILLCELL_X32 FILLER_88_664 ();
 FILLCELL_X32 FILLER_88_696 ();
 FILLCELL_X32 FILLER_88_728 ();
 FILLCELL_X32 FILLER_88_760 ();
 FILLCELL_X32 FILLER_88_792 ();
 FILLCELL_X32 FILLER_88_824 ();
 FILLCELL_X32 FILLER_88_856 ();
 FILLCELL_X32 FILLER_88_888 ();
 FILLCELL_X32 FILLER_88_920 ();
 FILLCELL_X32 FILLER_88_952 ();
 FILLCELL_X32 FILLER_88_984 ();
 FILLCELL_X32 FILLER_88_1016 ();
 FILLCELL_X32 FILLER_88_1048 ();
 FILLCELL_X32 FILLER_88_1080 ();
 FILLCELL_X32 FILLER_88_1112 ();
 FILLCELL_X32 FILLER_88_1144 ();
 FILLCELL_X32 FILLER_88_1176 ();
 FILLCELL_X32 FILLER_88_1208 ();
 FILLCELL_X32 FILLER_88_1240 ();
 FILLCELL_X32 FILLER_88_1272 ();
 FILLCELL_X32 FILLER_88_1304 ();
 FILLCELL_X32 FILLER_88_1336 ();
 FILLCELL_X32 FILLER_88_1368 ();
 FILLCELL_X32 FILLER_88_1400 ();
 FILLCELL_X32 FILLER_88_1432 ();
 FILLCELL_X32 FILLER_88_1464 ();
 FILLCELL_X32 FILLER_88_1496 ();
 FILLCELL_X32 FILLER_88_1528 ();
 FILLCELL_X32 FILLER_88_1560 ();
 FILLCELL_X32 FILLER_88_1592 ();
 FILLCELL_X32 FILLER_88_1624 ();
 FILLCELL_X32 FILLER_88_1656 ();
 FILLCELL_X32 FILLER_88_1688 ();
 FILLCELL_X32 FILLER_88_1720 ();
 FILLCELL_X32 FILLER_88_1752 ();
 FILLCELL_X32 FILLER_88_1784 ();
 FILLCELL_X32 FILLER_88_1816 ();
 FILLCELL_X32 FILLER_88_1848 ();
 FILLCELL_X8 FILLER_88_1880 ();
 FILLCELL_X4 FILLER_88_1888 ();
 FILLCELL_X2 FILLER_88_1892 ();
 FILLCELL_X32 FILLER_88_1895 ();
 FILLCELL_X32 FILLER_88_1927 ();
 FILLCELL_X32 FILLER_88_1959 ();
 FILLCELL_X32 FILLER_88_1991 ();
 FILLCELL_X32 FILLER_88_2023 ();
 FILLCELL_X32 FILLER_88_2055 ();
 FILLCELL_X32 FILLER_88_2087 ();
 FILLCELL_X32 FILLER_88_2119 ();
 FILLCELL_X32 FILLER_88_2151 ();
 FILLCELL_X32 FILLER_88_2183 ();
 FILLCELL_X32 FILLER_88_2215 ();
 FILLCELL_X32 FILLER_88_2247 ();
 FILLCELL_X32 FILLER_88_2279 ();
 FILLCELL_X32 FILLER_88_2311 ();
 FILLCELL_X32 FILLER_88_2343 ();
 FILLCELL_X32 FILLER_88_2375 ();
 FILLCELL_X32 FILLER_88_2407 ();
 FILLCELL_X32 FILLER_88_2439 ();
 FILLCELL_X32 FILLER_88_2471 ();
 FILLCELL_X32 FILLER_88_2503 ();
 FILLCELL_X32 FILLER_88_2535 ();
 FILLCELL_X32 FILLER_88_2567 ();
 FILLCELL_X32 FILLER_88_2599 ();
 FILLCELL_X32 FILLER_88_2631 ();
 FILLCELL_X32 FILLER_88_2663 ();
 FILLCELL_X32 FILLER_88_2695 ();
 FILLCELL_X32 FILLER_88_2727 ();
 FILLCELL_X32 FILLER_88_2759 ();
 FILLCELL_X32 FILLER_88_2791 ();
 FILLCELL_X32 FILLER_88_2823 ();
 FILLCELL_X32 FILLER_88_2855 ();
 FILLCELL_X32 FILLER_88_2887 ();
 FILLCELL_X32 FILLER_88_2919 ();
 FILLCELL_X32 FILLER_88_2951 ();
 FILLCELL_X32 FILLER_88_2983 ();
 FILLCELL_X32 FILLER_88_3015 ();
 FILLCELL_X32 FILLER_88_3047 ();
 FILLCELL_X32 FILLER_88_3079 ();
 FILLCELL_X32 FILLER_88_3111 ();
 FILLCELL_X8 FILLER_88_3143 ();
 FILLCELL_X4 FILLER_88_3151 ();
 FILLCELL_X2 FILLER_88_3155 ();
 FILLCELL_X32 FILLER_88_3158 ();
 FILLCELL_X32 FILLER_88_3190 ();
 FILLCELL_X32 FILLER_88_3222 ();
 FILLCELL_X32 FILLER_88_3254 ();
 FILLCELL_X32 FILLER_88_3286 ();
 FILLCELL_X32 FILLER_88_3318 ();
 FILLCELL_X32 FILLER_88_3350 ();
 FILLCELL_X32 FILLER_88_3382 ();
 FILLCELL_X32 FILLER_88_3414 ();
 FILLCELL_X32 FILLER_88_3446 ();
 FILLCELL_X32 FILLER_88_3478 ();
 FILLCELL_X32 FILLER_88_3510 ();
 FILLCELL_X32 FILLER_88_3542 ();
 FILLCELL_X32 FILLER_88_3574 ();
 FILLCELL_X32 FILLER_88_3606 ();
 FILLCELL_X32 FILLER_88_3638 ();
 FILLCELL_X32 FILLER_88_3670 ();
 FILLCELL_X32 FILLER_88_3702 ();
 FILLCELL_X4 FILLER_88_3734 ();
 FILLCELL_X32 FILLER_89_1 ();
 FILLCELL_X32 FILLER_89_33 ();
 FILLCELL_X32 FILLER_89_65 ();
 FILLCELL_X32 FILLER_89_97 ();
 FILLCELL_X32 FILLER_89_129 ();
 FILLCELL_X32 FILLER_89_161 ();
 FILLCELL_X32 FILLER_89_193 ();
 FILLCELL_X32 FILLER_89_225 ();
 FILLCELL_X32 FILLER_89_257 ();
 FILLCELL_X32 FILLER_89_289 ();
 FILLCELL_X32 FILLER_89_321 ();
 FILLCELL_X32 FILLER_89_353 ();
 FILLCELL_X32 FILLER_89_385 ();
 FILLCELL_X32 FILLER_89_417 ();
 FILLCELL_X32 FILLER_89_449 ();
 FILLCELL_X32 FILLER_89_481 ();
 FILLCELL_X32 FILLER_89_513 ();
 FILLCELL_X32 FILLER_89_545 ();
 FILLCELL_X32 FILLER_89_577 ();
 FILLCELL_X32 FILLER_89_609 ();
 FILLCELL_X32 FILLER_89_641 ();
 FILLCELL_X32 FILLER_89_673 ();
 FILLCELL_X32 FILLER_89_705 ();
 FILLCELL_X32 FILLER_89_737 ();
 FILLCELL_X32 FILLER_89_769 ();
 FILLCELL_X32 FILLER_89_801 ();
 FILLCELL_X32 FILLER_89_833 ();
 FILLCELL_X32 FILLER_89_865 ();
 FILLCELL_X32 FILLER_89_897 ();
 FILLCELL_X32 FILLER_89_929 ();
 FILLCELL_X32 FILLER_89_961 ();
 FILLCELL_X32 FILLER_89_993 ();
 FILLCELL_X32 FILLER_89_1025 ();
 FILLCELL_X32 FILLER_89_1057 ();
 FILLCELL_X32 FILLER_89_1089 ();
 FILLCELL_X32 FILLER_89_1121 ();
 FILLCELL_X32 FILLER_89_1153 ();
 FILLCELL_X32 FILLER_89_1185 ();
 FILLCELL_X32 FILLER_89_1217 ();
 FILLCELL_X8 FILLER_89_1249 ();
 FILLCELL_X4 FILLER_89_1257 ();
 FILLCELL_X2 FILLER_89_1261 ();
 FILLCELL_X32 FILLER_89_1264 ();
 FILLCELL_X32 FILLER_89_1296 ();
 FILLCELL_X32 FILLER_89_1328 ();
 FILLCELL_X32 FILLER_89_1360 ();
 FILLCELL_X32 FILLER_89_1392 ();
 FILLCELL_X32 FILLER_89_1424 ();
 FILLCELL_X32 FILLER_89_1456 ();
 FILLCELL_X32 FILLER_89_1488 ();
 FILLCELL_X32 FILLER_89_1520 ();
 FILLCELL_X32 FILLER_89_1552 ();
 FILLCELL_X32 FILLER_89_1584 ();
 FILLCELL_X32 FILLER_89_1616 ();
 FILLCELL_X32 FILLER_89_1648 ();
 FILLCELL_X32 FILLER_89_1680 ();
 FILLCELL_X32 FILLER_89_1712 ();
 FILLCELL_X32 FILLER_89_1744 ();
 FILLCELL_X32 FILLER_89_1776 ();
 FILLCELL_X32 FILLER_89_1808 ();
 FILLCELL_X32 FILLER_89_1840 ();
 FILLCELL_X32 FILLER_89_1872 ();
 FILLCELL_X32 FILLER_89_1904 ();
 FILLCELL_X32 FILLER_89_1936 ();
 FILLCELL_X32 FILLER_89_1968 ();
 FILLCELL_X32 FILLER_89_2000 ();
 FILLCELL_X32 FILLER_89_2032 ();
 FILLCELL_X32 FILLER_89_2064 ();
 FILLCELL_X32 FILLER_89_2096 ();
 FILLCELL_X32 FILLER_89_2128 ();
 FILLCELL_X32 FILLER_89_2160 ();
 FILLCELL_X32 FILLER_89_2192 ();
 FILLCELL_X32 FILLER_89_2224 ();
 FILLCELL_X32 FILLER_89_2256 ();
 FILLCELL_X32 FILLER_89_2288 ();
 FILLCELL_X32 FILLER_89_2320 ();
 FILLCELL_X32 FILLER_89_2352 ();
 FILLCELL_X32 FILLER_89_2384 ();
 FILLCELL_X32 FILLER_89_2416 ();
 FILLCELL_X32 FILLER_89_2448 ();
 FILLCELL_X32 FILLER_89_2480 ();
 FILLCELL_X8 FILLER_89_2512 ();
 FILLCELL_X4 FILLER_89_2520 ();
 FILLCELL_X2 FILLER_89_2524 ();
 FILLCELL_X32 FILLER_89_2527 ();
 FILLCELL_X32 FILLER_89_2559 ();
 FILLCELL_X32 FILLER_89_2591 ();
 FILLCELL_X32 FILLER_89_2623 ();
 FILLCELL_X32 FILLER_89_2655 ();
 FILLCELL_X32 FILLER_89_2687 ();
 FILLCELL_X32 FILLER_89_2719 ();
 FILLCELL_X32 FILLER_89_2751 ();
 FILLCELL_X32 FILLER_89_2783 ();
 FILLCELL_X32 FILLER_89_2815 ();
 FILLCELL_X32 FILLER_89_2847 ();
 FILLCELL_X32 FILLER_89_2879 ();
 FILLCELL_X32 FILLER_89_2911 ();
 FILLCELL_X32 FILLER_89_2943 ();
 FILLCELL_X32 FILLER_89_2975 ();
 FILLCELL_X32 FILLER_89_3007 ();
 FILLCELL_X32 FILLER_89_3039 ();
 FILLCELL_X32 FILLER_89_3071 ();
 FILLCELL_X32 FILLER_89_3103 ();
 FILLCELL_X32 FILLER_89_3135 ();
 FILLCELL_X32 FILLER_89_3167 ();
 FILLCELL_X32 FILLER_89_3199 ();
 FILLCELL_X32 FILLER_89_3231 ();
 FILLCELL_X32 FILLER_89_3263 ();
 FILLCELL_X32 FILLER_89_3295 ();
 FILLCELL_X32 FILLER_89_3327 ();
 FILLCELL_X32 FILLER_89_3359 ();
 FILLCELL_X32 FILLER_89_3391 ();
 FILLCELL_X32 FILLER_89_3423 ();
 FILLCELL_X32 FILLER_89_3455 ();
 FILLCELL_X32 FILLER_89_3487 ();
 FILLCELL_X32 FILLER_89_3519 ();
 FILLCELL_X32 FILLER_89_3551 ();
 FILLCELL_X32 FILLER_89_3583 ();
 FILLCELL_X32 FILLER_89_3615 ();
 FILLCELL_X32 FILLER_89_3647 ();
 FILLCELL_X32 FILLER_89_3679 ();
 FILLCELL_X16 FILLER_89_3711 ();
 FILLCELL_X8 FILLER_89_3727 ();
 FILLCELL_X2 FILLER_89_3735 ();
 FILLCELL_X1 FILLER_89_3737 ();
 FILLCELL_X32 FILLER_90_1 ();
 FILLCELL_X32 FILLER_90_33 ();
 FILLCELL_X32 FILLER_90_65 ();
 FILLCELL_X32 FILLER_90_97 ();
 FILLCELL_X32 FILLER_90_129 ();
 FILLCELL_X32 FILLER_90_161 ();
 FILLCELL_X32 FILLER_90_193 ();
 FILLCELL_X32 FILLER_90_225 ();
 FILLCELL_X32 FILLER_90_257 ();
 FILLCELL_X32 FILLER_90_289 ();
 FILLCELL_X32 FILLER_90_321 ();
 FILLCELL_X32 FILLER_90_353 ();
 FILLCELL_X32 FILLER_90_385 ();
 FILLCELL_X32 FILLER_90_417 ();
 FILLCELL_X32 FILLER_90_449 ();
 FILLCELL_X32 FILLER_90_481 ();
 FILLCELL_X32 FILLER_90_513 ();
 FILLCELL_X32 FILLER_90_545 ();
 FILLCELL_X32 FILLER_90_577 ();
 FILLCELL_X16 FILLER_90_609 ();
 FILLCELL_X4 FILLER_90_625 ();
 FILLCELL_X2 FILLER_90_629 ();
 FILLCELL_X32 FILLER_90_632 ();
 FILLCELL_X32 FILLER_90_664 ();
 FILLCELL_X32 FILLER_90_696 ();
 FILLCELL_X32 FILLER_90_728 ();
 FILLCELL_X32 FILLER_90_760 ();
 FILLCELL_X32 FILLER_90_792 ();
 FILLCELL_X32 FILLER_90_824 ();
 FILLCELL_X32 FILLER_90_856 ();
 FILLCELL_X32 FILLER_90_888 ();
 FILLCELL_X32 FILLER_90_920 ();
 FILLCELL_X32 FILLER_90_952 ();
 FILLCELL_X32 FILLER_90_984 ();
 FILLCELL_X32 FILLER_90_1016 ();
 FILLCELL_X32 FILLER_90_1048 ();
 FILLCELL_X32 FILLER_90_1080 ();
 FILLCELL_X32 FILLER_90_1112 ();
 FILLCELL_X32 FILLER_90_1144 ();
 FILLCELL_X32 FILLER_90_1176 ();
 FILLCELL_X32 FILLER_90_1208 ();
 FILLCELL_X32 FILLER_90_1240 ();
 FILLCELL_X32 FILLER_90_1272 ();
 FILLCELL_X32 FILLER_90_1304 ();
 FILLCELL_X32 FILLER_90_1336 ();
 FILLCELL_X32 FILLER_90_1368 ();
 FILLCELL_X32 FILLER_90_1400 ();
 FILLCELL_X32 FILLER_90_1432 ();
 FILLCELL_X32 FILLER_90_1464 ();
 FILLCELL_X32 FILLER_90_1496 ();
 FILLCELL_X32 FILLER_90_1528 ();
 FILLCELL_X32 FILLER_90_1560 ();
 FILLCELL_X32 FILLER_90_1592 ();
 FILLCELL_X32 FILLER_90_1624 ();
 FILLCELL_X32 FILLER_90_1656 ();
 FILLCELL_X32 FILLER_90_1688 ();
 FILLCELL_X32 FILLER_90_1720 ();
 FILLCELL_X32 FILLER_90_1752 ();
 FILLCELL_X32 FILLER_90_1784 ();
 FILLCELL_X32 FILLER_90_1816 ();
 FILLCELL_X32 FILLER_90_1848 ();
 FILLCELL_X8 FILLER_90_1880 ();
 FILLCELL_X4 FILLER_90_1888 ();
 FILLCELL_X2 FILLER_90_1892 ();
 FILLCELL_X32 FILLER_90_1895 ();
 FILLCELL_X32 FILLER_90_1927 ();
 FILLCELL_X32 FILLER_90_1959 ();
 FILLCELL_X32 FILLER_90_1991 ();
 FILLCELL_X32 FILLER_90_2023 ();
 FILLCELL_X32 FILLER_90_2055 ();
 FILLCELL_X32 FILLER_90_2087 ();
 FILLCELL_X32 FILLER_90_2119 ();
 FILLCELL_X32 FILLER_90_2151 ();
 FILLCELL_X32 FILLER_90_2183 ();
 FILLCELL_X32 FILLER_90_2215 ();
 FILLCELL_X32 FILLER_90_2247 ();
 FILLCELL_X32 FILLER_90_2279 ();
 FILLCELL_X32 FILLER_90_2311 ();
 FILLCELL_X32 FILLER_90_2343 ();
 FILLCELL_X32 FILLER_90_2375 ();
 FILLCELL_X32 FILLER_90_2407 ();
 FILLCELL_X32 FILLER_90_2439 ();
 FILLCELL_X32 FILLER_90_2471 ();
 FILLCELL_X32 FILLER_90_2503 ();
 FILLCELL_X32 FILLER_90_2535 ();
 FILLCELL_X32 FILLER_90_2567 ();
 FILLCELL_X32 FILLER_90_2599 ();
 FILLCELL_X32 FILLER_90_2631 ();
 FILLCELL_X32 FILLER_90_2663 ();
 FILLCELL_X32 FILLER_90_2695 ();
 FILLCELL_X32 FILLER_90_2727 ();
 FILLCELL_X32 FILLER_90_2759 ();
 FILLCELL_X32 FILLER_90_2791 ();
 FILLCELL_X32 FILLER_90_2823 ();
 FILLCELL_X32 FILLER_90_2855 ();
 FILLCELL_X32 FILLER_90_2887 ();
 FILLCELL_X32 FILLER_90_2919 ();
 FILLCELL_X32 FILLER_90_2951 ();
 FILLCELL_X32 FILLER_90_2983 ();
 FILLCELL_X32 FILLER_90_3015 ();
 FILLCELL_X32 FILLER_90_3047 ();
 FILLCELL_X32 FILLER_90_3079 ();
 FILLCELL_X32 FILLER_90_3111 ();
 FILLCELL_X8 FILLER_90_3143 ();
 FILLCELL_X4 FILLER_90_3151 ();
 FILLCELL_X2 FILLER_90_3155 ();
 FILLCELL_X32 FILLER_90_3158 ();
 FILLCELL_X32 FILLER_90_3190 ();
 FILLCELL_X32 FILLER_90_3222 ();
 FILLCELL_X32 FILLER_90_3254 ();
 FILLCELL_X32 FILLER_90_3286 ();
 FILLCELL_X32 FILLER_90_3318 ();
 FILLCELL_X32 FILLER_90_3350 ();
 FILLCELL_X32 FILLER_90_3382 ();
 FILLCELL_X32 FILLER_90_3414 ();
 FILLCELL_X32 FILLER_90_3446 ();
 FILLCELL_X32 FILLER_90_3478 ();
 FILLCELL_X32 FILLER_90_3510 ();
 FILLCELL_X32 FILLER_90_3542 ();
 FILLCELL_X32 FILLER_90_3574 ();
 FILLCELL_X32 FILLER_90_3606 ();
 FILLCELL_X32 FILLER_90_3638 ();
 FILLCELL_X32 FILLER_90_3670 ();
 FILLCELL_X32 FILLER_90_3702 ();
 FILLCELL_X4 FILLER_90_3734 ();
 FILLCELL_X32 FILLER_91_1 ();
 FILLCELL_X32 FILLER_91_33 ();
 FILLCELL_X32 FILLER_91_65 ();
 FILLCELL_X32 FILLER_91_97 ();
 FILLCELL_X32 FILLER_91_129 ();
 FILLCELL_X32 FILLER_91_161 ();
 FILLCELL_X32 FILLER_91_193 ();
 FILLCELL_X32 FILLER_91_225 ();
 FILLCELL_X32 FILLER_91_257 ();
 FILLCELL_X32 FILLER_91_289 ();
 FILLCELL_X32 FILLER_91_321 ();
 FILLCELL_X32 FILLER_91_353 ();
 FILLCELL_X32 FILLER_91_385 ();
 FILLCELL_X32 FILLER_91_417 ();
 FILLCELL_X32 FILLER_91_449 ();
 FILLCELL_X32 FILLER_91_481 ();
 FILLCELL_X32 FILLER_91_513 ();
 FILLCELL_X32 FILLER_91_545 ();
 FILLCELL_X32 FILLER_91_577 ();
 FILLCELL_X32 FILLER_91_609 ();
 FILLCELL_X32 FILLER_91_641 ();
 FILLCELL_X32 FILLER_91_673 ();
 FILLCELL_X32 FILLER_91_705 ();
 FILLCELL_X32 FILLER_91_737 ();
 FILLCELL_X32 FILLER_91_769 ();
 FILLCELL_X32 FILLER_91_801 ();
 FILLCELL_X32 FILLER_91_833 ();
 FILLCELL_X32 FILLER_91_865 ();
 FILLCELL_X32 FILLER_91_897 ();
 FILLCELL_X32 FILLER_91_929 ();
 FILLCELL_X32 FILLER_91_961 ();
 FILLCELL_X32 FILLER_91_993 ();
 FILLCELL_X32 FILLER_91_1025 ();
 FILLCELL_X32 FILLER_91_1057 ();
 FILLCELL_X32 FILLER_91_1089 ();
 FILLCELL_X32 FILLER_91_1121 ();
 FILLCELL_X32 FILLER_91_1153 ();
 FILLCELL_X32 FILLER_91_1185 ();
 FILLCELL_X32 FILLER_91_1217 ();
 FILLCELL_X8 FILLER_91_1249 ();
 FILLCELL_X4 FILLER_91_1257 ();
 FILLCELL_X2 FILLER_91_1261 ();
 FILLCELL_X32 FILLER_91_1264 ();
 FILLCELL_X32 FILLER_91_1296 ();
 FILLCELL_X32 FILLER_91_1328 ();
 FILLCELL_X32 FILLER_91_1360 ();
 FILLCELL_X32 FILLER_91_1392 ();
 FILLCELL_X32 FILLER_91_1424 ();
 FILLCELL_X32 FILLER_91_1456 ();
 FILLCELL_X32 FILLER_91_1488 ();
 FILLCELL_X32 FILLER_91_1520 ();
 FILLCELL_X32 FILLER_91_1552 ();
 FILLCELL_X32 FILLER_91_1584 ();
 FILLCELL_X32 FILLER_91_1616 ();
 FILLCELL_X32 FILLER_91_1648 ();
 FILLCELL_X32 FILLER_91_1680 ();
 FILLCELL_X32 FILLER_91_1712 ();
 FILLCELL_X32 FILLER_91_1744 ();
 FILLCELL_X32 FILLER_91_1776 ();
 FILLCELL_X32 FILLER_91_1808 ();
 FILLCELL_X32 FILLER_91_1840 ();
 FILLCELL_X32 FILLER_91_1872 ();
 FILLCELL_X32 FILLER_91_1904 ();
 FILLCELL_X32 FILLER_91_1936 ();
 FILLCELL_X32 FILLER_91_1968 ();
 FILLCELL_X32 FILLER_91_2000 ();
 FILLCELL_X32 FILLER_91_2032 ();
 FILLCELL_X32 FILLER_91_2064 ();
 FILLCELL_X32 FILLER_91_2096 ();
 FILLCELL_X32 FILLER_91_2128 ();
 FILLCELL_X32 FILLER_91_2160 ();
 FILLCELL_X32 FILLER_91_2192 ();
 FILLCELL_X32 FILLER_91_2224 ();
 FILLCELL_X32 FILLER_91_2256 ();
 FILLCELL_X32 FILLER_91_2288 ();
 FILLCELL_X32 FILLER_91_2320 ();
 FILLCELL_X32 FILLER_91_2352 ();
 FILLCELL_X32 FILLER_91_2384 ();
 FILLCELL_X32 FILLER_91_2416 ();
 FILLCELL_X32 FILLER_91_2448 ();
 FILLCELL_X32 FILLER_91_2480 ();
 FILLCELL_X8 FILLER_91_2512 ();
 FILLCELL_X4 FILLER_91_2520 ();
 FILLCELL_X2 FILLER_91_2524 ();
 FILLCELL_X32 FILLER_91_2527 ();
 FILLCELL_X32 FILLER_91_2559 ();
 FILLCELL_X32 FILLER_91_2591 ();
 FILLCELL_X32 FILLER_91_2623 ();
 FILLCELL_X32 FILLER_91_2655 ();
 FILLCELL_X32 FILLER_91_2687 ();
 FILLCELL_X32 FILLER_91_2719 ();
 FILLCELL_X32 FILLER_91_2751 ();
 FILLCELL_X32 FILLER_91_2783 ();
 FILLCELL_X32 FILLER_91_2815 ();
 FILLCELL_X32 FILLER_91_2847 ();
 FILLCELL_X32 FILLER_91_2879 ();
 FILLCELL_X32 FILLER_91_2911 ();
 FILLCELL_X32 FILLER_91_2943 ();
 FILLCELL_X32 FILLER_91_2975 ();
 FILLCELL_X32 FILLER_91_3007 ();
 FILLCELL_X32 FILLER_91_3039 ();
 FILLCELL_X32 FILLER_91_3071 ();
 FILLCELL_X32 FILLER_91_3103 ();
 FILLCELL_X32 FILLER_91_3135 ();
 FILLCELL_X32 FILLER_91_3167 ();
 FILLCELL_X32 FILLER_91_3199 ();
 FILLCELL_X32 FILLER_91_3231 ();
 FILLCELL_X32 FILLER_91_3263 ();
 FILLCELL_X32 FILLER_91_3295 ();
 FILLCELL_X32 FILLER_91_3327 ();
 FILLCELL_X32 FILLER_91_3359 ();
 FILLCELL_X32 FILLER_91_3391 ();
 FILLCELL_X32 FILLER_91_3423 ();
 FILLCELL_X32 FILLER_91_3455 ();
 FILLCELL_X32 FILLER_91_3487 ();
 FILLCELL_X32 FILLER_91_3519 ();
 FILLCELL_X32 FILLER_91_3551 ();
 FILLCELL_X32 FILLER_91_3583 ();
 FILLCELL_X32 FILLER_91_3615 ();
 FILLCELL_X32 FILLER_91_3647 ();
 FILLCELL_X32 FILLER_91_3679 ();
 FILLCELL_X16 FILLER_91_3711 ();
 FILLCELL_X8 FILLER_91_3727 ();
 FILLCELL_X2 FILLER_91_3735 ();
 FILLCELL_X1 FILLER_91_3737 ();
 FILLCELL_X32 FILLER_92_1 ();
 FILLCELL_X32 FILLER_92_33 ();
 FILLCELL_X32 FILLER_92_65 ();
 FILLCELL_X32 FILLER_92_97 ();
 FILLCELL_X32 FILLER_92_129 ();
 FILLCELL_X32 FILLER_92_161 ();
 FILLCELL_X32 FILLER_92_193 ();
 FILLCELL_X32 FILLER_92_225 ();
 FILLCELL_X32 FILLER_92_257 ();
 FILLCELL_X32 FILLER_92_289 ();
 FILLCELL_X32 FILLER_92_321 ();
 FILLCELL_X32 FILLER_92_353 ();
 FILLCELL_X32 FILLER_92_385 ();
 FILLCELL_X32 FILLER_92_417 ();
 FILLCELL_X32 FILLER_92_449 ();
 FILLCELL_X32 FILLER_92_481 ();
 FILLCELL_X32 FILLER_92_513 ();
 FILLCELL_X32 FILLER_92_545 ();
 FILLCELL_X32 FILLER_92_577 ();
 FILLCELL_X16 FILLER_92_609 ();
 FILLCELL_X4 FILLER_92_625 ();
 FILLCELL_X2 FILLER_92_629 ();
 FILLCELL_X32 FILLER_92_632 ();
 FILLCELL_X32 FILLER_92_664 ();
 FILLCELL_X32 FILLER_92_696 ();
 FILLCELL_X32 FILLER_92_728 ();
 FILLCELL_X32 FILLER_92_760 ();
 FILLCELL_X32 FILLER_92_792 ();
 FILLCELL_X32 FILLER_92_824 ();
 FILLCELL_X32 FILLER_92_856 ();
 FILLCELL_X32 FILLER_92_888 ();
 FILLCELL_X32 FILLER_92_920 ();
 FILLCELL_X32 FILLER_92_952 ();
 FILLCELL_X32 FILLER_92_984 ();
 FILLCELL_X32 FILLER_92_1016 ();
 FILLCELL_X32 FILLER_92_1048 ();
 FILLCELL_X32 FILLER_92_1080 ();
 FILLCELL_X32 FILLER_92_1112 ();
 FILLCELL_X32 FILLER_92_1144 ();
 FILLCELL_X32 FILLER_92_1176 ();
 FILLCELL_X32 FILLER_92_1208 ();
 FILLCELL_X32 FILLER_92_1240 ();
 FILLCELL_X32 FILLER_92_1272 ();
 FILLCELL_X32 FILLER_92_1304 ();
 FILLCELL_X32 FILLER_92_1336 ();
 FILLCELL_X32 FILLER_92_1368 ();
 FILLCELL_X32 FILLER_92_1400 ();
 FILLCELL_X32 FILLER_92_1432 ();
 FILLCELL_X32 FILLER_92_1464 ();
 FILLCELL_X32 FILLER_92_1496 ();
 FILLCELL_X32 FILLER_92_1528 ();
 FILLCELL_X32 FILLER_92_1560 ();
 FILLCELL_X32 FILLER_92_1592 ();
 FILLCELL_X32 FILLER_92_1624 ();
 FILLCELL_X32 FILLER_92_1656 ();
 FILLCELL_X32 FILLER_92_1688 ();
 FILLCELL_X32 FILLER_92_1720 ();
 FILLCELL_X32 FILLER_92_1752 ();
 FILLCELL_X32 FILLER_92_1784 ();
 FILLCELL_X32 FILLER_92_1816 ();
 FILLCELL_X32 FILLER_92_1848 ();
 FILLCELL_X8 FILLER_92_1880 ();
 FILLCELL_X4 FILLER_92_1888 ();
 FILLCELL_X2 FILLER_92_1892 ();
 FILLCELL_X32 FILLER_92_1895 ();
 FILLCELL_X32 FILLER_92_1927 ();
 FILLCELL_X32 FILLER_92_1959 ();
 FILLCELL_X32 FILLER_92_1991 ();
 FILLCELL_X32 FILLER_92_2023 ();
 FILLCELL_X32 FILLER_92_2055 ();
 FILLCELL_X32 FILLER_92_2087 ();
 FILLCELL_X32 FILLER_92_2119 ();
 FILLCELL_X32 FILLER_92_2151 ();
 FILLCELL_X32 FILLER_92_2183 ();
 FILLCELL_X32 FILLER_92_2215 ();
 FILLCELL_X32 FILLER_92_2247 ();
 FILLCELL_X32 FILLER_92_2279 ();
 FILLCELL_X32 FILLER_92_2311 ();
 FILLCELL_X32 FILLER_92_2343 ();
 FILLCELL_X32 FILLER_92_2375 ();
 FILLCELL_X32 FILLER_92_2407 ();
 FILLCELL_X32 FILLER_92_2439 ();
 FILLCELL_X32 FILLER_92_2471 ();
 FILLCELL_X32 FILLER_92_2503 ();
 FILLCELL_X32 FILLER_92_2535 ();
 FILLCELL_X32 FILLER_92_2567 ();
 FILLCELL_X32 FILLER_92_2599 ();
 FILLCELL_X32 FILLER_92_2631 ();
 FILLCELL_X32 FILLER_92_2663 ();
 FILLCELL_X32 FILLER_92_2695 ();
 FILLCELL_X32 FILLER_92_2727 ();
 FILLCELL_X32 FILLER_92_2759 ();
 FILLCELL_X32 FILLER_92_2791 ();
 FILLCELL_X32 FILLER_92_2823 ();
 FILLCELL_X32 FILLER_92_2855 ();
 FILLCELL_X32 FILLER_92_2887 ();
 FILLCELL_X32 FILLER_92_2919 ();
 FILLCELL_X32 FILLER_92_2951 ();
 FILLCELL_X32 FILLER_92_2983 ();
 FILLCELL_X32 FILLER_92_3015 ();
 FILLCELL_X32 FILLER_92_3047 ();
 FILLCELL_X32 FILLER_92_3079 ();
 FILLCELL_X32 FILLER_92_3111 ();
 FILLCELL_X8 FILLER_92_3143 ();
 FILLCELL_X4 FILLER_92_3151 ();
 FILLCELL_X2 FILLER_92_3155 ();
 FILLCELL_X32 FILLER_92_3158 ();
 FILLCELL_X32 FILLER_92_3190 ();
 FILLCELL_X32 FILLER_92_3222 ();
 FILLCELL_X32 FILLER_92_3254 ();
 FILLCELL_X32 FILLER_92_3286 ();
 FILLCELL_X32 FILLER_92_3318 ();
 FILLCELL_X32 FILLER_92_3350 ();
 FILLCELL_X32 FILLER_92_3382 ();
 FILLCELL_X32 FILLER_92_3414 ();
 FILLCELL_X32 FILLER_92_3446 ();
 FILLCELL_X32 FILLER_92_3478 ();
 FILLCELL_X32 FILLER_92_3510 ();
 FILLCELL_X32 FILLER_92_3542 ();
 FILLCELL_X32 FILLER_92_3574 ();
 FILLCELL_X32 FILLER_92_3606 ();
 FILLCELL_X32 FILLER_92_3638 ();
 FILLCELL_X32 FILLER_92_3670 ();
 FILLCELL_X32 FILLER_92_3702 ();
 FILLCELL_X4 FILLER_92_3734 ();
 FILLCELL_X32 FILLER_93_1 ();
 FILLCELL_X32 FILLER_93_33 ();
 FILLCELL_X32 FILLER_93_65 ();
 FILLCELL_X32 FILLER_93_97 ();
 FILLCELL_X32 FILLER_93_129 ();
 FILLCELL_X32 FILLER_93_161 ();
 FILLCELL_X32 FILLER_93_193 ();
 FILLCELL_X32 FILLER_93_225 ();
 FILLCELL_X32 FILLER_93_257 ();
 FILLCELL_X32 FILLER_93_289 ();
 FILLCELL_X32 FILLER_93_321 ();
 FILLCELL_X32 FILLER_93_353 ();
 FILLCELL_X32 FILLER_93_385 ();
 FILLCELL_X32 FILLER_93_417 ();
 FILLCELL_X32 FILLER_93_449 ();
 FILLCELL_X32 FILLER_93_481 ();
 FILLCELL_X32 FILLER_93_513 ();
 FILLCELL_X32 FILLER_93_545 ();
 FILLCELL_X32 FILLER_93_577 ();
 FILLCELL_X32 FILLER_93_609 ();
 FILLCELL_X32 FILLER_93_641 ();
 FILLCELL_X32 FILLER_93_673 ();
 FILLCELL_X32 FILLER_93_705 ();
 FILLCELL_X32 FILLER_93_737 ();
 FILLCELL_X32 FILLER_93_769 ();
 FILLCELL_X32 FILLER_93_801 ();
 FILLCELL_X32 FILLER_93_833 ();
 FILLCELL_X32 FILLER_93_865 ();
 FILLCELL_X32 FILLER_93_897 ();
 FILLCELL_X32 FILLER_93_929 ();
 FILLCELL_X32 FILLER_93_961 ();
 FILLCELL_X32 FILLER_93_993 ();
 FILLCELL_X32 FILLER_93_1025 ();
 FILLCELL_X32 FILLER_93_1057 ();
 FILLCELL_X32 FILLER_93_1089 ();
 FILLCELL_X32 FILLER_93_1121 ();
 FILLCELL_X32 FILLER_93_1153 ();
 FILLCELL_X32 FILLER_93_1185 ();
 FILLCELL_X32 FILLER_93_1217 ();
 FILLCELL_X8 FILLER_93_1249 ();
 FILLCELL_X4 FILLER_93_1257 ();
 FILLCELL_X2 FILLER_93_1261 ();
 FILLCELL_X32 FILLER_93_1264 ();
 FILLCELL_X32 FILLER_93_1296 ();
 FILLCELL_X32 FILLER_93_1328 ();
 FILLCELL_X32 FILLER_93_1360 ();
 FILLCELL_X32 FILLER_93_1392 ();
 FILLCELL_X32 FILLER_93_1424 ();
 FILLCELL_X32 FILLER_93_1456 ();
 FILLCELL_X32 FILLER_93_1488 ();
 FILLCELL_X32 FILLER_93_1520 ();
 FILLCELL_X32 FILLER_93_1552 ();
 FILLCELL_X32 FILLER_93_1584 ();
 FILLCELL_X32 FILLER_93_1616 ();
 FILLCELL_X32 FILLER_93_1648 ();
 FILLCELL_X32 FILLER_93_1680 ();
 FILLCELL_X32 FILLER_93_1712 ();
 FILLCELL_X32 FILLER_93_1744 ();
 FILLCELL_X32 FILLER_93_1776 ();
 FILLCELL_X32 FILLER_93_1808 ();
 FILLCELL_X32 FILLER_93_1840 ();
 FILLCELL_X32 FILLER_93_1872 ();
 FILLCELL_X32 FILLER_93_1904 ();
 FILLCELL_X32 FILLER_93_1936 ();
 FILLCELL_X32 FILLER_93_1968 ();
 FILLCELL_X32 FILLER_93_2000 ();
 FILLCELL_X32 FILLER_93_2032 ();
 FILLCELL_X32 FILLER_93_2064 ();
 FILLCELL_X32 FILLER_93_2096 ();
 FILLCELL_X32 FILLER_93_2128 ();
 FILLCELL_X32 FILLER_93_2160 ();
 FILLCELL_X32 FILLER_93_2192 ();
 FILLCELL_X32 FILLER_93_2224 ();
 FILLCELL_X32 FILLER_93_2256 ();
 FILLCELL_X32 FILLER_93_2288 ();
 FILLCELL_X32 FILLER_93_2320 ();
 FILLCELL_X32 FILLER_93_2352 ();
 FILLCELL_X32 FILLER_93_2384 ();
 FILLCELL_X32 FILLER_93_2416 ();
 FILLCELL_X32 FILLER_93_2448 ();
 FILLCELL_X32 FILLER_93_2480 ();
 FILLCELL_X8 FILLER_93_2512 ();
 FILLCELL_X4 FILLER_93_2520 ();
 FILLCELL_X2 FILLER_93_2524 ();
 FILLCELL_X32 FILLER_93_2527 ();
 FILLCELL_X32 FILLER_93_2559 ();
 FILLCELL_X32 FILLER_93_2591 ();
 FILLCELL_X32 FILLER_93_2623 ();
 FILLCELL_X32 FILLER_93_2655 ();
 FILLCELL_X32 FILLER_93_2687 ();
 FILLCELL_X32 FILLER_93_2719 ();
 FILLCELL_X32 FILLER_93_2751 ();
 FILLCELL_X32 FILLER_93_2783 ();
 FILLCELL_X32 FILLER_93_2815 ();
 FILLCELL_X32 FILLER_93_2847 ();
 FILLCELL_X32 FILLER_93_2879 ();
 FILLCELL_X32 FILLER_93_2911 ();
 FILLCELL_X32 FILLER_93_2943 ();
 FILLCELL_X32 FILLER_93_2975 ();
 FILLCELL_X32 FILLER_93_3007 ();
 FILLCELL_X32 FILLER_93_3039 ();
 FILLCELL_X32 FILLER_93_3071 ();
 FILLCELL_X32 FILLER_93_3103 ();
 FILLCELL_X32 FILLER_93_3135 ();
 FILLCELL_X32 FILLER_93_3167 ();
 FILLCELL_X32 FILLER_93_3199 ();
 FILLCELL_X32 FILLER_93_3231 ();
 FILLCELL_X32 FILLER_93_3263 ();
 FILLCELL_X32 FILLER_93_3295 ();
 FILLCELL_X32 FILLER_93_3327 ();
 FILLCELL_X32 FILLER_93_3359 ();
 FILLCELL_X32 FILLER_93_3391 ();
 FILLCELL_X32 FILLER_93_3423 ();
 FILLCELL_X32 FILLER_93_3455 ();
 FILLCELL_X32 FILLER_93_3487 ();
 FILLCELL_X32 FILLER_93_3519 ();
 FILLCELL_X32 FILLER_93_3551 ();
 FILLCELL_X32 FILLER_93_3583 ();
 FILLCELL_X32 FILLER_93_3615 ();
 FILLCELL_X32 FILLER_93_3647 ();
 FILLCELL_X32 FILLER_93_3679 ();
 FILLCELL_X16 FILLER_93_3711 ();
 FILLCELL_X8 FILLER_93_3727 ();
 FILLCELL_X2 FILLER_93_3735 ();
 FILLCELL_X1 FILLER_93_3737 ();
 FILLCELL_X32 FILLER_94_1 ();
 FILLCELL_X32 FILLER_94_33 ();
 FILLCELL_X32 FILLER_94_65 ();
 FILLCELL_X32 FILLER_94_97 ();
 FILLCELL_X32 FILLER_94_129 ();
 FILLCELL_X32 FILLER_94_161 ();
 FILLCELL_X32 FILLER_94_193 ();
 FILLCELL_X32 FILLER_94_225 ();
 FILLCELL_X32 FILLER_94_257 ();
 FILLCELL_X32 FILLER_94_289 ();
 FILLCELL_X32 FILLER_94_321 ();
 FILLCELL_X32 FILLER_94_353 ();
 FILLCELL_X32 FILLER_94_385 ();
 FILLCELL_X32 FILLER_94_417 ();
 FILLCELL_X32 FILLER_94_449 ();
 FILLCELL_X32 FILLER_94_481 ();
 FILLCELL_X32 FILLER_94_513 ();
 FILLCELL_X32 FILLER_94_545 ();
 FILLCELL_X32 FILLER_94_577 ();
 FILLCELL_X16 FILLER_94_609 ();
 FILLCELL_X4 FILLER_94_625 ();
 FILLCELL_X2 FILLER_94_629 ();
 FILLCELL_X32 FILLER_94_632 ();
 FILLCELL_X32 FILLER_94_664 ();
 FILLCELL_X32 FILLER_94_696 ();
 FILLCELL_X32 FILLER_94_728 ();
 FILLCELL_X32 FILLER_94_760 ();
 FILLCELL_X32 FILLER_94_792 ();
 FILLCELL_X32 FILLER_94_824 ();
 FILLCELL_X32 FILLER_94_856 ();
 FILLCELL_X32 FILLER_94_888 ();
 FILLCELL_X32 FILLER_94_920 ();
 FILLCELL_X32 FILLER_94_952 ();
 FILLCELL_X32 FILLER_94_984 ();
 FILLCELL_X32 FILLER_94_1016 ();
 FILLCELL_X32 FILLER_94_1048 ();
 FILLCELL_X32 FILLER_94_1080 ();
 FILLCELL_X32 FILLER_94_1112 ();
 FILLCELL_X32 FILLER_94_1144 ();
 FILLCELL_X32 FILLER_94_1176 ();
 FILLCELL_X32 FILLER_94_1208 ();
 FILLCELL_X32 FILLER_94_1240 ();
 FILLCELL_X32 FILLER_94_1272 ();
 FILLCELL_X32 FILLER_94_1304 ();
 FILLCELL_X32 FILLER_94_1336 ();
 FILLCELL_X32 FILLER_94_1368 ();
 FILLCELL_X32 FILLER_94_1400 ();
 FILLCELL_X32 FILLER_94_1432 ();
 FILLCELL_X32 FILLER_94_1464 ();
 FILLCELL_X32 FILLER_94_1496 ();
 FILLCELL_X32 FILLER_94_1528 ();
 FILLCELL_X32 FILLER_94_1560 ();
 FILLCELL_X32 FILLER_94_1592 ();
 FILLCELL_X32 FILLER_94_1624 ();
 FILLCELL_X32 FILLER_94_1656 ();
 FILLCELL_X32 FILLER_94_1688 ();
 FILLCELL_X32 FILLER_94_1720 ();
 FILLCELL_X32 FILLER_94_1752 ();
 FILLCELL_X32 FILLER_94_1784 ();
 FILLCELL_X32 FILLER_94_1816 ();
 FILLCELL_X32 FILLER_94_1848 ();
 FILLCELL_X8 FILLER_94_1880 ();
 FILLCELL_X4 FILLER_94_1888 ();
 FILLCELL_X2 FILLER_94_1892 ();
 FILLCELL_X32 FILLER_94_1895 ();
 FILLCELL_X32 FILLER_94_1927 ();
 FILLCELL_X32 FILLER_94_1959 ();
 FILLCELL_X32 FILLER_94_1991 ();
 FILLCELL_X32 FILLER_94_2023 ();
 FILLCELL_X32 FILLER_94_2055 ();
 FILLCELL_X32 FILLER_94_2087 ();
 FILLCELL_X32 FILLER_94_2119 ();
 FILLCELL_X32 FILLER_94_2151 ();
 FILLCELL_X32 FILLER_94_2183 ();
 FILLCELL_X32 FILLER_94_2215 ();
 FILLCELL_X32 FILLER_94_2247 ();
 FILLCELL_X32 FILLER_94_2279 ();
 FILLCELL_X32 FILLER_94_2311 ();
 FILLCELL_X32 FILLER_94_2343 ();
 FILLCELL_X32 FILLER_94_2375 ();
 FILLCELL_X32 FILLER_94_2407 ();
 FILLCELL_X32 FILLER_94_2439 ();
 FILLCELL_X32 FILLER_94_2471 ();
 FILLCELL_X32 FILLER_94_2503 ();
 FILLCELL_X32 FILLER_94_2535 ();
 FILLCELL_X32 FILLER_94_2567 ();
 FILLCELL_X32 FILLER_94_2599 ();
 FILLCELL_X32 FILLER_94_2631 ();
 FILLCELL_X32 FILLER_94_2663 ();
 FILLCELL_X32 FILLER_94_2695 ();
 FILLCELL_X32 FILLER_94_2727 ();
 FILLCELL_X32 FILLER_94_2759 ();
 FILLCELL_X32 FILLER_94_2791 ();
 FILLCELL_X32 FILLER_94_2823 ();
 FILLCELL_X32 FILLER_94_2855 ();
 FILLCELL_X32 FILLER_94_2887 ();
 FILLCELL_X32 FILLER_94_2919 ();
 FILLCELL_X32 FILLER_94_2951 ();
 FILLCELL_X32 FILLER_94_2983 ();
 FILLCELL_X32 FILLER_94_3015 ();
 FILLCELL_X32 FILLER_94_3047 ();
 FILLCELL_X32 FILLER_94_3079 ();
 FILLCELL_X32 FILLER_94_3111 ();
 FILLCELL_X8 FILLER_94_3143 ();
 FILLCELL_X4 FILLER_94_3151 ();
 FILLCELL_X2 FILLER_94_3155 ();
 FILLCELL_X32 FILLER_94_3158 ();
 FILLCELL_X32 FILLER_94_3190 ();
 FILLCELL_X32 FILLER_94_3222 ();
 FILLCELL_X32 FILLER_94_3254 ();
 FILLCELL_X32 FILLER_94_3286 ();
 FILLCELL_X32 FILLER_94_3318 ();
 FILLCELL_X32 FILLER_94_3350 ();
 FILLCELL_X32 FILLER_94_3382 ();
 FILLCELL_X32 FILLER_94_3414 ();
 FILLCELL_X32 FILLER_94_3446 ();
 FILLCELL_X32 FILLER_94_3478 ();
 FILLCELL_X32 FILLER_94_3510 ();
 FILLCELL_X32 FILLER_94_3542 ();
 FILLCELL_X32 FILLER_94_3574 ();
 FILLCELL_X32 FILLER_94_3606 ();
 FILLCELL_X32 FILLER_94_3638 ();
 FILLCELL_X32 FILLER_94_3670 ();
 FILLCELL_X32 FILLER_94_3702 ();
 FILLCELL_X4 FILLER_94_3734 ();
 FILLCELL_X32 FILLER_95_1 ();
 FILLCELL_X32 FILLER_95_33 ();
 FILLCELL_X32 FILLER_95_65 ();
 FILLCELL_X32 FILLER_95_97 ();
 FILLCELL_X32 FILLER_95_129 ();
 FILLCELL_X32 FILLER_95_161 ();
 FILLCELL_X32 FILLER_95_193 ();
 FILLCELL_X32 FILLER_95_225 ();
 FILLCELL_X32 FILLER_95_257 ();
 FILLCELL_X32 FILLER_95_289 ();
 FILLCELL_X32 FILLER_95_321 ();
 FILLCELL_X32 FILLER_95_353 ();
 FILLCELL_X32 FILLER_95_385 ();
 FILLCELL_X32 FILLER_95_417 ();
 FILLCELL_X32 FILLER_95_449 ();
 FILLCELL_X32 FILLER_95_481 ();
 FILLCELL_X32 FILLER_95_513 ();
 FILLCELL_X32 FILLER_95_545 ();
 FILLCELL_X32 FILLER_95_577 ();
 FILLCELL_X32 FILLER_95_609 ();
 FILLCELL_X32 FILLER_95_641 ();
 FILLCELL_X32 FILLER_95_673 ();
 FILLCELL_X32 FILLER_95_705 ();
 FILLCELL_X32 FILLER_95_737 ();
 FILLCELL_X32 FILLER_95_769 ();
 FILLCELL_X32 FILLER_95_801 ();
 FILLCELL_X32 FILLER_95_833 ();
 FILLCELL_X32 FILLER_95_865 ();
 FILLCELL_X32 FILLER_95_897 ();
 FILLCELL_X32 FILLER_95_929 ();
 FILLCELL_X32 FILLER_95_961 ();
 FILLCELL_X32 FILLER_95_993 ();
 FILLCELL_X32 FILLER_95_1025 ();
 FILLCELL_X32 FILLER_95_1057 ();
 FILLCELL_X32 FILLER_95_1089 ();
 FILLCELL_X32 FILLER_95_1121 ();
 FILLCELL_X32 FILLER_95_1153 ();
 FILLCELL_X32 FILLER_95_1185 ();
 FILLCELL_X32 FILLER_95_1217 ();
 FILLCELL_X8 FILLER_95_1249 ();
 FILLCELL_X4 FILLER_95_1257 ();
 FILLCELL_X2 FILLER_95_1261 ();
 FILLCELL_X32 FILLER_95_1264 ();
 FILLCELL_X32 FILLER_95_1296 ();
 FILLCELL_X32 FILLER_95_1328 ();
 FILLCELL_X32 FILLER_95_1360 ();
 FILLCELL_X32 FILLER_95_1392 ();
 FILLCELL_X32 FILLER_95_1424 ();
 FILLCELL_X32 FILLER_95_1456 ();
 FILLCELL_X32 FILLER_95_1488 ();
 FILLCELL_X32 FILLER_95_1520 ();
 FILLCELL_X32 FILLER_95_1552 ();
 FILLCELL_X32 FILLER_95_1584 ();
 FILLCELL_X32 FILLER_95_1616 ();
 FILLCELL_X32 FILLER_95_1648 ();
 FILLCELL_X32 FILLER_95_1680 ();
 FILLCELL_X32 FILLER_95_1712 ();
 FILLCELL_X32 FILLER_95_1744 ();
 FILLCELL_X32 FILLER_95_1776 ();
 FILLCELL_X32 FILLER_95_1808 ();
 FILLCELL_X32 FILLER_95_1840 ();
 FILLCELL_X32 FILLER_95_1872 ();
 FILLCELL_X32 FILLER_95_1904 ();
 FILLCELL_X32 FILLER_95_1936 ();
 FILLCELL_X32 FILLER_95_1968 ();
 FILLCELL_X32 FILLER_95_2000 ();
 FILLCELL_X32 FILLER_95_2032 ();
 FILLCELL_X32 FILLER_95_2064 ();
 FILLCELL_X32 FILLER_95_2096 ();
 FILLCELL_X32 FILLER_95_2128 ();
 FILLCELL_X32 FILLER_95_2160 ();
 FILLCELL_X32 FILLER_95_2192 ();
 FILLCELL_X32 FILLER_95_2224 ();
 FILLCELL_X32 FILLER_95_2256 ();
 FILLCELL_X32 FILLER_95_2288 ();
 FILLCELL_X32 FILLER_95_2320 ();
 FILLCELL_X32 FILLER_95_2352 ();
 FILLCELL_X32 FILLER_95_2384 ();
 FILLCELL_X32 FILLER_95_2416 ();
 FILLCELL_X32 FILLER_95_2448 ();
 FILLCELL_X32 FILLER_95_2480 ();
 FILLCELL_X8 FILLER_95_2512 ();
 FILLCELL_X4 FILLER_95_2520 ();
 FILLCELL_X2 FILLER_95_2524 ();
 FILLCELL_X32 FILLER_95_2527 ();
 FILLCELL_X32 FILLER_95_2559 ();
 FILLCELL_X32 FILLER_95_2591 ();
 FILLCELL_X32 FILLER_95_2623 ();
 FILLCELL_X32 FILLER_95_2655 ();
 FILLCELL_X32 FILLER_95_2687 ();
 FILLCELL_X32 FILLER_95_2719 ();
 FILLCELL_X32 FILLER_95_2751 ();
 FILLCELL_X32 FILLER_95_2783 ();
 FILLCELL_X32 FILLER_95_2815 ();
 FILLCELL_X32 FILLER_95_2847 ();
 FILLCELL_X32 FILLER_95_2879 ();
 FILLCELL_X32 FILLER_95_2911 ();
 FILLCELL_X32 FILLER_95_2943 ();
 FILLCELL_X32 FILLER_95_2975 ();
 FILLCELL_X32 FILLER_95_3007 ();
 FILLCELL_X32 FILLER_95_3039 ();
 FILLCELL_X32 FILLER_95_3071 ();
 FILLCELL_X32 FILLER_95_3103 ();
 FILLCELL_X32 FILLER_95_3135 ();
 FILLCELL_X32 FILLER_95_3167 ();
 FILLCELL_X32 FILLER_95_3199 ();
 FILLCELL_X32 FILLER_95_3231 ();
 FILLCELL_X32 FILLER_95_3263 ();
 FILLCELL_X32 FILLER_95_3295 ();
 FILLCELL_X32 FILLER_95_3327 ();
 FILLCELL_X32 FILLER_95_3359 ();
 FILLCELL_X32 FILLER_95_3391 ();
 FILLCELL_X32 FILLER_95_3423 ();
 FILLCELL_X32 FILLER_95_3455 ();
 FILLCELL_X32 FILLER_95_3487 ();
 FILLCELL_X32 FILLER_95_3519 ();
 FILLCELL_X32 FILLER_95_3551 ();
 FILLCELL_X32 FILLER_95_3583 ();
 FILLCELL_X32 FILLER_95_3615 ();
 FILLCELL_X32 FILLER_95_3647 ();
 FILLCELL_X32 FILLER_95_3679 ();
 FILLCELL_X16 FILLER_95_3711 ();
 FILLCELL_X8 FILLER_95_3727 ();
 FILLCELL_X2 FILLER_95_3735 ();
 FILLCELL_X1 FILLER_95_3737 ();
 FILLCELL_X32 FILLER_96_1 ();
 FILLCELL_X32 FILLER_96_33 ();
 FILLCELL_X32 FILLER_96_65 ();
 FILLCELL_X32 FILLER_96_97 ();
 FILLCELL_X32 FILLER_96_129 ();
 FILLCELL_X32 FILLER_96_161 ();
 FILLCELL_X32 FILLER_96_193 ();
 FILLCELL_X32 FILLER_96_225 ();
 FILLCELL_X32 FILLER_96_257 ();
 FILLCELL_X32 FILLER_96_289 ();
 FILLCELL_X32 FILLER_96_321 ();
 FILLCELL_X32 FILLER_96_353 ();
 FILLCELL_X32 FILLER_96_385 ();
 FILLCELL_X32 FILLER_96_417 ();
 FILLCELL_X32 FILLER_96_449 ();
 FILLCELL_X32 FILLER_96_481 ();
 FILLCELL_X32 FILLER_96_513 ();
 FILLCELL_X32 FILLER_96_545 ();
 FILLCELL_X32 FILLER_96_577 ();
 FILLCELL_X16 FILLER_96_609 ();
 FILLCELL_X4 FILLER_96_625 ();
 FILLCELL_X2 FILLER_96_629 ();
 FILLCELL_X32 FILLER_96_632 ();
 FILLCELL_X32 FILLER_96_664 ();
 FILLCELL_X32 FILLER_96_696 ();
 FILLCELL_X32 FILLER_96_728 ();
 FILLCELL_X32 FILLER_96_760 ();
 FILLCELL_X32 FILLER_96_792 ();
 FILLCELL_X32 FILLER_96_824 ();
 FILLCELL_X32 FILLER_96_856 ();
 FILLCELL_X32 FILLER_96_888 ();
 FILLCELL_X32 FILLER_96_920 ();
 FILLCELL_X32 FILLER_96_952 ();
 FILLCELL_X32 FILLER_96_984 ();
 FILLCELL_X32 FILLER_96_1016 ();
 FILLCELL_X32 FILLER_96_1048 ();
 FILLCELL_X32 FILLER_96_1080 ();
 FILLCELL_X32 FILLER_96_1112 ();
 FILLCELL_X32 FILLER_96_1144 ();
 FILLCELL_X32 FILLER_96_1176 ();
 FILLCELL_X32 FILLER_96_1208 ();
 FILLCELL_X32 FILLER_96_1240 ();
 FILLCELL_X32 FILLER_96_1272 ();
 FILLCELL_X32 FILLER_96_1304 ();
 FILLCELL_X32 FILLER_96_1336 ();
 FILLCELL_X32 FILLER_96_1368 ();
 FILLCELL_X32 FILLER_96_1400 ();
 FILLCELL_X32 FILLER_96_1432 ();
 FILLCELL_X32 FILLER_96_1464 ();
 FILLCELL_X32 FILLER_96_1496 ();
 FILLCELL_X32 FILLER_96_1528 ();
 FILLCELL_X32 FILLER_96_1560 ();
 FILLCELL_X32 FILLER_96_1592 ();
 FILLCELL_X32 FILLER_96_1624 ();
 FILLCELL_X32 FILLER_96_1656 ();
 FILLCELL_X32 FILLER_96_1688 ();
 FILLCELL_X32 FILLER_96_1720 ();
 FILLCELL_X32 FILLER_96_1752 ();
 FILLCELL_X32 FILLER_96_1784 ();
 FILLCELL_X32 FILLER_96_1816 ();
 FILLCELL_X32 FILLER_96_1848 ();
 FILLCELL_X8 FILLER_96_1880 ();
 FILLCELL_X4 FILLER_96_1888 ();
 FILLCELL_X2 FILLER_96_1892 ();
 FILLCELL_X32 FILLER_96_1895 ();
 FILLCELL_X32 FILLER_96_1927 ();
 FILLCELL_X32 FILLER_96_1959 ();
 FILLCELL_X32 FILLER_96_1991 ();
 FILLCELL_X32 FILLER_96_2023 ();
 FILLCELL_X32 FILLER_96_2055 ();
 FILLCELL_X32 FILLER_96_2087 ();
 FILLCELL_X32 FILLER_96_2119 ();
 FILLCELL_X32 FILLER_96_2151 ();
 FILLCELL_X32 FILLER_96_2183 ();
 FILLCELL_X32 FILLER_96_2215 ();
 FILLCELL_X32 FILLER_96_2247 ();
 FILLCELL_X32 FILLER_96_2279 ();
 FILLCELL_X32 FILLER_96_2311 ();
 FILLCELL_X32 FILLER_96_2343 ();
 FILLCELL_X32 FILLER_96_2375 ();
 FILLCELL_X32 FILLER_96_2407 ();
 FILLCELL_X32 FILLER_96_2439 ();
 FILLCELL_X32 FILLER_96_2471 ();
 FILLCELL_X32 FILLER_96_2503 ();
 FILLCELL_X32 FILLER_96_2535 ();
 FILLCELL_X32 FILLER_96_2567 ();
 FILLCELL_X32 FILLER_96_2599 ();
 FILLCELL_X32 FILLER_96_2631 ();
 FILLCELL_X32 FILLER_96_2663 ();
 FILLCELL_X32 FILLER_96_2695 ();
 FILLCELL_X32 FILLER_96_2727 ();
 FILLCELL_X32 FILLER_96_2759 ();
 FILLCELL_X32 FILLER_96_2791 ();
 FILLCELL_X32 FILLER_96_2823 ();
 FILLCELL_X32 FILLER_96_2855 ();
 FILLCELL_X32 FILLER_96_2887 ();
 FILLCELL_X32 FILLER_96_2919 ();
 FILLCELL_X32 FILLER_96_2951 ();
 FILLCELL_X32 FILLER_96_2983 ();
 FILLCELL_X32 FILLER_96_3015 ();
 FILLCELL_X32 FILLER_96_3047 ();
 FILLCELL_X32 FILLER_96_3079 ();
 FILLCELL_X32 FILLER_96_3111 ();
 FILLCELL_X8 FILLER_96_3143 ();
 FILLCELL_X4 FILLER_96_3151 ();
 FILLCELL_X2 FILLER_96_3155 ();
 FILLCELL_X32 FILLER_96_3158 ();
 FILLCELL_X32 FILLER_96_3190 ();
 FILLCELL_X32 FILLER_96_3222 ();
 FILLCELL_X32 FILLER_96_3254 ();
 FILLCELL_X32 FILLER_96_3286 ();
 FILLCELL_X32 FILLER_96_3318 ();
 FILLCELL_X32 FILLER_96_3350 ();
 FILLCELL_X32 FILLER_96_3382 ();
 FILLCELL_X32 FILLER_96_3414 ();
 FILLCELL_X32 FILLER_96_3446 ();
 FILLCELL_X32 FILLER_96_3478 ();
 FILLCELL_X32 FILLER_96_3510 ();
 FILLCELL_X32 FILLER_96_3542 ();
 FILLCELL_X32 FILLER_96_3574 ();
 FILLCELL_X32 FILLER_96_3606 ();
 FILLCELL_X32 FILLER_96_3638 ();
 FILLCELL_X32 FILLER_96_3670 ();
 FILLCELL_X32 FILLER_96_3702 ();
 FILLCELL_X4 FILLER_96_3734 ();
 FILLCELL_X32 FILLER_97_1 ();
 FILLCELL_X32 FILLER_97_33 ();
 FILLCELL_X32 FILLER_97_65 ();
 FILLCELL_X32 FILLER_97_97 ();
 FILLCELL_X32 FILLER_97_129 ();
 FILLCELL_X32 FILLER_97_161 ();
 FILLCELL_X32 FILLER_97_193 ();
 FILLCELL_X32 FILLER_97_225 ();
 FILLCELL_X32 FILLER_97_257 ();
 FILLCELL_X32 FILLER_97_289 ();
 FILLCELL_X32 FILLER_97_321 ();
 FILLCELL_X32 FILLER_97_353 ();
 FILLCELL_X32 FILLER_97_385 ();
 FILLCELL_X32 FILLER_97_417 ();
 FILLCELL_X32 FILLER_97_449 ();
 FILLCELL_X32 FILLER_97_481 ();
 FILLCELL_X32 FILLER_97_513 ();
 FILLCELL_X32 FILLER_97_545 ();
 FILLCELL_X32 FILLER_97_577 ();
 FILLCELL_X32 FILLER_97_609 ();
 FILLCELL_X32 FILLER_97_641 ();
 FILLCELL_X32 FILLER_97_673 ();
 FILLCELL_X32 FILLER_97_705 ();
 FILLCELL_X32 FILLER_97_737 ();
 FILLCELL_X32 FILLER_97_769 ();
 FILLCELL_X32 FILLER_97_801 ();
 FILLCELL_X32 FILLER_97_833 ();
 FILLCELL_X32 FILLER_97_865 ();
 FILLCELL_X32 FILLER_97_897 ();
 FILLCELL_X32 FILLER_97_929 ();
 FILLCELL_X32 FILLER_97_961 ();
 FILLCELL_X32 FILLER_97_993 ();
 FILLCELL_X32 FILLER_97_1025 ();
 FILLCELL_X32 FILLER_97_1057 ();
 FILLCELL_X32 FILLER_97_1089 ();
 FILLCELL_X32 FILLER_97_1121 ();
 FILLCELL_X32 FILLER_97_1153 ();
 FILLCELL_X32 FILLER_97_1185 ();
 FILLCELL_X32 FILLER_97_1217 ();
 FILLCELL_X8 FILLER_97_1249 ();
 FILLCELL_X4 FILLER_97_1257 ();
 FILLCELL_X2 FILLER_97_1261 ();
 FILLCELL_X32 FILLER_97_1264 ();
 FILLCELL_X32 FILLER_97_1296 ();
 FILLCELL_X32 FILLER_97_1328 ();
 FILLCELL_X32 FILLER_97_1360 ();
 FILLCELL_X32 FILLER_97_1392 ();
 FILLCELL_X32 FILLER_97_1424 ();
 FILLCELL_X32 FILLER_97_1456 ();
 FILLCELL_X32 FILLER_97_1488 ();
 FILLCELL_X32 FILLER_97_1520 ();
 FILLCELL_X32 FILLER_97_1552 ();
 FILLCELL_X32 FILLER_97_1584 ();
 FILLCELL_X32 FILLER_97_1616 ();
 FILLCELL_X32 FILLER_97_1648 ();
 FILLCELL_X32 FILLER_97_1680 ();
 FILLCELL_X32 FILLER_97_1712 ();
 FILLCELL_X32 FILLER_97_1744 ();
 FILLCELL_X32 FILLER_97_1776 ();
 FILLCELL_X32 FILLER_97_1808 ();
 FILLCELL_X32 FILLER_97_1840 ();
 FILLCELL_X32 FILLER_97_1872 ();
 FILLCELL_X32 FILLER_97_1904 ();
 FILLCELL_X32 FILLER_97_1936 ();
 FILLCELL_X32 FILLER_97_1968 ();
 FILLCELL_X32 FILLER_97_2000 ();
 FILLCELL_X32 FILLER_97_2032 ();
 FILLCELL_X32 FILLER_97_2064 ();
 FILLCELL_X32 FILLER_97_2096 ();
 FILLCELL_X32 FILLER_97_2128 ();
 FILLCELL_X32 FILLER_97_2160 ();
 FILLCELL_X32 FILLER_97_2192 ();
 FILLCELL_X32 FILLER_97_2224 ();
 FILLCELL_X32 FILLER_97_2256 ();
 FILLCELL_X32 FILLER_97_2288 ();
 FILLCELL_X32 FILLER_97_2320 ();
 FILLCELL_X32 FILLER_97_2352 ();
 FILLCELL_X32 FILLER_97_2384 ();
 FILLCELL_X32 FILLER_97_2416 ();
 FILLCELL_X32 FILLER_97_2448 ();
 FILLCELL_X32 FILLER_97_2480 ();
 FILLCELL_X8 FILLER_97_2512 ();
 FILLCELL_X4 FILLER_97_2520 ();
 FILLCELL_X2 FILLER_97_2524 ();
 FILLCELL_X32 FILLER_97_2527 ();
 FILLCELL_X32 FILLER_97_2559 ();
 FILLCELL_X32 FILLER_97_2591 ();
 FILLCELL_X32 FILLER_97_2623 ();
 FILLCELL_X32 FILLER_97_2655 ();
 FILLCELL_X32 FILLER_97_2687 ();
 FILLCELL_X32 FILLER_97_2719 ();
 FILLCELL_X32 FILLER_97_2751 ();
 FILLCELL_X32 FILLER_97_2783 ();
 FILLCELL_X32 FILLER_97_2815 ();
 FILLCELL_X32 FILLER_97_2847 ();
 FILLCELL_X32 FILLER_97_2879 ();
 FILLCELL_X32 FILLER_97_2911 ();
 FILLCELL_X32 FILLER_97_2943 ();
 FILLCELL_X32 FILLER_97_2975 ();
 FILLCELL_X32 FILLER_97_3007 ();
 FILLCELL_X32 FILLER_97_3039 ();
 FILLCELL_X32 FILLER_97_3071 ();
 FILLCELL_X32 FILLER_97_3103 ();
 FILLCELL_X32 FILLER_97_3135 ();
 FILLCELL_X32 FILLER_97_3167 ();
 FILLCELL_X32 FILLER_97_3199 ();
 FILLCELL_X32 FILLER_97_3231 ();
 FILLCELL_X32 FILLER_97_3263 ();
 FILLCELL_X32 FILLER_97_3295 ();
 FILLCELL_X32 FILLER_97_3327 ();
 FILLCELL_X32 FILLER_97_3359 ();
 FILLCELL_X32 FILLER_97_3391 ();
 FILLCELL_X32 FILLER_97_3423 ();
 FILLCELL_X32 FILLER_97_3455 ();
 FILLCELL_X32 FILLER_97_3487 ();
 FILLCELL_X32 FILLER_97_3519 ();
 FILLCELL_X32 FILLER_97_3551 ();
 FILLCELL_X32 FILLER_97_3583 ();
 FILLCELL_X32 FILLER_97_3615 ();
 FILLCELL_X32 FILLER_97_3647 ();
 FILLCELL_X32 FILLER_97_3679 ();
 FILLCELL_X16 FILLER_97_3711 ();
 FILLCELL_X8 FILLER_97_3727 ();
 FILLCELL_X2 FILLER_97_3735 ();
 FILLCELL_X1 FILLER_97_3737 ();
 FILLCELL_X32 FILLER_98_1 ();
 FILLCELL_X32 FILLER_98_33 ();
 FILLCELL_X32 FILLER_98_65 ();
 FILLCELL_X32 FILLER_98_97 ();
 FILLCELL_X32 FILLER_98_129 ();
 FILLCELL_X32 FILLER_98_161 ();
 FILLCELL_X32 FILLER_98_193 ();
 FILLCELL_X32 FILLER_98_225 ();
 FILLCELL_X32 FILLER_98_257 ();
 FILLCELL_X32 FILLER_98_289 ();
 FILLCELL_X32 FILLER_98_321 ();
 FILLCELL_X32 FILLER_98_353 ();
 FILLCELL_X32 FILLER_98_385 ();
 FILLCELL_X32 FILLER_98_417 ();
 FILLCELL_X32 FILLER_98_449 ();
 FILLCELL_X32 FILLER_98_481 ();
 FILLCELL_X32 FILLER_98_513 ();
 FILLCELL_X32 FILLER_98_545 ();
 FILLCELL_X32 FILLER_98_577 ();
 FILLCELL_X16 FILLER_98_609 ();
 FILLCELL_X4 FILLER_98_625 ();
 FILLCELL_X2 FILLER_98_629 ();
 FILLCELL_X32 FILLER_98_632 ();
 FILLCELL_X32 FILLER_98_664 ();
 FILLCELL_X32 FILLER_98_696 ();
 FILLCELL_X32 FILLER_98_728 ();
 FILLCELL_X32 FILLER_98_760 ();
 FILLCELL_X32 FILLER_98_792 ();
 FILLCELL_X32 FILLER_98_824 ();
 FILLCELL_X32 FILLER_98_856 ();
 FILLCELL_X32 FILLER_98_888 ();
 FILLCELL_X32 FILLER_98_920 ();
 FILLCELL_X32 FILLER_98_952 ();
 FILLCELL_X32 FILLER_98_984 ();
 FILLCELL_X32 FILLER_98_1016 ();
 FILLCELL_X32 FILLER_98_1048 ();
 FILLCELL_X32 FILLER_98_1080 ();
 FILLCELL_X32 FILLER_98_1112 ();
 FILLCELL_X32 FILLER_98_1144 ();
 FILLCELL_X32 FILLER_98_1176 ();
 FILLCELL_X32 FILLER_98_1208 ();
 FILLCELL_X32 FILLER_98_1240 ();
 FILLCELL_X32 FILLER_98_1272 ();
 FILLCELL_X32 FILLER_98_1304 ();
 FILLCELL_X32 FILLER_98_1336 ();
 FILLCELL_X32 FILLER_98_1368 ();
 FILLCELL_X32 FILLER_98_1400 ();
 FILLCELL_X32 FILLER_98_1432 ();
 FILLCELL_X32 FILLER_98_1464 ();
 FILLCELL_X32 FILLER_98_1496 ();
 FILLCELL_X32 FILLER_98_1528 ();
 FILLCELL_X32 FILLER_98_1560 ();
 FILLCELL_X32 FILLER_98_1592 ();
 FILLCELL_X32 FILLER_98_1624 ();
 FILLCELL_X32 FILLER_98_1656 ();
 FILLCELL_X32 FILLER_98_1688 ();
 FILLCELL_X32 FILLER_98_1720 ();
 FILLCELL_X32 FILLER_98_1752 ();
 FILLCELL_X32 FILLER_98_1784 ();
 FILLCELL_X32 FILLER_98_1816 ();
 FILLCELL_X32 FILLER_98_1848 ();
 FILLCELL_X8 FILLER_98_1880 ();
 FILLCELL_X4 FILLER_98_1888 ();
 FILLCELL_X2 FILLER_98_1892 ();
 FILLCELL_X32 FILLER_98_1895 ();
 FILLCELL_X32 FILLER_98_1927 ();
 FILLCELL_X32 FILLER_98_1959 ();
 FILLCELL_X32 FILLER_98_1991 ();
 FILLCELL_X32 FILLER_98_2023 ();
 FILLCELL_X32 FILLER_98_2055 ();
 FILLCELL_X32 FILLER_98_2087 ();
 FILLCELL_X32 FILLER_98_2119 ();
 FILLCELL_X32 FILLER_98_2151 ();
 FILLCELL_X32 FILLER_98_2183 ();
 FILLCELL_X32 FILLER_98_2215 ();
 FILLCELL_X32 FILLER_98_2247 ();
 FILLCELL_X32 FILLER_98_2279 ();
 FILLCELL_X32 FILLER_98_2311 ();
 FILLCELL_X32 FILLER_98_2343 ();
 FILLCELL_X32 FILLER_98_2375 ();
 FILLCELL_X32 FILLER_98_2407 ();
 FILLCELL_X32 FILLER_98_2439 ();
 FILLCELL_X32 FILLER_98_2471 ();
 FILLCELL_X32 FILLER_98_2503 ();
 FILLCELL_X32 FILLER_98_2535 ();
 FILLCELL_X32 FILLER_98_2567 ();
 FILLCELL_X32 FILLER_98_2599 ();
 FILLCELL_X32 FILLER_98_2631 ();
 FILLCELL_X32 FILLER_98_2663 ();
 FILLCELL_X32 FILLER_98_2695 ();
 FILLCELL_X32 FILLER_98_2727 ();
 FILLCELL_X32 FILLER_98_2759 ();
 FILLCELL_X32 FILLER_98_2791 ();
 FILLCELL_X32 FILLER_98_2823 ();
 FILLCELL_X32 FILLER_98_2855 ();
 FILLCELL_X32 FILLER_98_2887 ();
 FILLCELL_X32 FILLER_98_2919 ();
 FILLCELL_X32 FILLER_98_2951 ();
 FILLCELL_X32 FILLER_98_2983 ();
 FILLCELL_X32 FILLER_98_3015 ();
 FILLCELL_X32 FILLER_98_3047 ();
 FILLCELL_X32 FILLER_98_3079 ();
 FILLCELL_X32 FILLER_98_3111 ();
 FILLCELL_X8 FILLER_98_3143 ();
 FILLCELL_X4 FILLER_98_3151 ();
 FILLCELL_X2 FILLER_98_3155 ();
 FILLCELL_X32 FILLER_98_3158 ();
 FILLCELL_X32 FILLER_98_3190 ();
 FILLCELL_X32 FILLER_98_3222 ();
 FILLCELL_X32 FILLER_98_3254 ();
 FILLCELL_X32 FILLER_98_3286 ();
 FILLCELL_X32 FILLER_98_3318 ();
 FILLCELL_X32 FILLER_98_3350 ();
 FILLCELL_X32 FILLER_98_3382 ();
 FILLCELL_X32 FILLER_98_3414 ();
 FILLCELL_X32 FILLER_98_3446 ();
 FILLCELL_X32 FILLER_98_3478 ();
 FILLCELL_X32 FILLER_98_3510 ();
 FILLCELL_X32 FILLER_98_3542 ();
 FILLCELL_X32 FILLER_98_3574 ();
 FILLCELL_X32 FILLER_98_3606 ();
 FILLCELL_X32 FILLER_98_3638 ();
 FILLCELL_X32 FILLER_98_3670 ();
 FILLCELL_X32 FILLER_98_3702 ();
 FILLCELL_X4 FILLER_98_3734 ();
 FILLCELL_X32 FILLER_99_1 ();
 FILLCELL_X32 FILLER_99_33 ();
 FILLCELL_X32 FILLER_99_65 ();
 FILLCELL_X32 FILLER_99_97 ();
 FILLCELL_X32 FILLER_99_129 ();
 FILLCELL_X32 FILLER_99_161 ();
 FILLCELL_X32 FILLER_99_193 ();
 FILLCELL_X32 FILLER_99_225 ();
 FILLCELL_X32 FILLER_99_257 ();
 FILLCELL_X32 FILLER_99_289 ();
 FILLCELL_X32 FILLER_99_321 ();
 FILLCELL_X32 FILLER_99_353 ();
 FILLCELL_X32 FILLER_99_385 ();
 FILLCELL_X32 FILLER_99_417 ();
 FILLCELL_X32 FILLER_99_449 ();
 FILLCELL_X32 FILLER_99_481 ();
 FILLCELL_X32 FILLER_99_513 ();
 FILLCELL_X32 FILLER_99_545 ();
 FILLCELL_X32 FILLER_99_577 ();
 FILLCELL_X32 FILLER_99_609 ();
 FILLCELL_X32 FILLER_99_641 ();
 FILLCELL_X32 FILLER_99_673 ();
 FILLCELL_X32 FILLER_99_705 ();
 FILLCELL_X32 FILLER_99_737 ();
 FILLCELL_X32 FILLER_99_769 ();
 FILLCELL_X32 FILLER_99_801 ();
 FILLCELL_X32 FILLER_99_833 ();
 FILLCELL_X32 FILLER_99_865 ();
 FILLCELL_X32 FILLER_99_897 ();
 FILLCELL_X32 FILLER_99_929 ();
 FILLCELL_X32 FILLER_99_961 ();
 FILLCELL_X32 FILLER_99_993 ();
 FILLCELL_X32 FILLER_99_1025 ();
 FILLCELL_X32 FILLER_99_1057 ();
 FILLCELL_X32 FILLER_99_1089 ();
 FILLCELL_X32 FILLER_99_1121 ();
 FILLCELL_X32 FILLER_99_1153 ();
 FILLCELL_X32 FILLER_99_1185 ();
 FILLCELL_X32 FILLER_99_1217 ();
 FILLCELL_X8 FILLER_99_1249 ();
 FILLCELL_X4 FILLER_99_1257 ();
 FILLCELL_X2 FILLER_99_1261 ();
 FILLCELL_X32 FILLER_99_1264 ();
 FILLCELL_X32 FILLER_99_1296 ();
 FILLCELL_X32 FILLER_99_1328 ();
 FILLCELL_X32 FILLER_99_1360 ();
 FILLCELL_X32 FILLER_99_1392 ();
 FILLCELL_X32 FILLER_99_1424 ();
 FILLCELL_X32 FILLER_99_1456 ();
 FILLCELL_X32 FILLER_99_1488 ();
 FILLCELL_X32 FILLER_99_1520 ();
 FILLCELL_X32 FILLER_99_1552 ();
 FILLCELL_X32 FILLER_99_1584 ();
 FILLCELL_X32 FILLER_99_1616 ();
 FILLCELL_X32 FILLER_99_1648 ();
 FILLCELL_X32 FILLER_99_1680 ();
 FILLCELL_X32 FILLER_99_1712 ();
 FILLCELL_X32 FILLER_99_1744 ();
 FILLCELL_X32 FILLER_99_1776 ();
 FILLCELL_X32 FILLER_99_1808 ();
 FILLCELL_X32 FILLER_99_1840 ();
 FILLCELL_X32 FILLER_99_1872 ();
 FILLCELL_X32 FILLER_99_1904 ();
 FILLCELL_X32 FILLER_99_1936 ();
 FILLCELL_X32 FILLER_99_1968 ();
 FILLCELL_X32 FILLER_99_2000 ();
 FILLCELL_X32 FILLER_99_2032 ();
 FILLCELL_X32 FILLER_99_2064 ();
 FILLCELL_X32 FILLER_99_2096 ();
 FILLCELL_X32 FILLER_99_2128 ();
 FILLCELL_X32 FILLER_99_2160 ();
 FILLCELL_X32 FILLER_99_2192 ();
 FILLCELL_X32 FILLER_99_2224 ();
 FILLCELL_X32 FILLER_99_2256 ();
 FILLCELL_X32 FILLER_99_2288 ();
 FILLCELL_X32 FILLER_99_2320 ();
 FILLCELL_X32 FILLER_99_2352 ();
 FILLCELL_X32 FILLER_99_2384 ();
 FILLCELL_X32 FILLER_99_2416 ();
 FILLCELL_X32 FILLER_99_2448 ();
 FILLCELL_X32 FILLER_99_2480 ();
 FILLCELL_X8 FILLER_99_2512 ();
 FILLCELL_X4 FILLER_99_2520 ();
 FILLCELL_X2 FILLER_99_2524 ();
 FILLCELL_X32 FILLER_99_2527 ();
 FILLCELL_X32 FILLER_99_2559 ();
 FILLCELL_X32 FILLER_99_2591 ();
 FILLCELL_X32 FILLER_99_2623 ();
 FILLCELL_X32 FILLER_99_2655 ();
 FILLCELL_X32 FILLER_99_2687 ();
 FILLCELL_X32 FILLER_99_2719 ();
 FILLCELL_X32 FILLER_99_2751 ();
 FILLCELL_X32 FILLER_99_2783 ();
 FILLCELL_X32 FILLER_99_2815 ();
 FILLCELL_X32 FILLER_99_2847 ();
 FILLCELL_X32 FILLER_99_2879 ();
 FILLCELL_X32 FILLER_99_2911 ();
 FILLCELL_X32 FILLER_99_2943 ();
 FILLCELL_X32 FILLER_99_2975 ();
 FILLCELL_X32 FILLER_99_3007 ();
 FILLCELL_X32 FILLER_99_3039 ();
 FILLCELL_X32 FILLER_99_3071 ();
 FILLCELL_X32 FILLER_99_3103 ();
 FILLCELL_X32 FILLER_99_3135 ();
 FILLCELL_X32 FILLER_99_3167 ();
 FILLCELL_X32 FILLER_99_3199 ();
 FILLCELL_X32 FILLER_99_3231 ();
 FILLCELL_X32 FILLER_99_3263 ();
 FILLCELL_X32 FILLER_99_3295 ();
 FILLCELL_X32 FILLER_99_3327 ();
 FILLCELL_X32 FILLER_99_3359 ();
 FILLCELL_X32 FILLER_99_3391 ();
 FILLCELL_X32 FILLER_99_3423 ();
 FILLCELL_X32 FILLER_99_3455 ();
 FILLCELL_X32 FILLER_99_3487 ();
 FILLCELL_X32 FILLER_99_3519 ();
 FILLCELL_X32 FILLER_99_3551 ();
 FILLCELL_X32 FILLER_99_3583 ();
 FILLCELL_X32 FILLER_99_3615 ();
 FILLCELL_X32 FILLER_99_3647 ();
 FILLCELL_X32 FILLER_99_3679 ();
 FILLCELL_X16 FILLER_99_3711 ();
 FILLCELL_X8 FILLER_99_3727 ();
 FILLCELL_X2 FILLER_99_3735 ();
 FILLCELL_X1 FILLER_99_3737 ();
 FILLCELL_X32 FILLER_100_1 ();
 FILLCELL_X32 FILLER_100_33 ();
 FILLCELL_X32 FILLER_100_65 ();
 FILLCELL_X32 FILLER_100_97 ();
 FILLCELL_X32 FILLER_100_129 ();
 FILLCELL_X32 FILLER_100_161 ();
 FILLCELL_X32 FILLER_100_193 ();
 FILLCELL_X32 FILLER_100_225 ();
 FILLCELL_X32 FILLER_100_257 ();
 FILLCELL_X32 FILLER_100_289 ();
 FILLCELL_X32 FILLER_100_321 ();
 FILLCELL_X32 FILLER_100_353 ();
 FILLCELL_X32 FILLER_100_385 ();
 FILLCELL_X32 FILLER_100_417 ();
 FILLCELL_X32 FILLER_100_449 ();
 FILLCELL_X32 FILLER_100_481 ();
 FILLCELL_X32 FILLER_100_513 ();
 FILLCELL_X32 FILLER_100_545 ();
 FILLCELL_X32 FILLER_100_577 ();
 FILLCELL_X16 FILLER_100_609 ();
 FILLCELL_X4 FILLER_100_625 ();
 FILLCELL_X2 FILLER_100_629 ();
 FILLCELL_X32 FILLER_100_632 ();
 FILLCELL_X32 FILLER_100_664 ();
 FILLCELL_X32 FILLER_100_696 ();
 FILLCELL_X32 FILLER_100_728 ();
 FILLCELL_X32 FILLER_100_760 ();
 FILLCELL_X32 FILLER_100_792 ();
 FILLCELL_X32 FILLER_100_824 ();
 FILLCELL_X32 FILLER_100_856 ();
 FILLCELL_X32 FILLER_100_888 ();
 FILLCELL_X32 FILLER_100_920 ();
 FILLCELL_X32 FILLER_100_952 ();
 FILLCELL_X32 FILLER_100_984 ();
 FILLCELL_X32 FILLER_100_1016 ();
 FILLCELL_X32 FILLER_100_1048 ();
 FILLCELL_X32 FILLER_100_1080 ();
 FILLCELL_X32 FILLER_100_1112 ();
 FILLCELL_X32 FILLER_100_1144 ();
 FILLCELL_X32 FILLER_100_1176 ();
 FILLCELL_X32 FILLER_100_1208 ();
 FILLCELL_X32 FILLER_100_1240 ();
 FILLCELL_X32 FILLER_100_1272 ();
 FILLCELL_X32 FILLER_100_1304 ();
 FILLCELL_X32 FILLER_100_1336 ();
 FILLCELL_X32 FILLER_100_1368 ();
 FILLCELL_X32 FILLER_100_1400 ();
 FILLCELL_X32 FILLER_100_1432 ();
 FILLCELL_X32 FILLER_100_1464 ();
 FILLCELL_X32 FILLER_100_1496 ();
 FILLCELL_X32 FILLER_100_1528 ();
 FILLCELL_X32 FILLER_100_1560 ();
 FILLCELL_X32 FILLER_100_1592 ();
 FILLCELL_X32 FILLER_100_1624 ();
 FILLCELL_X32 FILLER_100_1656 ();
 FILLCELL_X32 FILLER_100_1688 ();
 FILLCELL_X32 FILLER_100_1720 ();
 FILLCELL_X32 FILLER_100_1752 ();
 FILLCELL_X32 FILLER_100_1784 ();
 FILLCELL_X32 FILLER_100_1816 ();
 FILLCELL_X32 FILLER_100_1848 ();
 FILLCELL_X8 FILLER_100_1880 ();
 FILLCELL_X4 FILLER_100_1888 ();
 FILLCELL_X2 FILLER_100_1892 ();
 FILLCELL_X32 FILLER_100_1895 ();
 FILLCELL_X32 FILLER_100_1927 ();
 FILLCELL_X32 FILLER_100_1959 ();
 FILLCELL_X32 FILLER_100_1991 ();
 FILLCELL_X32 FILLER_100_2023 ();
 FILLCELL_X32 FILLER_100_2055 ();
 FILLCELL_X32 FILLER_100_2087 ();
 FILLCELL_X32 FILLER_100_2119 ();
 FILLCELL_X32 FILLER_100_2151 ();
 FILLCELL_X32 FILLER_100_2183 ();
 FILLCELL_X32 FILLER_100_2215 ();
 FILLCELL_X32 FILLER_100_2247 ();
 FILLCELL_X32 FILLER_100_2279 ();
 FILLCELL_X32 FILLER_100_2311 ();
 FILLCELL_X32 FILLER_100_2343 ();
 FILLCELL_X32 FILLER_100_2375 ();
 FILLCELL_X32 FILLER_100_2407 ();
 FILLCELL_X32 FILLER_100_2439 ();
 FILLCELL_X32 FILLER_100_2471 ();
 FILLCELL_X32 FILLER_100_2503 ();
 FILLCELL_X32 FILLER_100_2535 ();
 FILLCELL_X32 FILLER_100_2567 ();
 FILLCELL_X32 FILLER_100_2599 ();
 FILLCELL_X32 FILLER_100_2631 ();
 FILLCELL_X32 FILLER_100_2663 ();
 FILLCELL_X32 FILLER_100_2695 ();
 FILLCELL_X32 FILLER_100_2727 ();
 FILLCELL_X32 FILLER_100_2759 ();
 FILLCELL_X32 FILLER_100_2791 ();
 FILLCELL_X32 FILLER_100_2823 ();
 FILLCELL_X32 FILLER_100_2855 ();
 FILLCELL_X32 FILLER_100_2887 ();
 FILLCELL_X32 FILLER_100_2919 ();
 FILLCELL_X32 FILLER_100_2951 ();
 FILLCELL_X32 FILLER_100_2983 ();
 FILLCELL_X32 FILLER_100_3015 ();
 FILLCELL_X32 FILLER_100_3047 ();
 FILLCELL_X32 FILLER_100_3079 ();
 FILLCELL_X32 FILLER_100_3111 ();
 FILLCELL_X8 FILLER_100_3143 ();
 FILLCELL_X4 FILLER_100_3151 ();
 FILLCELL_X2 FILLER_100_3155 ();
 FILLCELL_X32 FILLER_100_3158 ();
 FILLCELL_X32 FILLER_100_3190 ();
 FILLCELL_X32 FILLER_100_3222 ();
 FILLCELL_X32 FILLER_100_3254 ();
 FILLCELL_X32 FILLER_100_3286 ();
 FILLCELL_X32 FILLER_100_3318 ();
 FILLCELL_X32 FILLER_100_3350 ();
 FILLCELL_X32 FILLER_100_3382 ();
 FILLCELL_X32 FILLER_100_3414 ();
 FILLCELL_X32 FILLER_100_3446 ();
 FILLCELL_X32 FILLER_100_3478 ();
 FILLCELL_X32 FILLER_100_3510 ();
 FILLCELL_X32 FILLER_100_3542 ();
 FILLCELL_X32 FILLER_100_3574 ();
 FILLCELL_X32 FILLER_100_3606 ();
 FILLCELL_X32 FILLER_100_3638 ();
 FILLCELL_X32 FILLER_100_3670 ();
 FILLCELL_X32 FILLER_100_3702 ();
 FILLCELL_X4 FILLER_100_3734 ();
 FILLCELL_X32 FILLER_101_1 ();
 FILLCELL_X32 FILLER_101_33 ();
 FILLCELL_X32 FILLER_101_65 ();
 FILLCELL_X32 FILLER_101_97 ();
 FILLCELL_X32 FILLER_101_129 ();
 FILLCELL_X32 FILLER_101_161 ();
 FILLCELL_X32 FILLER_101_193 ();
 FILLCELL_X32 FILLER_101_225 ();
 FILLCELL_X32 FILLER_101_257 ();
 FILLCELL_X32 FILLER_101_289 ();
 FILLCELL_X32 FILLER_101_321 ();
 FILLCELL_X32 FILLER_101_353 ();
 FILLCELL_X32 FILLER_101_385 ();
 FILLCELL_X32 FILLER_101_417 ();
 FILLCELL_X32 FILLER_101_449 ();
 FILLCELL_X32 FILLER_101_481 ();
 FILLCELL_X32 FILLER_101_513 ();
 FILLCELL_X32 FILLER_101_545 ();
 FILLCELL_X32 FILLER_101_577 ();
 FILLCELL_X32 FILLER_101_609 ();
 FILLCELL_X32 FILLER_101_641 ();
 FILLCELL_X32 FILLER_101_673 ();
 FILLCELL_X32 FILLER_101_705 ();
 FILLCELL_X32 FILLER_101_737 ();
 FILLCELL_X32 FILLER_101_769 ();
 FILLCELL_X32 FILLER_101_801 ();
 FILLCELL_X32 FILLER_101_833 ();
 FILLCELL_X32 FILLER_101_865 ();
 FILLCELL_X32 FILLER_101_897 ();
 FILLCELL_X32 FILLER_101_929 ();
 FILLCELL_X32 FILLER_101_961 ();
 FILLCELL_X32 FILLER_101_993 ();
 FILLCELL_X32 FILLER_101_1025 ();
 FILLCELL_X32 FILLER_101_1057 ();
 FILLCELL_X32 FILLER_101_1089 ();
 FILLCELL_X32 FILLER_101_1121 ();
 FILLCELL_X32 FILLER_101_1153 ();
 FILLCELL_X32 FILLER_101_1185 ();
 FILLCELL_X32 FILLER_101_1217 ();
 FILLCELL_X8 FILLER_101_1249 ();
 FILLCELL_X4 FILLER_101_1257 ();
 FILLCELL_X2 FILLER_101_1261 ();
 FILLCELL_X32 FILLER_101_1264 ();
 FILLCELL_X32 FILLER_101_1296 ();
 FILLCELL_X32 FILLER_101_1328 ();
 FILLCELL_X32 FILLER_101_1360 ();
 FILLCELL_X32 FILLER_101_1392 ();
 FILLCELL_X32 FILLER_101_1424 ();
 FILLCELL_X32 FILLER_101_1456 ();
 FILLCELL_X32 FILLER_101_1488 ();
 FILLCELL_X32 FILLER_101_1520 ();
 FILLCELL_X32 FILLER_101_1552 ();
 FILLCELL_X32 FILLER_101_1584 ();
 FILLCELL_X32 FILLER_101_1616 ();
 FILLCELL_X32 FILLER_101_1648 ();
 FILLCELL_X32 FILLER_101_1680 ();
 FILLCELL_X32 FILLER_101_1712 ();
 FILLCELL_X32 FILLER_101_1744 ();
 FILLCELL_X32 FILLER_101_1776 ();
 FILLCELL_X32 FILLER_101_1808 ();
 FILLCELL_X32 FILLER_101_1840 ();
 FILLCELL_X32 FILLER_101_1872 ();
 FILLCELL_X32 FILLER_101_1904 ();
 FILLCELL_X32 FILLER_101_1936 ();
 FILLCELL_X32 FILLER_101_1968 ();
 FILLCELL_X32 FILLER_101_2000 ();
 FILLCELL_X32 FILLER_101_2032 ();
 FILLCELL_X32 FILLER_101_2064 ();
 FILLCELL_X32 FILLER_101_2096 ();
 FILLCELL_X32 FILLER_101_2128 ();
 FILLCELL_X32 FILLER_101_2160 ();
 FILLCELL_X32 FILLER_101_2192 ();
 FILLCELL_X32 FILLER_101_2224 ();
 FILLCELL_X32 FILLER_101_2256 ();
 FILLCELL_X32 FILLER_101_2288 ();
 FILLCELL_X32 FILLER_101_2320 ();
 FILLCELL_X32 FILLER_101_2352 ();
 FILLCELL_X32 FILLER_101_2384 ();
 FILLCELL_X32 FILLER_101_2416 ();
 FILLCELL_X32 FILLER_101_2448 ();
 FILLCELL_X32 FILLER_101_2480 ();
 FILLCELL_X8 FILLER_101_2512 ();
 FILLCELL_X4 FILLER_101_2520 ();
 FILLCELL_X2 FILLER_101_2524 ();
 FILLCELL_X32 FILLER_101_2527 ();
 FILLCELL_X32 FILLER_101_2559 ();
 FILLCELL_X32 FILLER_101_2591 ();
 FILLCELL_X32 FILLER_101_2623 ();
 FILLCELL_X32 FILLER_101_2655 ();
 FILLCELL_X32 FILLER_101_2687 ();
 FILLCELL_X32 FILLER_101_2719 ();
 FILLCELL_X32 FILLER_101_2751 ();
 FILLCELL_X32 FILLER_101_2783 ();
 FILLCELL_X32 FILLER_101_2815 ();
 FILLCELL_X32 FILLER_101_2847 ();
 FILLCELL_X32 FILLER_101_2879 ();
 FILLCELL_X32 FILLER_101_2911 ();
 FILLCELL_X32 FILLER_101_2943 ();
 FILLCELL_X32 FILLER_101_2975 ();
 FILLCELL_X32 FILLER_101_3007 ();
 FILLCELL_X32 FILLER_101_3039 ();
 FILLCELL_X32 FILLER_101_3071 ();
 FILLCELL_X32 FILLER_101_3103 ();
 FILLCELL_X32 FILLER_101_3135 ();
 FILLCELL_X32 FILLER_101_3167 ();
 FILLCELL_X32 FILLER_101_3199 ();
 FILLCELL_X32 FILLER_101_3231 ();
 FILLCELL_X32 FILLER_101_3263 ();
 FILLCELL_X32 FILLER_101_3295 ();
 FILLCELL_X32 FILLER_101_3327 ();
 FILLCELL_X32 FILLER_101_3359 ();
 FILLCELL_X32 FILLER_101_3391 ();
 FILLCELL_X32 FILLER_101_3423 ();
 FILLCELL_X32 FILLER_101_3455 ();
 FILLCELL_X32 FILLER_101_3487 ();
 FILLCELL_X32 FILLER_101_3519 ();
 FILLCELL_X32 FILLER_101_3551 ();
 FILLCELL_X32 FILLER_101_3583 ();
 FILLCELL_X32 FILLER_101_3615 ();
 FILLCELL_X32 FILLER_101_3647 ();
 FILLCELL_X32 FILLER_101_3679 ();
 FILLCELL_X16 FILLER_101_3711 ();
 FILLCELL_X8 FILLER_101_3727 ();
 FILLCELL_X2 FILLER_101_3735 ();
 FILLCELL_X1 FILLER_101_3737 ();
 FILLCELL_X32 FILLER_102_1 ();
 FILLCELL_X32 FILLER_102_33 ();
 FILLCELL_X32 FILLER_102_65 ();
 FILLCELL_X32 FILLER_102_97 ();
 FILLCELL_X32 FILLER_102_129 ();
 FILLCELL_X32 FILLER_102_161 ();
 FILLCELL_X32 FILLER_102_193 ();
 FILLCELL_X32 FILLER_102_225 ();
 FILLCELL_X32 FILLER_102_257 ();
 FILLCELL_X32 FILLER_102_289 ();
 FILLCELL_X32 FILLER_102_321 ();
 FILLCELL_X32 FILLER_102_353 ();
 FILLCELL_X32 FILLER_102_385 ();
 FILLCELL_X32 FILLER_102_417 ();
 FILLCELL_X32 FILLER_102_449 ();
 FILLCELL_X32 FILLER_102_481 ();
 FILLCELL_X32 FILLER_102_513 ();
 FILLCELL_X32 FILLER_102_545 ();
 FILLCELL_X32 FILLER_102_577 ();
 FILLCELL_X16 FILLER_102_609 ();
 FILLCELL_X4 FILLER_102_625 ();
 FILLCELL_X2 FILLER_102_629 ();
 FILLCELL_X32 FILLER_102_632 ();
 FILLCELL_X32 FILLER_102_664 ();
 FILLCELL_X32 FILLER_102_696 ();
 FILLCELL_X32 FILLER_102_728 ();
 FILLCELL_X32 FILLER_102_760 ();
 FILLCELL_X32 FILLER_102_792 ();
 FILLCELL_X32 FILLER_102_824 ();
 FILLCELL_X32 FILLER_102_856 ();
 FILLCELL_X32 FILLER_102_888 ();
 FILLCELL_X32 FILLER_102_920 ();
 FILLCELL_X32 FILLER_102_952 ();
 FILLCELL_X32 FILLER_102_984 ();
 FILLCELL_X32 FILLER_102_1016 ();
 FILLCELL_X32 FILLER_102_1048 ();
 FILLCELL_X32 FILLER_102_1080 ();
 FILLCELL_X32 FILLER_102_1112 ();
 FILLCELL_X32 FILLER_102_1144 ();
 FILLCELL_X32 FILLER_102_1176 ();
 FILLCELL_X32 FILLER_102_1208 ();
 FILLCELL_X32 FILLER_102_1240 ();
 FILLCELL_X32 FILLER_102_1272 ();
 FILLCELL_X32 FILLER_102_1304 ();
 FILLCELL_X32 FILLER_102_1336 ();
 FILLCELL_X32 FILLER_102_1368 ();
 FILLCELL_X32 FILLER_102_1400 ();
 FILLCELL_X32 FILLER_102_1432 ();
 FILLCELL_X32 FILLER_102_1464 ();
 FILLCELL_X32 FILLER_102_1496 ();
 FILLCELL_X32 FILLER_102_1528 ();
 FILLCELL_X32 FILLER_102_1560 ();
 FILLCELL_X32 FILLER_102_1592 ();
 FILLCELL_X32 FILLER_102_1624 ();
 FILLCELL_X32 FILLER_102_1656 ();
 FILLCELL_X32 FILLER_102_1688 ();
 FILLCELL_X32 FILLER_102_1720 ();
 FILLCELL_X32 FILLER_102_1752 ();
 FILLCELL_X32 FILLER_102_1784 ();
 FILLCELL_X32 FILLER_102_1816 ();
 FILLCELL_X32 FILLER_102_1848 ();
 FILLCELL_X8 FILLER_102_1880 ();
 FILLCELL_X4 FILLER_102_1888 ();
 FILLCELL_X2 FILLER_102_1892 ();
 FILLCELL_X32 FILLER_102_1895 ();
 FILLCELL_X32 FILLER_102_1927 ();
 FILLCELL_X32 FILLER_102_1959 ();
 FILLCELL_X32 FILLER_102_1991 ();
 FILLCELL_X32 FILLER_102_2023 ();
 FILLCELL_X32 FILLER_102_2055 ();
 FILLCELL_X32 FILLER_102_2087 ();
 FILLCELL_X32 FILLER_102_2119 ();
 FILLCELL_X32 FILLER_102_2151 ();
 FILLCELL_X32 FILLER_102_2183 ();
 FILLCELL_X32 FILLER_102_2215 ();
 FILLCELL_X32 FILLER_102_2247 ();
 FILLCELL_X32 FILLER_102_2279 ();
 FILLCELL_X32 FILLER_102_2311 ();
 FILLCELL_X32 FILLER_102_2343 ();
 FILLCELL_X32 FILLER_102_2375 ();
 FILLCELL_X32 FILLER_102_2407 ();
 FILLCELL_X32 FILLER_102_2439 ();
 FILLCELL_X32 FILLER_102_2471 ();
 FILLCELL_X32 FILLER_102_2503 ();
 FILLCELL_X32 FILLER_102_2535 ();
 FILLCELL_X32 FILLER_102_2567 ();
 FILLCELL_X32 FILLER_102_2599 ();
 FILLCELL_X32 FILLER_102_2631 ();
 FILLCELL_X32 FILLER_102_2663 ();
 FILLCELL_X32 FILLER_102_2695 ();
 FILLCELL_X32 FILLER_102_2727 ();
 FILLCELL_X32 FILLER_102_2759 ();
 FILLCELL_X32 FILLER_102_2791 ();
 FILLCELL_X32 FILLER_102_2823 ();
 FILLCELL_X32 FILLER_102_2855 ();
 FILLCELL_X32 FILLER_102_2887 ();
 FILLCELL_X32 FILLER_102_2919 ();
 FILLCELL_X32 FILLER_102_2951 ();
 FILLCELL_X32 FILLER_102_2983 ();
 FILLCELL_X32 FILLER_102_3015 ();
 FILLCELL_X32 FILLER_102_3047 ();
 FILLCELL_X32 FILLER_102_3079 ();
 FILLCELL_X32 FILLER_102_3111 ();
 FILLCELL_X8 FILLER_102_3143 ();
 FILLCELL_X4 FILLER_102_3151 ();
 FILLCELL_X2 FILLER_102_3155 ();
 FILLCELL_X32 FILLER_102_3158 ();
 FILLCELL_X32 FILLER_102_3190 ();
 FILLCELL_X32 FILLER_102_3222 ();
 FILLCELL_X32 FILLER_102_3254 ();
 FILLCELL_X32 FILLER_102_3286 ();
 FILLCELL_X32 FILLER_102_3318 ();
 FILLCELL_X32 FILLER_102_3350 ();
 FILLCELL_X32 FILLER_102_3382 ();
 FILLCELL_X32 FILLER_102_3414 ();
 FILLCELL_X32 FILLER_102_3446 ();
 FILLCELL_X32 FILLER_102_3478 ();
 FILLCELL_X32 FILLER_102_3510 ();
 FILLCELL_X32 FILLER_102_3542 ();
 FILLCELL_X32 FILLER_102_3574 ();
 FILLCELL_X32 FILLER_102_3606 ();
 FILLCELL_X32 FILLER_102_3638 ();
 FILLCELL_X32 FILLER_102_3670 ();
 FILLCELL_X32 FILLER_102_3702 ();
 FILLCELL_X4 FILLER_102_3734 ();
 FILLCELL_X32 FILLER_103_1 ();
 FILLCELL_X32 FILLER_103_33 ();
 FILLCELL_X32 FILLER_103_65 ();
 FILLCELL_X32 FILLER_103_97 ();
 FILLCELL_X32 FILLER_103_129 ();
 FILLCELL_X32 FILLER_103_161 ();
 FILLCELL_X32 FILLER_103_193 ();
 FILLCELL_X32 FILLER_103_225 ();
 FILLCELL_X32 FILLER_103_257 ();
 FILLCELL_X32 FILLER_103_289 ();
 FILLCELL_X32 FILLER_103_321 ();
 FILLCELL_X32 FILLER_103_353 ();
 FILLCELL_X32 FILLER_103_385 ();
 FILLCELL_X32 FILLER_103_417 ();
 FILLCELL_X32 FILLER_103_449 ();
 FILLCELL_X32 FILLER_103_481 ();
 FILLCELL_X32 FILLER_103_513 ();
 FILLCELL_X32 FILLER_103_545 ();
 FILLCELL_X32 FILLER_103_577 ();
 FILLCELL_X32 FILLER_103_609 ();
 FILLCELL_X32 FILLER_103_641 ();
 FILLCELL_X32 FILLER_103_673 ();
 FILLCELL_X32 FILLER_103_705 ();
 FILLCELL_X32 FILLER_103_737 ();
 FILLCELL_X32 FILLER_103_769 ();
 FILLCELL_X32 FILLER_103_801 ();
 FILLCELL_X32 FILLER_103_833 ();
 FILLCELL_X32 FILLER_103_865 ();
 FILLCELL_X32 FILLER_103_897 ();
 FILLCELL_X32 FILLER_103_929 ();
 FILLCELL_X32 FILLER_103_961 ();
 FILLCELL_X32 FILLER_103_993 ();
 FILLCELL_X32 FILLER_103_1025 ();
 FILLCELL_X32 FILLER_103_1057 ();
 FILLCELL_X32 FILLER_103_1089 ();
 FILLCELL_X32 FILLER_103_1121 ();
 FILLCELL_X32 FILLER_103_1153 ();
 FILLCELL_X32 FILLER_103_1185 ();
 FILLCELL_X32 FILLER_103_1217 ();
 FILLCELL_X8 FILLER_103_1249 ();
 FILLCELL_X4 FILLER_103_1257 ();
 FILLCELL_X2 FILLER_103_1261 ();
 FILLCELL_X32 FILLER_103_1264 ();
 FILLCELL_X32 FILLER_103_1296 ();
 FILLCELL_X32 FILLER_103_1328 ();
 FILLCELL_X32 FILLER_103_1360 ();
 FILLCELL_X32 FILLER_103_1392 ();
 FILLCELL_X32 FILLER_103_1424 ();
 FILLCELL_X32 FILLER_103_1456 ();
 FILLCELL_X32 FILLER_103_1488 ();
 FILLCELL_X32 FILLER_103_1520 ();
 FILLCELL_X32 FILLER_103_1552 ();
 FILLCELL_X32 FILLER_103_1584 ();
 FILLCELL_X32 FILLER_103_1616 ();
 FILLCELL_X32 FILLER_103_1648 ();
 FILLCELL_X32 FILLER_103_1680 ();
 FILLCELL_X32 FILLER_103_1712 ();
 FILLCELL_X32 FILLER_103_1744 ();
 FILLCELL_X32 FILLER_103_1776 ();
 FILLCELL_X32 FILLER_103_1808 ();
 FILLCELL_X32 FILLER_103_1840 ();
 FILLCELL_X32 FILLER_103_1872 ();
 FILLCELL_X32 FILLER_103_1904 ();
 FILLCELL_X32 FILLER_103_1936 ();
 FILLCELL_X32 FILLER_103_1968 ();
 FILLCELL_X32 FILLER_103_2000 ();
 FILLCELL_X32 FILLER_103_2032 ();
 FILLCELL_X32 FILLER_103_2064 ();
 FILLCELL_X32 FILLER_103_2096 ();
 FILLCELL_X32 FILLER_103_2128 ();
 FILLCELL_X32 FILLER_103_2160 ();
 FILLCELL_X32 FILLER_103_2192 ();
 FILLCELL_X32 FILLER_103_2224 ();
 FILLCELL_X32 FILLER_103_2256 ();
 FILLCELL_X32 FILLER_103_2288 ();
 FILLCELL_X32 FILLER_103_2320 ();
 FILLCELL_X32 FILLER_103_2352 ();
 FILLCELL_X32 FILLER_103_2384 ();
 FILLCELL_X32 FILLER_103_2416 ();
 FILLCELL_X32 FILLER_103_2448 ();
 FILLCELL_X32 FILLER_103_2480 ();
 FILLCELL_X8 FILLER_103_2512 ();
 FILLCELL_X4 FILLER_103_2520 ();
 FILLCELL_X2 FILLER_103_2524 ();
 FILLCELL_X32 FILLER_103_2527 ();
 FILLCELL_X32 FILLER_103_2559 ();
 FILLCELL_X32 FILLER_103_2591 ();
 FILLCELL_X32 FILLER_103_2623 ();
 FILLCELL_X32 FILLER_103_2655 ();
 FILLCELL_X32 FILLER_103_2687 ();
 FILLCELL_X32 FILLER_103_2719 ();
 FILLCELL_X32 FILLER_103_2751 ();
 FILLCELL_X32 FILLER_103_2783 ();
 FILLCELL_X32 FILLER_103_2815 ();
 FILLCELL_X32 FILLER_103_2847 ();
 FILLCELL_X32 FILLER_103_2879 ();
 FILLCELL_X32 FILLER_103_2911 ();
 FILLCELL_X32 FILLER_103_2943 ();
 FILLCELL_X32 FILLER_103_2975 ();
 FILLCELL_X32 FILLER_103_3007 ();
 FILLCELL_X32 FILLER_103_3039 ();
 FILLCELL_X32 FILLER_103_3071 ();
 FILLCELL_X32 FILLER_103_3103 ();
 FILLCELL_X32 FILLER_103_3135 ();
 FILLCELL_X32 FILLER_103_3167 ();
 FILLCELL_X32 FILLER_103_3199 ();
 FILLCELL_X32 FILLER_103_3231 ();
 FILLCELL_X32 FILLER_103_3263 ();
 FILLCELL_X32 FILLER_103_3295 ();
 FILLCELL_X32 FILLER_103_3327 ();
 FILLCELL_X32 FILLER_103_3359 ();
 FILLCELL_X32 FILLER_103_3391 ();
 FILLCELL_X32 FILLER_103_3423 ();
 FILLCELL_X32 FILLER_103_3455 ();
 FILLCELL_X32 FILLER_103_3487 ();
 FILLCELL_X32 FILLER_103_3519 ();
 FILLCELL_X32 FILLER_103_3551 ();
 FILLCELL_X32 FILLER_103_3583 ();
 FILLCELL_X32 FILLER_103_3615 ();
 FILLCELL_X32 FILLER_103_3647 ();
 FILLCELL_X32 FILLER_103_3679 ();
 FILLCELL_X16 FILLER_103_3711 ();
 FILLCELL_X8 FILLER_103_3727 ();
 FILLCELL_X2 FILLER_103_3735 ();
 FILLCELL_X1 FILLER_103_3737 ();
 FILLCELL_X32 FILLER_104_1 ();
 FILLCELL_X32 FILLER_104_33 ();
 FILLCELL_X32 FILLER_104_65 ();
 FILLCELL_X32 FILLER_104_97 ();
 FILLCELL_X32 FILLER_104_129 ();
 FILLCELL_X32 FILLER_104_161 ();
 FILLCELL_X32 FILLER_104_193 ();
 FILLCELL_X32 FILLER_104_225 ();
 FILLCELL_X32 FILLER_104_257 ();
 FILLCELL_X32 FILLER_104_289 ();
 FILLCELL_X32 FILLER_104_321 ();
 FILLCELL_X32 FILLER_104_353 ();
 FILLCELL_X32 FILLER_104_385 ();
 FILLCELL_X32 FILLER_104_417 ();
 FILLCELL_X32 FILLER_104_449 ();
 FILLCELL_X32 FILLER_104_481 ();
 FILLCELL_X32 FILLER_104_513 ();
 FILLCELL_X32 FILLER_104_545 ();
 FILLCELL_X32 FILLER_104_577 ();
 FILLCELL_X16 FILLER_104_609 ();
 FILLCELL_X4 FILLER_104_625 ();
 FILLCELL_X2 FILLER_104_629 ();
 FILLCELL_X32 FILLER_104_632 ();
 FILLCELL_X32 FILLER_104_664 ();
 FILLCELL_X32 FILLER_104_696 ();
 FILLCELL_X32 FILLER_104_728 ();
 FILLCELL_X32 FILLER_104_760 ();
 FILLCELL_X32 FILLER_104_792 ();
 FILLCELL_X32 FILLER_104_824 ();
 FILLCELL_X32 FILLER_104_856 ();
 FILLCELL_X32 FILLER_104_888 ();
 FILLCELL_X32 FILLER_104_920 ();
 FILLCELL_X32 FILLER_104_952 ();
 FILLCELL_X32 FILLER_104_984 ();
 FILLCELL_X32 FILLER_104_1016 ();
 FILLCELL_X32 FILLER_104_1048 ();
 FILLCELL_X32 FILLER_104_1080 ();
 FILLCELL_X32 FILLER_104_1112 ();
 FILLCELL_X32 FILLER_104_1144 ();
 FILLCELL_X32 FILLER_104_1176 ();
 FILLCELL_X32 FILLER_104_1208 ();
 FILLCELL_X32 FILLER_104_1240 ();
 FILLCELL_X32 FILLER_104_1272 ();
 FILLCELL_X32 FILLER_104_1304 ();
 FILLCELL_X32 FILLER_104_1336 ();
 FILLCELL_X32 FILLER_104_1368 ();
 FILLCELL_X32 FILLER_104_1400 ();
 FILLCELL_X32 FILLER_104_1432 ();
 FILLCELL_X32 FILLER_104_1464 ();
 FILLCELL_X32 FILLER_104_1496 ();
 FILLCELL_X32 FILLER_104_1528 ();
 FILLCELL_X32 FILLER_104_1560 ();
 FILLCELL_X32 FILLER_104_1592 ();
 FILLCELL_X32 FILLER_104_1624 ();
 FILLCELL_X32 FILLER_104_1656 ();
 FILLCELL_X32 FILLER_104_1688 ();
 FILLCELL_X32 FILLER_104_1720 ();
 FILLCELL_X32 FILLER_104_1752 ();
 FILLCELL_X32 FILLER_104_1784 ();
 FILLCELL_X32 FILLER_104_1816 ();
 FILLCELL_X32 FILLER_104_1848 ();
 FILLCELL_X8 FILLER_104_1880 ();
 FILLCELL_X4 FILLER_104_1888 ();
 FILLCELL_X2 FILLER_104_1892 ();
 FILLCELL_X32 FILLER_104_1895 ();
 FILLCELL_X32 FILLER_104_1927 ();
 FILLCELL_X32 FILLER_104_1959 ();
 FILLCELL_X32 FILLER_104_1991 ();
 FILLCELL_X32 FILLER_104_2023 ();
 FILLCELL_X32 FILLER_104_2055 ();
 FILLCELL_X32 FILLER_104_2087 ();
 FILLCELL_X32 FILLER_104_2119 ();
 FILLCELL_X32 FILLER_104_2151 ();
 FILLCELL_X32 FILLER_104_2183 ();
 FILLCELL_X32 FILLER_104_2215 ();
 FILLCELL_X32 FILLER_104_2247 ();
 FILLCELL_X32 FILLER_104_2279 ();
 FILLCELL_X32 FILLER_104_2311 ();
 FILLCELL_X32 FILLER_104_2343 ();
 FILLCELL_X32 FILLER_104_2375 ();
 FILLCELL_X32 FILLER_104_2407 ();
 FILLCELL_X32 FILLER_104_2439 ();
 FILLCELL_X32 FILLER_104_2471 ();
 FILLCELL_X32 FILLER_104_2503 ();
 FILLCELL_X32 FILLER_104_2535 ();
 FILLCELL_X32 FILLER_104_2567 ();
 FILLCELL_X32 FILLER_104_2599 ();
 FILLCELL_X32 FILLER_104_2631 ();
 FILLCELL_X32 FILLER_104_2663 ();
 FILLCELL_X32 FILLER_104_2695 ();
 FILLCELL_X32 FILLER_104_2727 ();
 FILLCELL_X32 FILLER_104_2759 ();
 FILLCELL_X32 FILLER_104_2791 ();
 FILLCELL_X32 FILLER_104_2823 ();
 FILLCELL_X32 FILLER_104_2855 ();
 FILLCELL_X32 FILLER_104_2887 ();
 FILLCELL_X32 FILLER_104_2919 ();
 FILLCELL_X32 FILLER_104_2951 ();
 FILLCELL_X32 FILLER_104_2983 ();
 FILLCELL_X32 FILLER_104_3015 ();
 FILLCELL_X32 FILLER_104_3047 ();
 FILLCELL_X32 FILLER_104_3079 ();
 FILLCELL_X32 FILLER_104_3111 ();
 FILLCELL_X8 FILLER_104_3143 ();
 FILLCELL_X4 FILLER_104_3151 ();
 FILLCELL_X2 FILLER_104_3155 ();
 FILLCELL_X32 FILLER_104_3158 ();
 FILLCELL_X32 FILLER_104_3190 ();
 FILLCELL_X32 FILLER_104_3222 ();
 FILLCELL_X32 FILLER_104_3254 ();
 FILLCELL_X32 FILLER_104_3286 ();
 FILLCELL_X32 FILLER_104_3318 ();
 FILLCELL_X32 FILLER_104_3350 ();
 FILLCELL_X32 FILLER_104_3382 ();
 FILLCELL_X32 FILLER_104_3414 ();
 FILLCELL_X32 FILLER_104_3446 ();
 FILLCELL_X32 FILLER_104_3478 ();
 FILLCELL_X32 FILLER_104_3510 ();
 FILLCELL_X32 FILLER_104_3542 ();
 FILLCELL_X32 FILLER_104_3574 ();
 FILLCELL_X32 FILLER_104_3606 ();
 FILLCELL_X32 FILLER_104_3638 ();
 FILLCELL_X32 FILLER_104_3670 ();
 FILLCELL_X32 FILLER_104_3702 ();
 FILLCELL_X4 FILLER_104_3734 ();
 FILLCELL_X32 FILLER_105_1 ();
 FILLCELL_X32 FILLER_105_33 ();
 FILLCELL_X32 FILLER_105_65 ();
 FILLCELL_X32 FILLER_105_97 ();
 FILLCELL_X32 FILLER_105_129 ();
 FILLCELL_X32 FILLER_105_161 ();
 FILLCELL_X32 FILLER_105_193 ();
 FILLCELL_X32 FILLER_105_225 ();
 FILLCELL_X32 FILLER_105_257 ();
 FILLCELL_X32 FILLER_105_289 ();
 FILLCELL_X32 FILLER_105_321 ();
 FILLCELL_X32 FILLER_105_353 ();
 FILLCELL_X32 FILLER_105_385 ();
 FILLCELL_X32 FILLER_105_417 ();
 FILLCELL_X32 FILLER_105_449 ();
 FILLCELL_X32 FILLER_105_481 ();
 FILLCELL_X32 FILLER_105_513 ();
 FILLCELL_X32 FILLER_105_545 ();
 FILLCELL_X32 FILLER_105_577 ();
 FILLCELL_X32 FILLER_105_609 ();
 FILLCELL_X32 FILLER_105_641 ();
 FILLCELL_X32 FILLER_105_673 ();
 FILLCELL_X32 FILLER_105_705 ();
 FILLCELL_X32 FILLER_105_737 ();
 FILLCELL_X32 FILLER_105_769 ();
 FILLCELL_X32 FILLER_105_801 ();
 FILLCELL_X32 FILLER_105_833 ();
 FILLCELL_X32 FILLER_105_865 ();
 FILLCELL_X32 FILLER_105_897 ();
 FILLCELL_X32 FILLER_105_929 ();
 FILLCELL_X32 FILLER_105_961 ();
 FILLCELL_X32 FILLER_105_993 ();
 FILLCELL_X32 FILLER_105_1025 ();
 FILLCELL_X32 FILLER_105_1057 ();
 FILLCELL_X32 FILLER_105_1089 ();
 FILLCELL_X32 FILLER_105_1121 ();
 FILLCELL_X32 FILLER_105_1153 ();
 FILLCELL_X32 FILLER_105_1185 ();
 FILLCELL_X32 FILLER_105_1217 ();
 FILLCELL_X8 FILLER_105_1249 ();
 FILLCELL_X4 FILLER_105_1257 ();
 FILLCELL_X2 FILLER_105_1261 ();
 FILLCELL_X32 FILLER_105_1264 ();
 FILLCELL_X32 FILLER_105_1296 ();
 FILLCELL_X32 FILLER_105_1328 ();
 FILLCELL_X32 FILLER_105_1360 ();
 FILLCELL_X32 FILLER_105_1392 ();
 FILLCELL_X32 FILLER_105_1424 ();
 FILLCELL_X32 FILLER_105_1456 ();
 FILLCELL_X32 FILLER_105_1488 ();
 FILLCELL_X32 FILLER_105_1520 ();
 FILLCELL_X32 FILLER_105_1552 ();
 FILLCELL_X32 FILLER_105_1584 ();
 FILLCELL_X32 FILLER_105_1616 ();
 FILLCELL_X32 FILLER_105_1648 ();
 FILLCELL_X32 FILLER_105_1680 ();
 FILLCELL_X32 FILLER_105_1712 ();
 FILLCELL_X32 FILLER_105_1744 ();
 FILLCELL_X32 FILLER_105_1776 ();
 FILLCELL_X32 FILLER_105_1808 ();
 FILLCELL_X32 FILLER_105_1840 ();
 FILLCELL_X32 FILLER_105_1872 ();
 FILLCELL_X32 FILLER_105_1904 ();
 FILLCELL_X32 FILLER_105_1936 ();
 FILLCELL_X32 FILLER_105_1968 ();
 FILLCELL_X32 FILLER_105_2000 ();
 FILLCELL_X32 FILLER_105_2032 ();
 FILLCELL_X32 FILLER_105_2064 ();
 FILLCELL_X32 FILLER_105_2096 ();
 FILLCELL_X32 FILLER_105_2128 ();
 FILLCELL_X32 FILLER_105_2160 ();
 FILLCELL_X32 FILLER_105_2192 ();
 FILLCELL_X32 FILLER_105_2224 ();
 FILLCELL_X32 FILLER_105_2256 ();
 FILLCELL_X32 FILLER_105_2288 ();
 FILLCELL_X32 FILLER_105_2320 ();
 FILLCELL_X32 FILLER_105_2352 ();
 FILLCELL_X32 FILLER_105_2384 ();
 FILLCELL_X32 FILLER_105_2416 ();
 FILLCELL_X32 FILLER_105_2448 ();
 FILLCELL_X32 FILLER_105_2480 ();
 FILLCELL_X8 FILLER_105_2512 ();
 FILLCELL_X4 FILLER_105_2520 ();
 FILLCELL_X2 FILLER_105_2524 ();
 FILLCELL_X32 FILLER_105_2527 ();
 FILLCELL_X32 FILLER_105_2559 ();
 FILLCELL_X32 FILLER_105_2591 ();
 FILLCELL_X32 FILLER_105_2623 ();
 FILLCELL_X32 FILLER_105_2655 ();
 FILLCELL_X32 FILLER_105_2687 ();
 FILLCELL_X32 FILLER_105_2719 ();
 FILLCELL_X32 FILLER_105_2751 ();
 FILLCELL_X32 FILLER_105_2783 ();
 FILLCELL_X32 FILLER_105_2815 ();
 FILLCELL_X32 FILLER_105_2847 ();
 FILLCELL_X32 FILLER_105_2879 ();
 FILLCELL_X32 FILLER_105_2911 ();
 FILLCELL_X32 FILLER_105_2943 ();
 FILLCELL_X32 FILLER_105_2975 ();
 FILLCELL_X32 FILLER_105_3007 ();
 FILLCELL_X32 FILLER_105_3039 ();
 FILLCELL_X32 FILLER_105_3071 ();
 FILLCELL_X32 FILLER_105_3103 ();
 FILLCELL_X32 FILLER_105_3135 ();
 FILLCELL_X32 FILLER_105_3167 ();
 FILLCELL_X32 FILLER_105_3199 ();
 FILLCELL_X32 FILLER_105_3231 ();
 FILLCELL_X32 FILLER_105_3263 ();
 FILLCELL_X32 FILLER_105_3295 ();
 FILLCELL_X32 FILLER_105_3327 ();
 FILLCELL_X32 FILLER_105_3359 ();
 FILLCELL_X32 FILLER_105_3391 ();
 FILLCELL_X32 FILLER_105_3423 ();
 FILLCELL_X32 FILLER_105_3455 ();
 FILLCELL_X32 FILLER_105_3487 ();
 FILLCELL_X32 FILLER_105_3519 ();
 FILLCELL_X32 FILLER_105_3551 ();
 FILLCELL_X32 FILLER_105_3583 ();
 FILLCELL_X32 FILLER_105_3615 ();
 FILLCELL_X32 FILLER_105_3647 ();
 FILLCELL_X32 FILLER_105_3679 ();
 FILLCELL_X16 FILLER_105_3711 ();
 FILLCELL_X8 FILLER_105_3727 ();
 FILLCELL_X2 FILLER_105_3735 ();
 FILLCELL_X1 FILLER_105_3737 ();
 FILLCELL_X32 FILLER_106_1 ();
 FILLCELL_X32 FILLER_106_33 ();
 FILLCELL_X32 FILLER_106_65 ();
 FILLCELL_X32 FILLER_106_97 ();
 FILLCELL_X32 FILLER_106_129 ();
 FILLCELL_X32 FILLER_106_161 ();
 FILLCELL_X32 FILLER_106_193 ();
 FILLCELL_X32 FILLER_106_225 ();
 FILLCELL_X32 FILLER_106_257 ();
 FILLCELL_X32 FILLER_106_289 ();
 FILLCELL_X32 FILLER_106_321 ();
 FILLCELL_X32 FILLER_106_353 ();
 FILLCELL_X32 FILLER_106_385 ();
 FILLCELL_X32 FILLER_106_417 ();
 FILLCELL_X32 FILLER_106_449 ();
 FILLCELL_X32 FILLER_106_481 ();
 FILLCELL_X32 FILLER_106_513 ();
 FILLCELL_X32 FILLER_106_545 ();
 FILLCELL_X32 FILLER_106_577 ();
 FILLCELL_X16 FILLER_106_609 ();
 FILLCELL_X4 FILLER_106_625 ();
 FILLCELL_X2 FILLER_106_629 ();
 FILLCELL_X32 FILLER_106_632 ();
 FILLCELL_X32 FILLER_106_664 ();
 FILLCELL_X32 FILLER_106_696 ();
 FILLCELL_X32 FILLER_106_728 ();
 FILLCELL_X32 FILLER_106_760 ();
 FILLCELL_X32 FILLER_106_792 ();
 FILLCELL_X32 FILLER_106_824 ();
 FILLCELL_X32 FILLER_106_856 ();
 FILLCELL_X32 FILLER_106_888 ();
 FILLCELL_X32 FILLER_106_920 ();
 FILLCELL_X32 FILLER_106_952 ();
 FILLCELL_X32 FILLER_106_984 ();
 FILLCELL_X32 FILLER_106_1016 ();
 FILLCELL_X32 FILLER_106_1048 ();
 FILLCELL_X32 FILLER_106_1080 ();
 FILLCELL_X32 FILLER_106_1112 ();
 FILLCELL_X32 FILLER_106_1144 ();
 FILLCELL_X32 FILLER_106_1176 ();
 FILLCELL_X32 FILLER_106_1208 ();
 FILLCELL_X32 FILLER_106_1240 ();
 FILLCELL_X32 FILLER_106_1272 ();
 FILLCELL_X32 FILLER_106_1304 ();
 FILLCELL_X32 FILLER_106_1336 ();
 FILLCELL_X32 FILLER_106_1368 ();
 FILLCELL_X32 FILLER_106_1400 ();
 FILLCELL_X32 FILLER_106_1432 ();
 FILLCELL_X32 FILLER_106_1464 ();
 FILLCELL_X32 FILLER_106_1496 ();
 FILLCELL_X32 FILLER_106_1528 ();
 FILLCELL_X32 FILLER_106_1560 ();
 FILLCELL_X32 FILLER_106_1592 ();
 FILLCELL_X32 FILLER_106_1624 ();
 FILLCELL_X32 FILLER_106_1656 ();
 FILLCELL_X32 FILLER_106_1688 ();
 FILLCELL_X32 FILLER_106_1720 ();
 FILLCELL_X32 FILLER_106_1752 ();
 FILLCELL_X32 FILLER_106_1784 ();
 FILLCELL_X32 FILLER_106_1816 ();
 FILLCELL_X32 FILLER_106_1848 ();
 FILLCELL_X8 FILLER_106_1880 ();
 FILLCELL_X4 FILLER_106_1888 ();
 FILLCELL_X2 FILLER_106_1892 ();
 FILLCELL_X32 FILLER_106_1895 ();
 FILLCELL_X32 FILLER_106_1927 ();
 FILLCELL_X32 FILLER_106_1959 ();
 FILLCELL_X32 FILLER_106_1991 ();
 FILLCELL_X32 FILLER_106_2023 ();
 FILLCELL_X32 FILLER_106_2055 ();
 FILLCELL_X32 FILLER_106_2087 ();
 FILLCELL_X32 FILLER_106_2119 ();
 FILLCELL_X32 FILLER_106_2151 ();
 FILLCELL_X32 FILLER_106_2183 ();
 FILLCELL_X32 FILLER_106_2215 ();
 FILLCELL_X32 FILLER_106_2247 ();
 FILLCELL_X32 FILLER_106_2279 ();
 FILLCELL_X32 FILLER_106_2311 ();
 FILLCELL_X32 FILLER_106_2343 ();
 FILLCELL_X32 FILLER_106_2375 ();
 FILLCELL_X32 FILLER_106_2407 ();
 FILLCELL_X32 FILLER_106_2439 ();
 FILLCELL_X32 FILLER_106_2471 ();
 FILLCELL_X32 FILLER_106_2503 ();
 FILLCELL_X32 FILLER_106_2535 ();
 FILLCELL_X32 FILLER_106_2567 ();
 FILLCELL_X32 FILLER_106_2599 ();
 FILLCELL_X32 FILLER_106_2631 ();
 FILLCELL_X32 FILLER_106_2663 ();
 FILLCELL_X32 FILLER_106_2695 ();
 FILLCELL_X32 FILLER_106_2727 ();
 FILLCELL_X32 FILLER_106_2759 ();
 FILLCELL_X32 FILLER_106_2791 ();
 FILLCELL_X32 FILLER_106_2823 ();
 FILLCELL_X32 FILLER_106_2855 ();
 FILLCELL_X32 FILLER_106_2887 ();
 FILLCELL_X32 FILLER_106_2919 ();
 FILLCELL_X32 FILLER_106_2951 ();
 FILLCELL_X32 FILLER_106_2983 ();
 FILLCELL_X32 FILLER_106_3015 ();
 FILLCELL_X32 FILLER_106_3047 ();
 FILLCELL_X32 FILLER_106_3079 ();
 FILLCELL_X32 FILLER_106_3111 ();
 FILLCELL_X8 FILLER_106_3143 ();
 FILLCELL_X4 FILLER_106_3151 ();
 FILLCELL_X2 FILLER_106_3155 ();
 FILLCELL_X32 FILLER_106_3158 ();
 FILLCELL_X32 FILLER_106_3190 ();
 FILLCELL_X32 FILLER_106_3222 ();
 FILLCELL_X32 FILLER_106_3254 ();
 FILLCELL_X32 FILLER_106_3286 ();
 FILLCELL_X32 FILLER_106_3318 ();
 FILLCELL_X32 FILLER_106_3350 ();
 FILLCELL_X32 FILLER_106_3382 ();
 FILLCELL_X32 FILLER_106_3414 ();
 FILLCELL_X32 FILLER_106_3446 ();
 FILLCELL_X32 FILLER_106_3478 ();
 FILLCELL_X32 FILLER_106_3510 ();
 FILLCELL_X32 FILLER_106_3542 ();
 FILLCELL_X32 FILLER_106_3574 ();
 FILLCELL_X32 FILLER_106_3606 ();
 FILLCELL_X32 FILLER_106_3638 ();
 FILLCELL_X32 FILLER_106_3670 ();
 FILLCELL_X32 FILLER_106_3702 ();
 FILLCELL_X4 FILLER_106_3734 ();
 FILLCELL_X32 FILLER_107_1 ();
 FILLCELL_X32 FILLER_107_33 ();
 FILLCELL_X32 FILLER_107_65 ();
 FILLCELL_X32 FILLER_107_97 ();
 FILLCELL_X32 FILLER_107_129 ();
 FILLCELL_X32 FILLER_107_161 ();
 FILLCELL_X32 FILLER_107_193 ();
 FILLCELL_X32 FILLER_107_225 ();
 FILLCELL_X32 FILLER_107_257 ();
 FILLCELL_X32 FILLER_107_289 ();
 FILLCELL_X32 FILLER_107_321 ();
 FILLCELL_X32 FILLER_107_353 ();
 FILLCELL_X32 FILLER_107_385 ();
 FILLCELL_X32 FILLER_107_417 ();
 FILLCELL_X32 FILLER_107_449 ();
 FILLCELL_X32 FILLER_107_481 ();
 FILLCELL_X32 FILLER_107_513 ();
 FILLCELL_X32 FILLER_107_545 ();
 FILLCELL_X32 FILLER_107_577 ();
 FILLCELL_X32 FILLER_107_609 ();
 FILLCELL_X32 FILLER_107_641 ();
 FILLCELL_X32 FILLER_107_673 ();
 FILLCELL_X32 FILLER_107_705 ();
 FILLCELL_X32 FILLER_107_737 ();
 FILLCELL_X32 FILLER_107_769 ();
 FILLCELL_X32 FILLER_107_801 ();
 FILLCELL_X32 FILLER_107_833 ();
 FILLCELL_X32 FILLER_107_865 ();
 FILLCELL_X32 FILLER_107_897 ();
 FILLCELL_X32 FILLER_107_929 ();
 FILLCELL_X32 FILLER_107_961 ();
 FILLCELL_X32 FILLER_107_993 ();
 FILLCELL_X32 FILLER_107_1025 ();
 FILLCELL_X32 FILLER_107_1057 ();
 FILLCELL_X32 FILLER_107_1089 ();
 FILLCELL_X32 FILLER_107_1121 ();
 FILLCELL_X32 FILLER_107_1153 ();
 FILLCELL_X32 FILLER_107_1185 ();
 FILLCELL_X32 FILLER_107_1217 ();
 FILLCELL_X8 FILLER_107_1249 ();
 FILLCELL_X4 FILLER_107_1257 ();
 FILLCELL_X2 FILLER_107_1261 ();
 FILLCELL_X32 FILLER_107_1264 ();
 FILLCELL_X32 FILLER_107_1296 ();
 FILLCELL_X32 FILLER_107_1328 ();
 FILLCELL_X32 FILLER_107_1360 ();
 FILLCELL_X32 FILLER_107_1392 ();
 FILLCELL_X32 FILLER_107_1424 ();
 FILLCELL_X32 FILLER_107_1456 ();
 FILLCELL_X32 FILLER_107_1488 ();
 FILLCELL_X32 FILLER_107_1520 ();
 FILLCELL_X32 FILLER_107_1552 ();
 FILLCELL_X32 FILLER_107_1584 ();
 FILLCELL_X32 FILLER_107_1616 ();
 FILLCELL_X32 FILLER_107_1648 ();
 FILLCELL_X32 FILLER_107_1680 ();
 FILLCELL_X32 FILLER_107_1712 ();
 FILLCELL_X32 FILLER_107_1744 ();
 FILLCELL_X32 FILLER_107_1776 ();
 FILLCELL_X32 FILLER_107_1808 ();
 FILLCELL_X32 FILLER_107_1840 ();
 FILLCELL_X32 FILLER_107_1872 ();
 FILLCELL_X32 FILLER_107_1904 ();
 FILLCELL_X32 FILLER_107_1936 ();
 FILLCELL_X32 FILLER_107_1968 ();
 FILLCELL_X32 FILLER_107_2000 ();
 FILLCELL_X32 FILLER_107_2032 ();
 FILLCELL_X32 FILLER_107_2064 ();
 FILLCELL_X32 FILLER_107_2096 ();
 FILLCELL_X32 FILLER_107_2128 ();
 FILLCELL_X32 FILLER_107_2160 ();
 FILLCELL_X32 FILLER_107_2192 ();
 FILLCELL_X32 FILLER_107_2224 ();
 FILLCELL_X32 FILLER_107_2256 ();
 FILLCELL_X32 FILLER_107_2288 ();
 FILLCELL_X32 FILLER_107_2320 ();
 FILLCELL_X32 FILLER_107_2352 ();
 FILLCELL_X32 FILLER_107_2384 ();
 FILLCELL_X32 FILLER_107_2416 ();
 FILLCELL_X32 FILLER_107_2448 ();
 FILLCELL_X32 FILLER_107_2480 ();
 FILLCELL_X8 FILLER_107_2512 ();
 FILLCELL_X4 FILLER_107_2520 ();
 FILLCELL_X2 FILLER_107_2524 ();
 FILLCELL_X32 FILLER_107_2527 ();
 FILLCELL_X32 FILLER_107_2559 ();
 FILLCELL_X32 FILLER_107_2591 ();
 FILLCELL_X32 FILLER_107_2623 ();
 FILLCELL_X32 FILLER_107_2655 ();
 FILLCELL_X32 FILLER_107_2687 ();
 FILLCELL_X32 FILLER_107_2719 ();
 FILLCELL_X32 FILLER_107_2751 ();
 FILLCELL_X32 FILLER_107_2783 ();
 FILLCELL_X32 FILLER_107_2815 ();
 FILLCELL_X32 FILLER_107_2847 ();
 FILLCELL_X32 FILLER_107_2879 ();
 FILLCELL_X32 FILLER_107_2911 ();
 FILLCELL_X32 FILLER_107_2943 ();
 FILLCELL_X32 FILLER_107_2975 ();
 FILLCELL_X32 FILLER_107_3007 ();
 FILLCELL_X32 FILLER_107_3039 ();
 FILLCELL_X32 FILLER_107_3071 ();
 FILLCELL_X32 FILLER_107_3103 ();
 FILLCELL_X32 FILLER_107_3135 ();
 FILLCELL_X32 FILLER_107_3167 ();
 FILLCELL_X32 FILLER_107_3199 ();
 FILLCELL_X32 FILLER_107_3231 ();
 FILLCELL_X32 FILLER_107_3263 ();
 FILLCELL_X32 FILLER_107_3295 ();
 FILLCELL_X32 FILLER_107_3327 ();
 FILLCELL_X32 FILLER_107_3359 ();
 FILLCELL_X32 FILLER_107_3391 ();
 FILLCELL_X32 FILLER_107_3423 ();
 FILLCELL_X32 FILLER_107_3455 ();
 FILLCELL_X32 FILLER_107_3487 ();
 FILLCELL_X32 FILLER_107_3519 ();
 FILLCELL_X32 FILLER_107_3551 ();
 FILLCELL_X32 FILLER_107_3583 ();
 FILLCELL_X32 FILLER_107_3615 ();
 FILLCELL_X32 FILLER_107_3647 ();
 FILLCELL_X32 FILLER_107_3679 ();
 FILLCELL_X16 FILLER_107_3711 ();
 FILLCELL_X8 FILLER_107_3727 ();
 FILLCELL_X2 FILLER_107_3735 ();
 FILLCELL_X1 FILLER_107_3737 ();
 FILLCELL_X32 FILLER_108_1 ();
 FILLCELL_X32 FILLER_108_33 ();
 FILLCELL_X32 FILLER_108_65 ();
 FILLCELL_X32 FILLER_108_97 ();
 FILLCELL_X32 FILLER_108_129 ();
 FILLCELL_X32 FILLER_108_161 ();
 FILLCELL_X32 FILLER_108_193 ();
 FILLCELL_X32 FILLER_108_225 ();
 FILLCELL_X32 FILLER_108_257 ();
 FILLCELL_X32 FILLER_108_289 ();
 FILLCELL_X32 FILLER_108_321 ();
 FILLCELL_X32 FILLER_108_353 ();
 FILLCELL_X32 FILLER_108_385 ();
 FILLCELL_X32 FILLER_108_417 ();
 FILLCELL_X32 FILLER_108_449 ();
 FILLCELL_X32 FILLER_108_481 ();
 FILLCELL_X32 FILLER_108_513 ();
 FILLCELL_X32 FILLER_108_545 ();
 FILLCELL_X32 FILLER_108_577 ();
 FILLCELL_X16 FILLER_108_609 ();
 FILLCELL_X4 FILLER_108_625 ();
 FILLCELL_X2 FILLER_108_629 ();
 FILLCELL_X32 FILLER_108_632 ();
 FILLCELL_X32 FILLER_108_664 ();
 FILLCELL_X32 FILLER_108_696 ();
 FILLCELL_X32 FILLER_108_728 ();
 FILLCELL_X32 FILLER_108_760 ();
 FILLCELL_X32 FILLER_108_792 ();
 FILLCELL_X32 FILLER_108_824 ();
 FILLCELL_X32 FILLER_108_856 ();
 FILLCELL_X32 FILLER_108_888 ();
 FILLCELL_X32 FILLER_108_920 ();
 FILLCELL_X32 FILLER_108_952 ();
 FILLCELL_X32 FILLER_108_984 ();
 FILLCELL_X32 FILLER_108_1016 ();
 FILLCELL_X32 FILLER_108_1048 ();
 FILLCELL_X32 FILLER_108_1080 ();
 FILLCELL_X32 FILLER_108_1112 ();
 FILLCELL_X32 FILLER_108_1144 ();
 FILLCELL_X32 FILLER_108_1176 ();
 FILLCELL_X32 FILLER_108_1208 ();
 FILLCELL_X32 FILLER_108_1240 ();
 FILLCELL_X32 FILLER_108_1272 ();
 FILLCELL_X32 FILLER_108_1304 ();
 FILLCELL_X32 FILLER_108_1336 ();
 FILLCELL_X32 FILLER_108_1368 ();
 FILLCELL_X32 FILLER_108_1400 ();
 FILLCELL_X32 FILLER_108_1432 ();
 FILLCELL_X32 FILLER_108_1464 ();
 FILLCELL_X32 FILLER_108_1496 ();
 FILLCELL_X32 FILLER_108_1528 ();
 FILLCELL_X32 FILLER_108_1560 ();
 FILLCELL_X32 FILLER_108_1592 ();
 FILLCELL_X32 FILLER_108_1624 ();
 FILLCELL_X32 FILLER_108_1656 ();
 FILLCELL_X32 FILLER_108_1688 ();
 FILLCELL_X32 FILLER_108_1720 ();
 FILLCELL_X32 FILLER_108_1752 ();
 FILLCELL_X32 FILLER_108_1784 ();
 FILLCELL_X32 FILLER_108_1816 ();
 FILLCELL_X32 FILLER_108_1848 ();
 FILLCELL_X8 FILLER_108_1880 ();
 FILLCELL_X4 FILLER_108_1888 ();
 FILLCELL_X2 FILLER_108_1892 ();
 FILLCELL_X32 FILLER_108_1895 ();
 FILLCELL_X32 FILLER_108_1927 ();
 FILLCELL_X32 FILLER_108_1959 ();
 FILLCELL_X32 FILLER_108_1991 ();
 FILLCELL_X32 FILLER_108_2023 ();
 FILLCELL_X32 FILLER_108_2055 ();
 FILLCELL_X32 FILLER_108_2087 ();
 FILLCELL_X32 FILLER_108_2119 ();
 FILLCELL_X32 FILLER_108_2151 ();
 FILLCELL_X32 FILLER_108_2183 ();
 FILLCELL_X32 FILLER_108_2215 ();
 FILLCELL_X32 FILLER_108_2247 ();
 FILLCELL_X32 FILLER_108_2279 ();
 FILLCELL_X32 FILLER_108_2311 ();
 FILLCELL_X32 FILLER_108_2343 ();
 FILLCELL_X32 FILLER_108_2375 ();
 FILLCELL_X32 FILLER_108_2407 ();
 FILLCELL_X32 FILLER_108_2439 ();
 FILLCELL_X32 FILLER_108_2471 ();
 FILLCELL_X32 FILLER_108_2503 ();
 FILLCELL_X32 FILLER_108_2535 ();
 FILLCELL_X32 FILLER_108_2567 ();
 FILLCELL_X32 FILLER_108_2599 ();
 FILLCELL_X32 FILLER_108_2631 ();
 FILLCELL_X32 FILLER_108_2663 ();
 FILLCELL_X32 FILLER_108_2695 ();
 FILLCELL_X32 FILLER_108_2727 ();
 FILLCELL_X32 FILLER_108_2759 ();
 FILLCELL_X32 FILLER_108_2791 ();
 FILLCELL_X32 FILLER_108_2823 ();
 FILLCELL_X32 FILLER_108_2855 ();
 FILLCELL_X32 FILLER_108_2887 ();
 FILLCELL_X32 FILLER_108_2919 ();
 FILLCELL_X32 FILLER_108_2951 ();
 FILLCELL_X32 FILLER_108_2983 ();
 FILLCELL_X32 FILLER_108_3015 ();
 FILLCELL_X32 FILLER_108_3047 ();
 FILLCELL_X32 FILLER_108_3079 ();
 FILLCELL_X32 FILLER_108_3111 ();
 FILLCELL_X8 FILLER_108_3143 ();
 FILLCELL_X4 FILLER_108_3151 ();
 FILLCELL_X2 FILLER_108_3155 ();
 FILLCELL_X32 FILLER_108_3158 ();
 FILLCELL_X32 FILLER_108_3190 ();
 FILLCELL_X32 FILLER_108_3222 ();
 FILLCELL_X32 FILLER_108_3254 ();
 FILLCELL_X32 FILLER_108_3286 ();
 FILLCELL_X32 FILLER_108_3318 ();
 FILLCELL_X32 FILLER_108_3350 ();
 FILLCELL_X32 FILLER_108_3382 ();
 FILLCELL_X32 FILLER_108_3414 ();
 FILLCELL_X32 FILLER_108_3446 ();
 FILLCELL_X32 FILLER_108_3478 ();
 FILLCELL_X32 FILLER_108_3510 ();
 FILLCELL_X32 FILLER_108_3542 ();
 FILLCELL_X32 FILLER_108_3574 ();
 FILLCELL_X32 FILLER_108_3606 ();
 FILLCELL_X32 FILLER_108_3638 ();
 FILLCELL_X32 FILLER_108_3670 ();
 FILLCELL_X32 FILLER_108_3702 ();
 FILLCELL_X4 FILLER_108_3734 ();
 FILLCELL_X32 FILLER_109_1 ();
 FILLCELL_X32 FILLER_109_33 ();
 FILLCELL_X32 FILLER_109_65 ();
 FILLCELL_X32 FILLER_109_97 ();
 FILLCELL_X32 FILLER_109_129 ();
 FILLCELL_X32 FILLER_109_161 ();
 FILLCELL_X32 FILLER_109_193 ();
 FILLCELL_X32 FILLER_109_225 ();
 FILLCELL_X32 FILLER_109_257 ();
 FILLCELL_X32 FILLER_109_289 ();
 FILLCELL_X32 FILLER_109_321 ();
 FILLCELL_X32 FILLER_109_353 ();
 FILLCELL_X32 FILLER_109_385 ();
 FILLCELL_X32 FILLER_109_417 ();
 FILLCELL_X32 FILLER_109_449 ();
 FILLCELL_X32 FILLER_109_481 ();
 FILLCELL_X32 FILLER_109_513 ();
 FILLCELL_X32 FILLER_109_545 ();
 FILLCELL_X32 FILLER_109_577 ();
 FILLCELL_X32 FILLER_109_609 ();
 FILLCELL_X32 FILLER_109_641 ();
 FILLCELL_X32 FILLER_109_673 ();
 FILLCELL_X32 FILLER_109_705 ();
 FILLCELL_X32 FILLER_109_737 ();
 FILLCELL_X32 FILLER_109_769 ();
 FILLCELL_X32 FILLER_109_801 ();
 FILLCELL_X32 FILLER_109_833 ();
 FILLCELL_X32 FILLER_109_865 ();
 FILLCELL_X32 FILLER_109_897 ();
 FILLCELL_X32 FILLER_109_929 ();
 FILLCELL_X32 FILLER_109_961 ();
 FILLCELL_X32 FILLER_109_993 ();
 FILLCELL_X32 FILLER_109_1025 ();
 FILLCELL_X32 FILLER_109_1057 ();
 FILLCELL_X32 FILLER_109_1089 ();
 FILLCELL_X32 FILLER_109_1121 ();
 FILLCELL_X32 FILLER_109_1153 ();
 FILLCELL_X32 FILLER_109_1185 ();
 FILLCELL_X32 FILLER_109_1217 ();
 FILLCELL_X8 FILLER_109_1249 ();
 FILLCELL_X4 FILLER_109_1257 ();
 FILLCELL_X2 FILLER_109_1261 ();
 FILLCELL_X32 FILLER_109_1264 ();
 FILLCELL_X32 FILLER_109_1296 ();
 FILLCELL_X32 FILLER_109_1328 ();
 FILLCELL_X32 FILLER_109_1360 ();
 FILLCELL_X32 FILLER_109_1392 ();
 FILLCELL_X32 FILLER_109_1424 ();
 FILLCELL_X32 FILLER_109_1456 ();
 FILLCELL_X32 FILLER_109_1488 ();
 FILLCELL_X32 FILLER_109_1520 ();
 FILLCELL_X32 FILLER_109_1552 ();
 FILLCELL_X32 FILLER_109_1584 ();
 FILLCELL_X32 FILLER_109_1616 ();
 FILLCELL_X32 FILLER_109_1648 ();
 FILLCELL_X32 FILLER_109_1680 ();
 FILLCELL_X32 FILLER_109_1712 ();
 FILLCELL_X32 FILLER_109_1744 ();
 FILLCELL_X32 FILLER_109_1776 ();
 FILLCELL_X32 FILLER_109_1808 ();
 FILLCELL_X32 FILLER_109_1840 ();
 FILLCELL_X32 FILLER_109_1872 ();
 FILLCELL_X32 FILLER_109_1904 ();
 FILLCELL_X32 FILLER_109_1936 ();
 FILLCELL_X32 FILLER_109_1968 ();
 FILLCELL_X32 FILLER_109_2000 ();
 FILLCELL_X32 FILLER_109_2032 ();
 FILLCELL_X32 FILLER_109_2064 ();
 FILLCELL_X32 FILLER_109_2096 ();
 FILLCELL_X32 FILLER_109_2128 ();
 FILLCELL_X32 FILLER_109_2160 ();
 FILLCELL_X32 FILLER_109_2192 ();
 FILLCELL_X32 FILLER_109_2224 ();
 FILLCELL_X32 FILLER_109_2256 ();
 FILLCELL_X32 FILLER_109_2288 ();
 FILLCELL_X32 FILLER_109_2320 ();
 FILLCELL_X32 FILLER_109_2352 ();
 FILLCELL_X32 FILLER_109_2384 ();
 FILLCELL_X32 FILLER_109_2416 ();
 FILLCELL_X32 FILLER_109_2448 ();
 FILLCELL_X32 FILLER_109_2480 ();
 FILLCELL_X8 FILLER_109_2512 ();
 FILLCELL_X4 FILLER_109_2520 ();
 FILLCELL_X2 FILLER_109_2524 ();
 FILLCELL_X32 FILLER_109_2527 ();
 FILLCELL_X32 FILLER_109_2559 ();
 FILLCELL_X32 FILLER_109_2591 ();
 FILLCELL_X32 FILLER_109_2623 ();
 FILLCELL_X32 FILLER_109_2655 ();
 FILLCELL_X32 FILLER_109_2687 ();
 FILLCELL_X32 FILLER_109_2719 ();
 FILLCELL_X32 FILLER_109_2751 ();
 FILLCELL_X32 FILLER_109_2783 ();
 FILLCELL_X32 FILLER_109_2815 ();
 FILLCELL_X32 FILLER_109_2847 ();
 FILLCELL_X32 FILLER_109_2879 ();
 FILLCELL_X32 FILLER_109_2911 ();
 FILLCELL_X32 FILLER_109_2943 ();
 FILLCELL_X32 FILLER_109_2975 ();
 FILLCELL_X32 FILLER_109_3007 ();
 FILLCELL_X32 FILLER_109_3039 ();
 FILLCELL_X32 FILLER_109_3071 ();
 FILLCELL_X32 FILLER_109_3103 ();
 FILLCELL_X32 FILLER_109_3135 ();
 FILLCELL_X32 FILLER_109_3167 ();
 FILLCELL_X32 FILLER_109_3199 ();
 FILLCELL_X32 FILLER_109_3231 ();
 FILLCELL_X32 FILLER_109_3263 ();
 FILLCELL_X32 FILLER_109_3295 ();
 FILLCELL_X32 FILLER_109_3327 ();
 FILLCELL_X32 FILLER_109_3359 ();
 FILLCELL_X32 FILLER_109_3391 ();
 FILLCELL_X32 FILLER_109_3423 ();
 FILLCELL_X32 FILLER_109_3455 ();
 FILLCELL_X32 FILLER_109_3487 ();
 FILLCELL_X32 FILLER_109_3519 ();
 FILLCELL_X32 FILLER_109_3551 ();
 FILLCELL_X32 FILLER_109_3583 ();
 FILLCELL_X32 FILLER_109_3615 ();
 FILLCELL_X32 FILLER_109_3647 ();
 FILLCELL_X32 FILLER_109_3679 ();
 FILLCELL_X16 FILLER_109_3711 ();
 FILLCELL_X8 FILLER_109_3727 ();
 FILLCELL_X2 FILLER_109_3735 ();
 FILLCELL_X1 FILLER_109_3737 ();
 FILLCELL_X32 FILLER_110_1 ();
 FILLCELL_X32 FILLER_110_33 ();
 FILLCELL_X32 FILLER_110_65 ();
 FILLCELL_X32 FILLER_110_97 ();
 FILLCELL_X32 FILLER_110_129 ();
 FILLCELL_X32 FILLER_110_161 ();
 FILLCELL_X32 FILLER_110_193 ();
 FILLCELL_X32 FILLER_110_225 ();
 FILLCELL_X32 FILLER_110_257 ();
 FILLCELL_X32 FILLER_110_289 ();
 FILLCELL_X32 FILLER_110_321 ();
 FILLCELL_X32 FILLER_110_353 ();
 FILLCELL_X32 FILLER_110_385 ();
 FILLCELL_X32 FILLER_110_417 ();
 FILLCELL_X32 FILLER_110_449 ();
 FILLCELL_X32 FILLER_110_481 ();
 FILLCELL_X32 FILLER_110_513 ();
 FILLCELL_X32 FILLER_110_545 ();
 FILLCELL_X32 FILLER_110_577 ();
 FILLCELL_X16 FILLER_110_609 ();
 FILLCELL_X4 FILLER_110_625 ();
 FILLCELL_X2 FILLER_110_629 ();
 FILLCELL_X32 FILLER_110_632 ();
 FILLCELL_X32 FILLER_110_664 ();
 FILLCELL_X32 FILLER_110_696 ();
 FILLCELL_X32 FILLER_110_728 ();
 FILLCELL_X32 FILLER_110_760 ();
 FILLCELL_X32 FILLER_110_792 ();
 FILLCELL_X32 FILLER_110_824 ();
 FILLCELL_X32 FILLER_110_856 ();
 FILLCELL_X32 FILLER_110_888 ();
 FILLCELL_X32 FILLER_110_920 ();
 FILLCELL_X32 FILLER_110_952 ();
 FILLCELL_X32 FILLER_110_984 ();
 FILLCELL_X32 FILLER_110_1016 ();
 FILLCELL_X32 FILLER_110_1048 ();
 FILLCELL_X32 FILLER_110_1080 ();
 FILLCELL_X32 FILLER_110_1112 ();
 FILLCELL_X32 FILLER_110_1144 ();
 FILLCELL_X32 FILLER_110_1176 ();
 FILLCELL_X32 FILLER_110_1208 ();
 FILLCELL_X32 FILLER_110_1240 ();
 FILLCELL_X32 FILLER_110_1272 ();
 FILLCELL_X32 FILLER_110_1304 ();
 FILLCELL_X32 FILLER_110_1336 ();
 FILLCELL_X32 FILLER_110_1368 ();
 FILLCELL_X32 FILLER_110_1400 ();
 FILLCELL_X32 FILLER_110_1432 ();
 FILLCELL_X32 FILLER_110_1464 ();
 FILLCELL_X32 FILLER_110_1496 ();
 FILLCELL_X32 FILLER_110_1528 ();
 FILLCELL_X32 FILLER_110_1560 ();
 FILLCELL_X32 FILLER_110_1592 ();
 FILLCELL_X32 FILLER_110_1624 ();
 FILLCELL_X32 FILLER_110_1656 ();
 FILLCELL_X32 FILLER_110_1688 ();
 FILLCELL_X32 FILLER_110_1720 ();
 FILLCELL_X32 FILLER_110_1752 ();
 FILLCELL_X32 FILLER_110_1784 ();
 FILLCELL_X32 FILLER_110_1816 ();
 FILLCELL_X32 FILLER_110_1848 ();
 FILLCELL_X8 FILLER_110_1880 ();
 FILLCELL_X4 FILLER_110_1888 ();
 FILLCELL_X2 FILLER_110_1892 ();
 FILLCELL_X32 FILLER_110_1895 ();
 FILLCELL_X32 FILLER_110_1927 ();
 FILLCELL_X32 FILLER_110_1959 ();
 FILLCELL_X32 FILLER_110_1991 ();
 FILLCELL_X32 FILLER_110_2023 ();
 FILLCELL_X32 FILLER_110_2055 ();
 FILLCELL_X32 FILLER_110_2087 ();
 FILLCELL_X32 FILLER_110_2119 ();
 FILLCELL_X32 FILLER_110_2151 ();
 FILLCELL_X32 FILLER_110_2183 ();
 FILLCELL_X32 FILLER_110_2215 ();
 FILLCELL_X32 FILLER_110_2247 ();
 FILLCELL_X32 FILLER_110_2279 ();
 FILLCELL_X32 FILLER_110_2311 ();
 FILLCELL_X32 FILLER_110_2343 ();
 FILLCELL_X32 FILLER_110_2375 ();
 FILLCELL_X32 FILLER_110_2407 ();
 FILLCELL_X32 FILLER_110_2439 ();
 FILLCELL_X32 FILLER_110_2471 ();
 FILLCELL_X32 FILLER_110_2503 ();
 FILLCELL_X32 FILLER_110_2535 ();
 FILLCELL_X32 FILLER_110_2567 ();
 FILLCELL_X32 FILLER_110_2599 ();
 FILLCELL_X32 FILLER_110_2631 ();
 FILLCELL_X32 FILLER_110_2663 ();
 FILLCELL_X32 FILLER_110_2695 ();
 FILLCELL_X32 FILLER_110_2727 ();
 FILLCELL_X32 FILLER_110_2759 ();
 FILLCELL_X32 FILLER_110_2791 ();
 FILLCELL_X32 FILLER_110_2823 ();
 FILLCELL_X32 FILLER_110_2855 ();
 FILLCELL_X32 FILLER_110_2887 ();
 FILLCELL_X32 FILLER_110_2919 ();
 FILLCELL_X32 FILLER_110_2951 ();
 FILLCELL_X32 FILLER_110_2983 ();
 FILLCELL_X32 FILLER_110_3015 ();
 FILLCELL_X32 FILLER_110_3047 ();
 FILLCELL_X32 FILLER_110_3079 ();
 FILLCELL_X32 FILLER_110_3111 ();
 FILLCELL_X8 FILLER_110_3143 ();
 FILLCELL_X4 FILLER_110_3151 ();
 FILLCELL_X2 FILLER_110_3155 ();
 FILLCELL_X32 FILLER_110_3158 ();
 FILLCELL_X32 FILLER_110_3190 ();
 FILLCELL_X32 FILLER_110_3222 ();
 FILLCELL_X32 FILLER_110_3254 ();
 FILLCELL_X32 FILLER_110_3286 ();
 FILLCELL_X32 FILLER_110_3318 ();
 FILLCELL_X32 FILLER_110_3350 ();
 FILLCELL_X32 FILLER_110_3382 ();
 FILLCELL_X32 FILLER_110_3414 ();
 FILLCELL_X32 FILLER_110_3446 ();
 FILLCELL_X32 FILLER_110_3478 ();
 FILLCELL_X32 FILLER_110_3510 ();
 FILLCELL_X32 FILLER_110_3542 ();
 FILLCELL_X32 FILLER_110_3574 ();
 FILLCELL_X32 FILLER_110_3606 ();
 FILLCELL_X32 FILLER_110_3638 ();
 FILLCELL_X32 FILLER_110_3670 ();
 FILLCELL_X32 FILLER_110_3702 ();
 FILLCELL_X4 FILLER_110_3734 ();
 FILLCELL_X32 FILLER_111_1 ();
 FILLCELL_X32 FILLER_111_33 ();
 FILLCELL_X32 FILLER_111_65 ();
 FILLCELL_X32 FILLER_111_97 ();
 FILLCELL_X32 FILLER_111_129 ();
 FILLCELL_X32 FILLER_111_161 ();
 FILLCELL_X32 FILLER_111_193 ();
 FILLCELL_X32 FILLER_111_225 ();
 FILLCELL_X32 FILLER_111_257 ();
 FILLCELL_X32 FILLER_111_289 ();
 FILLCELL_X32 FILLER_111_321 ();
 FILLCELL_X32 FILLER_111_353 ();
 FILLCELL_X32 FILLER_111_385 ();
 FILLCELL_X32 FILLER_111_417 ();
 FILLCELL_X32 FILLER_111_449 ();
 FILLCELL_X32 FILLER_111_481 ();
 FILLCELL_X32 FILLER_111_513 ();
 FILLCELL_X32 FILLER_111_545 ();
 FILLCELL_X32 FILLER_111_577 ();
 FILLCELL_X32 FILLER_111_609 ();
 FILLCELL_X32 FILLER_111_641 ();
 FILLCELL_X32 FILLER_111_673 ();
 FILLCELL_X32 FILLER_111_705 ();
 FILLCELL_X32 FILLER_111_737 ();
 FILLCELL_X32 FILLER_111_769 ();
 FILLCELL_X32 FILLER_111_801 ();
 FILLCELL_X32 FILLER_111_833 ();
 FILLCELL_X32 FILLER_111_865 ();
 FILLCELL_X32 FILLER_111_897 ();
 FILLCELL_X32 FILLER_111_929 ();
 FILLCELL_X32 FILLER_111_961 ();
 FILLCELL_X32 FILLER_111_993 ();
 FILLCELL_X32 FILLER_111_1025 ();
 FILLCELL_X32 FILLER_111_1057 ();
 FILLCELL_X32 FILLER_111_1089 ();
 FILLCELL_X32 FILLER_111_1121 ();
 FILLCELL_X32 FILLER_111_1153 ();
 FILLCELL_X32 FILLER_111_1185 ();
 FILLCELL_X32 FILLER_111_1217 ();
 FILLCELL_X8 FILLER_111_1249 ();
 FILLCELL_X4 FILLER_111_1257 ();
 FILLCELL_X2 FILLER_111_1261 ();
 FILLCELL_X32 FILLER_111_1264 ();
 FILLCELL_X32 FILLER_111_1296 ();
 FILLCELL_X32 FILLER_111_1328 ();
 FILLCELL_X32 FILLER_111_1360 ();
 FILLCELL_X32 FILLER_111_1392 ();
 FILLCELL_X32 FILLER_111_1424 ();
 FILLCELL_X32 FILLER_111_1456 ();
 FILLCELL_X32 FILLER_111_1488 ();
 FILLCELL_X32 FILLER_111_1520 ();
 FILLCELL_X32 FILLER_111_1552 ();
 FILLCELL_X32 FILLER_111_1584 ();
 FILLCELL_X32 FILLER_111_1616 ();
 FILLCELL_X32 FILLER_111_1648 ();
 FILLCELL_X32 FILLER_111_1680 ();
 FILLCELL_X32 FILLER_111_1712 ();
 FILLCELL_X32 FILLER_111_1744 ();
 FILLCELL_X32 FILLER_111_1776 ();
 FILLCELL_X32 FILLER_111_1808 ();
 FILLCELL_X32 FILLER_111_1840 ();
 FILLCELL_X32 FILLER_111_1872 ();
 FILLCELL_X32 FILLER_111_1904 ();
 FILLCELL_X32 FILLER_111_1936 ();
 FILLCELL_X32 FILLER_111_1968 ();
 FILLCELL_X32 FILLER_111_2000 ();
 FILLCELL_X32 FILLER_111_2032 ();
 FILLCELL_X32 FILLER_111_2064 ();
 FILLCELL_X32 FILLER_111_2096 ();
 FILLCELL_X32 FILLER_111_2128 ();
 FILLCELL_X32 FILLER_111_2160 ();
 FILLCELL_X32 FILLER_111_2192 ();
 FILLCELL_X32 FILLER_111_2224 ();
 FILLCELL_X32 FILLER_111_2256 ();
 FILLCELL_X32 FILLER_111_2288 ();
 FILLCELL_X32 FILLER_111_2320 ();
 FILLCELL_X32 FILLER_111_2352 ();
 FILLCELL_X32 FILLER_111_2384 ();
 FILLCELL_X32 FILLER_111_2416 ();
 FILLCELL_X32 FILLER_111_2448 ();
 FILLCELL_X32 FILLER_111_2480 ();
 FILLCELL_X8 FILLER_111_2512 ();
 FILLCELL_X4 FILLER_111_2520 ();
 FILLCELL_X2 FILLER_111_2524 ();
 FILLCELL_X32 FILLER_111_2527 ();
 FILLCELL_X32 FILLER_111_2559 ();
 FILLCELL_X32 FILLER_111_2591 ();
 FILLCELL_X32 FILLER_111_2623 ();
 FILLCELL_X32 FILLER_111_2655 ();
 FILLCELL_X32 FILLER_111_2687 ();
 FILLCELL_X32 FILLER_111_2719 ();
 FILLCELL_X32 FILLER_111_2751 ();
 FILLCELL_X32 FILLER_111_2783 ();
 FILLCELL_X32 FILLER_111_2815 ();
 FILLCELL_X32 FILLER_111_2847 ();
 FILLCELL_X32 FILLER_111_2879 ();
 FILLCELL_X32 FILLER_111_2911 ();
 FILLCELL_X32 FILLER_111_2943 ();
 FILLCELL_X32 FILLER_111_2975 ();
 FILLCELL_X32 FILLER_111_3007 ();
 FILLCELL_X32 FILLER_111_3039 ();
 FILLCELL_X32 FILLER_111_3071 ();
 FILLCELL_X32 FILLER_111_3103 ();
 FILLCELL_X32 FILLER_111_3135 ();
 FILLCELL_X32 FILLER_111_3167 ();
 FILLCELL_X32 FILLER_111_3199 ();
 FILLCELL_X32 FILLER_111_3231 ();
 FILLCELL_X32 FILLER_111_3263 ();
 FILLCELL_X32 FILLER_111_3295 ();
 FILLCELL_X32 FILLER_111_3327 ();
 FILLCELL_X32 FILLER_111_3359 ();
 FILLCELL_X32 FILLER_111_3391 ();
 FILLCELL_X32 FILLER_111_3423 ();
 FILLCELL_X32 FILLER_111_3455 ();
 FILLCELL_X32 FILLER_111_3487 ();
 FILLCELL_X32 FILLER_111_3519 ();
 FILLCELL_X32 FILLER_111_3551 ();
 FILLCELL_X32 FILLER_111_3583 ();
 FILLCELL_X32 FILLER_111_3615 ();
 FILLCELL_X32 FILLER_111_3647 ();
 FILLCELL_X32 FILLER_111_3679 ();
 FILLCELL_X16 FILLER_111_3711 ();
 FILLCELL_X8 FILLER_111_3727 ();
 FILLCELL_X2 FILLER_111_3735 ();
 FILLCELL_X1 FILLER_111_3737 ();
 FILLCELL_X32 FILLER_112_1 ();
 FILLCELL_X32 FILLER_112_33 ();
 FILLCELL_X32 FILLER_112_65 ();
 FILLCELL_X32 FILLER_112_97 ();
 FILLCELL_X32 FILLER_112_129 ();
 FILLCELL_X32 FILLER_112_161 ();
 FILLCELL_X32 FILLER_112_193 ();
 FILLCELL_X32 FILLER_112_225 ();
 FILLCELL_X32 FILLER_112_257 ();
 FILLCELL_X32 FILLER_112_289 ();
 FILLCELL_X32 FILLER_112_321 ();
 FILLCELL_X32 FILLER_112_353 ();
 FILLCELL_X32 FILLER_112_385 ();
 FILLCELL_X32 FILLER_112_417 ();
 FILLCELL_X32 FILLER_112_449 ();
 FILLCELL_X32 FILLER_112_481 ();
 FILLCELL_X32 FILLER_112_513 ();
 FILLCELL_X32 FILLER_112_545 ();
 FILLCELL_X32 FILLER_112_577 ();
 FILLCELL_X16 FILLER_112_609 ();
 FILLCELL_X4 FILLER_112_625 ();
 FILLCELL_X2 FILLER_112_629 ();
 FILLCELL_X32 FILLER_112_632 ();
 FILLCELL_X32 FILLER_112_664 ();
 FILLCELL_X32 FILLER_112_696 ();
 FILLCELL_X32 FILLER_112_728 ();
 FILLCELL_X32 FILLER_112_760 ();
 FILLCELL_X32 FILLER_112_792 ();
 FILLCELL_X32 FILLER_112_824 ();
 FILLCELL_X32 FILLER_112_856 ();
 FILLCELL_X32 FILLER_112_888 ();
 FILLCELL_X32 FILLER_112_920 ();
 FILLCELL_X32 FILLER_112_952 ();
 FILLCELL_X32 FILLER_112_984 ();
 FILLCELL_X32 FILLER_112_1016 ();
 FILLCELL_X32 FILLER_112_1048 ();
 FILLCELL_X32 FILLER_112_1080 ();
 FILLCELL_X32 FILLER_112_1112 ();
 FILLCELL_X32 FILLER_112_1144 ();
 FILLCELL_X32 FILLER_112_1176 ();
 FILLCELL_X32 FILLER_112_1208 ();
 FILLCELL_X32 FILLER_112_1240 ();
 FILLCELL_X32 FILLER_112_1272 ();
 FILLCELL_X32 FILLER_112_1304 ();
 FILLCELL_X32 FILLER_112_1336 ();
 FILLCELL_X32 FILLER_112_1368 ();
 FILLCELL_X32 FILLER_112_1400 ();
 FILLCELL_X32 FILLER_112_1432 ();
 FILLCELL_X32 FILLER_112_1464 ();
 FILLCELL_X32 FILLER_112_1496 ();
 FILLCELL_X32 FILLER_112_1528 ();
 FILLCELL_X32 FILLER_112_1560 ();
 FILLCELL_X32 FILLER_112_1592 ();
 FILLCELL_X32 FILLER_112_1624 ();
 FILLCELL_X32 FILLER_112_1656 ();
 FILLCELL_X32 FILLER_112_1688 ();
 FILLCELL_X32 FILLER_112_1720 ();
 FILLCELL_X32 FILLER_112_1752 ();
 FILLCELL_X32 FILLER_112_1784 ();
 FILLCELL_X32 FILLER_112_1816 ();
 FILLCELL_X32 FILLER_112_1848 ();
 FILLCELL_X8 FILLER_112_1880 ();
 FILLCELL_X4 FILLER_112_1888 ();
 FILLCELL_X2 FILLER_112_1892 ();
 FILLCELL_X32 FILLER_112_1895 ();
 FILLCELL_X32 FILLER_112_1927 ();
 FILLCELL_X32 FILLER_112_1959 ();
 FILLCELL_X32 FILLER_112_1991 ();
 FILLCELL_X32 FILLER_112_2023 ();
 FILLCELL_X32 FILLER_112_2055 ();
 FILLCELL_X32 FILLER_112_2087 ();
 FILLCELL_X32 FILLER_112_2119 ();
 FILLCELL_X32 FILLER_112_2151 ();
 FILLCELL_X32 FILLER_112_2183 ();
 FILLCELL_X32 FILLER_112_2215 ();
 FILLCELL_X32 FILLER_112_2247 ();
 FILLCELL_X32 FILLER_112_2279 ();
 FILLCELL_X32 FILLER_112_2311 ();
 FILLCELL_X32 FILLER_112_2343 ();
 FILLCELL_X32 FILLER_112_2375 ();
 FILLCELL_X32 FILLER_112_2407 ();
 FILLCELL_X32 FILLER_112_2439 ();
 FILLCELL_X32 FILLER_112_2471 ();
 FILLCELL_X32 FILLER_112_2503 ();
 FILLCELL_X32 FILLER_112_2535 ();
 FILLCELL_X32 FILLER_112_2567 ();
 FILLCELL_X32 FILLER_112_2599 ();
 FILLCELL_X32 FILLER_112_2631 ();
 FILLCELL_X32 FILLER_112_2663 ();
 FILLCELL_X32 FILLER_112_2695 ();
 FILLCELL_X32 FILLER_112_2727 ();
 FILLCELL_X32 FILLER_112_2759 ();
 FILLCELL_X32 FILLER_112_2791 ();
 FILLCELL_X32 FILLER_112_2823 ();
 FILLCELL_X32 FILLER_112_2855 ();
 FILLCELL_X32 FILLER_112_2887 ();
 FILLCELL_X32 FILLER_112_2919 ();
 FILLCELL_X32 FILLER_112_2951 ();
 FILLCELL_X32 FILLER_112_2983 ();
 FILLCELL_X32 FILLER_112_3015 ();
 FILLCELL_X32 FILLER_112_3047 ();
 FILLCELL_X32 FILLER_112_3079 ();
 FILLCELL_X32 FILLER_112_3111 ();
 FILLCELL_X8 FILLER_112_3143 ();
 FILLCELL_X4 FILLER_112_3151 ();
 FILLCELL_X2 FILLER_112_3155 ();
 FILLCELL_X32 FILLER_112_3158 ();
 FILLCELL_X32 FILLER_112_3190 ();
 FILLCELL_X32 FILLER_112_3222 ();
 FILLCELL_X32 FILLER_112_3254 ();
 FILLCELL_X32 FILLER_112_3286 ();
 FILLCELL_X32 FILLER_112_3318 ();
 FILLCELL_X32 FILLER_112_3350 ();
 FILLCELL_X32 FILLER_112_3382 ();
 FILLCELL_X32 FILLER_112_3414 ();
 FILLCELL_X32 FILLER_112_3446 ();
 FILLCELL_X32 FILLER_112_3478 ();
 FILLCELL_X32 FILLER_112_3510 ();
 FILLCELL_X32 FILLER_112_3542 ();
 FILLCELL_X32 FILLER_112_3574 ();
 FILLCELL_X32 FILLER_112_3606 ();
 FILLCELL_X32 FILLER_112_3638 ();
 FILLCELL_X32 FILLER_112_3670 ();
 FILLCELL_X32 FILLER_112_3702 ();
 FILLCELL_X4 FILLER_112_3734 ();
 FILLCELL_X32 FILLER_113_1 ();
 FILLCELL_X32 FILLER_113_33 ();
 FILLCELL_X32 FILLER_113_65 ();
 FILLCELL_X32 FILLER_113_97 ();
 FILLCELL_X32 FILLER_113_129 ();
 FILLCELL_X32 FILLER_113_161 ();
 FILLCELL_X32 FILLER_113_193 ();
 FILLCELL_X32 FILLER_113_225 ();
 FILLCELL_X32 FILLER_113_257 ();
 FILLCELL_X32 FILLER_113_289 ();
 FILLCELL_X32 FILLER_113_321 ();
 FILLCELL_X32 FILLER_113_353 ();
 FILLCELL_X32 FILLER_113_385 ();
 FILLCELL_X32 FILLER_113_417 ();
 FILLCELL_X32 FILLER_113_449 ();
 FILLCELL_X32 FILLER_113_481 ();
 FILLCELL_X32 FILLER_113_513 ();
 FILLCELL_X32 FILLER_113_545 ();
 FILLCELL_X32 FILLER_113_577 ();
 FILLCELL_X32 FILLER_113_609 ();
 FILLCELL_X32 FILLER_113_641 ();
 FILLCELL_X32 FILLER_113_673 ();
 FILLCELL_X32 FILLER_113_705 ();
 FILLCELL_X32 FILLER_113_737 ();
 FILLCELL_X32 FILLER_113_769 ();
 FILLCELL_X32 FILLER_113_801 ();
 FILLCELL_X32 FILLER_113_833 ();
 FILLCELL_X32 FILLER_113_865 ();
 FILLCELL_X32 FILLER_113_897 ();
 FILLCELL_X32 FILLER_113_929 ();
 FILLCELL_X32 FILLER_113_961 ();
 FILLCELL_X32 FILLER_113_993 ();
 FILLCELL_X32 FILLER_113_1025 ();
 FILLCELL_X32 FILLER_113_1057 ();
 FILLCELL_X32 FILLER_113_1089 ();
 FILLCELL_X32 FILLER_113_1121 ();
 FILLCELL_X32 FILLER_113_1153 ();
 FILLCELL_X32 FILLER_113_1185 ();
 FILLCELL_X32 FILLER_113_1217 ();
 FILLCELL_X8 FILLER_113_1249 ();
 FILLCELL_X4 FILLER_113_1257 ();
 FILLCELL_X2 FILLER_113_1261 ();
 FILLCELL_X32 FILLER_113_1264 ();
 FILLCELL_X32 FILLER_113_1296 ();
 FILLCELL_X32 FILLER_113_1328 ();
 FILLCELL_X32 FILLER_113_1360 ();
 FILLCELL_X32 FILLER_113_1392 ();
 FILLCELL_X32 FILLER_113_1424 ();
 FILLCELL_X32 FILLER_113_1456 ();
 FILLCELL_X32 FILLER_113_1488 ();
 FILLCELL_X32 FILLER_113_1520 ();
 FILLCELL_X32 FILLER_113_1552 ();
 FILLCELL_X32 FILLER_113_1584 ();
 FILLCELL_X32 FILLER_113_1616 ();
 FILLCELL_X32 FILLER_113_1648 ();
 FILLCELL_X32 FILLER_113_1680 ();
 FILLCELL_X32 FILLER_113_1712 ();
 FILLCELL_X32 FILLER_113_1744 ();
 FILLCELL_X32 FILLER_113_1776 ();
 FILLCELL_X32 FILLER_113_1808 ();
 FILLCELL_X32 FILLER_113_1840 ();
 FILLCELL_X32 FILLER_113_1872 ();
 FILLCELL_X32 FILLER_113_1904 ();
 FILLCELL_X32 FILLER_113_1936 ();
 FILLCELL_X32 FILLER_113_1968 ();
 FILLCELL_X32 FILLER_113_2000 ();
 FILLCELL_X32 FILLER_113_2032 ();
 FILLCELL_X32 FILLER_113_2064 ();
 FILLCELL_X32 FILLER_113_2096 ();
 FILLCELL_X32 FILLER_113_2128 ();
 FILLCELL_X32 FILLER_113_2160 ();
 FILLCELL_X32 FILLER_113_2192 ();
 FILLCELL_X32 FILLER_113_2224 ();
 FILLCELL_X32 FILLER_113_2256 ();
 FILLCELL_X32 FILLER_113_2288 ();
 FILLCELL_X32 FILLER_113_2320 ();
 FILLCELL_X32 FILLER_113_2352 ();
 FILLCELL_X32 FILLER_113_2384 ();
 FILLCELL_X32 FILLER_113_2416 ();
 FILLCELL_X32 FILLER_113_2448 ();
 FILLCELL_X32 FILLER_113_2480 ();
 FILLCELL_X8 FILLER_113_2512 ();
 FILLCELL_X4 FILLER_113_2520 ();
 FILLCELL_X2 FILLER_113_2524 ();
 FILLCELL_X32 FILLER_113_2527 ();
 FILLCELL_X32 FILLER_113_2559 ();
 FILLCELL_X32 FILLER_113_2591 ();
 FILLCELL_X32 FILLER_113_2623 ();
 FILLCELL_X32 FILLER_113_2655 ();
 FILLCELL_X32 FILLER_113_2687 ();
 FILLCELL_X32 FILLER_113_2719 ();
 FILLCELL_X32 FILLER_113_2751 ();
 FILLCELL_X32 FILLER_113_2783 ();
 FILLCELL_X32 FILLER_113_2815 ();
 FILLCELL_X32 FILLER_113_2847 ();
 FILLCELL_X32 FILLER_113_2879 ();
 FILLCELL_X32 FILLER_113_2911 ();
 FILLCELL_X32 FILLER_113_2943 ();
 FILLCELL_X32 FILLER_113_2975 ();
 FILLCELL_X32 FILLER_113_3007 ();
 FILLCELL_X32 FILLER_113_3039 ();
 FILLCELL_X32 FILLER_113_3071 ();
 FILLCELL_X32 FILLER_113_3103 ();
 FILLCELL_X32 FILLER_113_3135 ();
 FILLCELL_X32 FILLER_113_3167 ();
 FILLCELL_X32 FILLER_113_3199 ();
 FILLCELL_X32 FILLER_113_3231 ();
 FILLCELL_X32 FILLER_113_3263 ();
 FILLCELL_X32 FILLER_113_3295 ();
 FILLCELL_X32 FILLER_113_3327 ();
 FILLCELL_X32 FILLER_113_3359 ();
 FILLCELL_X32 FILLER_113_3391 ();
 FILLCELL_X32 FILLER_113_3423 ();
 FILLCELL_X32 FILLER_113_3455 ();
 FILLCELL_X32 FILLER_113_3487 ();
 FILLCELL_X32 FILLER_113_3519 ();
 FILLCELL_X32 FILLER_113_3551 ();
 FILLCELL_X32 FILLER_113_3583 ();
 FILLCELL_X32 FILLER_113_3615 ();
 FILLCELL_X32 FILLER_113_3647 ();
 FILLCELL_X32 FILLER_113_3679 ();
 FILLCELL_X16 FILLER_113_3711 ();
 FILLCELL_X8 FILLER_113_3727 ();
 FILLCELL_X2 FILLER_113_3735 ();
 FILLCELL_X1 FILLER_113_3737 ();
 FILLCELL_X32 FILLER_114_1 ();
 FILLCELL_X32 FILLER_114_33 ();
 FILLCELL_X32 FILLER_114_65 ();
 FILLCELL_X32 FILLER_114_97 ();
 FILLCELL_X32 FILLER_114_129 ();
 FILLCELL_X32 FILLER_114_161 ();
 FILLCELL_X32 FILLER_114_193 ();
 FILLCELL_X32 FILLER_114_225 ();
 FILLCELL_X32 FILLER_114_257 ();
 FILLCELL_X32 FILLER_114_289 ();
 FILLCELL_X32 FILLER_114_321 ();
 FILLCELL_X32 FILLER_114_353 ();
 FILLCELL_X32 FILLER_114_385 ();
 FILLCELL_X32 FILLER_114_417 ();
 FILLCELL_X32 FILLER_114_449 ();
 FILLCELL_X32 FILLER_114_481 ();
 FILLCELL_X32 FILLER_114_513 ();
 FILLCELL_X32 FILLER_114_545 ();
 FILLCELL_X32 FILLER_114_577 ();
 FILLCELL_X16 FILLER_114_609 ();
 FILLCELL_X4 FILLER_114_625 ();
 FILLCELL_X2 FILLER_114_629 ();
 FILLCELL_X32 FILLER_114_632 ();
 FILLCELL_X32 FILLER_114_664 ();
 FILLCELL_X32 FILLER_114_696 ();
 FILLCELL_X32 FILLER_114_728 ();
 FILLCELL_X32 FILLER_114_760 ();
 FILLCELL_X32 FILLER_114_792 ();
 FILLCELL_X32 FILLER_114_824 ();
 FILLCELL_X32 FILLER_114_856 ();
 FILLCELL_X32 FILLER_114_888 ();
 FILLCELL_X32 FILLER_114_920 ();
 FILLCELL_X32 FILLER_114_952 ();
 FILLCELL_X32 FILLER_114_984 ();
 FILLCELL_X32 FILLER_114_1016 ();
 FILLCELL_X32 FILLER_114_1048 ();
 FILLCELL_X32 FILLER_114_1080 ();
 FILLCELL_X32 FILLER_114_1112 ();
 FILLCELL_X32 FILLER_114_1144 ();
 FILLCELL_X32 FILLER_114_1176 ();
 FILLCELL_X32 FILLER_114_1208 ();
 FILLCELL_X32 FILLER_114_1240 ();
 FILLCELL_X32 FILLER_114_1272 ();
 FILLCELL_X32 FILLER_114_1304 ();
 FILLCELL_X32 FILLER_114_1336 ();
 FILLCELL_X32 FILLER_114_1368 ();
 FILLCELL_X32 FILLER_114_1400 ();
 FILLCELL_X32 FILLER_114_1432 ();
 FILLCELL_X32 FILLER_114_1464 ();
 FILLCELL_X32 FILLER_114_1496 ();
 FILLCELL_X32 FILLER_114_1528 ();
 FILLCELL_X32 FILLER_114_1560 ();
 FILLCELL_X32 FILLER_114_1592 ();
 FILLCELL_X32 FILLER_114_1624 ();
 FILLCELL_X32 FILLER_114_1656 ();
 FILLCELL_X32 FILLER_114_1688 ();
 FILLCELL_X32 FILLER_114_1720 ();
 FILLCELL_X32 FILLER_114_1752 ();
 FILLCELL_X32 FILLER_114_1784 ();
 FILLCELL_X32 FILLER_114_1816 ();
 FILLCELL_X32 FILLER_114_1848 ();
 FILLCELL_X8 FILLER_114_1880 ();
 FILLCELL_X4 FILLER_114_1888 ();
 FILLCELL_X2 FILLER_114_1892 ();
 FILLCELL_X32 FILLER_114_1895 ();
 FILLCELL_X32 FILLER_114_1927 ();
 FILLCELL_X32 FILLER_114_1959 ();
 FILLCELL_X32 FILLER_114_1991 ();
 FILLCELL_X32 FILLER_114_2023 ();
 FILLCELL_X32 FILLER_114_2055 ();
 FILLCELL_X32 FILLER_114_2087 ();
 FILLCELL_X32 FILLER_114_2119 ();
 FILLCELL_X32 FILLER_114_2151 ();
 FILLCELL_X32 FILLER_114_2183 ();
 FILLCELL_X32 FILLER_114_2215 ();
 FILLCELL_X32 FILLER_114_2247 ();
 FILLCELL_X32 FILLER_114_2279 ();
 FILLCELL_X32 FILLER_114_2311 ();
 FILLCELL_X32 FILLER_114_2343 ();
 FILLCELL_X32 FILLER_114_2375 ();
 FILLCELL_X32 FILLER_114_2407 ();
 FILLCELL_X32 FILLER_114_2439 ();
 FILLCELL_X32 FILLER_114_2471 ();
 FILLCELL_X32 FILLER_114_2503 ();
 FILLCELL_X32 FILLER_114_2535 ();
 FILLCELL_X32 FILLER_114_2567 ();
 FILLCELL_X32 FILLER_114_2599 ();
 FILLCELL_X32 FILLER_114_2631 ();
 FILLCELL_X32 FILLER_114_2663 ();
 FILLCELL_X32 FILLER_114_2695 ();
 FILLCELL_X32 FILLER_114_2727 ();
 FILLCELL_X32 FILLER_114_2759 ();
 FILLCELL_X32 FILLER_114_2791 ();
 FILLCELL_X32 FILLER_114_2823 ();
 FILLCELL_X32 FILLER_114_2855 ();
 FILLCELL_X32 FILLER_114_2887 ();
 FILLCELL_X32 FILLER_114_2919 ();
 FILLCELL_X32 FILLER_114_2951 ();
 FILLCELL_X32 FILLER_114_2983 ();
 FILLCELL_X32 FILLER_114_3015 ();
 FILLCELL_X32 FILLER_114_3047 ();
 FILLCELL_X32 FILLER_114_3079 ();
 FILLCELL_X32 FILLER_114_3111 ();
 FILLCELL_X8 FILLER_114_3143 ();
 FILLCELL_X4 FILLER_114_3151 ();
 FILLCELL_X2 FILLER_114_3155 ();
 FILLCELL_X32 FILLER_114_3158 ();
 FILLCELL_X32 FILLER_114_3190 ();
 FILLCELL_X32 FILLER_114_3222 ();
 FILLCELL_X32 FILLER_114_3254 ();
 FILLCELL_X32 FILLER_114_3286 ();
 FILLCELL_X32 FILLER_114_3318 ();
 FILLCELL_X32 FILLER_114_3350 ();
 FILLCELL_X32 FILLER_114_3382 ();
 FILLCELL_X32 FILLER_114_3414 ();
 FILLCELL_X32 FILLER_114_3446 ();
 FILLCELL_X32 FILLER_114_3478 ();
 FILLCELL_X32 FILLER_114_3510 ();
 FILLCELL_X32 FILLER_114_3542 ();
 FILLCELL_X32 FILLER_114_3574 ();
 FILLCELL_X32 FILLER_114_3606 ();
 FILLCELL_X32 FILLER_114_3638 ();
 FILLCELL_X32 FILLER_114_3670 ();
 FILLCELL_X32 FILLER_114_3702 ();
 FILLCELL_X4 FILLER_114_3734 ();
 FILLCELL_X32 FILLER_115_1 ();
 FILLCELL_X32 FILLER_115_33 ();
 FILLCELL_X32 FILLER_115_65 ();
 FILLCELL_X32 FILLER_115_97 ();
 FILLCELL_X32 FILLER_115_129 ();
 FILLCELL_X32 FILLER_115_161 ();
 FILLCELL_X32 FILLER_115_193 ();
 FILLCELL_X32 FILLER_115_225 ();
 FILLCELL_X32 FILLER_115_257 ();
 FILLCELL_X32 FILLER_115_289 ();
 FILLCELL_X32 FILLER_115_321 ();
 FILLCELL_X32 FILLER_115_353 ();
 FILLCELL_X32 FILLER_115_385 ();
 FILLCELL_X32 FILLER_115_417 ();
 FILLCELL_X32 FILLER_115_449 ();
 FILLCELL_X32 FILLER_115_481 ();
 FILLCELL_X32 FILLER_115_513 ();
 FILLCELL_X32 FILLER_115_545 ();
 FILLCELL_X32 FILLER_115_577 ();
 FILLCELL_X32 FILLER_115_609 ();
 FILLCELL_X32 FILLER_115_641 ();
 FILLCELL_X32 FILLER_115_673 ();
 FILLCELL_X32 FILLER_115_705 ();
 FILLCELL_X32 FILLER_115_737 ();
 FILLCELL_X32 FILLER_115_769 ();
 FILLCELL_X32 FILLER_115_801 ();
 FILLCELL_X32 FILLER_115_833 ();
 FILLCELL_X32 FILLER_115_865 ();
 FILLCELL_X32 FILLER_115_897 ();
 FILLCELL_X32 FILLER_115_929 ();
 FILLCELL_X32 FILLER_115_961 ();
 FILLCELL_X32 FILLER_115_993 ();
 FILLCELL_X32 FILLER_115_1025 ();
 FILLCELL_X32 FILLER_115_1057 ();
 FILLCELL_X32 FILLER_115_1089 ();
 FILLCELL_X32 FILLER_115_1121 ();
 FILLCELL_X32 FILLER_115_1153 ();
 FILLCELL_X32 FILLER_115_1185 ();
 FILLCELL_X32 FILLER_115_1217 ();
 FILLCELL_X8 FILLER_115_1249 ();
 FILLCELL_X4 FILLER_115_1257 ();
 FILLCELL_X2 FILLER_115_1261 ();
 FILLCELL_X32 FILLER_115_1264 ();
 FILLCELL_X32 FILLER_115_1296 ();
 FILLCELL_X32 FILLER_115_1328 ();
 FILLCELL_X32 FILLER_115_1360 ();
 FILLCELL_X32 FILLER_115_1392 ();
 FILLCELL_X32 FILLER_115_1424 ();
 FILLCELL_X32 FILLER_115_1456 ();
 FILLCELL_X32 FILLER_115_1488 ();
 FILLCELL_X32 FILLER_115_1520 ();
 FILLCELL_X32 FILLER_115_1552 ();
 FILLCELL_X32 FILLER_115_1584 ();
 FILLCELL_X32 FILLER_115_1616 ();
 FILLCELL_X32 FILLER_115_1648 ();
 FILLCELL_X32 FILLER_115_1680 ();
 FILLCELL_X32 FILLER_115_1712 ();
 FILLCELL_X32 FILLER_115_1744 ();
 FILLCELL_X32 FILLER_115_1776 ();
 FILLCELL_X32 FILLER_115_1808 ();
 FILLCELL_X32 FILLER_115_1840 ();
 FILLCELL_X32 FILLER_115_1872 ();
 FILLCELL_X32 FILLER_115_1904 ();
 FILLCELL_X32 FILLER_115_1936 ();
 FILLCELL_X32 FILLER_115_1968 ();
 FILLCELL_X32 FILLER_115_2000 ();
 FILLCELL_X32 FILLER_115_2032 ();
 FILLCELL_X32 FILLER_115_2064 ();
 FILLCELL_X32 FILLER_115_2096 ();
 FILLCELL_X32 FILLER_115_2128 ();
 FILLCELL_X32 FILLER_115_2160 ();
 FILLCELL_X32 FILLER_115_2192 ();
 FILLCELL_X32 FILLER_115_2224 ();
 FILLCELL_X32 FILLER_115_2256 ();
 FILLCELL_X32 FILLER_115_2288 ();
 FILLCELL_X32 FILLER_115_2320 ();
 FILLCELL_X32 FILLER_115_2352 ();
 FILLCELL_X32 FILLER_115_2384 ();
 FILLCELL_X32 FILLER_115_2416 ();
 FILLCELL_X32 FILLER_115_2448 ();
 FILLCELL_X32 FILLER_115_2480 ();
 FILLCELL_X8 FILLER_115_2512 ();
 FILLCELL_X4 FILLER_115_2520 ();
 FILLCELL_X2 FILLER_115_2524 ();
 FILLCELL_X32 FILLER_115_2527 ();
 FILLCELL_X32 FILLER_115_2559 ();
 FILLCELL_X32 FILLER_115_2591 ();
 FILLCELL_X32 FILLER_115_2623 ();
 FILLCELL_X32 FILLER_115_2655 ();
 FILLCELL_X32 FILLER_115_2687 ();
 FILLCELL_X32 FILLER_115_2719 ();
 FILLCELL_X32 FILLER_115_2751 ();
 FILLCELL_X32 FILLER_115_2783 ();
 FILLCELL_X32 FILLER_115_2815 ();
 FILLCELL_X32 FILLER_115_2847 ();
 FILLCELL_X32 FILLER_115_2879 ();
 FILLCELL_X32 FILLER_115_2911 ();
 FILLCELL_X32 FILLER_115_2943 ();
 FILLCELL_X32 FILLER_115_2975 ();
 FILLCELL_X32 FILLER_115_3007 ();
 FILLCELL_X32 FILLER_115_3039 ();
 FILLCELL_X32 FILLER_115_3071 ();
 FILLCELL_X32 FILLER_115_3103 ();
 FILLCELL_X32 FILLER_115_3135 ();
 FILLCELL_X32 FILLER_115_3167 ();
 FILLCELL_X32 FILLER_115_3199 ();
 FILLCELL_X32 FILLER_115_3231 ();
 FILLCELL_X32 FILLER_115_3263 ();
 FILLCELL_X32 FILLER_115_3295 ();
 FILLCELL_X32 FILLER_115_3327 ();
 FILLCELL_X32 FILLER_115_3359 ();
 FILLCELL_X32 FILLER_115_3391 ();
 FILLCELL_X32 FILLER_115_3423 ();
 FILLCELL_X32 FILLER_115_3455 ();
 FILLCELL_X32 FILLER_115_3487 ();
 FILLCELL_X32 FILLER_115_3519 ();
 FILLCELL_X32 FILLER_115_3551 ();
 FILLCELL_X32 FILLER_115_3583 ();
 FILLCELL_X32 FILLER_115_3615 ();
 FILLCELL_X32 FILLER_115_3647 ();
 FILLCELL_X32 FILLER_115_3679 ();
 FILLCELL_X16 FILLER_115_3711 ();
 FILLCELL_X8 FILLER_115_3727 ();
 FILLCELL_X2 FILLER_115_3735 ();
 FILLCELL_X1 FILLER_115_3737 ();
 FILLCELL_X32 FILLER_116_1 ();
 FILLCELL_X32 FILLER_116_33 ();
 FILLCELL_X32 FILLER_116_65 ();
 FILLCELL_X32 FILLER_116_97 ();
 FILLCELL_X32 FILLER_116_129 ();
 FILLCELL_X32 FILLER_116_161 ();
 FILLCELL_X32 FILLER_116_193 ();
 FILLCELL_X32 FILLER_116_225 ();
 FILLCELL_X32 FILLER_116_257 ();
 FILLCELL_X32 FILLER_116_289 ();
 FILLCELL_X32 FILLER_116_321 ();
 FILLCELL_X32 FILLER_116_353 ();
 FILLCELL_X32 FILLER_116_385 ();
 FILLCELL_X32 FILLER_116_417 ();
 FILLCELL_X32 FILLER_116_449 ();
 FILLCELL_X32 FILLER_116_481 ();
 FILLCELL_X32 FILLER_116_513 ();
 FILLCELL_X32 FILLER_116_545 ();
 FILLCELL_X32 FILLER_116_577 ();
 FILLCELL_X16 FILLER_116_609 ();
 FILLCELL_X4 FILLER_116_625 ();
 FILLCELL_X2 FILLER_116_629 ();
 FILLCELL_X32 FILLER_116_632 ();
 FILLCELL_X32 FILLER_116_664 ();
 FILLCELL_X32 FILLER_116_696 ();
 FILLCELL_X32 FILLER_116_728 ();
 FILLCELL_X32 FILLER_116_760 ();
 FILLCELL_X32 FILLER_116_792 ();
 FILLCELL_X32 FILLER_116_824 ();
 FILLCELL_X32 FILLER_116_856 ();
 FILLCELL_X32 FILLER_116_888 ();
 FILLCELL_X32 FILLER_116_920 ();
 FILLCELL_X32 FILLER_116_952 ();
 FILLCELL_X32 FILLER_116_984 ();
 FILLCELL_X32 FILLER_116_1016 ();
 FILLCELL_X32 FILLER_116_1048 ();
 FILLCELL_X32 FILLER_116_1080 ();
 FILLCELL_X32 FILLER_116_1112 ();
 FILLCELL_X32 FILLER_116_1144 ();
 FILLCELL_X32 FILLER_116_1176 ();
 FILLCELL_X32 FILLER_116_1208 ();
 FILLCELL_X32 FILLER_116_1240 ();
 FILLCELL_X32 FILLER_116_1272 ();
 FILLCELL_X32 FILLER_116_1304 ();
 FILLCELL_X32 FILLER_116_1336 ();
 FILLCELL_X32 FILLER_116_1368 ();
 FILLCELL_X32 FILLER_116_1400 ();
 FILLCELL_X32 FILLER_116_1432 ();
 FILLCELL_X32 FILLER_116_1464 ();
 FILLCELL_X32 FILLER_116_1496 ();
 FILLCELL_X32 FILLER_116_1528 ();
 FILLCELL_X32 FILLER_116_1560 ();
 FILLCELL_X32 FILLER_116_1592 ();
 FILLCELL_X32 FILLER_116_1624 ();
 FILLCELL_X32 FILLER_116_1656 ();
 FILLCELL_X32 FILLER_116_1688 ();
 FILLCELL_X32 FILLER_116_1720 ();
 FILLCELL_X32 FILLER_116_1752 ();
 FILLCELL_X32 FILLER_116_1784 ();
 FILLCELL_X32 FILLER_116_1816 ();
 FILLCELL_X32 FILLER_116_1848 ();
 FILLCELL_X8 FILLER_116_1880 ();
 FILLCELL_X4 FILLER_116_1888 ();
 FILLCELL_X2 FILLER_116_1892 ();
 FILLCELL_X32 FILLER_116_1895 ();
 FILLCELL_X32 FILLER_116_1927 ();
 FILLCELL_X32 FILLER_116_1959 ();
 FILLCELL_X32 FILLER_116_1991 ();
 FILLCELL_X32 FILLER_116_2023 ();
 FILLCELL_X32 FILLER_116_2055 ();
 FILLCELL_X32 FILLER_116_2087 ();
 FILLCELL_X32 FILLER_116_2119 ();
 FILLCELL_X32 FILLER_116_2151 ();
 FILLCELL_X32 FILLER_116_2183 ();
 FILLCELL_X32 FILLER_116_2215 ();
 FILLCELL_X32 FILLER_116_2247 ();
 FILLCELL_X32 FILLER_116_2279 ();
 FILLCELL_X32 FILLER_116_2311 ();
 FILLCELL_X32 FILLER_116_2343 ();
 FILLCELL_X32 FILLER_116_2375 ();
 FILLCELL_X32 FILLER_116_2407 ();
 FILLCELL_X32 FILLER_116_2439 ();
 FILLCELL_X32 FILLER_116_2471 ();
 FILLCELL_X32 FILLER_116_2503 ();
 FILLCELL_X32 FILLER_116_2535 ();
 FILLCELL_X32 FILLER_116_2567 ();
 FILLCELL_X32 FILLER_116_2599 ();
 FILLCELL_X32 FILLER_116_2631 ();
 FILLCELL_X32 FILLER_116_2663 ();
 FILLCELL_X32 FILLER_116_2695 ();
 FILLCELL_X32 FILLER_116_2727 ();
 FILLCELL_X32 FILLER_116_2759 ();
 FILLCELL_X32 FILLER_116_2791 ();
 FILLCELL_X32 FILLER_116_2823 ();
 FILLCELL_X32 FILLER_116_2855 ();
 FILLCELL_X32 FILLER_116_2887 ();
 FILLCELL_X32 FILLER_116_2919 ();
 FILLCELL_X32 FILLER_116_2951 ();
 FILLCELL_X32 FILLER_116_2983 ();
 FILLCELL_X32 FILLER_116_3015 ();
 FILLCELL_X32 FILLER_116_3047 ();
 FILLCELL_X32 FILLER_116_3079 ();
 FILLCELL_X32 FILLER_116_3111 ();
 FILLCELL_X8 FILLER_116_3143 ();
 FILLCELL_X4 FILLER_116_3151 ();
 FILLCELL_X2 FILLER_116_3155 ();
 FILLCELL_X32 FILLER_116_3158 ();
 FILLCELL_X32 FILLER_116_3190 ();
 FILLCELL_X32 FILLER_116_3222 ();
 FILLCELL_X32 FILLER_116_3254 ();
 FILLCELL_X32 FILLER_116_3286 ();
 FILLCELL_X32 FILLER_116_3318 ();
 FILLCELL_X32 FILLER_116_3350 ();
 FILLCELL_X32 FILLER_116_3382 ();
 FILLCELL_X32 FILLER_116_3414 ();
 FILLCELL_X32 FILLER_116_3446 ();
 FILLCELL_X32 FILLER_116_3478 ();
 FILLCELL_X32 FILLER_116_3510 ();
 FILLCELL_X32 FILLER_116_3542 ();
 FILLCELL_X32 FILLER_116_3574 ();
 FILLCELL_X32 FILLER_116_3606 ();
 FILLCELL_X32 FILLER_116_3638 ();
 FILLCELL_X32 FILLER_116_3670 ();
 FILLCELL_X32 FILLER_116_3702 ();
 FILLCELL_X4 FILLER_116_3734 ();
 FILLCELL_X32 FILLER_117_1 ();
 FILLCELL_X32 FILLER_117_33 ();
 FILLCELL_X32 FILLER_117_65 ();
 FILLCELL_X32 FILLER_117_97 ();
 FILLCELL_X32 FILLER_117_129 ();
 FILLCELL_X32 FILLER_117_161 ();
 FILLCELL_X32 FILLER_117_193 ();
 FILLCELL_X32 FILLER_117_225 ();
 FILLCELL_X32 FILLER_117_257 ();
 FILLCELL_X32 FILLER_117_289 ();
 FILLCELL_X32 FILLER_117_321 ();
 FILLCELL_X32 FILLER_117_353 ();
 FILLCELL_X32 FILLER_117_385 ();
 FILLCELL_X32 FILLER_117_417 ();
 FILLCELL_X32 FILLER_117_449 ();
 FILLCELL_X32 FILLER_117_481 ();
 FILLCELL_X32 FILLER_117_513 ();
 FILLCELL_X32 FILLER_117_545 ();
 FILLCELL_X32 FILLER_117_577 ();
 FILLCELL_X32 FILLER_117_609 ();
 FILLCELL_X32 FILLER_117_641 ();
 FILLCELL_X32 FILLER_117_673 ();
 FILLCELL_X32 FILLER_117_705 ();
 FILLCELL_X32 FILLER_117_737 ();
 FILLCELL_X32 FILLER_117_769 ();
 FILLCELL_X32 FILLER_117_801 ();
 FILLCELL_X32 FILLER_117_833 ();
 FILLCELL_X32 FILLER_117_865 ();
 FILLCELL_X32 FILLER_117_897 ();
 FILLCELL_X32 FILLER_117_929 ();
 FILLCELL_X32 FILLER_117_961 ();
 FILLCELL_X32 FILLER_117_993 ();
 FILLCELL_X32 FILLER_117_1025 ();
 FILLCELL_X32 FILLER_117_1057 ();
 FILLCELL_X32 FILLER_117_1089 ();
 FILLCELL_X32 FILLER_117_1121 ();
 FILLCELL_X32 FILLER_117_1153 ();
 FILLCELL_X32 FILLER_117_1185 ();
 FILLCELL_X32 FILLER_117_1217 ();
 FILLCELL_X8 FILLER_117_1249 ();
 FILLCELL_X4 FILLER_117_1257 ();
 FILLCELL_X2 FILLER_117_1261 ();
 FILLCELL_X32 FILLER_117_1264 ();
 FILLCELL_X32 FILLER_117_1296 ();
 FILLCELL_X32 FILLER_117_1328 ();
 FILLCELL_X32 FILLER_117_1360 ();
 FILLCELL_X32 FILLER_117_1392 ();
 FILLCELL_X32 FILLER_117_1424 ();
 FILLCELL_X32 FILLER_117_1456 ();
 FILLCELL_X32 FILLER_117_1488 ();
 FILLCELL_X32 FILLER_117_1520 ();
 FILLCELL_X32 FILLER_117_1552 ();
 FILLCELL_X32 FILLER_117_1584 ();
 FILLCELL_X32 FILLER_117_1616 ();
 FILLCELL_X32 FILLER_117_1648 ();
 FILLCELL_X32 FILLER_117_1680 ();
 FILLCELL_X32 FILLER_117_1712 ();
 FILLCELL_X32 FILLER_117_1744 ();
 FILLCELL_X32 FILLER_117_1776 ();
 FILLCELL_X32 FILLER_117_1808 ();
 FILLCELL_X32 FILLER_117_1840 ();
 FILLCELL_X32 FILLER_117_1872 ();
 FILLCELL_X32 FILLER_117_1904 ();
 FILLCELL_X32 FILLER_117_1936 ();
 FILLCELL_X32 FILLER_117_1968 ();
 FILLCELL_X32 FILLER_117_2000 ();
 FILLCELL_X32 FILLER_117_2032 ();
 FILLCELL_X32 FILLER_117_2064 ();
 FILLCELL_X32 FILLER_117_2096 ();
 FILLCELL_X32 FILLER_117_2128 ();
 FILLCELL_X32 FILLER_117_2160 ();
 FILLCELL_X32 FILLER_117_2192 ();
 FILLCELL_X32 FILLER_117_2224 ();
 FILLCELL_X32 FILLER_117_2256 ();
 FILLCELL_X32 FILLER_117_2288 ();
 FILLCELL_X32 FILLER_117_2320 ();
 FILLCELL_X32 FILLER_117_2352 ();
 FILLCELL_X32 FILLER_117_2384 ();
 FILLCELL_X32 FILLER_117_2416 ();
 FILLCELL_X32 FILLER_117_2448 ();
 FILLCELL_X32 FILLER_117_2480 ();
 FILLCELL_X8 FILLER_117_2512 ();
 FILLCELL_X4 FILLER_117_2520 ();
 FILLCELL_X2 FILLER_117_2524 ();
 FILLCELL_X32 FILLER_117_2527 ();
 FILLCELL_X32 FILLER_117_2559 ();
 FILLCELL_X32 FILLER_117_2591 ();
 FILLCELL_X32 FILLER_117_2623 ();
 FILLCELL_X32 FILLER_117_2655 ();
 FILLCELL_X32 FILLER_117_2687 ();
 FILLCELL_X32 FILLER_117_2719 ();
 FILLCELL_X32 FILLER_117_2751 ();
 FILLCELL_X32 FILLER_117_2783 ();
 FILLCELL_X32 FILLER_117_2815 ();
 FILLCELL_X32 FILLER_117_2847 ();
 FILLCELL_X32 FILLER_117_2879 ();
 FILLCELL_X32 FILLER_117_2911 ();
 FILLCELL_X32 FILLER_117_2943 ();
 FILLCELL_X32 FILLER_117_2975 ();
 FILLCELL_X32 FILLER_117_3007 ();
 FILLCELL_X32 FILLER_117_3039 ();
 FILLCELL_X32 FILLER_117_3071 ();
 FILLCELL_X32 FILLER_117_3103 ();
 FILLCELL_X32 FILLER_117_3135 ();
 FILLCELL_X32 FILLER_117_3167 ();
 FILLCELL_X32 FILLER_117_3199 ();
 FILLCELL_X32 FILLER_117_3231 ();
 FILLCELL_X32 FILLER_117_3263 ();
 FILLCELL_X32 FILLER_117_3295 ();
 FILLCELL_X32 FILLER_117_3327 ();
 FILLCELL_X32 FILLER_117_3359 ();
 FILLCELL_X32 FILLER_117_3391 ();
 FILLCELL_X32 FILLER_117_3423 ();
 FILLCELL_X32 FILLER_117_3455 ();
 FILLCELL_X32 FILLER_117_3487 ();
 FILLCELL_X32 FILLER_117_3519 ();
 FILLCELL_X32 FILLER_117_3551 ();
 FILLCELL_X32 FILLER_117_3583 ();
 FILLCELL_X32 FILLER_117_3615 ();
 FILLCELL_X32 FILLER_117_3647 ();
 FILLCELL_X32 FILLER_117_3679 ();
 FILLCELL_X16 FILLER_117_3711 ();
 FILLCELL_X8 FILLER_117_3727 ();
 FILLCELL_X2 FILLER_117_3735 ();
 FILLCELL_X1 FILLER_117_3737 ();
 FILLCELL_X32 FILLER_118_1 ();
 FILLCELL_X32 FILLER_118_33 ();
 FILLCELL_X32 FILLER_118_65 ();
 FILLCELL_X32 FILLER_118_97 ();
 FILLCELL_X32 FILLER_118_129 ();
 FILLCELL_X32 FILLER_118_161 ();
 FILLCELL_X32 FILLER_118_193 ();
 FILLCELL_X32 FILLER_118_225 ();
 FILLCELL_X32 FILLER_118_257 ();
 FILLCELL_X32 FILLER_118_289 ();
 FILLCELL_X32 FILLER_118_321 ();
 FILLCELL_X32 FILLER_118_353 ();
 FILLCELL_X32 FILLER_118_385 ();
 FILLCELL_X32 FILLER_118_417 ();
 FILLCELL_X32 FILLER_118_449 ();
 FILLCELL_X32 FILLER_118_481 ();
 FILLCELL_X32 FILLER_118_513 ();
 FILLCELL_X32 FILLER_118_545 ();
 FILLCELL_X32 FILLER_118_577 ();
 FILLCELL_X16 FILLER_118_609 ();
 FILLCELL_X4 FILLER_118_625 ();
 FILLCELL_X2 FILLER_118_629 ();
 FILLCELL_X32 FILLER_118_632 ();
 FILLCELL_X32 FILLER_118_664 ();
 FILLCELL_X32 FILLER_118_696 ();
 FILLCELL_X32 FILLER_118_728 ();
 FILLCELL_X32 FILLER_118_760 ();
 FILLCELL_X32 FILLER_118_792 ();
 FILLCELL_X32 FILLER_118_824 ();
 FILLCELL_X32 FILLER_118_856 ();
 FILLCELL_X32 FILLER_118_888 ();
 FILLCELL_X32 FILLER_118_920 ();
 FILLCELL_X32 FILLER_118_952 ();
 FILLCELL_X32 FILLER_118_984 ();
 FILLCELL_X32 FILLER_118_1016 ();
 FILLCELL_X32 FILLER_118_1048 ();
 FILLCELL_X32 FILLER_118_1080 ();
 FILLCELL_X32 FILLER_118_1112 ();
 FILLCELL_X32 FILLER_118_1144 ();
 FILLCELL_X32 FILLER_118_1176 ();
 FILLCELL_X32 FILLER_118_1208 ();
 FILLCELL_X32 FILLER_118_1240 ();
 FILLCELL_X32 FILLER_118_1272 ();
 FILLCELL_X32 FILLER_118_1304 ();
 FILLCELL_X32 FILLER_118_1336 ();
 FILLCELL_X32 FILLER_118_1368 ();
 FILLCELL_X32 FILLER_118_1400 ();
 FILLCELL_X32 FILLER_118_1432 ();
 FILLCELL_X32 FILLER_118_1464 ();
 FILLCELL_X32 FILLER_118_1496 ();
 FILLCELL_X32 FILLER_118_1528 ();
 FILLCELL_X32 FILLER_118_1560 ();
 FILLCELL_X32 FILLER_118_1592 ();
 FILLCELL_X32 FILLER_118_1624 ();
 FILLCELL_X32 FILLER_118_1656 ();
 FILLCELL_X32 FILLER_118_1688 ();
 FILLCELL_X32 FILLER_118_1720 ();
 FILLCELL_X32 FILLER_118_1752 ();
 FILLCELL_X32 FILLER_118_1784 ();
 FILLCELL_X32 FILLER_118_1816 ();
 FILLCELL_X32 FILLER_118_1848 ();
 FILLCELL_X8 FILLER_118_1880 ();
 FILLCELL_X4 FILLER_118_1888 ();
 FILLCELL_X2 FILLER_118_1892 ();
 FILLCELL_X32 FILLER_118_1895 ();
 FILLCELL_X32 FILLER_118_1927 ();
 FILLCELL_X32 FILLER_118_1959 ();
 FILLCELL_X32 FILLER_118_1991 ();
 FILLCELL_X32 FILLER_118_2023 ();
 FILLCELL_X32 FILLER_118_2055 ();
 FILLCELL_X32 FILLER_118_2087 ();
 FILLCELL_X32 FILLER_118_2119 ();
 FILLCELL_X32 FILLER_118_2151 ();
 FILLCELL_X32 FILLER_118_2183 ();
 FILLCELL_X32 FILLER_118_2215 ();
 FILLCELL_X32 FILLER_118_2247 ();
 FILLCELL_X32 FILLER_118_2279 ();
 FILLCELL_X32 FILLER_118_2311 ();
 FILLCELL_X32 FILLER_118_2343 ();
 FILLCELL_X32 FILLER_118_2375 ();
 FILLCELL_X32 FILLER_118_2407 ();
 FILLCELL_X32 FILLER_118_2439 ();
 FILLCELL_X32 FILLER_118_2471 ();
 FILLCELL_X32 FILLER_118_2503 ();
 FILLCELL_X32 FILLER_118_2535 ();
 FILLCELL_X32 FILLER_118_2567 ();
 FILLCELL_X32 FILLER_118_2599 ();
 FILLCELL_X32 FILLER_118_2631 ();
 FILLCELL_X32 FILLER_118_2663 ();
 FILLCELL_X32 FILLER_118_2695 ();
 FILLCELL_X32 FILLER_118_2727 ();
 FILLCELL_X32 FILLER_118_2759 ();
 FILLCELL_X32 FILLER_118_2791 ();
 FILLCELL_X32 FILLER_118_2823 ();
 FILLCELL_X32 FILLER_118_2855 ();
 FILLCELL_X32 FILLER_118_2887 ();
 FILLCELL_X32 FILLER_118_2919 ();
 FILLCELL_X32 FILLER_118_2951 ();
 FILLCELL_X32 FILLER_118_2983 ();
 FILLCELL_X32 FILLER_118_3015 ();
 FILLCELL_X32 FILLER_118_3047 ();
 FILLCELL_X32 FILLER_118_3079 ();
 FILLCELL_X32 FILLER_118_3111 ();
 FILLCELL_X8 FILLER_118_3143 ();
 FILLCELL_X4 FILLER_118_3151 ();
 FILLCELL_X2 FILLER_118_3155 ();
 FILLCELL_X32 FILLER_118_3158 ();
 FILLCELL_X32 FILLER_118_3190 ();
 FILLCELL_X32 FILLER_118_3222 ();
 FILLCELL_X32 FILLER_118_3254 ();
 FILLCELL_X32 FILLER_118_3286 ();
 FILLCELL_X32 FILLER_118_3318 ();
 FILLCELL_X32 FILLER_118_3350 ();
 FILLCELL_X32 FILLER_118_3382 ();
 FILLCELL_X32 FILLER_118_3414 ();
 FILLCELL_X32 FILLER_118_3446 ();
 FILLCELL_X32 FILLER_118_3478 ();
 FILLCELL_X32 FILLER_118_3510 ();
 FILLCELL_X32 FILLER_118_3542 ();
 FILLCELL_X32 FILLER_118_3574 ();
 FILLCELL_X32 FILLER_118_3606 ();
 FILLCELL_X32 FILLER_118_3638 ();
 FILLCELL_X32 FILLER_118_3670 ();
 FILLCELL_X32 FILLER_118_3702 ();
 FILLCELL_X4 FILLER_118_3734 ();
 FILLCELL_X32 FILLER_119_1 ();
 FILLCELL_X32 FILLER_119_33 ();
 FILLCELL_X32 FILLER_119_65 ();
 FILLCELL_X32 FILLER_119_97 ();
 FILLCELL_X32 FILLER_119_129 ();
 FILLCELL_X32 FILLER_119_161 ();
 FILLCELL_X32 FILLER_119_193 ();
 FILLCELL_X32 FILLER_119_225 ();
 FILLCELL_X32 FILLER_119_257 ();
 FILLCELL_X32 FILLER_119_289 ();
 FILLCELL_X32 FILLER_119_321 ();
 FILLCELL_X32 FILLER_119_353 ();
 FILLCELL_X32 FILLER_119_385 ();
 FILLCELL_X32 FILLER_119_417 ();
 FILLCELL_X32 FILLER_119_449 ();
 FILLCELL_X32 FILLER_119_481 ();
 FILLCELL_X32 FILLER_119_513 ();
 FILLCELL_X32 FILLER_119_545 ();
 FILLCELL_X32 FILLER_119_577 ();
 FILLCELL_X32 FILLER_119_609 ();
 FILLCELL_X32 FILLER_119_641 ();
 FILLCELL_X32 FILLER_119_673 ();
 FILLCELL_X32 FILLER_119_705 ();
 FILLCELL_X32 FILLER_119_737 ();
 FILLCELL_X32 FILLER_119_769 ();
 FILLCELL_X32 FILLER_119_801 ();
 FILLCELL_X32 FILLER_119_833 ();
 FILLCELL_X32 FILLER_119_865 ();
 FILLCELL_X32 FILLER_119_897 ();
 FILLCELL_X32 FILLER_119_929 ();
 FILLCELL_X32 FILLER_119_961 ();
 FILLCELL_X32 FILLER_119_993 ();
 FILLCELL_X32 FILLER_119_1025 ();
 FILLCELL_X32 FILLER_119_1057 ();
 FILLCELL_X32 FILLER_119_1089 ();
 FILLCELL_X32 FILLER_119_1121 ();
 FILLCELL_X32 FILLER_119_1153 ();
 FILLCELL_X32 FILLER_119_1185 ();
 FILLCELL_X32 FILLER_119_1217 ();
 FILLCELL_X8 FILLER_119_1249 ();
 FILLCELL_X4 FILLER_119_1257 ();
 FILLCELL_X2 FILLER_119_1261 ();
 FILLCELL_X32 FILLER_119_1264 ();
 FILLCELL_X32 FILLER_119_1296 ();
 FILLCELL_X32 FILLER_119_1328 ();
 FILLCELL_X32 FILLER_119_1360 ();
 FILLCELL_X32 FILLER_119_1392 ();
 FILLCELL_X32 FILLER_119_1424 ();
 FILLCELL_X32 FILLER_119_1456 ();
 FILLCELL_X32 FILLER_119_1488 ();
 FILLCELL_X32 FILLER_119_1520 ();
 FILLCELL_X32 FILLER_119_1552 ();
 FILLCELL_X32 FILLER_119_1584 ();
 FILLCELL_X32 FILLER_119_1616 ();
 FILLCELL_X32 FILLER_119_1648 ();
 FILLCELL_X32 FILLER_119_1680 ();
 FILLCELL_X32 FILLER_119_1712 ();
 FILLCELL_X32 FILLER_119_1744 ();
 FILLCELL_X32 FILLER_119_1776 ();
 FILLCELL_X32 FILLER_119_1808 ();
 FILLCELL_X32 FILLER_119_1840 ();
 FILLCELL_X32 FILLER_119_1872 ();
 FILLCELL_X32 FILLER_119_1904 ();
 FILLCELL_X32 FILLER_119_1936 ();
 FILLCELL_X32 FILLER_119_1968 ();
 FILLCELL_X32 FILLER_119_2000 ();
 FILLCELL_X32 FILLER_119_2032 ();
 FILLCELL_X32 FILLER_119_2064 ();
 FILLCELL_X32 FILLER_119_2096 ();
 FILLCELL_X32 FILLER_119_2128 ();
 FILLCELL_X32 FILLER_119_2160 ();
 FILLCELL_X32 FILLER_119_2192 ();
 FILLCELL_X32 FILLER_119_2224 ();
 FILLCELL_X32 FILLER_119_2256 ();
 FILLCELL_X32 FILLER_119_2288 ();
 FILLCELL_X32 FILLER_119_2320 ();
 FILLCELL_X32 FILLER_119_2352 ();
 FILLCELL_X32 FILLER_119_2384 ();
 FILLCELL_X32 FILLER_119_2416 ();
 FILLCELL_X32 FILLER_119_2448 ();
 FILLCELL_X32 FILLER_119_2480 ();
 FILLCELL_X8 FILLER_119_2512 ();
 FILLCELL_X4 FILLER_119_2520 ();
 FILLCELL_X2 FILLER_119_2524 ();
 FILLCELL_X32 FILLER_119_2527 ();
 FILLCELL_X32 FILLER_119_2559 ();
 FILLCELL_X32 FILLER_119_2591 ();
 FILLCELL_X32 FILLER_119_2623 ();
 FILLCELL_X32 FILLER_119_2655 ();
 FILLCELL_X32 FILLER_119_2687 ();
 FILLCELL_X32 FILLER_119_2719 ();
 FILLCELL_X32 FILLER_119_2751 ();
 FILLCELL_X32 FILLER_119_2783 ();
 FILLCELL_X32 FILLER_119_2815 ();
 FILLCELL_X32 FILLER_119_2847 ();
 FILLCELL_X32 FILLER_119_2879 ();
 FILLCELL_X32 FILLER_119_2911 ();
 FILLCELL_X32 FILLER_119_2943 ();
 FILLCELL_X32 FILLER_119_2975 ();
 FILLCELL_X32 FILLER_119_3007 ();
 FILLCELL_X32 FILLER_119_3039 ();
 FILLCELL_X32 FILLER_119_3071 ();
 FILLCELL_X32 FILLER_119_3103 ();
 FILLCELL_X32 FILLER_119_3135 ();
 FILLCELL_X32 FILLER_119_3167 ();
 FILLCELL_X32 FILLER_119_3199 ();
 FILLCELL_X32 FILLER_119_3231 ();
 FILLCELL_X32 FILLER_119_3263 ();
 FILLCELL_X32 FILLER_119_3295 ();
 FILLCELL_X32 FILLER_119_3327 ();
 FILLCELL_X32 FILLER_119_3359 ();
 FILLCELL_X32 FILLER_119_3391 ();
 FILLCELL_X32 FILLER_119_3423 ();
 FILLCELL_X32 FILLER_119_3455 ();
 FILLCELL_X32 FILLER_119_3487 ();
 FILLCELL_X32 FILLER_119_3519 ();
 FILLCELL_X32 FILLER_119_3551 ();
 FILLCELL_X32 FILLER_119_3583 ();
 FILLCELL_X32 FILLER_119_3615 ();
 FILLCELL_X32 FILLER_119_3647 ();
 FILLCELL_X32 FILLER_119_3679 ();
 FILLCELL_X16 FILLER_119_3711 ();
 FILLCELL_X8 FILLER_119_3727 ();
 FILLCELL_X2 FILLER_119_3735 ();
 FILLCELL_X1 FILLER_119_3737 ();
 FILLCELL_X32 FILLER_120_1 ();
 FILLCELL_X32 FILLER_120_33 ();
 FILLCELL_X32 FILLER_120_65 ();
 FILLCELL_X32 FILLER_120_97 ();
 FILLCELL_X32 FILLER_120_129 ();
 FILLCELL_X32 FILLER_120_161 ();
 FILLCELL_X32 FILLER_120_193 ();
 FILLCELL_X32 FILLER_120_225 ();
 FILLCELL_X32 FILLER_120_257 ();
 FILLCELL_X32 FILLER_120_289 ();
 FILLCELL_X32 FILLER_120_321 ();
 FILLCELL_X32 FILLER_120_353 ();
 FILLCELL_X32 FILLER_120_385 ();
 FILLCELL_X32 FILLER_120_417 ();
 FILLCELL_X32 FILLER_120_449 ();
 FILLCELL_X32 FILLER_120_481 ();
 FILLCELL_X32 FILLER_120_513 ();
 FILLCELL_X32 FILLER_120_545 ();
 FILLCELL_X32 FILLER_120_577 ();
 FILLCELL_X16 FILLER_120_609 ();
 FILLCELL_X4 FILLER_120_625 ();
 FILLCELL_X2 FILLER_120_629 ();
 FILLCELL_X32 FILLER_120_632 ();
 FILLCELL_X32 FILLER_120_664 ();
 FILLCELL_X32 FILLER_120_696 ();
 FILLCELL_X32 FILLER_120_728 ();
 FILLCELL_X32 FILLER_120_760 ();
 FILLCELL_X32 FILLER_120_792 ();
 FILLCELL_X32 FILLER_120_824 ();
 FILLCELL_X32 FILLER_120_856 ();
 FILLCELL_X32 FILLER_120_888 ();
 FILLCELL_X32 FILLER_120_920 ();
 FILLCELL_X32 FILLER_120_952 ();
 FILLCELL_X32 FILLER_120_984 ();
 FILLCELL_X32 FILLER_120_1016 ();
 FILLCELL_X32 FILLER_120_1048 ();
 FILLCELL_X32 FILLER_120_1080 ();
 FILLCELL_X32 FILLER_120_1112 ();
 FILLCELL_X32 FILLER_120_1144 ();
 FILLCELL_X32 FILLER_120_1176 ();
 FILLCELL_X32 FILLER_120_1208 ();
 FILLCELL_X32 FILLER_120_1240 ();
 FILLCELL_X32 FILLER_120_1272 ();
 FILLCELL_X32 FILLER_120_1304 ();
 FILLCELL_X32 FILLER_120_1336 ();
 FILLCELL_X32 FILLER_120_1368 ();
 FILLCELL_X32 FILLER_120_1400 ();
 FILLCELL_X32 FILLER_120_1432 ();
 FILLCELL_X32 FILLER_120_1464 ();
 FILLCELL_X32 FILLER_120_1496 ();
 FILLCELL_X32 FILLER_120_1528 ();
 FILLCELL_X32 FILLER_120_1560 ();
 FILLCELL_X32 FILLER_120_1592 ();
 FILLCELL_X32 FILLER_120_1624 ();
 FILLCELL_X32 FILLER_120_1656 ();
 FILLCELL_X32 FILLER_120_1688 ();
 FILLCELL_X32 FILLER_120_1720 ();
 FILLCELL_X32 FILLER_120_1752 ();
 FILLCELL_X32 FILLER_120_1784 ();
 FILLCELL_X32 FILLER_120_1816 ();
 FILLCELL_X32 FILLER_120_1848 ();
 FILLCELL_X8 FILLER_120_1880 ();
 FILLCELL_X4 FILLER_120_1888 ();
 FILLCELL_X2 FILLER_120_1892 ();
 FILLCELL_X32 FILLER_120_1895 ();
 FILLCELL_X32 FILLER_120_1927 ();
 FILLCELL_X32 FILLER_120_1959 ();
 FILLCELL_X32 FILLER_120_1991 ();
 FILLCELL_X32 FILLER_120_2023 ();
 FILLCELL_X32 FILLER_120_2055 ();
 FILLCELL_X32 FILLER_120_2087 ();
 FILLCELL_X32 FILLER_120_2119 ();
 FILLCELL_X32 FILLER_120_2151 ();
 FILLCELL_X32 FILLER_120_2183 ();
 FILLCELL_X32 FILLER_120_2215 ();
 FILLCELL_X32 FILLER_120_2247 ();
 FILLCELL_X32 FILLER_120_2279 ();
 FILLCELL_X32 FILLER_120_2311 ();
 FILLCELL_X32 FILLER_120_2343 ();
 FILLCELL_X32 FILLER_120_2375 ();
 FILLCELL_X32 FILLER_120_2407 ();
 FILLCELL_X32 FILLER_120_2439 ();
 FILLCELL_X32 FILLER_120_2471 ();
 FILLCELL_X32 FILLER_120_2503 ();
 FILLCELL_X32 FILLER_120_2535 ();
 FILLCELL_X32 FILLER_120_2567 ();
 FILLCELL_X32 FILLER_120_2599 ();
 FILLCELL_X32 FILLER_120_2631 ();
 FILLCELL_X32 FILLER_120_2663 ();
 FILLCELL_X32 FILLER_120_2695 ();
 FILLCELL_X32 FILLER_120_2727 ();
 FILLCELL_X32 FILLER_120_2759 ();
 FILLCELL_X32 FILLER_120_2791 ();
 FILLCELL_X32 FILLER_120_2823 ();
 FILLCELL_X32 FILLER_120_2855 ();
 FILLCELL_X32 FILLER_120_2887 ();
 FILLCELL_X32 FILLER_120_2919 ();
 FILLCELL_X32 FILLER_120_2951 ();
 FILLCELL_X32 FILLER_120_2983 ();
 FILLCELL_X32 FILLER_120_3015 ();
 FILLCELL_X32 FILLER_120_3047 ();
 FILLCELL_X32 FILLER_120_3079 ();
 FILLCELL_X32 FILLER_120_3111 ();
 FILLCELL_X8 FILLER_120_3143 ();
 FILLCELL_X4 FILLER_120_3151 ();
 FILLCELL_X2 FILLER_120_3155 ();
 FILLCELL_X32 FILLER_120_3158 ();
 FILLCELL_X32 FILLER_120_3190 ();
 FILLCELL_X32 FILLER_120_3222 ();
 FILLCELL_X32 FILLER_120_3254 ();
 FILLCELL_X32 FILLER_120_3286 ();
 FILLCELL_X32 FILLER_120_3318 ();
 FILLCELL_X32 FILLER_120_3350 ();
 FILLCELL_X32 FILLER_120_3382 ();
 FILLCELL_X32 FILLER_120_3414 ();
 FILLCELL_X32 FILLER_120_3446 ();
 FILLCELL_X32 FILLER_120_3478 ();
 FILLCELL_X32 FILLER_120_3510 ();
 FILLCELL_X32 FILLER_120_3542 ();
 FILLCELL_X32 FILLER_120_3574 ();
 FILLCELL_X32 FILLER_120_3606 ();
 FILLCELL_X32 FILLER_120_3638 ();
 FILLCELL_X32 FILLER_120_3670 ();
 FILLCELL_X32 FILLER_120_3702 ();
 FILLCELL_X4 FILLER_120_3734 ();
 FILLCELL_X32 FILLER_121_1 ();
 FILLCELL_X32 FILLER_121_33 ();
 FILLCELL_X32 FILLER_121_65 ();
 FILLCELL_X32 FILLER_121_97 ();
 FILLCELL_X32 FILLER_121_129 ();
 FILLCELL_X32 FILLER_121_161 ();
 FILLCELL_X32 FILLER_121_193 ();
 FILLCELL_X32 FILLER_121_225 ();
 FILLCELL_X32 FILLER_121_257 ();
 FILLCELL_X32 FILLER_121_289 ();
 FILLCELL_X32 FILLER_121_321 ();
 FILLCELL_X32 FILLER_121_353 ();
 FILLCELL_X32 FILLER_121_385 ();
 FILLCELL_X32 FILLER_121_417 ();
 FILLCELL_X32 FILLER_121_449 ();
 FILLCELL_X32 FILLER_121_481 ();
 FILLCELL_X32 FILLER_121_513 ();
 FILLCELL_X32 FILLER_121_545 ();
 FILLCELL_X32 FILLER_121_577 ();
 FILLCELL_X32 FILLER_121_609 ();
 FILLCELL_X32 FILLER_121_641 ();
 FILLCELL_X32 FILLER_121_673 ();
 FILLCELL_X32 FILLER_121_705 ();
 FILLCELL_X32 FILLER_121_737 ();
 FILLCELL_X32 FILLER_121_769 ();
 FILLCELL_X32 FILLER_121_801 ();
 FILLCELL_X32 FILLER_121_833 ();
 FILLCELL_X32 FILLER_121_865 ();
 FILLCELL_X32 FILLER_121_897 ();
 FILLCELL_X32 FILLER_121_929 ();
 FILLCELL_X32 FILLER_121_961 ();
 FILLCELL_X32 FILLER_121_993 ();
 FILLCELL_X32 FILLER_121_1025 ();
 FILLCELL_X32 FILLER_121_1057 ();
 FILLCELL_X32 FILLER_121_1089 ();
 FILLCELL_X32 FILLER_121_1121 ();
 FILLCELL_X32 FILLER_121_1153 ();
 FILLCELL_X32 FILLER_121_1185 ();
 FILLCELL_X32 FILLER_121_1217 ();
 FILLCELL_X8 FILLER_121_1249 ();
 FILLCELL_X4 FILLER_121_1257 ();
 FILLCELL_X2 FILLER_121_1261 ();
 FILLCELL_X32 FILLER_121_1264 ();
 FILLCELL_X32 FILLER_121_1296 ();
 FILLCELL_X32 FILLER_121_1328 ();
 FILLCELL_X32 FILLER_121_1360 ();
 FILLCELL_X32 FILLER_121_1392 ();
 FILLCELL_X32 FILLER_121_1424 ();
 FILLCELL_X32 FILLER_121_1456 ();
 FILLCELL_X32 FILLER_121_1488 ();
 FILLCELL_X32 FILLER_121_1520 ();
 FILLCELL_X32 FILLER_121_1552 ();
 FILLCELL_X32 FILLER_121_1584 ();
 FILLCELL_X32 FILLER_121_1616 ();
 FILLCELL_X32 FILLER_121_1648 ();
 FILLCELL_X32 FILLER_121_1680 ();
 FILLCELL_X32 FILLER_121_1712 ();
 FILLCELL_X32 FILLER_121_1744 ();
 FILLCELL_X32 FILLER_121_1776 ();
 FILLCELL_X32 FILLER_121_1808 ();
 FILLCELL_X32 FILLER_121_1840 ();
 FILLCELL_X32 FILLER_121_1872 ();
 FILLCELL_X32 FILLER_121_1904 ();
 FILLCELL_X32 FILLER_121_1936 ();
 FILLCELL_X32 FILLER_121_1968 ();
 FILLCELL_X32 FILLER_121_2000 ();
 FILLCELL_X32 FILLER_121_2032 ();
 FILLCELL_X32 FILLER_121_2064 ();
 FILLCELL_X32 FILLER_121_2096 ();
 FILLCELL_X32 FILLER_121_2128 ();
 FILLCELL_X32 FILLER_121_2160 ();
 FILLCELL_X32 FILLER_121_2192 ();
 FILLCELL_X32 FILLER_121_2224 ();
 FILLCELL_X32 FILLER_121_2256 ();
 FILLCELL_X32 FILLER_121_2288 ();
 FILLCELL_X32 FILLER_121_2320 ();
 FILLCELL_X32 FILLER_121_2352 ();
 FILLCELL_X32 FILLER_121_2384 ();
 FILLCELL_X32 FILLER_121_2416 ();
 FILLCELL_X32 FILLER_121_2448 ();
 FILLCELL_X32 FILLER_121_2480 ();
 FILLCELL_X8 FILLER_121_2512 ();
 FILLCELL_X4 FILLER_121_2520 ();
 FILLCELL_X2 FILLER_121_2524 ();
 FILLCELL_X32 FILLER_121_2527 ();
 FILLCELL_X32 FILLER_121_2559 ();
 FILLCELL_X32 FILLER_121_2591 ();
 FILLCELL_X32 FILLER_121_2623 ();
 FILLCELL_X32 FILLER_121_2655 ();
 FILLCELL_X32 FILLER_121_2687 ();
 FILLCELL_X32 FILLER_121_2719 ();
 FILLCELL_X32 FILLER_121_2751 ();
 FILLCELL_X32 FILLER_121_2783 ();
 FILLCELL_X32 FILLER_121_2815 ();
 FILLCELL_X32 FILLER_121_2847 ();
 FILLCELL_X32 FILLER_121_2879 ();
 FILLCELL_X32 FILLER_121_2911 ();
 FILLCELL_X32 FILLER_121_2943 ();
 FILLCELL_X32 FILLER_121_2975 ();
 FILLCELL_X32 FILLER_121_3007 ();
 FILLCELL_X32 FILLER_121_3039 ();
 FILLCELL_X32 FILLER_121_3071 ();
 FILLCELL_X32 FILLER_121_3103 ();
 FILLCELL_X32 FILLER_121_3135 ();
 FILLCELL_X32 FILLER_121_3167 ();
 FILLCELL_X32 FILLER_121_3199 ();
 FILLCELL_X32 FILLER_121_3231 ();
 FILLCELL_X32 FILLER_121_3263 ();
 FILLCELL_X32 FILLER_121_3295 ();
 FILLCELL_X32 FILLER_121_3327 ();
 FILLCELL_X32 FILLER_121_3359 ();
 FILLCELL_X32 FILLER_121_3391 ();
 FILLCELL_X32 FILLER_121_3423 ();
 FILLCELL_X32 FILLER_121_3455 ();
 FILLCELL_X32 FILLER_121_3487 ();
 FILLCELL_X32 FILLER_121_3519 ();
 FILLCELL_X32 FILLER_121_3551 ();
 FILLCELL_X32 FILLER_121_3583 ();
 FILLCELL_X32 FILLER_121_3615 ();
 FILLCELL_X32 FILLER_121_3647 ();
 FILLCELL_X32 FILLER_121_3679 ();
 FILLCELL_X16 FILLER_121_3711 ();
 FILLCELL_X8 FILLER_121_3727 ();
 FILLCELL_X2 FILLER_121_3735 ();
 FILLCELL_X1 FILLER_121_3737 ();
 FILLCELL_X32 FILLER_122_1 ();
 FILLCELL_X32 FILLER_122_33 ();
 FILLCELL_X32 FILLER_122_65 ();
 FILLCELL_X32 FILLER_122_97 ();
 FILLCELL_X32 FILLER_122_129 ();
 FILLCELL_X32 FILLER_122_161 ();
 FILLCELL_X32 FILLER_122_193 ();
 FILLCELL_X32 FILLER_122_225 ();
 FILLCELL_X32 FILLER_122_257 ();
 FILLCELL_X32 FILLER_122_289 ();
 FILLCELL_X32 FILLER_122_321 ();
 FILLCELL_X32 FILLER_122_353 ();
 FILLCELL_X32 FILLER_122_385 ();
 FILLCELL_X32 FILLER_122_417 ();
 FILLCELL_X32 FILLER_122_449 ();
 FILLCELL_X32 FILLER_122_481 ();
 FILLCELL_X32 FILLER_122_513 ();
 FILLCELL_X32 FILLER_122_545 ();
 FILLCELL_X32 FILLER_122_577 ();
 FILLCELL_X16 FILLER_122_609 ();
 FILLCELL_X4 FILLER_122_625 ();
 FILLCELL_X2 FILLER_122_629 ();
 FILLCELL_X32 FILLER_122_632 ();
 FILLCELL_X32 FILLER_122_664 ();
 FILLCELL_X32 FILLER_122_696 ();
 FILLCELL_X32 FILLER_122_728 ();
 FILLCELL_X32 FILLER_122_760 ();
 FILLCELL_X32 FILLER_122_792 ();
 FILLCELL_X32 FILLER_122_824 ();
 FILLCELL_X32 FILLER_122_856 ();
 FILLCELL_X32 FILLER_122_888 ();
 FILLCELL_X32 FILLER_122_920 ();
 FILLCELL_X32 FILLER_122_952 ();
 FILLCELL_X32 FILLER_122_984 ();
 FILLCELL_X32 FILLER_122_1016 ();
 FILLCELL_X32 FILLER_122_1048 ();
 FILLCELL_X32 FILLER_122_1080 ();
 FILLCELL_X32 FILLER_122_1112 ();
 FILLCELL_X32 FILLER_122_1144 ();
 FILLCELL_X32 FILLER_122_1176 ();
 FILLCELL_X32 FILLER_122_1208 ();
 FILLCELL_X32 FILLER_122_1240 ();
 FILLCELL_X32 FILLER_122_1272 ();
 FILLCELL_X32 FILLER_122_1304 ();
 FILLCELL_X32 FILLER_122_1336 ();
 FILLCELL_X32 FILLER_122_1368 ();
 FILLCELL_X32 FILLER_122_1400 ();
 FILLCELL_X32 FILLER_122_1432 ();
 FILLCELL_X32 FILLER_122_1464 ();
 FILLCELL_X32 FILLER_122_1496 ();
 FILLCELL_X32 FILLER_122_1528 ();
 FILLCELL_X32 FILLER_122_1560 ();
 FILLCELL_X32 FILLER_122_1592 ();
 FILLCELL_X32 FILLER_122_1624 ();
 FILLCELL_X32 FILLER_122_1656 ();
 FILLCELL_X32 FILLER_122_1688 ();
 FILLCELL_X32 FILLER_122_1720 ();
 FILLCELL_X32 FILLER_122_1752 ();
 FILLCELL_X32 FILLER_122_1784 ();
 FILLCELL_X32 FILLER_122_1816 ();
 FILLCELL_X32 FILLER_122_1848 ();
 FILLCELL_X8 FILLER_122_1880 ();
 FILLCELL_X4 FILLER_122_1888 ();
 FILLCELL_X2 FILLER_122_1892 ();
 FILLCELL_X32 FILLER_122_1895 ();
 FILLCELL_X32 FILLER_122_1927 ();
 FILLCELL_X32 FILLER_122_1959 ();
 FILLCELL_X32 FILLER_122_1991 ();
 FILLCELL_X32 FILLER_122_2023 ();
 FILLCELL_X32 FILLER_122_2055 ();
 FILLCELL_X32 FILLER_122_2087 ();
 FILLCELL_X32 FILLER_122_2119 ();
 FILLCELL_X32 FILLER_122_2151 ();
 FILLCELL_X32 FILLER_122_2183 ();
 FILLCELL_X32 FILLER_122_2215 ();
 FILLCELL_X32 FILLER_122_2247 ();
 FILLCELL_X32 FILLER_122_2279 ();
 FILLCELL_X32 FILLER_122_2311 ();
 FILLCELL_X32 FILLER_122_2343 ();
 FILLCELL_X32 FILLER_122_2375 ();
 FILLCELL_X32 FILLER_122_2407 ();
 FILLCELL_X32 FILLER_122_2439 ();
 FILLCELL_X32 FILLER_122_2471 ();
 FILLCELL_X32 FILLER_122_2503 ();
 FILLCELL_X32 FILLER_122_2535 ();
 FILLCELL_X32 FILLER_122_2567 ();
 FILLCELL_X32 FILLER_122_2599 ();
 FILLCELL_X32 FILLER_122_2631 ();
 FILLCELL_X32 FILLER_122_2663 ();
 FILLCELL_X32 FILLER_122_2695 ();
 FILLCELL_X32 FILLER_122_2727 ();
 FILLCELL_X32 FILLER_122_2759 ();
 FILLCELL_X32 FILLER_122_2791 ();
 FILLCELL_X32 FILLER_122_2823 ();
 FILLCELL_X32 FILLER_122_2855 ();
 FILLCELL_X32 FILLER_122_2887 ();
 FILLCELL_X32 FILLER_122_2919 ();
 FILLCELL_X32 FILLER_122_2951 ();
 FILLCELL_X32 FILLER_122_2983 ();
 FILLCELL_X32 FILLER_122_3015 ();
 FILLCELL_X32 FILLER_122_3047 ();
 FILLCELL_X32 FILLER_122_3079 ();
 FILLCELL_X32 FILLER_122_3111 ();
 FILLCELL_X8 FILLER_122_3143 ();
 FILLCELL_X4 FILLER_122_3151 ();
 FILLCELL_X2 FILLER_122_3155 ();
 FILLCELL_X32 FILLER_122_3158 ();
 FILLCELL_X32 FILLER_122_3190 ();
 FILLCELL_X32 FILLER_122_3222 ();
 FILLCELL_X32 FILLER_122_3254 ();
 FILLCELL_X32 FILLER_122_3286 ();
 FILLCELL_X32 FILLER_122_3318 ();
 FILLCELL_X32 FILLER_122_3350 ();
 FILLCELL_X32 FILLER_122_3382 ();
 FILLCELL_X32 FILLER_122_3414 ();
 FILLCELL_X32 FILLER_122_3446 ();
 FILLCELL_X32 FILLER_122_3478 ();
 FILLCELL_X32 FILLER_122_3510 ();
 FILLCELL_X32 FILLER_122_3542 ();
 FILLCELL_X32 FILLER_122_3574 ();
 FILLCELL_X32 FILLER_122_3606 ();
 FILLCELL_X32 FILLER_122_3638 ();
 FILLCELL_X32 FILLER_122_3670 ();
 FILLCELL_X32 FILLER_122_3702 ();
 FILLCELL_X4 FILLER_122_3734 ();
 FILLCELL_X32 FILLER_123_1 ();
 FILLCELL_X32 FILLER_123_33 ();
 FILLCELL_X32 FILLER_123_65 ();
 FILLCELL_X32 FILLER_123_97 ();
 FILLCELL_X32 FILLER_123_129 ();
 FILLCELL_X32 FILLER_123_161 ();
 FILLCELL_X32 FILLER_123_193 ();
 FILLCELL_X32 FILLER_123_225 ();
 FILLCELL_X32 FILLER_123_257 ();
 FILLCELL_X32 FILLER_123_289 ();
 FILLCELL_X32 FILLER_123_321 ();
 FILLCELL_X32 FILLER_123_353 ();
 FILLCELL_X32 FILLER_123_385 ();
 FILLCELL_X32 FILLER_123_417 ();
 FILLCELL_X32 FILLER_123_449 ();
 FILLCELL_X32 FILLER_123_481 ();
 FILLCELL_X32 FILLER_123_513 ();
 FILLCELL_X32 FILLER_123_545 ();
 FILLCELL_X32 FILLER_123_577 ();
 FILLCELL_X32 FILLER_123_609 ();
 FILLCELL_X32 FILLER_123_641 ();
 FILLCELL_X32 FILLER_123_673 ();
 FILLCELL_X32 FILLER_123_705 ();
 FILLCELL_X32 FILLER_123_737 ();
 FILLCELL_X32 FILLER_123_769 ();
 FILLCELL_X32 FILLER_123_801 ();
 FILLCELL_X32 FILLER_123_833 ();
 FILLCELL_X32 FILLER_123_865 ();
 FILLCELL_X32 FILLER_123_897 ();
 FILLCELL_X32 FILLER_123_929 ();
 FILLCELL_X32 FILLER_123_961 ();
 FILLCELL_X32 FILLER_123_993 ();
 FILLCELL_X32 FILLER_123_1025 ();
 FILLCELL_X32 FILLER_123_1057 ();
 FILLCELL_X32 FILLER_123_1089 ();
 FILLCELL_X32 FILLER_123_1121 ();
 FILLCELL_X32 FILLER_123_1153 ();
 FILLCELL_X32 FILLER_123_1185 ();
 FILLCELL_X32 FILLER_123_1217 ();
 FILLCELL_X8 FILLER_123_1249 ();
 FILLCELL_X4 FILLER_123_1257 ();
 FILLCELL_X2 FILLER_123_1261 ();
 FILLCELL_X32 FILLER_123_1264 ();
 FILLCELL_X32 FILLER_123_1296 ();
 FILLCELL_X32 FILLER_123_1328 ();
 FILLCELL_X32 FILLER_123_1360 ();
 FILLCELL_X32 FILLER_123_1392 ();
 FILLCELL_X32 FILLER_123_1424 ();
 FILLCELL_X32 FILLER_123_1456 ();
 FILLCELL_X32 FILLER_123_1488 ();
 FILLCELL_X32 FILLER_123_1520 ();
 FILLCELL_X32 FILLER_123_1552 ();
 FILLCELL_X32 FILLER_123_1584 ();
 FILLCELL_X32 FILLER_123_1616 ();
 FILLCELL_X32 FILLER_123_1648 ();
 FILLCELL_X32 FILLER_123_1680 ();
 FILLCELL_X32 FILLER_123_1712 ();
 FILLCELL_X32 FILLER_123_1744 ();
 FILLCELL_X32 FILLER_123_1776 ();
 FILLCELL_X32 FILLER_123_1808 ();
 FILLCELL_X32 FILLER_123_1840 ();
 FILLCELL_X32 FILLER_123_1872 ();
 FILLCELL_X32 FILLER_123_1904 ();
 FILLCELL_X32 FILLER_123_1936 ();
 FILLCELL_X32 FILLER_123_1968 ();
 FILLCELL_X32 FILLER_123_2000 ();
 FILLCELL_X32 FILLER_123_2032 ();
 FILLCELL_X32 FILLER_123_2064 ();
 FILLCELL_X32 FILLER_123_2096 ();
 FILLCELL_X32 FILLER_123_2128 ();
 FILLCELL_X32 FILLER_123_2160 ();
 FILLCELL_X32 FILLER_123_2192 ();
 FILLCELL_X32 FILLER_123_2224 ();
 FILLCELL_X32 FILLER_123_2256 ();
 FILLCELL_X32 FILLER_123_2288 ();
 FILLCELL_X32 FILLER_123_2320 ();
 FILLCELL_X32 FILLER_123_2352 ();
 FILLCELL_X32 FILLER_123_2384 ();
 FILLCELL_X32 FILLER_123_2416 ();
 FILLCELL_X32 FILLER_123_2448 ();
 FILLCELL_X32 FILLER_123_2480 ();
 FILLCELL_X8 FILLER_123_2512 ();
 FILLCELL_X4 FILLER_123_2520 ();
 FILLCELL_X2 FILLER_123_2524 ();
 FILLCELL_X32 FILLER_123_2527 ();
 FILLCELL_X32 FILLER_123_2559 ();
 FILLCELL_X32 FILLER_123_2591 ();
 FILLCELL_X32 FILLER_123_2623 ();
 FILLCELL_X32 FILLER_123_2655 ();
 FILLCELL_X32 FILLER_123_2687 ();
 FILLCELL_X32 FILLER_123_2719 ();
 FILLCELL_X32 FILLER_123_2751 ();
 FILLCELL_X32 FILLER_123_2783 ();
 FILLCELL_X32 FILLER_123_2815 ();
 FILLCELL_X32 FILLER_123_2847 ();
 FILLCELL_X32 FILLER_123_2879 ();
 FILLCELL_X32 FILLER_123_2911 ();
 FILLCELL_X32 FILLER_123_2943 ();
 FILLCELL_X32 FILLER_123_2975 ();
 FILLCELL_X32 FILLER_123_3007 ();
 FILLCELL_X32 FILLER_123_3039 ();
 FILLCELL_X32 FILLER_123_3071 ();
 FILLCELL_X32 FILLER_123_3103 ();
 FILLCELL_X32 FILLER_123_3135 ();
 FILLCELL_X32 FILLER_123_3167 ();
 FILLCELL_X32 FILLER_123_3199 ();
 FILLCELL_X32 FILLER_123_3231 ();
 FILLCELL_X32 FILLER_123_3263 ();
 FILLCELL_X32 FILLER_123_3295 ();
 FILLCELL_X32 FILLER_123_3327 ();
 FILLCELL_X32 FILLER_123_3359 ();
 FILLCELL_X32 FILLER_123_3391 ();
 FILLCELL_X32 FILLER_123_3423 ();
 FILLCELL_X32 FILLER_123_3455 ();
 FILLCELL_X32 FILLER_123_3487 ();
 FILLCELL_X32 FILLER_123_3519 ();
 FILLCELL_X32 FILLER_123_3551 ();
 FILLCELL_X32 FILLER_123_3583 ();
 FILLCELL_X32 FILLER_123_3615 ();
 FILLCELL_X32 FILLER_123_3647 ();
 FILLCELL_X32 FILLER_123_3679 ();
 FILLCELL_X16 FILLER_123_3711 ();
 FILLCELL_X8 FILLER_123_3727 ();
 FILLCELL_X2 FILLER_123_3735 ();
 FILLCELL_X1 FILLER_123_3737 ();
 FILLCELL_X32 FILLER_124_1 ();
 FILLCELL_X32 FILLER_124_33 ();
 FILLCELL_X32 FILLER_124_65 ();
 FILLCELL_X32 FILLER_124_97 ();
 FILLCELL_X32 FILLER_124_129 ();
 FILLCELL_X32 FILLER_124_161 ();
 FILLCELL_X32 FILLER_124_193 ();
 FILLCELL_X32 FILLER_124_225 ();
 FILLCELL_X32 FILLER_124_257 ();
 FILLCELL_X32 FILLER_124_289 ();
 FILLCELL_X32 FILLER_124_321 ();
 FILLCELL_X32 FILLER_124_353 ();
 FILLCELL_X32 FILLER_124_385 ();
 FILLCELL_X32 FILLER_124_417 ();
 FILLCELL_X32 FILLER_124_449 ();
 FILLCELL_X32 FILLER_124_481 ();
 FILLCELL_X32 FILLER_124_513 ();
 FILLCELL_X32 FILLER_124_545 ();
 FILLCELL_X32 FILLER_124_577 ();
 FILLCELL_X16 FILLER_124_609 ();
 FILLCELL_X4 FILLER_124_625 ();
 FILLCELL_X2 FILLER_124_629 ();
 FILLCELL_X32 FILLER_124_632 ();
 FILLCELL_X32 FILLER_124_664 ();
 FILLCELL_X32 FILLER_124_696 ();
 FILLCELL_X32 FILLER_124_728 ();
 FILLCELL_X32 FILLER_124_760 ();
 FILLCELL_X32 FILLER_124_792 ();
 FILLCELL_X32 FILLER_124_824 ();
 FILLCELL_X32 FILLER_124_856 ();
 FILLCELL_X32 FILLER_124_888 ();
 FILLCELL_X32 FILLER_124_920 ();
 FILLCELL_X32 FILLER_124_952 ();
 FILLCELL_X32 FILLER_124_984 ();
 FILLCELL_X32 FILLER_124_1016 ();
 FILLCELL_X32 FILLER_124_1048 ();
 FILLCELL_X32 FILLER_124_1080 ();
 FILLCELL_X32 FILLER_124_1112 ();
 FILLCELL_X32 FILLER_124_1144 ();
 FILLCELL_X32 FILLER_124_1176 ();
 FILLCELL_X32 FILLER_124_1208 ();
 FILLCELL_X32 FILLER_124_1240 ();
 FILLCELL_X32 FILLER_124_1272 ();
 FILLCELL_X32 FILLER_124_1304 ();
 FILLCELL_X32 FILLER_124_1336 ();
 FILLCELL_X32 FILLER_124_1368 ();
 FILLCELL_X32 FILLER_124_1400 ();
 FILLCELL_X32 FILLER_124_1432 ();
 FILLCELL_X32 FILLER_124_1464 ();
 FILLCELL_X32 FILLER_124_1496 ();
 FILLCELL_X32 FILLER_124_1528 ();
 FILLCELL_X32 FILLER_124_1560 ();
 FILLCELL_X32 FILLER_124_1592 ();
 FILLCELL_X32 FILLER_124_1624 ();
 FILLCELL_X32 FILLER_124_1656 ();
 FILLCELL_X32 FILLER_124_1688 ();
 FILLCELL_X32 FILLER_124_1720 ();
 FILLCELL_X32 FILLER_124_1752 ();
 FILLCELL_X32 FILLER_124_1784 ();
 FILLCELL_X32 FILLER_124_1816 ();
 FILLCELL_X32 FILLER_124_1848 ();
 FILLCELL_X8 FILLER_124_1880 ();
 FILLCELL_X4 FILLER_124_1888 ();
 FILLCELL_X2 FILLER_124_1892 ();
 FILLCELL_X32 FILLER_124_1895 ();
 FILLCELL_X32 FILLER_124_1927 ();
 FILLCELL_X32 FILLER_124_1959 ();
 FILLCELL_X32 FILLER_124_1991 ();
 FILLCELL_X32 FILLER_124_2023 ();
 FILLCELL_X32 FILLER_124_2055 ();
 FILLCELL_X32 FILLER_124_2087 ();
 FILLCELL_X32 FILLER_124_2119 ();
 FILLCELL_X32 FILLER_124_2151 ();
 FILLCELL_X32 FILLER_124_2183 ();
 FILLCELL_X32 FILLER_124_2215 ();
 FILLCELL_X32 FILLER_124_2247 ();
 FILLCELL_X32 FILLER_124_2279 ();
 FILLCELL_X32 FILLER_124_2311 ();
 FILLCELL_X32 FILLER_124_2343 ();
 FILLCELL_X32 FILLER_124_2375 ();
 FILLCELL_X32 FILLER_124_2407 ();
 FILLCELL_X32 FILLER_124_2439 ();
 FILLCELL_X32 FILLER_124_2471 ();
 FILLCELL_X32 FILLER_124_2503 ();
 FILLCELL_X32 FILLER_124_2535 ();
 FILLCELL_X32 FILLER_124_2567 ();
 FILLCELL_X32 FILLER_124_2599 ();
 FILLCELL_X32 FILLER_124_2631 ();
 FILLCELL_X32 FILLER_124_2663 ();
 FILLCELL_X32 FILLER_124_2695 ();
 FILLCELL_X32 FILLER_124_2727 ();
 FILLCELL_X32 FILLER_124_2759 ();
 FILLCELL_X32 FILLER_124_2791 ();
 FILLCELL_X32 FILLER_124_2823 ();
 FILLCELL_X32 FILLER_124_2855 ();
 FILLCELL_X32 FILLER_124_2887 ();
 FILLCELL_X32 FILLER_124_2919 ();
 FILLCELL_X32 FILLER_124_2951 ();
 FILLCELL_X32 FILLER_124_2983 ();
 FILLCELL_X32 FILLER_124_3015 ();
 FILLCELL_X32 FILLER_124_3047 ();
 FILLCELL_X32 FILLER_124_3079 ();
 FILLCELL_X32 FILLER_124_3111 ();
 FILLCELL_X8 FILLER_124_3143 ();
 FILLCELL_X4 FILLER_124_3151 ();
 FILLCELL_X2 FILLER_124_3155 ();
 FILLCELL_X32 FILLER_124_3158 ();
 FILLCELL_X32 FILLER_124_3190 ();
 FILLCELL_X32 FILLER_124_3222 ();
 FILLCELL_X32 FILLER_124_3254 ();
 FILLCELL_X32 FILLER_124_3286 ();
 FILLCELL_X32 FILLER_124_3318 ();
 FILLCELL_X32 FILLER_124_3350 ();
 FILLCELL_X32 FILLER_124_3382 ();
 FILLCELL_X32 FILLER_124_3414 ();
 FILLCELL_X32 FILLER_124_3446 ();
 FILLCELL_X32 FILLER_124_3478 ();
 FILLCELL_X32 FILLER_124_3510 ();
 FILLCELL_X32 FILLER_124_3542 ();
 FILLCELL_X32 FILLER_124_3574 ();
 FILLCELL_X32 FILLER_124_3606 ();
 FILLCELL_X32 FILLER_124_3638 ();
 FILLCELL_X32 FILLER_124_3670 ();
 FILLCELL_X32 FILLER_124_3702 ();
 FILLCELL_X4 FILLER_124_3734 ();
 FILLCELL_X32 FILLER_125_1 ();
 FILLCELL_X32 FILLER_125_33 ();
 FILLCELL_X32 FILLER_125_65 ();
 FILLCELL_X32 FILLER_125_97 ();
 FILLCELL_X32 FILLER_125_129 ();
 FILLCELL_X32 FILLER_125_161 ();
 FILLCELL_X32 FILLER_125_193 ();
 FILLCELL_X32 FILLER_125_225 ();
 FILLCELL_X32 FILLER_125_257 ();
 FILLCELL_X32 FILLER_125_289 ();
 FILLCELL_X32 FILLER_125_321 ();
 FILLCELL_X32 FILLER_125_353 ();
 FILLCELL_X32 FILLER_125_385 ();
 FILLCELL_X32 FILLER_125_417 ();
 FILLCELL_X32 FILLER_125_449 ();
 FILLCELL_X32 FILLER_125_481 ();
 FILLCELL_X32 FILLER_125_513 ();
 FILLCELL_X32 FILLER_125_545 ();
 FILLCELL_X32 FILLER_125_577 ();
 FILLCELL_X32 FILLER_125_609 ();
 FILLCELL_X32 FILLER_125_641 ();
 FILLCELL_X32 FILLER_125_673 ();
 FILLCELL_X32 FILLER_125_705 ();
 FILLCELL_X32 FILLER_125_737 ();
 FILLCELL_X32 FILLER_125_769 ();
 FILLCELL_X32 FILLER_125_801 ();
 FILLCELL_X32 FILLER_125_833 ();
 FILLCELL_X32 FILLER_125_865 ();
 FILLCELL_X32 FILLER_125_897 ();
 FILLCELL_X32 FILLER_125_929 ();
 FILLCELL_X32 FILLER_125_961 ();
 FILLCELL_X32 FILLER_125_993 ();
 FILLCELL_X32 FILLER_125_1025 ();
 FILLCELL_X32 FILLER_125_1057 ();
 FILLCELL_X32 FILLER_125_1089 ();
 FILLCELL_X32 FILLER_125_1121 ();
 FILLCELL_X32 FILLER_125_1153 ();
 FILLCELL_X32 FILLER_125_1185 ();
 FILLCELL_X32 FILLER_125_1217 ();
 FILLCELL_X8 FILLER_125_1249 ();
 FILLCELL_X4 FILLER_125_1257 ();
 FILLCELL_X2 FILLER_125_1261 ();
 FILLCELL_X32 FILLER_125_1264 ();
 FILLCELL_X32 FILLER_125_1296 ();
 FILLCELL_X32 FILLER_125_1328 ();
 FILLCELL_X32 FILLER_125_1360 ();
 FILLCELL_X32 FILLER_125_1392 ();
 FILLCELL_X32 FILLER_125_1424 ();
 FILLCELL_X32 FILLER_125_1456 ();
 FILLCELL_X32 FILLER_125_1488 ();
 FILLCELL_X32 FILLER_125_1520 ();
 FILLCELL_X32 FILLER_125_1552 ();
 FILLCELL_X32 FILLER_125_1584 ();
 FILLCELL_X32 FILLER_125_1616 ();
 FILLCELL_X32 FILLER_125_1648 ();
 FILLCELL_X32 FILLER_125_1680 ();
 FILLCELL_X32 FILLER_125_1712 ();
 FILLCELL_X32 FILLER_125_1744 ();
 FILLCELL_X32 FILLER_125_1776 ();
 FILLCELL_X32 FILLER_125_1808 ();
 FILLCELL_X32 FILLER_125_1840 ();
 FILLCELL_X32 FILLER_125_1872 ();
 FILLCELL_X32 FILLER_125_1904 ();
 FILLCELL_X32 FILLER_125_1936 ();
 FILLCELL_X32 FILLER_125_1968 ();
 FILLCELL_X32 FILLER_125_2000 ();
 FILLCELL_X32 FILLER_125_2032 ();
 FILLCELL_X32 FILLER_125_2064 ();
 FILLCELL_X32 FILLER_125_2096 ();
 FILLCELL_X32 FILLER_125_2128 ();
 FILLCELL_X32 FILLER_125_2160 ();
 FILLCELL_X32 FILLER_125_2192 ();
 FILLCELL_X32 FILLER_125_2224 ();
 FILLCELL_X32 FILLER_125_2256 ();
 FILLCELL_X32 FILLER_125_2288 ();
 FILLCELL_X32 FILLER_125_2320 ();
 FILLCELL_X32 FILLER_125_2352 ();
 FILLCELL_X32 FILLER_125_2384 ();
 FILLCELL_X32 FILLER_125_2416 ();
 FILLCELL_X32 FILLER_125_2448 ();
 FILLCELL_X32 FILLER_125_2480 ();
 FILLCELL_X8 FILLER_125_2512 ();
 FILLCELL_X4 FILLER_125_2520 ();
 FILLCELL_X2 FILLER_125_2524 ();
 FILLCELL_X32 FILLER_125_2527 ();
 FILLCELL_X32 FILLER_125_2559 ();
 FILLCELL_X32 FILLER_125_2591 ();
 FILLCELL_X32 FILLER_125_2623 ();
 FILLCELL_X32 FILLER_125_2655 ();
 FILLCELL_X32 FILLER_125_2687 ();
 FILLCELL_X32 FILLER_125_2719 ();
 FILLCELL_X32 FILLER_125_2751 ();
 FILLCELL_X32 FILLER_125_2783 ();
 FILLCELL_X32 FILLER_125_2815 ();
 FILLCELL_X32 FILLER_125_2847 ();
 FILLCELL_X32 FILLER_125_2879 ();
 FILLCELL_X32 FILLER_125_2911 ();
 FILLCELL_X32 FILLER_125_2943 ();
 FILLCELL_X32 FILLER_125_2975 ();
 FILLCELL_X32 FILLER_125_3007 ();
 FILLCELL_X32 FILLER_125_3039 ();
 FILLCELL_X32 FILLER_125_3071 ();
 FILLCELL_X32 FILLER_125_3103 ();
 FILLCELL_X32 FILLER_125_3135 ();
 FILLCELL_X32 FILLER_125_3167 ();
 FILLCELL_X32 FILLER_125_3199 ();
 FILLCELL_X32 FILLER_125_3231 ();
 FILLCELL_X32 FILLER_125_3263 ();
 FILLCELL_X32 FILLER_125_3295 ();
 FILLCELL_X32 FILLER_125_3327 ();
 FILLCELL_X32 FILLER_125_3359 ();
 FILLCELL_X32 FILLER_125_3391 ();
 FILLCELL_X32 FILLER_125_3423 ();
 FILLCELL_X32 FILLER_125_3455 ();
 FILLCELL_X32 FILLER_125_3487 ();
 FILLCELL_X32 FILLER_125_3519 ();
 FILLCELL_X32 FILLER_125_3551 ();
 FILLCELL_X32 FILLER_125_3583 ();
 FILLCELL_X32 FILLER_125_3615 ();
 FILLCELL_X32 FILLER_125_3647 ();
 FILLCELL_X32 FILLER_125_3679 ();
 FILLCELL_X16 FILLER_125_3711 ();
 FILLCELL_X8 FILLER_125_3727 ();
 FILLCELL_X2 FILLER_125_3735 ();
 FILLCELL_X1 FILLER_125_3737 ();
 FILLCELL_X32 FILLER_126_1 ();
 FILLCELL_X32 FILLER_126_33 ();
 FILLCELL_X32 FILLER_126_65 ();
 FILLCELL_X32 FILLER_126_97 ();
 FILLCELL_X32 FILLER_126_129 ();
 FILLCELL_X32 FILLER_126_161 ();
 FILLCELL_X32 FILLER_126_193 ();
 FILLCELL_X32 FILLER_126_225 ();
 FILLCELL_X32 FILLER_126_257 ();
 FILLCELL_X32 FILLER_126_289 ();
 FILLCELL_X32 FILLER_126_321 ();
 FILLCELL_X32 FILLER_126_353 ();
 FILLCELL_X32 FILLER_126_385 ();
 FILLCELL_X32 FILLER_126_417 ();
 FILLCELL_X32 FILLER_126_449 ();
 FILLCELL_X32 FILLER_126_481 ();
 FILLCELL_X32 FILLER_126_513 ();
 FILLCELL_X32 FILLER_126_545 ();
 FILLCELL_X32 FILLER_126_577 ();
 FILLCELL_X16 FILLER_126_609 ();
 FILLCELL_X4 FILLER_126_625 ();
 FILLCELL_X2 FILLER_126_629 ();
 FILLCELL_X32 FILLER_126_632 ();
 FILLCELL_X32 FILLER_126_664 ();
 FILLCELL_X32 FILLER_126_696 ();
 FILLCELL_X32 FILLER_126_728 ();
 FILLCELL_X32 FILLER_126_760 ();
 FILLCELL_X32 FILLER_126_792 ();
 FILLCELL_X32 FILLER_126_824 ();
 FILLCELL_X32 FILLER_126_856 ();
 FILLCELL_X32 FILLER_126_888 ();
 FILLCELL_X32 FILLER_126_920 ();
 FILLCELL_X32 FILLER_126_952 ();
 FILLCELL_X32 FILLER_126_984 ();
 FILLCELL_X32 FILLER_126_1016 ();
 FILLCELL_X32 FILLER_126_1048 ();
 FILLCELL_X32 FILLER_126_1080 ();
 FILLCELL_X32 FILLER_126_1112 ();
 FILLCELL_X32 FILLER_126_1144 ();
 FILLCELL_X32 FILLER_126_1176 ();
 FILLCELL_X32 FILLER_126_1208 ();
 FILLCELL_X32 FILLER_126_1240 ();
 FILLCELL_X32 FILLER_126_1272 ();
 FILLCELL_X32 FILLER_126_1304 ();
 FILLCELL_X32 FILLER_126_1336 ();
 FILLCELL_X32 FILLER_126_1368 ();
 FILLCELL_X32 FILLER_126_1400 ();
 FILLCELL_X32 FILLER_126_1432 ();
 FILLCELL_X32 FILLER_126_1464 ();
 FILLCELL_X32 FILLER_126_1496 ();
 FILLCELL_X32 FILLER_126_1528 ();
 FILLCELL_X32 FILLER_126_1560 ();
 FILLCELL_X32 FILLER_126_1592 ();
 FILLCELL_X32 FILLER_126_1624 ();
 FILLCELL_X32 FILLER_126_1656 ();
 FILLCELL_X32 FILLER_126_1688 ();
 FILLCELL_X32 FILLER_126_1720 ();
 FILLCELL_X32 FILLER_126_1752 ();
 FILLCELL_X32 FILLER_126_1784 ();
 FILLCELL_X32 FILLER_126_1816 ();
 FILLCELL_X32 FILLER_126_1848 ();
 FILLCELL_X8 FILLER_126_1880 ();
 FILLCELL_X4 FILLER_126_1888 ();
 FILLCELL_X2 FILLER_126_1892 ();
 FILLCELL_X32 FILLER_126_1895 ();
 FILLCELL_X32 FILLER_126_1927 ();
 FILLCELL_X32 FILLER_126_1959 ();
 FILLCELL_X32 FILLER_126_1991 ();
 FILLCELL_X32 FILLER_126_2023 ();
 FILLCELL_X32 FILLER_126_2055 ();
 FILLCELL_X32 FILLER_126_2087 ();
 FILLCELL_X32 FILLER_126_2119 ();
 FILLCELL_X32 FILLER_126_2151 ();
 FILLCELL_X32 FILLER_126_2183 ();
 FILLCELL_X32 FILLER_126_2215 ();
 FILLCELL_X32 FILLER_126_2247 ();
 FILLCELL_X32 FILLER_126_2279 ();
 FILLCELL_X32 FILLER_126_2311 ();
 FILLCELL_X32 FILLER_126_2343 ();
 FILLCELL_X32 FILLER_126_2375 ();
 FILLCELL_X32 FILLER_126_2407 ();
 FILLCELL_X32 FILLER_126_2439 ();
 FILLCELL_X32 FILLER_126_2471 ();
 FILLCELL_X32 FILLER_126_2503 ();
 FILLCELL_X32 FILLER_126_2535 ();
 FILLCELL_X32 FILLER_126_2567 ();
 FILLCELL_X32 FILLER_126_2599 ();
 FILLCELL_X32 FILLER_126_2631 ();
 FILLCELL_X32 FILLER_126_2663 ();
 FILLCELL_X32 FILLER_126_2695 ();
 FILLCELL_X32 FILLER_126_2727 ();
 FILLCELL_X32 FILLER_126_2759 ();
 FILLCELL_X32 FILLER_126_2791 ();
 FILLCELL_X32 FILLER_126_2823 ();
 FILLCELL_X32 FILLER_126_2855 ();
 FILLCELL_X32 FILLER_126_2887 ();
 FILLCELL_X32 FILLER_126_2919 ();
 FILLCELL_X32 FILLER_126_2951 ();
 FILLCELL_X32 FILLER_126_2983 ();
 FILLCELL_X32 FILLER_126_3015 ();
 FILLCELL_X32 FILLER_126_3047 ();
 FILLCELL_X32 FILLER_126_3079 ();
 FILLCELL_X32 FILLER_126_3111 ();
 FILLCELL_X8 FILLER_126_3143 ();
 FILLCELL_X4 FILLER_126_3151 ();
 FILLCELL_X2 FILLER_126_3155 ();
 FILLCELL_X32 FILLER_126_3158 ();
 FILLCELL_X32 FILLER_126_3190 ();
 FILLCELL_X32 FILLER_126_3222 ();
 FILLCELL_X32 FILLER_126_3254 ();
 FILLCELL_X32 FILLER_126_3286 ();
 FILLCELL_X32 FILLER_126_3318 ();
 FILLCELL_X32 FILLER_126_3350 ();
 FILLCELL_X32 FILLER_126_3382 ();
 FILLCELL_X32 FILLER_126_3414 ();
 FILLCELL_X32 FILLER_126_3446 ();
 FILLCELL_X32 FILLER_126_3478 ();
 FILLCELL_X32 FILLER_126_3510 ();
 FILLCELL_X32 FILLER_126_3542 ();
 FILLCELL_X32 FILLER_126_3574 ();
 FILLCELL_X32 FILLER_126_3606 ();
 FILLCELL_X32 FILLER_126_3638 ();
 FILLCELL_X32 FILLER_126_3670 ();
 FILLCELL_X32 FILLER_126_3702 ();
 FILLCELL_X4 FILLER_126_3734 ();
 FILLCELL_X32 FILLER_127_1 ();
 FILLCELL_X32 FILLER_127_33 ();
 FILLCELL_X32 FILLER_127_65 ();
 FILLCELL_X32 FILLER_127_97 ();
 FILLCELL_X32 FILLER_127_129 ();
 FILLCELL_X32 FILLER_127_161 ();
 FILLCELL_X32 FILLER_127_193 ();
 FILLCELL_X32 FILLER_127_225 ();
 FILLCELL_X32 FILLER_127_257 ();
 FILLCELL_X32 FILLER_127_289 ();
 FILLCELL_X32 FILLER_127_321 ();
 FILLCELL_X32 FILLER_127_353 ();
 FILLCELL_X32 FILLER_127_385 ();
 FILLCELL_X32 FILLER_127_417 ();
 FILLCELL_X32 FILLER_127_449 ();
 FILLCELL_X32 FILLER_127_481 ();
 FILLCELL_X32 FILLER_127_513 ();
 FILLCELL_X32 FILLER_127_545 ();
 FILLCELL_X32 FILLER_127_577 ();
 FILLCELL_X32 FILLER_127_609 ();
 FILLCELL_X32 FILLER_127_641 ();
 FILLCELL_X32 FILLER_127_673 ();
 FILLCELL_X32 FILLER_127_705 ();
 FILLCELL_X32 FILLER_127_737 ();
 FILLCELL_X32 FILLER_127_769 ();
 FILLCELL_X32 FILLER_127_801 ();
 FILLCELL_X32 FILLER_127_833 ();
 FILLCELL_X32 FILLER_127_865 ();
 FILLCELL_X32 FILLER_127_897 ();
 FILLCELL_X32 FILLER_127_929 ();
 FILLCELL_X32 FILLER_127_961 ();
 FILLCELL_X32 FILLER_127_993 ();
 FILLCELL_X32 FILLER_127_1025 ();
 FILLCELL_X32 FILLER_127_1057 ();
 FILLCELL_X32 FILLER_127_1089 ();
 FILLCELL_X32 FILLER_127_1121 ();
 FILLCELL_X32 FILLER_127_1153 ();
 FILLCELL_X32 FILLER_127_1185 ();
 FILLCELL_X32 FILLER_127_1217 ();
 FILLCELL_X8 FILLER_127_1249 ();
 FILLCELL_X4 FILLER_127_1257 ();
 FILLCELL_X2 FILLER_127_1261 ();
 FILLCELL_X32 FILLER_127_1264 ();
 FILLCELL_X32 FILLER_127_1296 ();
 FILLCELL_X32 FILLER_127_1328 ();
 FILLCELL_X32 FILLER_127_1360 ();
 FILLCELL_X32 FILLER_127_1392 ();
 FILLCELL_X32 FILLER_127_1424 ();
 FILLCELL_X32 FILLER_127_1456 ();
 FILLCELL_X32 FILLER_127_1488 ();
 FILLCELL_X32 FILLER_127_1520 ();
 FILLCELL_X32 FILLER_127_1552 ();
 FILLCELL_X32 FILLER_127_1584 ();
 FILLCELL_X32 FILLER_127_1616 ();
 FILLCELL_X32 FILLER_127_1648 ();
 FILLCELL_X32 FILLER_127_1680 ();
 FILLCELL_X32 FILLER_127_1712 ();
 FILLCELL_X32 FILLER_127_1744 ();
 FILLCELL_X32 FILLER_127_1776 ();
 FILLCELL_X32 FILLER_127_1808 ();
 FILLCELL_X32 FILLER_127_1840 ();
 FILLCELL_X32 FILLER_127_1872 ();
 FILLCELL_X32 FILLER_127_1904 ();
 FILLCELL_X32 FILLER_127_1936 ();
 FILLCELL_X32 FILLER_127_1968 ();
 FILLCELL_X32 FILLER_127_2000 ();
 FILLCELL_X32 FILLER_127_2032 ();
 FILLCELL_X32 FILLER_127_2064 ();
 FILLCELL_X32 FILLER_127_2096 ();
 FILLCELL_X32 FILLER_127_2128 ();
 FILLCELL_X32 FILLER_127_2160 ();
 FILLCELL_X32 FILLER_127_2192 ();
 FILLCELL_X32 FILLER_127_2224 ();
 FILLCELL_X32 FILLER_127_2256 ();
 FILLCELL_X32 FILLER_127_2288 ();
 FILLCELL_X32 FILLER_127_2320 ();
 FILLCELL_X32 FILLER_127_2352 ();
 FILLCELL_X32 FILLER_127_2384 ();
 FILLCELL_X32 FILLER_127_2416 ();
 FILLCELL_X32 FILLER_127_2448 ();
 FILLCELL_X32 FILLER_127_2480 ();
 FILLCELL_X8 FILLER_127_2512 ();
 FILLCELL_X4 FILLER_127_2520 ();
 FILLCELL_X2 FILLER_127_2524 ();
 FILLCELL_X32 FILLER_127_2527 ();
 FILLCELL_X32 FILLER_127_2559 ();
 FILLCELL_X32 FILLER_127_2591 ();
 FILLCELL_X32 FILLER_127_2623 ();
 FILLCELL_X32 FILLER_127_2655 ();
 FILLCELL_X32 FILLER_127_2687 ();
 FILLCELL_X32 FILLER_127_2719 ();
 FILLCELL_X32 FILLER_127_2751 ();
 FILLCELL_X32 FILLER_127_2783 ();
 FILLCELL_X32 FILLER_127_2815 ();
 FILLCELL_X32 FILLER_127_2847 ();
 FILLCELL_X32 FILLER_127_2879 ();
 FILLCELL_X32 FILLER_127_2911 ();
 FILLCELL_X32 FILLER_127_2943 ();
 FILLCELL_X32 FILLER_127_2975 ();
 FILLCELL_X32 FILLER_127_3007 ();
 FILLCELL_X32 FILLER_127_3039 ();
 FILLCELL_X32 FILLER_127_3071 ();
 FILLCELL_X32 FILLER_127_3103 ();
 FILLCELL_X32 FILLER_127_3135 ();
 FILLCELL_X32 FILLER_127_3167 ();
 FILLCELL_X32 FILLER_127_3199 ();
 FILLCELL_X32 FILLER_127_3231 ();
 FILLCELL_X32 FILLER_127_3263 ();
 FILLCELL_X32 FILLER_127_3295 ();
 FILLCELL_X32 FILLER_127_3327 ();
 FILLCELL_X32 FILLER_127_3359 ();
 FILLCELL_X32 FILLER_127_3391 ();
 FILLCELL_X32 FILLER_127_3423 ();
 FILLCELL_X32 FILLER_127_3455 ();
 FILLCELL_X32 FILLER_127_3487 ();
 FILLCELL_X32 FILLER_127_3519 ();
 FILLCELL_X32 FILLER_127_3551 ();
 FILLCELL_X32 FILLER_127_3583 ();
 FILLCELL_X32 FILLER_127_3615 ();
 FILLCELL_X32 FILLER_127_3647 ();
 FILLCELL_X32 FILLER_127_3679 ();
 FILLCELL_X16 FILLER_127_3711 ();
 FILLCELL_X8 FILLER_127_3727 ();
 FILLCELL_X2 FILLER_127_3735 ();
 FILLCELL_X1 FILLER_127_3737 ();
 FILLCELL_X32 FILLER_128_1 ();
 FILLCELL_X32 FILLER_128_33 ();
 FILLCELL_X32 FILLER_128_65 ();
 FILLCELL_X32 FILLER_128_97 ();
 FILLCELL_X32 FILLER_128_129 ();
 FILLCELL_X32 FILLER_128_161 ();
 FILLCELL_X32 FILLER_128_193 ();
 FILLCELL_X32 FILLER_128_225 ();
 FILLCELL_X32 FILLER_128_257 ();
 FILLCELL_X32 FILLER_128_289 ();
 FILLCELL_X32 FILLER_128_321 ();
 FILLCELL_X32 FILLER_128_353 ();
 FILLCELL_X32 FILLER_128_385 ();
 FILLCELL_X32 FILLER_128_417 ();
 FILLCELL_X32 FILLER_128_449 ();
 FILLCELL_X32 FILLER_128_481 ();
 FILLCELL_X32 FILLER_128_513 ();
 FILLCELL_X32 FILLER_128_545 ();
 FILLCELL_X32 FILLER_128_577 ();
 FILLCELL_X16 FILLER_128_609 ();
 FILLCELL_X4 FILLER_128_625 ();
 FILLCELL_X2 FILLER_128_629 ();
 FILLCELL_X32 FILLER_128_632 ();
 FILLCELL_X32 FILLER_128_664 ();
 FILLCELL_X32 FILLER_128_696 ();
 FILLCELL_X32 FILLER_128_728 ();
 FILLCELL_X32 FILLER_128_760 ();
 FILLCELL_X32 FILLER_128_792 ();
 FILLCELL_X32 FILLER_128_824 ();
 FILLCELL_X32 FILLER_128_856 ();
 FILLCELL_X32 FILLER_128_888 ();
 FILLCELL_X32 FILLER_128_920 ();
 FILLCELL_X32 FILLER_128_952 ();
 FILLCELL_X32 FILLER_128_984 ();
 FILLCELL_X32 FILLER_128_1016 ();
 FILLCELL_X32 FILLER_128_1048 ();
 FILLCELL_X32 FILLER_128_1080 ();
 FILLCELL_X32 FILLER_128_1112 ();
 FILLCELL_X32 FILLER_128_1144 ();
 FILLCELL_X32 FILLER_128_1176 ();
 FILLCELL_X32 FILLER_128_1208 ();
 FILLCELL_X32 FILLER_128_1240 ();
 FILLCELL_X32 FILLER_128_1272 ();
 FILLCELL_X32 FILLER_128_1304 ();
 FILLCELL_X32 FILLER_128_1336 ();
 FILLCELL_X32 FILLER_128_1368 ();
 FILLCELL_X32 FILLER_128_1400 ();
 FILLCELL_X32 FILLER_128_1432 ();
 FILLCELL_X32 FILLER_128_1464 ();
 FILLCELL_X32 FILLER_128_1496 ();
 FILLCELL_X32 FILLER_128_1528 ();
 FILLCELL_X32 FILLER_128_1560 ();
 FILLCELL_X32 FILLER_128_1592 ();
 FILLCELL_X32 FILLER_128_1624 ();
 FILLCELL_X32 FILLER_128_1656 ();
 FILLCELL_X32 FILLER_128_1688 ();
 FILLCELL_X32 FILLER_128_1720 ();
 FILLCELL_X32 FILLER_128_1752 ();
 FILLCELL_X32 FILLER_128_1784 ();
 FILLCELL_X32 FILLER_128_1816 ();
 FILLCELL_X32 FILLER_128_1848 ();
 FILLCELL_X8 FILLER_128_1880 ();
 FILLCELL_X4 FILLER_128_1888 ();
 FILLCELL_X2 FILLER_128_1892 ();
 FILLCELL_X32 FILLER_128_1895 ();
 FILLCELL_X32 FILLER_128_1927 ();
 FILLCELL_X32 FILLER_128_1959 ();
 FILLCELL_X32 FILLER_128_1991 ();
 FILLCELL_X32 FILLER_128_2023 ();
 FILLCELL_X32 FILLER_128_2055 ();
 FILLCELL_X32 FILLER_128_2087 ();
 FILLCELL_X32 FILLER_128_2119 ();
 FILLCELL_X32 FILLER_128_2151 ();
 FILLCELL_X32 FILLER_128_2183 ();
 FILLCELL_X32 FILLER_128_2215 ();
 FILLCELL_X32 FILLER_128_2247 ();
 FILLCELL_X32 FILLER_128_2279 ();
 FILLCELL_X32 FILLER_128_2311 ();
 FILLCELL_X32 FILLER_128_2343 ();
 FILLCELL_X32 FILLER_128_2375 ();
 FILLCELL_X32 FILLER_128_2407 ();
 FILLCELL_X32 FILLER_128_2439 ();
 FILLCELL_X32 FILLER_128_2471 ();
 FILLCELL_X32 FILLER_128_2503 ();
 FILLCELL_X32 FILLER_128_2535 ();
 FILLCELL_X32 FILLER_128_2567 ();
 FILLCELL_X32 FILLER_128_2599 ();
 FILLCELL_X32 FILLER_128_2631 ();
 FILLCELL_X32 FILLER_128_2663 ();
 FILLCELL_X32 FILLER_128_2695 ();
 FILLCELL_X32 FILLER_128_2727 ();
 FILLCELL_X32 FILLER_128_2759 ();
 FILLCELL_X32 FILLER_128_2791 ();
 FILLCELL_X32 FILLER_128_2823 ();
 FILLCELL_X32 FILLER_128_2855 ();
 FILLCELL_X32 FILLER_128_2887 ();
 FILLCELL_X32 FILLER_128_2919 ();
 FILLCELL_X32 FILLER_128_2951 ();
 FILLCELL_X32 FILLER_128_2983 ();
 FILLCELL_X32 FILLER_128_3015 ();
 FILLCELL_X32 FILLER_128_3047 ();
 FILLCELL_X32 FILLER_128_3079 ();
 FILLCELL_X32 FILLER_128_3111 ();
 FILLCELL_X8 FILLER_128_3143 ();
 FILLCELL_X4 FILLER_128_3151 ();
 FILLCELL_X2 FILLER_128_3155 ();
 FILLCELL_X32 FILLER_128_3158 ();
 FILLCELL_X32 FILLER_128_3190 ();
 FILLCELL_X32 FILLER_128_3222 ();
 FILLCELL_X32 FILLER_128_3254 ();
 FILLCELL_X32 FILLER_128_3286 ();
 FILLCELL_X32 FILLER_128_3318 ();
 FILLCELL_X32 FILLER_128_3350 ();
 FILLCELL_X32 FILLER_128_3382 ();
 FILLCELL_X32 FILLER_128_3414 ();
 FILLCELL_X32 FILLER_128_3446 ();
 FILLCELL_X32 FILLER_128_3478 ();
 FILLCELL_X32 FILLER_128_3510 ();
 FILLCELL_X32 FILLER_128_3542 ();
 FILLCELL_X32 FILLER_128_3574 ();
 FILLCELL_X32 FILLER_128_3606 ();
 FILLCELL_X32 FILLER_128_3638 ();
 FILLCELL_X32 FILLER_128_3670 ();
 FILLCELL_X32 FILLER_128_3702 ();
 FILLCELL_X4 FILLER_128_3734 ();
 FILLCELL_X32 FILLER_129_1 ();
 FILLCELL_X32 FILLER_129_33 ();
 FILLCELL_X32 FILLER_129_65 ();
 FILLCELL_X32 FILLER_129_97 ();
 FILLCELL_X32 FILLER_129_129 ();
 FILLCELL_X32 FILLER_129_161 ();
 FILLCELL_X32 FILLER_129_193 ();
 FILLCELL_X32 FILLER_129_225 ();
 FILLCELL_X32 FILLER_129_257 ();
 FILLCELL_X32 FILLER_129_289 ();
 FILLCELL_X32 FILLER_129_321 ();
 FILLCELL_X32 FILLER_129_353 ();
 FILLCELL_X32 FILLER_129_385 ();
 FILLCELL_X32 FILLER_129_417 ();
 FILLCELL_X32 FILLER_129_449 ();
 FILLCELL_X32 FILLER_129_481 ();
 FILLCELL_X32 FILLER_129_513 ();
 FILLCELL_X32 FILLER_129_545 ();
 FILLCELL_X32 FILLER_129_577 ();
 FILLCELL_X32 FILLER_129_609 ();
 FILLCELL_X32 FILLER_129_641 ();
 FILLCELL_X32 FILLER_129_673 ();
 FILLCELL_X32 FILLER_129_705 ();
 FILLCELL_X32 FILLER_129_737 ();
 FILLCELL_X32 FILLER_129_769 ();
 FILLCELL_X32 FILLER_129_801 ();
 FILLCELL_X32 FILLER_129_833 ();
 FILLCELL_X32 FILLER_129_865 ();
 FILLCELL_X32 FILLER_129_897 ();
 FILLCELL_X32 FILLER_129_929 ();
 FILLCELL_X32 FILLER_129_961 ();
 FILLCELL_X32 FILLER_129_993 ();
 FILLCELL_X32 FILLER_129_1025 ();
 FILLCELL_X32 FILLER_129_1057 ();
 FILLCELL_X32 FILLER_129_1089 ();
 FILLCELL_X32 FILLER_129_1121 ();
 FILLCELL_X32 FILLER_129_1153 ();
 FILLCELL_X32 FILLER_129_1185 ();
 FILLCELL_X32 FILLER_129_1217 ();
 FILLCELL_X8 FILLER_129_1249 ();
 FILLCELL_X4 FILLER_129_1257 ();
 FILLCELL_X2 FILLER_129_1261 ();
 FILLCELL_X32 FILLER_129_1264 ();
 FILLCELL_X32 FILLER_129_1296 ();
 FILLCELL_X32 FILLER_129_1328 ();
 FILLCELL_X32 FILLER_129_1360 ();
 FILLCELL_X32 FILLER_129_1392 ();
 FILLCELL_X32 FILLER_129_1424 ();
 FILLCELL_X32 FILLER_129_1456 ();
 FILLCELL_X32 FILLER_129_1488 ();
 FILLCELL_X32 FILLER_129_1520 ();
 FILLCELL_X32 FILLER_129_1552 ();
 FILLCELL_X32 FILLER_129_1584 ();
 FILLCELL_X32 FILLER_129_1616 ();
 FILLCELL_X32 FILLER_129_1648 ();
 FILLCELL_X32 FILLER_129_1680 ();
 FILLCELL_X32 FILLER_129_1712 ();
 FILLCELL_X32 FILLER_129_1744 ();
 FILLCELL_X32 FILLER_129_1776 ();
 FILLCELL_X32 FILLER_129_1808 ();
 FILLCELL_X32 FILLER_129_1840 ();
 FILLCELL_X32 FILLER_129_1872 ();
 FILLCELL_X32 FILLER_129_1904 ();
 FILLCELL_X32 FILLER_129_1936 ();
 FILLCELL_X32 FILLER_129_1968 ();
 FILLCELL_X32 FILLER_129_2000 ();
 FILLCELL_X32 FILLER_129_2032 ();
 FILLCELL_X32 FILLER_129_2064 ();
 FILLCELL_X32 FILLER_129_2096 ();
 FILLCELL_X32 FILLER_129_2128 ();
 FILLCELL_X32 FILLER_129_2160 ();
 FILLCELL_X32 FILLER_129_2192 ();
 FILLCELL_X32 FILLER_129_2224 ();
 FILLCELL_X32 FILLER_129_2256 ();
 FILLCELL_X32 FILLER_129_2288 ();
 FILLCELL_X32 FILLER_129_2320 ();
 FILLCELL_X32 FILLER_129_2352 ();
 FILLCELL_X32 FILLER_129_2384 ();
 FILLCELL_X32 FILLER_129_2416 ();
 FILLCELL_X32 FILLER_129_2448 ();
 FILLCELL_X32 FILLER_129_2480 ();
 FILLCELL_X8 FILLER_129_2512 ();
 FILLCELL_X4 FILLER_129_2520 ();
 FILLCELL_X2 FILLER_129_2524 ();
 FILLCELL_X32 FILLER_129_2527 ();
 FILLCELL_X32 FILLER_129_2559 ();
 FILLCELL_X32 FILLER_129_2591 ();
 FILLCELL_X32 FILLER_129_2623 ();
 FILLCELL_X32 FILLER_129_2655 ();
 FILLCELL_X32 FILLER_129_2687 ();
 FILLCELL_X32 FILLER_129_2719 ();
 FILLCELL_X32 FILLER_129_2751 ();
 FILLCELL_X32 FILLER_129_2783 ();
 FILLCELL_X32 FILLER_129_2815 ();
 FILLCELL_X32 FILLER_129_2847 ();
 FILLCELL_X32 FILLER_129_2879 ();
 FILLCELL_X32 FILLER_129_2911 ();
 FILLCELL_X32 FILLER_129_2943 ();
 FILLCELL_X32 FILLER_129_2975 ();
 FILLCELL_X32 FILLER_129_3007 ();
 FILLCELL_X32 FILLER_129_3039 ();
 FILLCELL_X32 FILLER_129_3071 ();
 FILLCELL_X32 FILLER_129_3103 ();
 FILLCELL_X32 FILLER_129_3135 ();
 FILLCELL_X32 FILLER_129_3167 ();
 FILLCELL_X32 FILLER_129_3199 ();
 FILLCELL_X32 FILLER_129_3231 ();
 FILLCELL_X32 FILLER_129_3263 ();
 FILLCELL_X32 FILLER_129_3295 ();
 FILLCELL_X32 FILLER_129_3327 ();
 FILLCELL_X32 FILLER_129_3359 ();
 FILLCELL_X32 FILLER_129_3391 ();
 FILLCELL_X32 FILLER_129_3423 ();
 FILLCELL_X32 FILLER_129_3455 ();
 FILLCELL_X32 FILLER_129_3487 ();
 FILLCELL_X32 FILLER_129_3519 ();
 FILLCELL_X32 FILLER_129_3551 ();
 FILLCELL_X32 FILLER_129_3583 ();
 FILLCELL_X32 FILLER_129_3615 ();
 FILLCELL_X32 FILLER_129_3647 ();
 FILLCELL_X32 FILLER_129_3679 ();
 FILLCELL_X16 FILLER_129_3711 ();
 FILLCELL_X8 FILLER_129_3727 ();
 FILLCELL_X2 FILLER_129_3735 ();
 FILLCELL_X1 FILLER_129_3737 ();
 FILLCELL_X32 FILLER_130_1 ();
 FILLCELL_X32 FILLER_130_33 ();
 FILLCELL_X32 FILLER_130_65 ();
 FILLCELL_X32 FILLER_130_97 ();
 FILLCELL_X32 FILLER_130_129 ();
 FILLCELL_X32 FILLER_130_161 ();
 FILLCELL_X32 FILLER_130_193 ();
 FILLCELL_X32 FILLER_130_225 ();
 FILLCELL_X32 FILLER_130_257 ();
 FILLCELL_X32 FILLER_130_289 ();
 FILLCELL_X32 FILLER_130_321 ();
 FILLCELL_X32 FILLER_130_353 ();
 FILLCELL_X32 FILLER_130_385 ();
 FILLCELL_X32 FILLER_130_417 ();
 FILLCELL_X32 FILLER_130_449 ();
 FILLCELL_X32 FILLER_130_481 ();
 FILLCELL_X32 FILLER_130_513 ();
 FILLCELL_X32 FILLER_130_545 ();
 FILLCELL_X32 FILLER_130_577 ();
 FILLCELL_X16 FILLER_130_609 ();
 FILLCELL_X4 FILLER_130_625 ();
 FILLCELL_X2 FILLER_130_629 ();
 FILLCELL_X32 FILLER_130_632 ();
 FILLCELL_X32 FILLER_130_664 ();
 FILLCELL_X32 FILLER_130_696 ();
 FILLCELL_X32 FILLER_130_728 ();
 FILLCELL_X32 FILLER_130_760 ();
 FILLCELL_X32 FILLER_130_792 ();
 FILLCELL_X32 FILLER_130_824 ();
 FILLCELL_X32 FILLER_130_856 ();
 FILLCELL_X32 FILLER_130_888 ();
 FILLCELL_X32 FILLER_130_920 ();
 FILLCELL_X32 FILLER_130_952 ();
 FILLCELL_X32 FILLER_130_984 ();
 FILLCELL_X32 FILLER_130_1016 ();
 FILLCELL_X32 FILLER_130_1048 ();
 FILLCELL_X32 FILLER_130_1080 ();
 FILLCELL_X32 FILLER_130_1112 ();
 FILLCELL_X32 FILLER_130_1144 ();
 FILLCELL_X32 FILLER_130_1176 ();
 FILLCELL_X32 FILLER_130_1208 ();
 FILLCELL_X32 FILLER_130_1240 ();
 FILLCELL_X32 FILLER_130_1272 ();
 FILLCELL_X32 FILLER_130_1304 ();
 FILLCELL_X32 FILLER_130_1336 ();
 FILLCELL_X32 FILLER_130_1368 ();
 FILLCELL_X32 FILLER_130_1400 ();
 FILLCELL_X32 FILLER_130_1432 ();
 FILLCELL_X32 FILLER_130_1464 ();
 FILLCELL_X32 FILLER_130_1496 ();
 FILLCELL_X32 FILLER_130_1528 ();
 FILLCELL_X32 FILLER_130_1560 ();
 FILLCELL_X32 FILLER_130_1592 ();
 FILLCELL_X32 FILLER_130_1624 ();
 FILLCELL_X32 FILLER_130_1656 ();
 FILLCELL_X32 FILLER_130_1688 ();
 FILLCELL_X32 FILLER_130_1720 ();
 FILLCELL_X32 FILLER_130_1752 ();
 FILLCELL_X32 FILLER_130_1784 ();
 FILLCELL_X32 FILLER_130_1816 ();
 FILLCELL_X32 FILLER_130_1848 ();
 FILLCELL_X8 FILLER_130_1880 ();
 FILLCELL_X4 FILLER_130_1888 ();
 FILLCELL_X2 FILLER_130_1892 ();
 FILLCELL_X32 FILLER_130_1895 ();
 FILLCELL_X32 FILLER_130_1927 ();
 FILLCELL_X32 FILLER_130_1959 ();
 FILLCELL_X32 FILLER_130_1991 ();
 FILLCELL_X32 FILLER_130_2023 ();
 FILLCELL_X32 FILLER_130_2055 ();
 FILLCELL_X32 FILLER_130_2087 ();
 FILLCELL_X32 FILLER_130_2119 ();
 FILLCELL_X32 FILLER_130_2151 ();
 FILLCELL_X32 FILLER_130_2183 ();
 FILLCELL_X32 FILLER_130_2215 ();
 FILLCELL_X32 FILLER_130_2247 ();
 FILLCELL_X32 FILLER_130_2279 ();
 FILLCELL_X32 FILLER_130_2311 ();
 FILLCELL_X32 FILLER_130_2343 ();
 FILLCELL_X32 FILLER_130_2375 ();
 FILLCELL_X32 FILLER_130_2407 ();
 FILLCELL_X32 FILLER_130_2439 ();
 FILLCELL_X32 FILLER_130_2471 ();
 FILLCELL_X32 FILLER_130_2503 ();
 FILLCELL_X32 FILLER_130_2535 ();
 FILLCELL_X32 FILLER_130_2567 ();
 FILLCELL_X32 FILLER_130_2599 ();
 FILLCELL_X32 FILLER_130_2631 ();
 FILLCELL_X32 FILLER_130_2663 ();
 FILLCELL_X32 FILLER_130_2695 ();
 FILLCELL_X32 FILLER_130_2727 ();
 FILLCELL_X32 FILLER_130_2759 ();
 FILLCELL_X32 FILLER_130_2791 ();
 FILLCELL_X32 FILLER_130_2823 ();
 FILLCELL_X32 FILLER_130_2855 ();
 FILLCELL_X32 FILLER_130_2887 ();
 FILLCELL_X32 FILLER_130_2919 ();
 FILLCELL_X32 FILLER_130_2951 ();
 FILLCELL_X32 FILLER_130_2983 ();
 FILLCELL_X32 FILLER_130_3015 ();
 FILLCELL_X32 FILLER_130_3047 ();
 FILLCELL_X32 FILLER_130_3079 ();
 FILLCELL_X32 FILLER_130_3111 ();
 FILLCELL_X8 FILLER_130_3143 ();
 FILLCELL_X4 FILLER_130_3151 ();
 FILLCELL_X2 FILLER_130_3155 ();
 FILLCELL_X32 FILLER_130_3158 ();
 FILLCELL_X32 FILLER_130_3190 ();
 FILLCELL_X32 FILLER_130_3222 ();
 FILLCELL_X32 FILLER_130_3254 ();
 FILLCELL_X32 FILLER_130_3286 ();
 FILLCELL_X32 FILLER_130_3318 ();
 FILLCELL_X32 FILLER_130_3350 ();
 FILLCELL_X32 FILLER_130_3382 ();
 FILLCELL_X32 FILLER_130_3414 ();
 FILLCELL_X32 FILLER_130_3446 ();
 FILLCELL_X32 FILLER_130_3478 ();
 FILLCELL_X32 FILLER_130_3510 ();
 FILLCELL_X32 FILLER_130_3542 ();
 FILLCELL_X32 FILLER_130_3574 ();
 FILLCELL_X32 FILLER_130_3606 ();
 FILLCELL_X32 FILLER_130_3638 ();
 FILLCELL_X32 FILLER_130_3670 ();
 FILLCELL_X32 FILLER_130_3702 ();
 FILLCELL_X4 FILLER_130_3734 ();
 FILLCELL_X32 FILLER_131_1 ();
 FILLCELL_X32 FILLER_131_33 ();
 FILLCELL_X32 FILLER_131_65 ();
 FILLCELL_X32 FILLER_131_97 ();
 FILLCELL_X32 FILLER_131_129 ();
 FILLCELL_X32 FILLER_131_161 ();
 FILLCELL_X32 FILLER_131_193 ();
 FILLCELL_X32 FILLER_131_225 ();
 FILLCELL_X32 FILLER_131_257 ();
 FILLCELL_X32 FILLER_131_289 ();
 FILLCELL_X32 FILLER_131_321 ();
 FILLCELL_X32 FILLER_131_353 ();
 FILLCELL_X32 FILLER_131_385 ();
 FILLCELL_X32 FILLER_131_417 ();
 FILLCELL_X32 FILLER_131_449 ();
 FILLCELL_X32 FILLER_131_481 ();
 FILLCELL_X32 FILLER_131_513 ();
 FILLCELL_X32 FILLER_131_545 ();
 FILLCELL_X32 FILLER_131_577 ();
 FILLCELL_X32 FILLER_131_609 ();
 FILLCELL_X32 FILLER_131_641 ();
 FILLCELL_X32 FILLER_131_673 ();
 FILLCELL_X32 FILLER_131_705 ();
 FILLCELL_X32 FILLER_131_737 ();
 FILLCELL_X32 FILLER_131_769 ();
 FILLCELL_X32 FILLER_131_801 ();
 FILLCELL_X32 FILLER_131_833 ();
 FILLCELL_X32 FILLER_131_865 ();
 FILLCELL_X32 FILLER_131_897 ();
 FILLCELL_X32 FILLER_131_929 ();
 FILLCELL_X32 FILLER_131_961 ();
 FILLCELL_X32 FILLER_131_993 ();
 FILLCELL_X32 FILLER_131_1025 ();
 FILLCELL_X32 FILLER_131_1057 ();
 FILLCELL_X32 FILLER_131_1089 ();
 FILLCELL_X32 FILLER_131_1121 ();
 FILLCELL_X32 FILLER_131_1153 ();
 FILLCELL_X32 FILLER_131_1185 ();
 FILLCELL_X32 FILLER_131_1217 ();
 FILLCELL_X8 FILLER_131_1249 ();
 FILLCELL_X4 FILLER_131_1257 ();
 FILLCELL_X2 FILLER_131_1261 ();
 FILLCELL_X32 FILLER_131_1264 ();
 FILLCELL_X32 FILLER_131_1296 ();
 FILLCELL_X32 FILLER_131_1328 ();
 FILLCELL_X32 FILLER_131_1360 ();
 FILLCELL_X32 FILLER_131_1392 ();
 FILLCELL_X32 FILLER_131_1424 ();
 FILLCELL_X32 FILLER_131_1456 ();
 FILLCELL_X32 FILLER_131_1488 ();
 FILLCELL_X32 FILLER_131_1520 ();
 FILLCELL_X32 FILLER_131_1552 ();
 FILLCELL_X32 FILLER_131_1584 ();
 FILLCELL_X32 FILLER_131_1616 ();
 FILLCELL_X32 FILLER_131_1648 ();
 FILLCELL_X32 FILLER_131_1680 ();
 FILLCELL_X32 FILLER_131_1712 ();
 FILLCELL_X32 FILLER_131_1744 ();
 FILLCELL_X32 FILLER_131_1776 ();
 FILLCELL_X32 FILLER_131_1808 ();
 FILLCELL_X32 FILLER_131_1840 ();
 FILLCELL_X32 FILLER_131_1872 ();
 FILLCELL_X32 FILLER_131_1904 ();
 FILLCELL_X32 FILLER_131_1936 ();
 FILLCELL_X32 FILLER_131_1968 ();
 FILLCELL_X32 FILLER_131_2000 ();
 FILLCELL_X32 FILLER_131_2032 ();
 FILLCELL_X32 FILLER_131_2064 ();
 FILLCELL_X32 FILLER_131_2096 ();
 FILLCELL_X32 FILLER_131_2128 ();
 FILLCELL_X32 FILLER_131_2160 ();
 FILLCELL_X32 FILLER_131_2192 ();
 FILLCELL_X32 FILLER_131_2224 ();
 FILLCELL_X32 FILLER_131_2256 ();
 FILLCELL_X32 FILLER_131_2288 ();
 FILLCELL_X32 FILLER_131_2320 ();
 FILLCELL_X32 FILLER_131_2352 ();
 FILLCELL_X32 FILLER_131_2384 ();
 FILLCELL_X32 FILLER_131_2416 ();
 FILLCELL_X32 FILLER_131_2448 ();
 FILLCELL_X32 FILLER_131_2480 ();
 FILLCELL_X8 FILLER_131_2512 ();
 FILLCELL_X4 FILLER_131_2520 ();
 FILLCELL_X2 FILLER_131_2524 ();
 FILLCELL_X32 FILLER_131_2527 ();
 FILLCELL_X32 FILLER_131_2559 ();
 FILLCELL_X32 FILLER_131_2591 ();
 FILLCELL_X32 FILLER_131_2623 ();
 FILLCELL_X32 FILLER_131_2655 ();
 FILLCELL_X32 FILLER_131_2687 ();
 FILLCELL_X32 FILLER_131_2719 ();
 FILLCELL_X32 FILLER_131_2751 ();
 FILLCELL_X32 FILLER_131_2783 ();
 FILLCELL_X32 FILLER_131_2815 ();
 FILLCELL_X32 FILLER_131_2847 ();
 FILLCELL_X32 FILLER_131_2879 ();
 FILLCELL_X32 FILLER_131_2911 ();
 FILLCELL_X32 FILLER_131_2943 ();
 FILLCELL_X32 FILLER_131_2975 ();
 FILLCELL_X32 FILLER_131_3007 ();
 FILLCELL_X32 FILLER_131_3039 ();
 FILLCELL_X32 FILLER_131_3071 ();
 FILLCELL_X32 FILLER_131_3103 ();
 FILLCELL_X32 FILLER_131_3135 ();
 FILLCELL_X32 FILLER_131_3167 ();
 FILLCELL_X32 FILLER_131_3199 ();
 FILLCELL_X32 FILLER_131_3231 ();
 FILLCELL_X32 FILLER_131_3263 ();
 FILLCELL_X32 FILLER_131_3295 ();
 FILLCELL_X32 FILLER_131_3327 ();
 FILLCELL_X32 FILLER_131_3359 ();
 FILLCELL_X32 FILLER_131_3391 ();
 FILLCELL_X32 FILLER_131_3423 ();
 FILLCELL_X32 FILLER_131_3455 ();
 FILLCELL_X32 FILLER_131_3487 ();
 FILLCELL_X32 FILLER_131_3519 ();
 FILLCELL_X32 FILLER_131_3551 ();
 FILLCELL_X32 FILLER_131_3583 ();
 FILLCELL_X32 FILLER_131_3615 ();
 FILLCELL_X32 FILLER_131_3647 ();
 FILLCELL_X32 FILLER_131_3679 ();
 FILLCELL_X16 FILLER_131_3711 ();
 FILLCELL_X8 FILLER_131_3727 ();
 FILLCELL_X2 FILLER_131_3735 ();
 FILLCELL_X1 FILLER_131_3737 ();
 FILLCELL_X32 FILLER_132_1 ();
 FILLCELL_X32 FILLER_132_33 ();
 FILLCELL_X32 FILLER_132_65 ();
 FILLCELL_X32 FILLER_132_97 ();
 FILLCELL_X32 FILLER_132_129 ();
 FILLCELL_X32 FILLER_132_161 ();
 FILLCELL_X32 FILLER_132_193 ();
 FILLCELL_X32 FILLER_132_225 ();
 FILLCELL_X32 FILLER_132_257 ();
 FILLCELL_X32 FILLER_132_289 ();
 FILLCELL_X32 FILLER_132_321 ();
 FILLCELL_X32 FILLER_132_353 ();
 FILLCELL_X32 FILLER_132_385 ();
 FILLCELL_X32 FILLER_132_417 ();
 FILLCELL_X32 FILLER_132_449 ();
 FILLCELL_X32 FILLER_132_481 ();
 FILLCELL_X32 FILLER_132_513 ();
 FILLCELL_X32 FILLER_132_545 ();
 FILLCELL_X32 FILLER_132_577 ();
 FILLCELL_X16 FILLER_132_609 ();
 FILLCELL_X4 FILLER_132_625 ();
 FILLCELL_X2 FILLER_132_629 ();
 FILLCELL_X32 FILLER_132_632 ();
 FILLCELL_X32 FILLER_132_664 ();
 FILLCELL_X32 FILLER_132_696 ();
 FILLCELL_X32 FILLER_132_728 ();
 FILLCELL_X32 FILLER_132_760 ();
 FILLCELL_X32 FILLER_132_792 ();
 FILLCELL_X32 FILLER_132_824 ();
 FILLCELL_X32 FILLER_132_856 ();
 FILLCELL_X32 FILLER_132_888 ();
 FILLCELL_X32 FILLER_132_920 ();
 FILLCELL_X32 FILLER_132_952 ();
 FILLCELL_X32 FILLER_132_984 ();
 FILLCELL_X32 FILLER_132_1016 ();
 FILLCELL_X32 FILLER_132_1048 ();
 FILLCELL_X32 FILLER_132_1080 ();
 FILLCELL_X32 FILLER_132_1112 ();
 FILLCELL_X32 FILLER_132_1144 ();
 FILLCELL_X32 FILLER_132_1176 ();
 FILLCELL_X32 FILLER_132_1208 ();
 FILLCELL_X32 FILLER_132_1240 ();
 FILLCELL_X32 FILLER_132_1272 ();
 FILLCELL_X32 FILLER_132_1304 ();
 FILLCELL_X32 FILLER_132_1336 ();
 FILLCELL_X32 FILLER_132_1368 ();
 FILLCELL_X32 FILLER_132_1400 ();
 FILLCELL_X32 FILLER_132_1432 ();
 FILLCELL_X32 FILLER_132_1464 ();
 FILLCELL_X32 FILLER_132_1496 ();
 FILLCELL_X32 FILLER_132_1528 ();
 FILLCELL_X32 FILLER_132_1560 ();
 FILLCELL_X32 FILLER_132_1592 ();
 FILLCELL_X32 FILLER_132_1624 ();
 FILLCELL_X32 FILLER_132_1656 ();
 FILLCELL_X32 FILLER_132_1688 ();
 FILLCELL_X32 FILLER_132_1720 ();
 FILLCELL_X32 FILLER_132_1752 ();
 FILLCELL_X32 FILLER_132_1784 ();
 FILLCELL_X32 FILLER_132_1816 ();
 FILLCELL_X32 FILLER_132_1848 ();
 FILLCELL_X8 FILLER_132_1880 ();
 FILLCELL_X4 FILLER_132_1888 ();
 FILLCELL_X2 FILLER_132_1892 ();
 FILLCELL_X32 FILLER_132_1895 ();
 FILLCELL_X32 FILLER_132_1927 ();
 FILLCELL_X32 FILLER_132_1959 ();
 FILLCELL_X32 FILLER_132_1991 ();
 FILLCELL_X32 FILLER_132_2023 ();
 FILLCELL_X32 FILLER_132_2055 ();
 FILLCELL_X32 FILLER_132_2087 ();
 FILLCELL_X32 FILLER_132_2119 ();
 FILLCELL_X32 FILLER_132_2151 ();
 FILLCELL_X32 FILLER_132_2183 ();
 FILLCELL_X32 FILLER_132_2215 ();
 FILLCELL_X32 FILLER_132_2247 ();
 FILLCELL_X32 FILLER_132_2279 ();
 FILLCELL_X32 FILLER_132_2311 ();
 FILLCELL_X32 FILLER_132_2343 ();
 FILLCELL_X32 FILLER_132_2375 ();
 FILLCELL_X32 FILLER_132_2407 ();
 FILLCELL_X32 FILLER_132_2439 ();
 FILLCELL_X32 FILLER_132_2471 ();
 FILLCELL_X32 FILLER_132_2503 ();
 FILLCELL_X32 FILLER_132_2535 ();
 FILLCELL_X32 FILLER_132_2567 ();
 FILLCELL_X32 FILLER_132_2599 ();
 FILLCELL_X32 FILLER_132_2631 ();
 FILLCELL_X32 FILLER_132_2663 ();
 FILLCELL_X32 FILLER_132_2695 ();
 FILLCELL_X32 FILLER_132_2727 ();
 FILLCELL_X32 FILLER_132_2759 ();
 FILLCELL_X32 FILLER_132_2791 ();
 FILLCELL_X32 FILLER_132_2823 ();
 FILLCELL_X32 FILLER_132_2855 ();
 FILLCELL_X32 FILLER_132_2887 ();
 FILLCELL_X32 FILLER_132_2919 ();
 FILLCELL_X32 FILLER_132_2951 ();
 FILLCELL_X32 FILLER_132_2983 ();
 FILLCELL_X32 FILLER_132_3015 ();
 FILLCELL_X32 FILLER_132_3047 ();
 FILLCELL_X32 FILLER_132_3079 ();
 FILLCELL_X32 FILLER_132_3111 ();
 FILLCELL_X8 FILLER_132_3143 ();
 FILLCELL_X4 FILLER_132_3151 ();
 FILLCELL_X2 FILLER_132_3155 ();
 FILLCELL_X32 FILLER_132_3158 ();
 FILLCELL_X32 FILLER_132_3190 ();
 FILLCELL_X32 FILLER_132_3222 ();
 FILLCELL_X32 FILLER_132_3254 ();
 FILLCELL_X32 FILLER_132_3286 ();
 FILLCELL_X32 FILLER_132_3318 ();
 FILLCELL_X32 FILLER_132_3350 ();
 FILLCELL_X32 FILLER_132_3382 ();
 FILLCELL_X32 FILLER_132_3414 ();
 FILLCELL_X32 FILLER_132_3446 ();
 FILLCELL_X32 FILLER_132_3478 ();
 FILLCELL_X32 FILLER_132_3510 ();
 FILLCELL_X32 FILLER_132_3542 ();
 FILLCELL_X32 FILLER_132_3574 ();
 FILLCELL_X32 FILLER_132_3606 ();
 FILLCELL_X32 FILLER_132_3638 ();
 FILLCELL_X32 FILLER_132_3670 ();
 FILLCELL_X32 FILLER_132_3702 ();
 FILLCELL_X4 FILLER_132_3734 ();
 FILLCELL_X32 FILLER_133_1 ();
 FILLCELL_X32 FILLER_133_33 ();
 FILLCELL_X32 FILLER_133_65 ();
 FILLCELL_X32 FILLER_133_97 ();
 FILLCELL_X32 FILLER_133_129 ();
 FILLCELL_X32 FILLER_133_161 ();
 FILLCELL_X32 FILLER_133_193 ();
 FILLCELL_X32 FILLER_133_225 ();
 FILLCELL_X32 FILLER_133_257 ();
 FILLCELL_X32 FILLER_133_289 ();
 FILLCELL_X32 FILLER_133_321 ();
 FILLCELL_X32 FILLER_133_353 ();
 FILLCELL_X32 FILLER_133_385 ();
 FILLCELL_X32 FILLER_133_417 ();
 FILLCELL_X32 FILLER_133_449 ();
 FILLCELL_X32 FILLER_133_481 ();
 FILLCELL_X32 FILLER_133_513 ();
 FILLCELL_X32 FILLER_133_545 ();
 FILLCELL_X32 FILLER_133_577 ();
 FILLCELL_X32 FILLER_133_609 ();
 FILLCELL_X32 FILLER_133_641 ();
 FILLCELL_X32 FILLER_133_673 ();
 FILLCELL_X32 FILLER_133_705 ();
 FILLCELL_X32 FILLER_133_737 ();
 FILLCELL_X32 FILLER_133_769 ();
 FILLCELL_X32 FILLER_133_801 ();
 FILLCELL_X32 FILLER_133_833 ();
 FILLCELL_X32 FILLER_133_865 ();
 FILLCELL_X32 FILLER_133_897 ();
 FILLCELL_X32 FILLER_133_929 ();
 FILLCELL_X32 FILLER_133_961 ();
 FILLCELL_X32 FILLER_133_993 ();
 FILLCELL_X32 FILLER_133_1025 ();
 FILLCELL_X32 FILLER_133_1057 ();
 FILLCELL_X32 FILLER_133_1089 ();
 FILLCELL_X32 FILLER_133_1121 ();
 FILLCELL_X32 FILLER_133_1153 ();
 FILLCELL_X32 FILLER_133_1185 ();
 FILLCELL_X32 FILLER_133_1217 ();
 FILLCELL_X8 FILLER_133_1249 ();
 FILLCELL_X4 FILLER_133_1257 ();
 FILLCELL_X2 FILLER_133_1261 ();
 FILLCELL_X32 FILLER_133_1264 ();
 FILLCELL_X32 FILLER_133_1296 ();
 FILLCELL_X32 FILLER_133_1328 ();
 FILLCELL_X32 FILLER_133_1360 ();
 FILLCELL_X32 FILLER_133_1392 ();
 FILLCELL_X32 FILLER_133_1424 ();
 FILLCELL_X32 FILLER_133_1456 ();
 FILLCELL_X32 FILLER_133_1488 ();
 FILLCELL_X32 FILLER_133_1520 ();
 FILLCELL_X32 FILLER_133_1552 ();
 FILLCELL_X32 FILLER_133_1584 ();
 FILLCELL_X32 FILLER_133_1616 ();
 FILLCELL_X32 FILLER_133_1648 ();
 FILLCELL_X32 FILLER_133_1680 ();
 FILLCELL_X32 FILLER_133_1712 ();
 FILLCELL_X32 FILLER_133_1744 ();
 FILLCELL_X32 FILLER_133_1776 ();
 FILLCELL_X32 FILLER_133_1808 ();
 FILLCELL_X32 FILLER_133_1840 ();
 FILLCELL_X32 FILLER_133_1872 ();
 FILLCELL_X32 FILLER_133_1904 ();
 FILLCELL_X32 FILLER_133_1936 ();
 FILLCELL_X32 FILLER_133_1968 ();
 FILLCELL_X32 FILLER_133_2000 ();
 FILLCELL_X32 FILLER_133_2032 ();
 FILLCELL_X32 FILLER_133_2064 ();
 FILLCELL_X32 FILLER_133_2096 ();
 FILLCELL_X32 FILLER_133_2128 ();
 FILLCELL_X32 FILLER_133_2160 ();
 FILLCELL_X32 FILLER_133_2192 ();
 FILLCELL_X32 FILLER_133_2224 ();
 FILLCELL_X32 FILLER_133_2256 ();
 FILLCELL_X32 FILLER_133_2288 ();
 FILLCELL_X32 FILLER_133_2320 ();
 FILLCELL_X32 FILLER_133_2352 ();
 FILLCELL_X32 FILLER_133_2384 ();
 FILLCELL_X32 FILLER_133_2416 ();
 FILLCELL_X32 FILLER_133_2448 ();
 FILLCELL_X32 FILLER_133_2480 ();
 FILLCELL_X8 FILLER_133_2512 ();
 FILLCELL_X4 FILLER_133_2520 ();
 FILLCELL_X2 FILLER_133_2524 ();
 FILLCELL_X32 FILLER_133_2527 ();
 FILLCELL_X32 FILLER_133_2559 ();
 FILLCELL_X32 FILLER_133_2591 ();
 FILLCELL_X32 FILLER_133_2623 ();
 FILLCELL_X32 FILLER_133_2655 ();
 FILLCELL_X32 FILLER_133_2687 ();
 FILLCELL_X32 FILLER_133_2719 ();
 FILLCELL_X32 FILLER_133_2751 ();
 FILLCELL_X32 FILLER_133_2783 ();
 FILLCELL_X32 FILLER_133_2815 ();
 FILLCELL_X32 FILLER_133_2847 ();
 FILLCELL_X32 FILLER_133_2879 ();
 FILLCELL_X32 FILLER_133_2911 ();
 FILLCELL_X32 FILLER_133_2943 ();
 FILLCELL_X32 FILLER_133_2975 ();
 FILLCELL_X32 FILLER_133_3007 ();
 FILLCELL_X32 FILLER_133_3039 ();
 FILLCELL_X32 FILLER_133_3071 ();
 FILLCELL_X32 FILLER_133_3103 ();
 FILLCELL_X32 FILLER_133_3135 ();
 FILLCELL_X32 FILLER_133_3167 ();
 FILLCELL_X32 FILLER_133_3199 ();
 FILLCELL_X32 FILLER_133_3231 ();
 FILLCELL_X32 FILLER_133_3263 ();
 FILLCELL_X32 FILLER_133_3295 ();
 FILLCELL_X32 FILLER_133_3327 ();
 FILLCELL_X32 FILLER_133_3359 ();
 FILLCELL_X32 FILLER_133_3391 ();
 FILLCELL_X32 FILLER_133_3423 ();
 FILLCELL_X32 FILLER_133_3455 ();
 FILLCELL_X32 FILLER_133_3487 ();
 FILLCELL_X32 FILLER_133_3519 ();
 FILLCELL_X32 FILLER_133_3551 ();
 FILLCELL_X32 FILLER_133_3583 ();
 FILLCELL_X32 FILLER_133_3615 ();
 FILLCELL_X32 FILLER_133_3647 ();
 FILLCELL_X32 FILLER_133_3679 ();
 FILLCELL_X16 FILLER_133_3711 ();
 FILLCELL_X8 FILLER_133_3727 ();
 FILLCELL_X2 FILLER_133_3735 ();
 FILLCELL_X1 FILLER_133_3737 ();
 FILLCELL_X32 FILLER_134_1 ();
 FILLCELL_X32 FILLER_134_33 ();
 FILLCELL_X32 FILLER_134_65 ();
 FILLCELL_X32 FILLER_134_97 ();
 FILLCELL_X32 FILLER_134_129 ();
 FILLCELL_X32 FILLER_134_161 ();
 FILLCELL_X32 FILLER_134_193 ();
 FILLCELL_X32 FILLER_134_225 ();
 FILLCELL_X32 FILLER_134_257 ();
 FILLCELL_X32 FILLER_134_289 ();
 FILLCELL_X32 FILLER_134_321 ();
 FILLCELL_X32 FILLER_134_353 ();
 FILLCELL_X32 FILLER_134_385 ();
 FILLCELL_X32 FILLER_134_417 ();
 FILLCELL_X32 FILLER_134_449 ();
 FILLCELL_X32 FILLER_134_481 ();
 FILLCELL_X32 FILLER_134_513 ();
 FILLCELL_X32 FILLER_134_545 ();
 FILLCELL_X32 FILLER_134_577 ();
 FILLCELL_X16 FILLER_134_609 ();
 FILLCELL_X4 FILLER_134_625 ();
 FILLCELL_X2 FILLER_134_629 ();
 FILLCELL_X32 FILLER_134_632 ();
 FILLCELL_X32 FILLER_134_664 ();
 FILLCELL_X32 FILLER_134_696 ();
 FILLCELL_X32 FILLER_134_728 ();
 FILLCELL_X32 FILLER_134_760 ();
 FILLCELL_X32 FILLER_134_792 ();
 FILLCELL_X32 FILLER_134_824 ();
 FILLCELL_X32 FILLER_134_856 ();
 FILLCELL_X32 FILLER_134_888 ();
 FILLCELL_X32 FILLER_134_920 ();
 FILLCELL_X32 FILLER_134_952 ();
 FILLCELL_X32 FILLER_134_984 ();
 FILLCELL_X32 FILLER_134_1016 ();
 FILLCELL_X32 FILLER_134_1048 ();
 FILLCELL_X32 FILLER_134_1080 ();
 FILLCELL_X32 FILLER_134_1112 ();
 FILLCELL_X32 FILLER_134_1144 ();
 FILLCELL_X32 FILLER_134_1176 ();
 FILLCELL_X32 FILLER_134_1208 ();
 FILLCELL_X32 FILLER_134_1240 ();
 FILLCELL_X32 FILLER_134_1272 ();
 FILLCELL_X32 FILLER_134_1304 ();
 FILLCELL_X32 FILLER_134_1336 ();
 FILLCELL_X32 FILLER_134_1368 ();
 FILLCELL_X32 FILLER_134_1400 ();
 FILLCELL_X32 FILLER_134_1432 ();
 FILLCELL_X32 FILLER_134_1464 ();
 FILLCELL_X32 FILLER_134_1496 ();
 FILLCELL_X32 FILLER_134_1528 ();
 FILLCELL_X32 FILLER_134_1560 ();
 FILLCELL_X32 FILLER_134_1592 ();
 FILLCELL_X32 FILLER_134_1624 ();
 FILLCELL_X32 FILLER_134_1656 ();
 FILLCELL_X32 FILLER_134_1688 ();
 FILLCELL_X32 FILLER_134_1720 ();
 FILLCELL_X32 FILLER_134_1752 ();
 FILLCELL_X32 FILLER_134_1784 ();
 FILLCELL_X32 FILLER_134_1816 ();
 FILLCELL_X32 FILLER_134_1848 ();
 FILLCELL_X8 FILLER_134_1880 ();
 FILLCELL_X4 FILLER_134_1888 ();
 FILLCELL_X2 FILLER_134_1892 ();
 FILLCELL_X32 FILLER_134_1895 ();
 FILLCELL_X32 FILLER_134_1927 ();
 FILLCELL_X32 FILLER_134_1959 ();
 FILLCELL_X32 FILLER_134_1991 ();
 FILLCELL_X32 FILLER_134_2023 ();
 FILLCELL_X32 FILLER_134_2055 ();
 FILLCELL_X32 FILLER_134_2087 ();
 FILLCELL_X32 FILLER_134_2119 ();
 FILLCELL_X32 FILLER_134_2151 ();
 FILLCELL_X32 FILLER_134_2183 ();
 FILLCELL_X32 FILLER_134_2215 ();
 FILLCELL_X32 FILLER_134_2247 ();
 FILLCELL_X32 FILLER_134_2279 ();
 FILLCELL_X32 FILLER_134_2311 ();
 FILLCELL_X32 FILLER_134_2343 ();
 FILLCELL_X32 FILLER_134_2375 ();
 FILLCELL_X32 FILLER_134_2407 ();
 FILLCELL_X32 FILLER_134_2439 ();
 FILLCELL_X32 FILLER_134_2471 ();
 FILLCELL_X32 FILLER_134_2503 ();
 FILLCELL_X32 FILLER_134_2535 ();
 FILLCELL_X32 FILLER_134_2567 ();
 FILLCELL_X32 FILLER_134_2599 ();
 FILLCELL_X32 FILLER_134_2631 ();
 FILLCELL_X32 FILLER_134_2663 ();
 FILLCELL_X32 FILLER_134_2695 ();
 FILLCELL_X32 FILLER_134_2727 ();
 FILLCELL_X32 FILLER_134_2759 ();
 FILLCELL_X32 FILLER_134_2791 ();
 FILLCELL_X32 FILLER_134_2823 ();
 FILLCELL_X32 FILLER_134_2855 ();
 FILLCELL_X32 FILLER_134_2887 ();
 FILLCELL_X32 FILLER_134_2919 ();
 FILLCELL_X32 FILLER_134_2951 ();
 FILLCELL_X32 FILLER_134_2983 ();
 FILLCELL_X32 FILLER_134_3015 ();
 FILLCELL_X32 FILLER_134_3047 ();
 FILLCELL_X32 FILLER_134_3079 ();
 FILLCELL_X32 FILLER_134_3111 ();
 FILLCELL_X8 FILLER_134_3143 ();
 FILLCELL_X4 FILLER_134_3151 ();
 FILLCELL_X2 FILLER_134_3155 ();
 FILLCELL_X32 FILLER_134_3158 ();
 FILLCELL_X32 FILLER_134_3190 ();
 FILLCELL_X32 FILLER_134_3222 ();
 FILLCELL_X32 FILLER_134_3254 ();
 FILLCELL_X32 FILLER_134_3286 ();
 FILLCELL_X32 FILLER_134_3318 ();
 FILLCELL_X32 FILLER_134_3350 ();
 FILLCELL_X32 FILLER_134_3382 ();
 FILLCELL_X32 FILLER_134_3414 ();
 FILLCELL_X32 FILLER_134_3446 ();
 FILLCELL_X32 FILLER_134_3478 ();
 FILLCELL_X32 FILLER_134_3510 ();
 FILLCELL_X32 FILLER_134_3542 ();
 FILLCELL_X32 FILLER_134_3574 ();
 FILLCELL_X32 FILLER_134_3606 ();
 FILLCELL_X32 FILLER_134_3638 ();
 FILLCELL_X32 FILLER_134_3670 ();
 FILLCELL_X32 FILLER_134_3702 ();
 FILLCELL_X4 FILLER_134_3734 ();
 FILLCELL_X32 FILLER_135_1 ();
 FILLCELL_X32 FILLER_135_33 ();
 FILLCELL_X32 FILLER_135_65 ();
 FILLCELL_X32 FILLER_135_97 ();
 FILLCELL_X32 FILLER_135_129 ();
 FILLCELL_X32 FILLER_135_161 ();
 FILLCELL_X32 FILLER_135_193 ();
 FILLCELL_X32 FILLER_135_225 ();
 FILLCELL_X32 FILLER_135_257 ();
 FILLCELL_X32 FILLER_135_289 ();
 FILLCELL_X32 FILLER_135_321 ();
 FILLCELL_X32 FILLER_135_353 ();
 FILLCELL_X32 FILLER_135_385 ();
 FILLCELL_X32 FILLER_135_417 ();
 FILLCELL_X32 FILLER_135_449 ();
 FILLCELL_X32 FILLER_135_481 ();
 FILLCELL_X32 FILLER_135_513 ();
 FILLCELL_X32 FILLER_135_545 ();
 FILLCELL_X32 FILLER_135_577 ();
 FILLCELL_X32 FILLER_135_609 ();
 FILLCELL_X32 FILLER_135_641 ();
 FILLCELL_X32 FILLER_135_673 ();
 FILLCELL_X32 FILLER_135_705 ();
 FILLCELL_X32 FILLER_135_737 ();
 FILLCELL_X32 FILLER_135_769 ();
 FILLCELL_X32 FILLER_135_801 ();
 FILLCELL_X32 FILLER_135_833 ();
 FILLCELL_X32 FILLER_135_865 ();
 FILLCELL_X32 FILLER_135_897 ();
 FILLCELL_X32 FILLER_135_929 ();
 FILLCELL_X32 FILLER_135_961 ();
 FILLCELL_X32 FILLER_135_993 ();
 FILLCELL_X32 FILLER_135_1025 ();
 FILLCELL_X32 FILLER_135_1057 ();
 FILLCELL_X32 FILLER_135_1089 ();
 FILLCELL_X32 FILLER_135_1121 ();
 FILLCELL_X32 FILLER_135_1153 ();
 FILLCELL_X32 FILLER_135_1185 ();
 FILLCELL_X32 FILLER_135_1217 ();
 FILLCELL_X8 FILLER_135_1249 ();
 FILLCELL_X4 FILLER_135_1257 ();
 FILLCELL_X2 FILLER_135_1261 ();
 FILLCELL_X32 FILLER_135_1264 ();
 FILLCELL_X32 FILLER_135_1296 ();
 FILLCELL_X32 FILLER_135_1328 ();
 FILLCELL_X32 FILLER_135_1360 ();
 FILLCELL_X32 FILLER_135_1392 ();
 FILLCELL_X32 FILLER_135_1424 ();
 FILLCELL_X32 FILLER_135_1456 ();
 FILLCELL_X32 FILLER_135_1488 ();
 FILLCELL_X32 FILLER_135_1520 ();
 FILLCELL_X32 FILLER_135_1552 ();
 FILLCELL_X32 FILLER_135_1584 ();
 FILLCELL_X32 FILLER_135_1616 ();
 FILLCELL_X32 FILLER_135_1648 ();
 FILLCELL_X32 FILLER_135_1680 ();
 FILLCELL_X32 FILLER_135_1712 ();
 FILLCELL_X32 FILLER_135_1744 ();
 FILLCELL_X32 FILLER_135_1776 ();
 FILLCELL_X32 FILLER_135_1808 ();
 FILLCELL_X32 FILLER_135_1840 ();
 FILLCELL_X32 FILLER_135_1872 ();
 FILLCELL_X32 FILLER_135_1904 ();
 FILLCELL_X32 FILLER_135_1936 ();
 FILLCELL_X32 FILLER_135_1968 ();
 FILLCELL_X32 FILLER_135_2000 ();
 FILLCELL_X32 FILLER_135_2032 ();
 FILLCELL_X32 FILLER_135_2064 ();
 FILLCELL_X32 FILLER_135_2096 ();
 FILLCELL_X32 FILLER_135_2128 ();
 FILLCELL_X32 FILLER_135_2160 ();
 FILLCELL_X32 FILLER_135_2192 ();
 FILLCELL_X32 FILLER_135_2224 ();
 FILLCELL_X32 FILLER_135_2256 ();
 FILLCELL_X32 FILLER_135_2288 ();
 FILLCELL_X32 FILLER_135_2320 ();
 FILLCELL_X32 FILLER_135_2352 ();
 FILLCELL_X32 FILLER_135_2384 ();
 FILLCELL_X32 FILLER_135_2416 ();
 FILLCELL_X32 FILLER_135_2448 ();
 FILLCELL_X32 FILLER_135_2480 ();
 FILLCELL_X8 FILLER_135_2512 ();
 FILLCELL_X4 FILLER_135_2520 ();
 FILLCELL_X2 FILLER_135_2524 ();
 FILLCELL_X32 FILLER_135_2527 ();
 FILLCELL_X32 FILLER_135_2559 ();
 FILLCELL_X32 FILLER_135_2591 ();
 FILLCELL_X32 FILLER_135_2623 ();
 FILLCELL_X32 FILLER_135_2655 ();
 FILLCELL_X32 FILLER_135_2687 ();
 FILLCELL_X32 FILLER_135_2719 ();
 FILLCELL_X32 FILLER_135_2751 ();
 FILLCELL_X32 FILLER_135_2783 ();
 FILLCELL_X32 FILLER_135_2815 ();
 FILLCELL_X32 FILLER_135_2847 ();
 FILLCELL_X32 FILLER_135_2879 ();
 FILLCELL_X32 FILLER_135_2911 ();
 FILLCELL_X32 FILLER_135_2943 ();
 FILLCELL_X32 FILLER_135_2975 ();
 FILLCELL_X32 FILLER_135_3007 ();
 FILLCELL_X32 FILLER_135_3039 ();
 FILLCELL_X32 FILLER_135_3071 ();
 FILLCELL_X32 FILLER_135_3103 ();
 FILLCELL_X32 FILLER_135_3135 ();
 FILLCELL_X32 FILLER_135_3167 ();
 FILLCELL_X32 FILLER_135_3199 ();
 FILLCELL_X32 FILLER_135_3231 ();
 FILLCELL_X32 FILLER_135_3263 ();
 FILLCELL_X32 FILLER_135_3295 ();
 FILLCELL_X32 FILLER_135_3327 ();
 FILLCELL_X32 FILLER_135_3359 ();
 FILLCELL_X32 FILLER_135_3391 ();
 FILLCELL_X32 FILLER_135_3423 ();
 FILLCELL_X32 FILLER_135_3455 ();
 FILLCELL_X32 FILLER_135_3487 ();
 FILLCELL_X32 FILLER_135_3519 ();
 FILLCELL_X32 FILLER_135_3551 ();
 FILLCELL_X32 FILLER_135_3583 ();
 FILLCELL_X32 FILLER_135_3615 ();
 FILLCELL_X32 FILLER_135_3647 ();
 FILLCELL_X32 FILLER_135_3679 ();
 FILLCELL_X16 FILLER_135_3711 ();
 FILLCELL_X8 FILLER_135_3727 ();
 FILLCELL_X2 FILLER_135_3735 ();
 FILLCELL_X1 FILLER_135_3737 ();
 FILLCELL_X32 FILLER_136_1 ();
 FILLCELL_X32 FILLER_136_33 ();
 FILLCELL_X32 FILLER_136_65 ();
 FILLCELL_X32 FILLER_136_97 ();
 FILLCELL_X32 FILLER_136_129 ();
 FILLCELL_X32 FILLER_136_161 ();
 FILLCELL_X32 FILLER_136_193 ();
 FILLCELL_X32 FILLER_136_225 ();
 FILLCELL_X32 FILLER_136_257 ();
 FILLCELL_X32 FILLER_136_289 ();
 FILLCELL_X32 FILLER_136_321 ();
 FILLCELL_X32 FILLER_136_353 ();
 FILLCELL_X32 FILLER_136_385 ();
 FILLCELL_X32 FILLER_136_417 ();
 FILLCELL_X32 FILLER_136_449 ();
 FILLCELL_X32 FILLER_136_481 ();
 FILLCELL_X32 FILLER_136_513 ();
 FILLCELL_X32 FILLER_136_545 ();
 FILLCELL_X32 FILLER_136_577 ();
 FILLCELL_X16 FILLER_136_609 ();
 FILLCELL_X4 FILLER_136_625 ();
 FILLCELL_X2 FILLER_136_629 ();
 FILLCELL_X32 FILLER_136_632 ();
 FILLCELL_X32 FILLER_136_664 ();
 FILLCELL_X32 FILLER_136_696 ();
 FILLCELL_X32 FILLER_136_728 ();
 FILLCELL_X32 FILLER_136_760 ();
 FILLCELL_X32 FILLER_136_792 ();
 FILLCELL_X32 FILLER_136_824 ();
 FILLCELL_X32 FILLER_136_856 ();
 FILLCELL_X32 FILLER_136_888 ();
 FILLCELL_X32 FILLER_136_920 ();
 FILLCELL_X32 FILLER_136_952 ();
 FILLCELL_X32 FILLER_136_984 ();
 FILLCELL_X32 FILLER_136_1016 ();
 FILLCELL_X32 FILLER_136_1048 ();
 FILLCELL_X32 FILLER_136_1080 ();
 FILLCELL_X32 FILLER_136_1112 ();
 FILLCELL_X32 FILLER_136_1144 ();
 FILLCELL_X32 FILLER_136_1176 ();
 FILLCELL_X32 FILLER_136_1208 ();
 FILLCELL_X32 FILLER_136_1240 ();
 FILLCELL_X32 FILLER_136_1272 ();
 FILLCELL_X32 FILLER_136_1304 ();
 FILLCELL_X32 FILLER_136_1336 ();
 FILLCELL_X32 FILLER_136_1368 ();
 FILLCELL_X32 FILLER_136_1400 ();
 FILLCELL_X32 FILLER_136_1432 ();
 FILLCELL_X32 FILLER_136_1464 ();
 FILLCELL_X32 FILLER_136_1496 ();
 FILLCELL_X32 FILLER_136_1528 ();
 FILLCELL_X32 FILLER_136_1560 ();
 FILLCELL_X32 FILLER_136_1592 ();
 FILLCELL_X32 FILLER_136_1624 ();
 FILLCELL_X32 FILLER_136_1656 ();
 FILLCELL_X32 FILLER_136_1688 ();
 FILLCELL_X32 FILLER_136_1720 ();
 FILLCELL_X32 FILLER_136_1752 ();
 FILLCELL_X32 FILLER_136_1784 ();
 FILLCELL_X32 FILLER_136_1816 ();
 FILLCELL_X32 FILLER_136_1848 ();
 FILLCELL_X8 FILLER_136_1880 ();
 FILLCELL_X4 FILLER_136_1888 ();
 FILLCELL_X2 FILLER_136_1892 ();
 FILLCELL_X32 FILLER_136_1895 ();
 FILLCELL_X32 FILLER_136_1927 ();
 FILLCELL_X32 FILLER_136_1959 ();
 FILLCELL_X32 FILLER_136_1991 ();
 FILLCELL_X32 FILLER_136_2023 ();
 FILLCELL_X32 FILLER_136_2055 ();
 FILLCELL_X32 FILLER_136_2087 ();
 FILLCELL_X32 FILLER_136_2119 ();
 FILLCELL_X32 FILLER_136_2151 ();
 FILLCELL_X32 FILLER_136_2183 ();
 FILLCELL_X32 FILLER_136_2215 ();
 FILLCELL_X32 FILLER_136_2247 ();
 FILLCELL_X32 FILLER_136_2279 ();
 FILLCELL_X32 FILLER_136_2311 ();
 FILLCELL_X32 FILLER_136_2343 ();
 FILLCELL_X32 FILLER_136_2375 ();
 FILLCELL_X32 FILLER_136_2407 ();
 FILLCELL_X32 FILLER_136_2439 ();
 FILLCELL_X32 FILLER_136_2471 ();
 FILLCELL_X32 FILLER_136_2503 ();
 FILLCELL_X32 FILLER_136_2535 ();
 FILLCELL_X32 FILLER_136_2567 ();
 FILLCELL_X32 FILLER_136_2599 ();
 FILLCELL_X32 FILLER_136_2631 ();
 FILLCELL_X32 FILLER_136_2663 ();
 FILLCELL_X32 FILLER_136_2695 ();
 FILLCELL_X32 FILLER_136_2727 ();
 FILLCELL_X32 FILLER_136_2759 ();
 FILLCELL_X32 FILLER_136_2791 ();
 FILLCELL_X32 FILLER_136_2823 ();
 FILLCELL_X32 FILLER_136_2855 ();
 FILLCELL_X32 FILLER_136_2887 ();
 FILLCELL_X32 FILLER_136_2919 ();
 FILLCELL_X32 FILLER_136_2951 ();
 FILLCELL_X32 FILLER_136_2983 ();
 FILLCELL_X32 FILLER_136_3015 ();
 FILLCELL_X32 FILLER_136_3047 ();
 FILLCELL_X32 FILLER_136_3079 ();
 FILLCELL_X32 FILLER_136_3111 ();
 FILLCELL_X8 FILLER_136_3143 ();
 FILLCELL_X4 FILLER_136_3151 ();
 FILLCELL_X2 FILLER_136_3155 ();
 FILLCELL_X32 FILLER_136_3158 ();
 FILLCELL_X32 FILLER_136_3190 ();
 FILLCELL_X32 FILLER_136_3222 ();
 FILLCELL_X32 FILLER_136_3254 ();
 FILLCELL_X32 FILLER_136_3286 ();
 FILLCELL_X32 FILLER_136_3318 ();
 FILLCELL_X32 FILLER_136_3350 ();
 FILLCELL_X32 FILLER_136_3382 ();
 FILLCELL_X32 FILLER_136_3414 ();
 FILLCELL_X32 FILLER_136_3446 ();
 FILLCELL_X32 FILLER_136_3478 ();
 FILLCELL_X32 FILLER_136_3510 ();
 FILLCELL_X32 FILLER_136_3542 ();
 FILLCELL_X32 FILLER_136_3574 ();
 FILLCELL_X32 FILLER_136_3606 ();
 FILLCELL_X32 FILLER_136_3638 ();
 FILLCELL_X32 FILLER_136_3670 ();
 FILLCELL_X32 FILLER_136_3702 ();
 FILLCELL_X4 FILLER_136_3734 ();
 FILLCELL_X32 FILLER_137_1 ();
 FILLCELL_X32 FILLER_137_33 ();
 FILLCELL_X32 FILLER_137_65 ();
 FILLCELL_X32 FILLER_137_97 ();
 FILLCELL_X32 FILLER_137_129 ();
 FILLCELL_X32 FILLER_137_161 ();
 FILLCELL_X32 FILLER_137_193 ();
 FILLCELL_X32 FILLER_137_225 ();
 FILLCELL_X32 FILLER_137_257 ();
 FILLCELL_X32 FILLER_137_289 ();
 FILLCELL_X32 FILLER_137_321 ();
 FILLCELL_X32 FILLER_137_353 ();
 FILLCELL_X32 FILLER_137_385 ();
 FILLCELL_X32 FILLER_137_417 ();
 FILLCELL_X32 FILLER_137_449 ();
 FILLCELL_X32 FILLER_137_481 ();
 FILLCELL_X32 FILLER_137_513 ();
 FILLCELL_X32 FILLER_137_545 ();
 FILLCELL_X32 FILLER_137_577 ();
 FILLCELL_X32 FILLER_137_609 ();
 FILLCELL_X32 FILLER_137_641 ();
 FILLCELL_X32 FILLER_137_673 ();
 FILLCELL_X32 FILLER_137_705 ();
 FILLCELL_X32 FILLER_137_737 ();
 FILLCELL_X32 FILLER_137_769 ();
 FILLCELL_X32 FILLER_137_801 ();
 FILLCELL_X32 FILLER_137_833 ();
 FILLCELL_X32 FILLER_137_865 ();
 FILLCELL_X32 FILLER_137_897 ();
 FILLCELL_X32 FILLER_137_929 ();
 FILLCELL_X32 FILLER_137_961 ();
 FILLCELL_X32 FILLER_137_993 ();
 FILLCELL_X32 FILLER_137_1025 ();
 FILLCELL_X32 FILLER_137_1057 ();
 FILLCELL_X32 FILLER_137_1089 ();
 FILLCELL_X32 FILLER_137_1121 ();
 FILLCELL_X32 FILLER_137_1153 ();
 FILLCELL_X32 FILLER_137_1185 ();
 FILLCELL_X32 FILLER_137_1217 ();
 FILLCELL_X8 FILLER_137_1249 ();
 FILLCELL_X4 FILLER_137_1257 ();
 FILLCELL_X2 FILLER_137_1261 ();
 FILLCELL_X32 FILLER_137_1264 ();
 FILLCELL_X32 FILLER_137_1296 ();
 FILLCELL_X32 FILLER_137_1328 ();
 FILLCELL_X32 FILLER_137_1360 ();
 FILLCELL_X32 FILLER_137_1392 ();
 FILLCELL_X32 FILLER_137_1424 ();
 FILLCELL_X32 FILLER_137_1456 ();
 FILLCELL_X32 FILLER_137_1488 ();
 FILLCELL_X32 FILLER_137_1520 ();
 FILLCELL_X32 FILLER_137_1552 ();
 FILLCELL_X32 FILLER_137_1584 ();
 FILLCELL_X32 FILLER_137_1616 ();
 FILLCELL_X32 FILLER_137_1648 ();
 FILLCELL_X32 FILLER_137_1680 ();
 FILLCELL_X32 FILLER_137_1712 ();
 FILLCELL_X32 FILLER_137_1744 ();
 FILLCELL_X32 FILLER_137_1776 ();
 FILLCELL_X32 FILLER_137_1808 ();
 FILLCELL_X32 FILLER_137_1840 ();
 FILLCELL_X32 FILLER_137_1872 ();
 FILLCELL_X32 FILLER_137_1904 ();
 FILLCELL_X32 FILLER_137_1936 ();
 FILLCELL_X32 FILLER_137_1968 ();
 FILLCELL_X32 FILLER_137_2000 ();
 FILLCELL_X32 FILLER_137_2032 ();
 FILLCELL_X32 FILLER_137_2064 ();
 FILLCELL_X32 FILLER_137_2096 ();
 FILLCELL_X32 FILLER_137_2128 ();
 FILLCELL_X32 FILLER_137_2160 ();
 FILLCELL_X32 FILLER_137_2192 ();
 FILLCELL_X32 FILLER_137_2224 ();
 FILLCELL_X32 FILLER_137_2256 ();
 FILLCELL_X32 FILLER_137_2288 ();
 FILLCELL_X32 FILLER_137_2320 ();
 FILLCELL_X32 FILLER_137_2352 ();
 FILLCELL_X32 FILLER_137_2384 ();
 FILLCELL_X32 FILLER_137_2416 ();
 FILLCELL_X32 FILLER_137_2448 ();
 FILLCELL_X32 FILLER_137_2480 ();
 FILLCELL_X8 FILLER_137_2512 ();
 FILLCELL_X4 FILLER_137_2520 ();
 FILLCELL_X2 FILLER_137_2524 ();
 FILLCELL_X32 FILLER_137_2527 ();
 FILLCELL_X32 FILLER_137_2559 ();
 FILLCELL_X32 FILLER_137_2591 ();
 FILLCELL_X32 FILLER_137_2623 ();
 FILLCELL_X32 FILLER_137_2655 ();
 FILLCELL_X32 FILLER_137_2687 ();
 FILLCELL_X32 FILLER_137_2719 ();
 FILLCELL_X32 FILLER_137_2751 ();
 FILLCELL_X32 FILLER_137_2783 ();
 FILLCELL_X32 FILLER_137_2815 ();
 FILLCELL_X32 FILLER_137_2847 ();
 FILLCELL_X32 FILLER_137_2879 ();
 FILLCELL_X32 FILLER_137_2911 ();
 FILLCELL_X32 FILLER_137_2943 ();
 FILLCELL_X32 FILLER_137_2975 ();
 FILLCELL_X32 FILLER_137_3007 ();
 FILLCELL_X32 FILLER_137_3039 ();
 FILLCELL_X32 FILLER_137_3071 ();
 FILLCELL_X32 FILLER_137_3103 ();
 FILLCELL_X32 FILLER_137_3135 ();
 FILLCELL_X32 FILLER_137_3167 ();
 FILLCELL_X32 FILLER_137_3199 ();
 FILLCELL_X32 FILLER_137_3231 ();
 FILLCELL_X32 FILLER_137_3263 ();
 FILLCELL_X32 FILLER_137_3295 ();
 FILLCELL_X32 FILLER_137_3327 ();
 FILLCELL_X32 FILLER_137_3359 ();
 FILLCELL_X32 FILLER_137_3391 ();
 FILLCELL_X32 FILLER_137_3423 ();
 FILLCELL_X32 FILLER_137_3455 ();
 FILLCELL_X32 FILLER_137_3487 ();
 FILLCELL_X32 FILLER_137_3519 ();
 FILLCELL_X32 FILLER_137_3551 ();
 FILLCELL_X32 FILLER_137_3583 ();
 FILLCELL_X32 FILLER_137_3615 ();
 FILLCELL_X32 FILLER_137_3647 ();
 FILLCELL_X32 FILLER_137_3679 ();
 FILLCELL_X16 FILLER_137_3711 ();
 FILLCELL_X8 FILLER_137_3727 ();
 FILLCELL_X2 FILLER_137_3735 ();
 FILLCELL_X1 FILLER_137_3737 ();
 FILLCELL_X32 FILLER_138_1 ();
 FILLCELL_X32 FILLER_138_33 ();
 FILLCELL_X32 FILLER_138_65 ();
 FILLCELL_X32 FILLER_138_97 ();
 FILLCELL_X32 FILLER_138_129 ();
 FILLCELL_X32 FILLER_138_161 ();
 FILLCELL_X32 FILLER_138_193 ();
 FILLCELL_X32 FILLER_138_225 ();
 FILLCELL_X32 FILLER_138_257 ();
 FILLCELL_X32 FILLER_138_289 ();
 FILLCELL_X32 FILLER_138_321 ();
 FILLCELL_X32 FILLER_138_353 ();
 FILLCELL_X32 FILLER_138_385 ();
 FILLCELL_X32 FILLER_138_417 ();
 FILLCELL_X32 FILLER_138_449 ();
 FILLCELL_X32 FILLER_138_481 ();
 FILLCELL_X32 FILLER_138_513 ();
 FILLCELL_X32 FILLER_138_545 ();
 FILLCELL_X32 FILLER_138_577 ();
 FILLCELL_X16 FILLER_138_609 ();
 FILLCELL_X4 FILLER_138_625 ();
 FILLCELL_X2 FILLER_138_629 ();
 FILLCELL_X32 FILLER_138_632 ();
 FILLCELL_X32 FILLER_138_664 ();
 FILLCELL_X32 FILLER_138_696 ();
 FILLCELL_X32 FILLER_138_728 ();
 FILLCELL_X32 FILLER_138_760 ();
 FILLCELL_X32 FILLER_138_792 ();
 FILLCELL_X32 FILLER_138_824 ();
 FILLCELL_X32 FILLER_138_856 ();
 FILLCELL_X32 FILLER_138_888 ();
 FILLCELL_X32 FILLER_138_920 ();
 FILLCELL_X32 FILLER_138_952 ();
 FILLCELL_X32 FILLER_138_984 ();
 FILLCELL_X32 FILLER_138_1016 ();
 FILLCELL_X32 FILLER_138_1048 ();
 FILLCELL_X32 FILLER_138_1080 ();
 FILLCELL_X32 FILLER_138_1112 ();
 FILLCELL_X32 FILLER_138_1144 ();
 FILLCELL_X32 FILLER_138_1176 ();
 FILLCELL_X32 FILLER_138_1208 ();
 FILLCELL_X32 FILLER_138_1240 ();
 FILLCELL_X32 FILLER_138_1272 ();
 FILLCELL_X32 FILLER_138_1304 ();
 FILLCELL_X32 FILLER_138_1336 ();
 FILLCELL_X32 FILLER_138_1368 ();
 FILLCELL_X32 FILLER_138_1400 ();
 FILLCELL_X32 FILLER_138_1432 ();
 FILLCELL_X32 FILLER_138_1464 ();
 FILLCELL_X32 FILLER_138_1496 ();
 FILLCELL_X32 FILLER_138_1528 ();
 FILLCELL_X32 FILLER_138_1560 ();
 FILLCELL_X32 FILLER_138_1592 ();
 FILLCELL_X32 FILLER_138_1624 ();
 FILLCELL_X32 FILLER_138_1656 ();
 FILLCELL_X32 FILLER_138_1688 ();
 FILLCELL_X32 FILLER_138_1720 ();
 FILLCELL_X32 FILLER_138_1752 ();
 FILLCELL_X32 FILLER_138_1784 ();
 FILLCELL_X32 FILLER_138_1816 ();
 FILLCELL_X32 FILLER_138_1848 ();
 FILLCELL_X8 FILLER_138_1880 ();
 FILLCELL_X4 FILLER_138_1888 ();
 FILLCELL_X2 FILLER_138_1892 ();
 FILLCELL_X32 FILLER_138_1895 ();
 FILLCELL_X32 FILLER_138_1927 ();
 FILLCELL_X32 FILLER_138_1959 ();
 FILLCELL_X32 FILLER_138_1991 ();
 FILLCELL_X32 FILLER_138_2023 ();
 FILLCELL_X32 FILLER_138_2055 ();
 FILLCELL_X32 FILLER_138_2087 ();
 FILLCELL_X32 FILLER_138_2119 ();
 FILLCELL_X32 FILLER_138_2151 ();
 FILLCELL_X32 FILLER_138_2183 ();
 FILLCELL_X32 FILLER_138_2215 ();
 FILLCELL_X32 FILLER_138_2247 ();
 FILLCELL_X32 FILLER_138_2279 ();
 FILLCELL_X32 FILLER_138_2311 ();
 FILLCELL_X32 FILLER_138_2343 ();
 FILLCELL_X32 FILLER_138_2375 ();
 FILLCELL_X32 FILLER_138_2407 ();
 FILLCELL_X32 FILLER_138_2439 ();
 FILLCELL_X32 FILLER_138_2471 ();
 FILLCELL_X32 FILLER_138_2503 ();
 FILLCELL_X32 FILLER_138_2535 ();
 FILLCELL_X32 FILLER_138_2567 ();
 FILLCELL_X32 FILLER_138_2599 ();
 FILLCELL_X32 FILLER_138_2631 ();
 FILLCELL_X32 FILLER_138_2663 ();
 FILLCELL_X32 FILLER_138_2695 ();
 FILLCELL_X32 FILLER_138_2727 ();
 FILLCELL_X32 FILLER_138_2759 ();
 FILLCELL_X32 FILLER_138_2791 ();
 FILLCELL_X32 FILLER_138_2823 ();
 FILLCELL_X32 FILLER_138_2855 ();
 FILLCELL_X32 FILLER_138_2887 ();
 FILLCELL_X32 FILLER_138_2919 ();
 FILLCELL_X32 FILLER_138_2951 ();
 FILLCELL_X32 FILLER_138_2983 ();
 FILLCELL_X32 FILLER_138_3015 ();
 FILLCELL_X32 FILLER_138_3047 ();
 FILLCELL_X32 FILLER_138_3079 ();
 FILLCELL_X32 FILLER_138_3111 ();
 FILLCELL_X8 FILLER_138_3143 ();
 FILLCELL_X4 FILLER_138_3151 ();
 FILLCELL_X2 FILLER_138_3155 ();
 FILLCELL_X32 FILLER_138_3158 ();
 FILLCELL_X32 FILLER_138_3190 ();
 FILLCELL_X32 FILLER_138_3222 ();
 FILLCELL_X32 FILLER_138_3254 ();
 FILLCELL_X32 FILLER_138_3286 ();
 FILLCELL_X32 FILLER_138_3318 ();
 FILLCELL_X32 FILLER_138_3350 ();
 FILLCELL_X32 FILLER_138_3382 ();
 FILLCELL_X32 FILLER_138_3414 ();
 FILLCELL_X32 FILLER_138_3446 ();
 FILLCELL_X32 FILLER_138_3478 ();
 FILLCELL_X32 FILLER_138_3510 ();
 FILLCELL_X32 FILLER_138_3542 ();
 FILLCELL_X32 FILLER_138_3574 ();
 FILLCELL_X32 FILLER_138_3606 ();
 FILLCELL_X32 FILLER_138_3638 ();
 FILLCELL_X32 FILLER_138_3670 ();
 FILLCELL_X32 FILLER_138_3702 ();
 FILLCELL_X4 FILLER_138_3734 ();
 FILLCELL_X32 FILLER_139_1 ();
 FILLCELL_X32 FILLER_139_33 ();
 FILLCELL_X32 FILLER_139_65 ();
 FILLCELL_X32 FILLER_139_97 ();
 FILLCELL_X32 FILLER_139_129 ();
 FILLCELL_X32 FILLER_139_161 ();
 FILLCELL_X32 FILLER_139_193 ();
 FILLCELL_X32 FILLER_139_225 ();
 FILLCELL_X32 FILLER_139_257 ();
 FILLCELL_X32 FILLER_139_289 ();
 FILLCELL_X32 FILLER_139_321 ();
 FILLCELL_X32 FILLER_139_353 ();
 FILLCELL_X32 FILLER_139_385 ();
 FILLCELL_X32 FILLER_139_417 ();
 FILLCELL_X32 FILLER_139_449 ();
 FILLCELL_X32 FILLER_139_481 ();
 FILLCELL_X32 FILLER_139_513 ();
 FILLCELL_X32 FILLER_139_545 ();
 FILLCELL_X32 FILLER_139_577 ();
 FILLCELL_X32 FILLER_139_609 ();
 FILLCELL_X32 FILLER_139_641 ();
 FILLCELL_X32 FILLER_139_673 ();
 FILLCELL_X32 FILLER_139_705 ();
 FILLCELL_X32 FILLER_139_737 ();
 FILLCELL_X32 FILLER_139_769 ();
 FILLCELL_X32 FILLER_139_801 ();
 FILLCELL_X32 FILLER_139_833 ();
 FILLCELL_X32 FILLER_139_865 ();
 FILLCELL_X32 FILLER_139_897 ();
 FILLCELL_X32 FILLER_139_929 ();
 FILLCELL_X32 FILLER_139_961 ();
 FILLCELL_X32 FILLER_139_993 ();
 FILLCELL_X32 FILLER_139_1025 ();
 FILLCELL_X32 FILLER_139_1057 ();
 FILLCELL_X32 FILLER_139_1089 ();
 FILLCELL_X32 FILLER_139_1121 ();
 FILLCELL_X32 FILLER_139_1153 ();
 FILLCELL_X32 FILLER_139_1185 ();
 FILLCELL_X32 FILLER_139_1217 ();
 FILLCELL_X8 FILLER_139_1249 ();
 FILLCELL_X4 FILLER_139_1257 ();
 FILLCELL_X2 FILLER_139_1261 ();
 FILLCELL_X32 FILLER_139_1264 ();
 FILLCELL_X32 FILLER_139_1296 ();
 FILLCELL_X32 FILLER_139_1328 ();
 FILLCELL_X32 FILLER_139_1360 ();
 FILLCELL_X32 FILLER_139_1392 ();
 FILLCELL_X32 FILLER_139_1424 ();
 FILLCELL_X32 FILLER_139_1456 ();
 FILLCELL_X32 FILLER_139_1488 ();
 FILLCELL_X32 FILLER_139_1520 ();
 FILLCELL_X32 FILLER_139_1552 ();
 FILLCELL_X32 FILLER_139_1584 ();
 FILLCELL_X32 FILLER_139_1616 ();
 FILLCELL_X32 FILLER_139_1648 ();
 FILLCELL_X32 FILLER_139_1680 ();
 FILLCELL_X32 FILLER_139_1712 ();
 FILLCELL_X32 FILLER_139_1744 ();
 FILLCELL_X32 FILLER_139_1776 ();
 FILLCELL_X32 FILLER_139_1808 ();
 FILLCELL_X32 FILLER_139_1840 ();
 FILLCELL_X32 FILLER_139_1872 ();
 FILLCELL_X32 FILLER_139_1904 ();
 FILLCELL_X32 FILLER_139_1936 ();
 FILLCELL_X32 FILLER_139_1968 ();
 FILLCELL_X32 FILLER_139_2000 ();
 FILLCELL_X32 FILLER_139_2032 ();
 FILLCELL_X32 FILLER_139_2064 ();
 FILLCELL_X32 FILLER_139_2096 ();
 FILLCELL_X32 FILLER_139_2128 ();
 FILLCELL_X32 FILLER_139_2160 ();
 FILLCELL_X32 FILLER_139_2192 ();
 FILLCELL_X32 FILLER_139_2224 ();
 FILLCELL_X32 FILLER_139_2256 ();
 FILLCELL_X32 FILLER_139_2288 ();
 FILLCELL_X32 FILLER_139_2320 ();
 FILLCELL_X32 FILLER_139_2352 ();
 FILLCELL_X32 FILLER_139_2384 ();
 FILLCELL_X32 FILLER_139_2416 ();
 FILLCELL_X32 FILLER_139_2448 ();
 FILLCELL_X32 FILLER_139_2480 ();
 FILLCELL_X8 FILLER_139_2512 ();
 FILLCELL_X4 FILLER_139_2520 ();
 FILLCELL_X2 FILLER_139_2524 ();
 FILLCELL_X32 FILLER_139_2527 ();
 FILLCELL_X32 FILLER_139_2559 ();
 FILLCELL_X32 FILLER_139_2591 ();
 FILLCELL_X32 FILLER_139_2623 ();
 FILLCELL_X32 FILLER_139_2655 ();
 FILLCELL_X32 FILLER_139_2687 ();
 FILLCELL_X32 FILLER_139_2719 ();
 FILLCELL_X32 FILLER_139_2751 ();
 FILLCELL_X32 FILLER_139_2783 ();
 FILLCELL_X32 FILLER_139_2815 ();
 FILLCELL_X32 FILLER_139_2847 ();
 FILLCELL_X32 FILLER_139_2879 ();
 FILLCELL_X32 FILLER_139_2911 ();
 FILLCELL_X32 FILLER_139_2943 ();
 FILLCELL_X32 FILLER_139_2975 ();
 FILLCELL_X32 FILLER_139_3007 ();
 FILLCELL_X32 FILLER_139_3039 ();
 FILLCELL_X32 FILLER_139_3071 ();
 FILLCELL_X32 FILLER_139_3103 ();
 FILLCELL_X32 FILLER_139_3135 ();
 FILLCELL_X32 FILLER_139_3167 ();
 FILLCELL_X32 FILLER_139_3199 ();
 FILLCELL_X32 FILLER_139_3231 ();
 FILLCELL_X32 FILLER_139_3263 ();
 FILLCELL_X32 FILLER_139_3295 ();
 FILLCELL_X32 FILLER_139_3327 ();
 FILLCELL_X32 FILLER_139_3359 ();
 FILLCELL_X32 FILLER_139_3391 ();
 FILLCELL_X32 FILLER_139_3423 ();
 FILLCELL_X32 FILLER_139_3455 ();
 FILLCELL_X32 FILLER_139_3487 ();
 FILLCELL_X32 FILLER_139_3519 ();
 FILLCELL_X32 FILLER_139_3551 ();
 FILLCELL_X32 FILLER_139_3583 ();
 FILLCELL_X32 FILLER_139_3615 ();
 FILLCELL_X32 FILLER_139_3647 ();
 FILLCELL_X32 FILLER_139_3679 ();
 FILLCELL_X16 FILLER_139_3711 ();
 FILLCELL_X8 FILLER_139_3727 ();
 FILLCELL_X2 FILLER_139_3735 ();
 FILLCELL_X1 FILLER_139_3737 ();
 FILLCELL_X32 FILLER_140_1 ();
 FILLCELL_X32 FILLER_140_33 ();
 FILLCELL_X32 FILLER_140_65 ();
 FILLCELL_X32 FILLER_140_97 ();
 FILLCELL_X32 FILLER_140_129 ();
 FILLCELL_X32 FILLER_140_161 ();
 FILLCELL_X32 FILLER_140_193 ();
 FILLCELL_X32 FILLER_140_225 ();
 FILLCELL_X32 FILLER_140_257 ();
 FILLCELL_X32 FILLER_140_289 ();
 FILLCELL_X32 FILLER_140_321 ();
 FILLCELL_X32 FILLER_140_353 ();
 FILLCELL_X32 FILLER_140_385 ();
 FILLCELL_X32 FILLER_140_417 ();
 FILLCELL_X32 FILLER_140_449 ();
 FILLCELL_X32 FILLER_140_481 ();
 FILLCELL_X32 FILLER_140_513 ();
 FILLCELL_X32 FILLER_140_545 ();
 FILLCELL_X32 FILLER_140_577 ();
 FILLCELL_X16 FILLER_140_609 ();
 FILLCELL_X4 FILLER_140_625 ();
 FILLCELL_X2 FILLER_140_629 ();
 FILLCELL_X32 FILLER_140_632 ();
 FILLCELL_X32 FILLER_140_664 ();
 FILLCELL_X32 FILLER_140_696 ();
 FILLCELL_X32 FILLER_140_728 ();
 FILLCELL_X32 FILLER_140_760 ();
 FILLCELL_X32 FILLER_140_792 ();
 FILLCELL_X32 FILLER_140_824 ();
 FILLCELL_X32 FILLER_140_856 ();
 FILLCELL_X32 FILLER_140_888 ();
 FILLCELL_X32 FILLER_140_920 ();
 FILLCELL_X32 FILLER_140_952 ();
 FILLCELL_X32 FILLER_140_984 ();
 FILLCELL_X32 FILLER_140_1016 ();
 FILLCELL_X32 FILLER_140_1048 ();
 FILLCELL_X32 FILLER_140_1080 ();
 FILLCELL_X32 FILLER_140_1112 ();
 FILLCELL_X32 FILLER_140_1144 ();
 FILLCELL_X32 FILLER_140_1176 ();
 FILLCELL_X32 FILLER_140_1208 ();
 FILLCELL_X32 FILLER_140_1240 ();
 FILLCELL_X32 FILLER_140_1272 ();
 FILLCELL_X32 FILLER_140_1304 ();
 FILLCELL_X32 FILLER_140_1336 ();
 FILLCELL_X32 FILLER_140_1368 ();
 FILLCELL_X32 FILLER_140_1400 ();
 FILLCELL_X32 FILLER_140_1432 ();
 FILLCELL_X32 FILLER_140_1464 ();
 FILLCELL_X32 FILLER_140_1496 ();
 FILLCELL_X32 FILLER_140_1528 ();
 FILLCELL_X32 FILLER_140_1560 ();
 FILLCELL_X32 FILLER_140_1592 ();
 FILLCELL_X32 FILLER_140_1624 ();
 FILLCELL_X32 FILLER_140_1656 ();
 FILLCELL_X32 FILLER_140_1688 ();
 FILLCELL_X32 FILLER_140_1720 ();
 FILLCELL_X32 FILLER_140_1752 ();
 FILLCELL_X32 FILLER_140_1784 ();
 FILLCELL_X32 FILLER_140_1816 ();
 FILLCELL_X32 FILLER_140_1848 ();
 FILLCELL_X8 FILLER_140_1880 ();
 FILLCELL_X4 FILLER_140_1888 ();
 FILLCELL_X2 FILLER_140_1892 ();
 FILLCELL_X32 FILLER_140_1895 ();
 FILLCELL_X32 FILLER_140_1927 ();
 FILLCELL_X32 FILLER_140_1959 ();
 FILLCELL_X32 FILLER_140_1991 ();
 FILLCELL_X32 FILLER_140_2023 ();
 FILLCELL_X32 FILLER_140_2055 ();
 FILLCELL_X32 FILLER_140_2087 ();
 FILLCELL_X32 FILLER_140_2119 ();
 FILLCELL_X32 FILLER_140_2151 ();
 FILLCELL_X32 FILLER_140_2183 ();
 FILLCELL_X32 FILLER_140_2215 ();
 FILLCELL_X32 FILLER_140_2247 ();
 FILLCELL_X32 FILLER_140_2279 ();
 FILLCELL_X32 FILLER_140_2311 ();
 FILLCELL_X32 FILLER_140_2343 ();
 FILLCELL_X32 FILLER_140_2375 ();
 FILLCELL_X32 FILLER_140_2407 ();
 FILLCELL_X32 FILLER_140_2439 ();
 FILLCELL_X32 FILLER_140_2471 ();
 FILLCELL_X32 FILLER_140_2503 ();
 FILLCELL_X32 FILLER_140_2535 ();
 FILLCELL_X32 FILLER_140_2567 ();
 FILLCELL_X32 FILLER_140_2599 ();
 FILLCELL_X32 FILLER_140_2631 ();
 FILLCELL_X32 FILLER_140_2663 ();
 FILLCELL_X32 FILLER_140_2695 ();
 FILLCELL_X32 FILLER_140_2727 ();
 FILLCELL_X32 FILLER_140_2759 ();
 FILLCELL_X32 FILLER_140_2791 ();
 FILLCELL_X32 FILLER_140_2823 ();
 FILLCELL_X32 FILLER_140_2855 ();
 FILLCELL_X32 FILLER_140_2887 ();
 FILLCELL_X32 FILLER_140_2919 ();
 FILLCELL_X32 FILLER_140_2951 ();
 FILLCELL_X32 FILLER_140_2983 ();
 FILLCELL_X32 FILLER_140_3015 ();
 FILLCELL_X32 FILLER_140_3047 ();
 FILLCELL_X32 FILLER_140_3079 ();
 FILLCELL_X32 FILLER_140_3111 ();
 FILLCELL_X8 FILLER_140_3143 ();
 FILLCELL_X4 FILLER_140_3151 ();
 FILLCELL_X2 FILLER_140_3155 ();
 FILLCELL_X32 FILLER_140_3158 ();
 FILLCELL_X32 FILLER_140_3190 ();
 FILLCELL_X32 FILLER_140_3222 ();
 FILLCELL_X32 FILLER_140_3254 ();
 FILLCELL_X32 FILLER_140_3286 ();
 FILLCELL_X32 FILLER_140_3318 ();
 FILLCELL_X32 FILLER_140_3350 ();
 FILLCELL_X32 FILLER_140_3382 ();
 FILLCELL_X32 FILLER_140_3414 ();
 FILLCELL_X32 FILLER_140_3446 ();
 FILLCELL_X32 FILLER_140_3478 ();
 FILLCELL_X32 FILLER_140_3510 ();
 FILLCELL_X32 FILLER_140_3542 ();
 FILLCELL_X32 FILLER_140_3574 ();
 FILLCELL_X32 FILLER_140_3606 ();
 FILLCELL_X32 FILLER_140_3638 ();
 FILLCELL_X32 FILLER_140_3670 ();
 FILLCELL_X32 FILLER_140_3702 ();
 FILLCELL_X4 FILLER_140_3734 ();
 FILLCELL_X32 FILLER_141_1 ();
 FILLCELL_X32 FILLER_141_33 ();
 FILLCELL_X32 FILLER_141_65 ();
 FILLCELL_X32 FILLER_141_97 ();
 FILLCELL_X32 FILLER_141_129 ();
 FILLCELL_X32 FILLER_141_161 ();
 FILLCELL_X32 FILLER_141_193 ();
 FILLCELL_X32 FILLER_141_225 ();
 FILLCELL_X32 FILLER_141_257 ();
 FILLCELL_X32 FILLER_141_289 ();
 FILLCELL_X32 FILLER_141_321 ();
 FILLCELL_X32 FILLER_141_353 ();
 FILLCELL_X32 FILLER_141_385 ();
 FILLCELL_X32 FILLER_141_417 ();
 FILLCELL_X32 FILLER_141_449 ();
 FILLCELL_X32 FILLER_141_481 ();
 FILLCELL_X32 FILLER_141_513 ();
 FILLCELL_X32 FILLER_141_545 ();
 FILLCELL_X32 FILLER_141_577 ();
 FILLCELL_X32 FILLER_141_609 ();
 FILLCELL_X32 FILLER_141_641 ();
 FILLCELL_X32 FILLER_141_673 ();
 FILLCELL_X32 FILLER_141_705 ();
 FILLCELL_X32 FILLER_141_737 ();
 FILLCELL_X32 FILLER_141_769 ();
 FILLCELL_X32 FILLER_141_801 ();
 FILLCELL_X32 FILLER_141_833 ();
 FILLCELL_X32 FILLER_141_865 ();
 FILLCELL_X32 FILLER_141_897 ();
 FILLCELL_X32 FILLER_141_929 ();
 FILLCELL_X32 FILLER_141_961 ();
 FILLCELL_X32 FILLER_141_993 ();
 FILLCELL_X32 FILLER_141_1025 ();
 FILLCELL_X32 FILLER_141_1057 ();
 FILLCELL_X32 FILLER_141_1089 ();
 FILLCELL_X32 FILLER_141_1121 ();
 FILLCELL_X32 FILLER_141_1153 ();
 FILLCELL_X32 FILLER_141_1185 ();
 FILLCELL_X32 FILLER_141_1217 ();
 FILLCELL_X8 FILLER_141_1249 ();
 FILLCELL_X4 FILLER_141_1257 ();
 FILLCELL_X2 FILLER_141_1261 ();
 FILLCELL_X32 FILLER_141_1264 ();
 FILLCELL_X32 FILLER_141_1296 ();
 FILLCELL_X32 FILLER_141_1328 ();
 FILLCELL_X32 FILLER_141_1360 ();
 FILLCELL_X32 FILLER_141_1392 ();
 FILLCELL_X32 FILLER_141_1424 ();
 FILLCELL_X32 FILLER_141_1456 ();
 FILLCELL_X32 FILLER_141_1488 ();
 FILLCELL_X32 FILLER_141_1520 ();
 FILLCELL_X32 FILLER_141_1552 ();
 FILLCELL_X32 FILLER_141_1584 ();
 FILLCELL_X32 FILLER_141_1616 ();
 FILLCELL_X32 FILLER_141_1648 ();
 FILLCELL_X32 FILLER_141_1680 ();
 FILLCELL_X32 FILLER_141_1712 ();
 FILLCELL_X32 FILLER_141_1744 ();
 FILLCELL_X32 FILLER_141_1776 ();
 FILLCELL_X32 FILLER_141_1808 ();
 FILLCELL_X32 FILLER_141_1840 ();
 FILLCELL_X32 FILLER_141_1872 ();
 FILLCELL_X32 FILLER_141_1904 ();
 FILLCELL_X32 FILLER_141_1936 ();
 FILLCELL_X32 FILLER_141_1968 ();
 FILLCELL_X32 FILLER_141_2000 ();
 FILLCELL_X32 FILLER_141_2032 ();
 FILLCELL_X32 FILLER_141_2064 ();
 FILLCELL_X32 FILLER_141_2096 ();
 FILLCELL_X32 FILLER_141_2128 ();
 FILLCELL_X32 FILLER_141_2160 ();
 FILLCELL_X32 FILLER_141_2192 ();
 FILLCELL_X32 FILLER_141_2224 ();
 FILLCELL_X32 FILLER_141_2256 ();
 FILLCELL_X32 FILLER_141_2288 ();
 FILLCELL_X32 FILLER_141_2320 ();
 FILLCELL_X32 FILLER_141_2352 ();
 FILLCELL_X32 FILLER_141_2384 ();
 FILLCELL_X32 FILLER_141_2416 ();
 FILLCELL_X32 FILLER_141_2448 ();
 FILLCELL_X32 FILLER_141_2480 ();
 FILLCELL_X8 FILLER_141_2512 ();
 FILLCELL_X4 FILLER_141_2520 ();
 FILLCELL_X2 FILLER_141_2524 ();
 FILLCELL_X32 FILLER_141_2527 ();
 FILLCELL_X32 FILLER_141_2559 ();
 FILLCELL_X32 FILLER_141_2591 ();
 FILLCELL_X32 FILLER_141_2623 ();
 FILLCELL_X32 FILLER_141_2655 ();
 FILLCELL_X32 FILLER_141_2687 ();
 FILLCELL_X32 FILLER_141_2719 ();
 FILLCELL_X32 FILLER_141_2751 ();
 FILLCELL_X32 FILLER_141_2783 ();
 FILLCELL_X32 FILLER_141_2815 ();
 FILLCELL_X32 FILLER_141_2847 ();
 FILLCELL_X32 FILLER_141_2879 ();
 FILLCELL_X32 FILLER_141_2911 ();
 FILLCELL_X32 FILLER_141_2943 ();
 FILLCELL_X32 FILLER_141_2975 ();
 FILLCELL_X32 FILLER_141_3007 ();
 FILLCELL_X32 FILLER_141_3039 ();
 FILLCELL_X32 FILLER_141_3071 ();
 FILLCELL_X32 FILLER_141_3103 ();
 FILLCELL_X32 FILLER_141_3135 ();
 FILLCELL_X32 FILLER_141_3167 ();
 FILLCELL_X32 FILLER_141_3199 ();
 FILLCELL_X32 FILLER_141_3231 ();
 FILLCELL_X32 FILLER_141_3263 ();
 FILLCELL_X32 FILLER_141_3295 ();
 FILLCELL_X32 FILLER_141_3327 ();
 FILLCELL_X32 FILLER_141_3359 ();
 FILLCELL_X32 FILLER_141_3391 ();
 FILLCELL_X32 FILLER_141_3423 ();
 FILLCELL_X32 FILLER_141_3455 ();
 FILLCELL_X32 FILLER_141_3487 ();
 FILLCELL_X32 FILLER_141_3519 ();
 FILLCELL_X32 FILLER_141_3551 ();
 FILLCELL_X32 FILLER_141_3583 ();
 FILLCELL_X32 FILLER_141_3615 ();
 FILLCELL_X32 FILLER_141_3647 ();
 FILLCELL_X32 FILLER_141_3679 ();
 FILLCELL_X16 FILLER_141_3711 ();
 FILLCELL_X8 FILLER_141_3727 ();
 FILLCELL_X2 FILLER_141_3735 ();
 FILLCELL_X1 FILLER_141_3737 ();
 FILLCELL_X32 FILLER_142_1 ();
 FILLCELL_X32 FILLER_142_33 ();
 FILLCELL_X32 FILLER_142_65 ();
 FILLCELL_X32 FILLER_142_97 ();
 FILLCELL_X32 FILLER_142_129 ();
 FILLCELL_X32 FILLER_142_161 ();
 FILLCELL_X32 FILLER_142_193 ();
 FILLCELL_X32 FILLER_142_225 ();
 FILLCELL_X32 FILLER_142_257 ();
 FILLCELL_X32 FILLER_142_289 ();
 FILLCELL_X32 FILLER_142_321 ();
 FILLCELL_X32 FILLER_142_353 ();
 FILLCELL_X32 FILLER_142_385 ();
 FILLCELL_X32 FILLER_142_417 ();
 FILLCELL_X32 FILLER_142_449 ();
 FILLCELL_X32 FILLER_142_481 ();
 FILLCELL_X32 FILLER_142_513 ();
 FILLCELL_X32 FILLER_142_545 ();
 FILLCELL_X32 FILLER_142_577 ();
 FILLCELL_X16 FILLER_142_609 ();
 FILLCELL_X4 FILLER_142_625 ();
 FILLCELL_X2 FILLER_142_629 ();
 FILLCELL_X32 FILLER_142_632 ();
 FILLCELL_X32 FILLER_142_664 ();
 FILLCELL_X32 FILLER_142_696 ();
 FILLCELL_X32 FILLER_142_728 ();
 FILLCELL_X32 FILLER_142_760 ();
 FILLCELL_X32 FILLER_142_792 ();
 FILLCELL_X32 FILLER_142_824 ();
 FILLCELL_X32 FILLER_142_856 ();
 FILLCELL_X32 FILLER_142_888 ();
 FILLCELL_X32 FILLER_142_920 ();
 FILLCELL_X32 FILLER_142_952 ();
 FILLCELL_X32 FILLER_142_984 ();
 FILLCELL_X32 FILLER_142_1016 ();
 FILLCELL_X32 FILLER_142_1048 ();
 FILLCELL_X32 FILLER_142_1080 ();
 FILLCELL_X32 FILLER_142_1112 ();
 FILLCELL_X32 FILLER_142_1144 ();
 FILLCELL_X32 FILLER_142_1176 ();
 FILLCELL_X32 FILLER_142_1208 ();
 FILLCELL_X32 FILLER_142_1240 ();
 FILLCELL_X32 FILLER_142_1272 ();
 FILLCELL_X32 FILLER_142_1304 ();
 FILLCELL_X32 FILLER_142_1336 ();
 FILLCELL_X32 FILLER_142_1368 ();
 FILLCELL_X32 FILLER_142_1400 ();
 FILLCELL_X32 FILLER_142_1432 ();
 FILLCELL_X32 FILLER_142_1464 ();
 FILLCELL_X32 FILLER_142_1496 ();
 FILLCELL_X32 FILLER_142_1528 ();
 FILLCELL_X32 FILLER_142_1560 ();
 FILLCELL_X32 FILLER_142_1592 ();
 FILLCELL_X32 FILLER_142_1624 ();
 FILLCELL_X32 FILLER_142_1656 ();
 FILLCELL_X32 FILLER_142_1688 ();
 FILLCELL_X32 FILLER_142_1720 ();
 FILLCELL_X32 FILLER_142_1752 ();
 FILLCELL_X32 FILLER_142_1784 ();
 FILLCELL_X32 FILLER_142_1816 ();
 FILLCELL_X32 FILLER_142_1848 ();
 FILLCELL_X8 FILLER_142_1880 ();
 FILLCELL_X4 FILLER_142_1888 ();
 FILLCELL_X2 FILLER_142_1892 ();
 FILLCELL_X32 FILLER_142_1895 ();
 FILLCELL_X32 FILLER_142_1927 ();
 FILLCELL_X32 FILLER_142_1959 ();
 FILLCELL_X32 FILLER_142_1991 ();
 FILLCELL_X32 FILLER_142_2023 ();
 FILLCELL_X32 FILLER_142_2055 ();
 FILLCELL_X32 FILLER_142_2087 ();
 FILLCELL_X32 FILLER_142_2119 ();
 FILLCELL_X32 FILLER_142_2151 ();
 FILLCELL_X32 FILLER_142_2183 ();
 FILLCELL_X32 FILLER_142_2215 ();
 FILLCELL_X32 FILLER_142_2247 ();
 FILLCELL_X32 FILLER_142_2279 ();
 FILLCELL_X32 FILLER_142_2311 ();
 FILLCELL_X32 FILLER_142_2343 ();
 FILLCELL_X32 FILLER_142_2375 ();
 FILLCELL_X32 FILLER_142_2407 ();
 FILLCELL_X32 FILLER_142_2439 ();
 FILLCELL_X32 FILLER_142_2471 ();
 FILLCELL_X32 FILLER_142_2503 ();
 FILLCELL_X32 FILLER_142_2535 ();
 FILLCELL_X32 FILLER_142_2567 ();
 FILLCELL_X32 FILLER_142_2599 ();
 FILLCELL_X32 FILLER_142_2631 ();
 FILLCELL_X32 FILLER_142_2663 ();
 FILLCELL_X32 FILLER_142_2695 ();
 FILLCELL_X32 FILLER_142_2727 ();
 FILLCELL_X32 FILLER_142_2759 ();
 FILLCELL_X32 FILLER_142_2791 ();
 FILLCELL_X32 FILLER_142_2823 ();
 FILLCELL_X32 FILLER_142_2855 ();
 FILLCELL_X32 FILLER_142_2887 ();
 FILLCELL_X32 FILLER_142_2919 ();
 FILLCELL_X32 FILLER_142_2951 ();
 FILLCELL_X32 FILLER_142_2983 ();
 FILLCELL_X32 FILLER_142_3015 ();
 FILLCELL_X32 FILLER_142_3047 ();
 FILLCELL_X32 FILLER_142_3079 ();
 FILLCELL_X32 FILLER_142_3111 ();
 FILLCELL_X8 FILLER_142_3143 ();
 FILLCELL_X4 FILLER_142_3151 ();
 FILLCELL_X2 FILLER_142_3155 ();
 FILLCELL_X32 FILLER_142_3158 ();
 FILLCELL_X32 FILLER_142_3190 ();
 FILLCELL_X32 FILLER_142_3222 ();
 FILLCELL_X32 FILLER_142_3254 ();
 FILLCELL_X32 FILLER_142_3286 ();
 FILLCELL_X32 FILLER_142_3318 ();
 FILLCELL_X32 FILLER_142_3350 ();
 FILLCELL_X32 FILLER_142_3382 ();
 FILLCELL_X32 FILLER_142_3414 ();
 FILLCELL_X32 FILLER_142_3446 ();
 FILLCELL_X32 FILLER_142_3478 ();
 FILLCELL_X32 FILLER_142_3510 ();
 FILLCELL_X32 FILLER_142_3542 ();
 FILLCELL_X32 FILLER_142_3574 ();
 FILLCELL_X32 FILLER_142_3606 ();
 FILLCELL_X32 FILLER_142_3638 ();
 FILLCELL_X32 FILLER_142_3670 ();
 FILLCELL_X32 FILLER_142_3702 ();
 FILLCELL_X4 FILLER_142_3734 ();
 FILLCELL_X32 FILLER_143_1 ();
 FILLCELL_X32 FILLER_143_33 ();
 FILLCELL_X32 FILLER_143_65 ();
 FILLCELL_X32 FILLER_143_97 ();
 FILLCELL_X32 FILLER_143_129 ();
 FILLCELL_X32 FILLER_143_161 ();
 FILLCELL_X32 FILLER_143_193 ();
 FILLCELL_X32 FILLER_143_225 ();
 FILLCELL_X32 FILLER_143_257 ();
 FILLCELL_X32 FILLER_143_289 ();
 FILLCELL_X32 FILLER_143_321 ();
 FILLCELL_X32 FILLER_143_353 ();
 FILLCELL_X32 FILLER_143_385 ();
 FILLCELL_X32 FILLER_143_417 ();
 FILLCELL_X32 FILLER_143_449 ();
 FILLCELL_X32 FILLER_143_481 ();
 FILLCELL_X32 FILLER_143_513 ();
 FILLCELL_X32 FILLER_143_545 ();
 FILLCELL_X32 FILLER_143_577 ();
 FILLCELL_X32 FILLER_143_609 ();
 FILLCELL_X32 FILLER_143_641 ();
 FILLCELL_X32 FILLER_143_673 ();
 FILLCELL_X32 FILLER_143_705 ();
 FILLCELL_X32 FILLER_143_737 ();
 FILLCELL_X32 FILLER_143_769 ();
 FILLCELL_X32 FILLER_143_801 ();
 FILLCELL_X32 FILLER_143_833 ();
 FILLCELL_X32 FILLER_143_865 ();
 FILLCELL_X32 FILLER_143_897 ();
 FILLCELL_X32 FILLER_143_929 ();
 FILLCELL_X32 FILLER_143_961 ();
 FILLCELL_X32 FILLER_143_993 ();
 FILLCELL_X32 FILLER_143_1025 ();
 FILLCELL_X32 FILLER_143_1057 ();
 FILLCELL_X32 FILLER_143_1089 ();
 FILLCELL_X32 FILLER_143_1121 ();
 FILLCELL_X32 FILLER_143_1153 ();
 FILLCELL_X32 FILLER_143_1185 ();
 FILLCELL_X32 FILLER_143_1217 ();
 FILLCELL_X8 FILLER_143_1249 ();
 FILLCELL_X4 FILLER_143_1257 ();
 FILLCELL_X2 FILLER_143_1261 ();
 FILLCELL_X32 FILLER_143_1264 ();
 FILLCELL_X32 FILLER_143_1296 ();
 FILLCELL_X32 FILLER_143_1328 ();
 FILLCELL_X32 FILLER_143_1360 ();
 FILLCELL_X32 FILLER_143_1392 ();
 FILLCELL_X32 FILLER_143_1424 ();
 FILLCELL_X32 FILLER_143_1456 ();
 FILLCELL_X32 FILLER_143_1488 ();
 FILLCELL_X32 FILLER_143_1520 ();
 FILLCELL_X32 FILLER_143_1552 ();
 FILLCELL_X32 FILLER_143_1584 ();
 FILLCELL_X32 FILLER_143_1616 ();
 FILLCELL_X32 FILLER_143_1648 ();
 FILLCELL_X32 FILLER_143_1680 ();
 FILLCELL_X32 FILLER_143_1712 ();
 FILLCELL_X32 FILLER_143_1744 ();
 FILLCELL_X32 FILLER_143_1776 ();
 FILLCELL_X32 FILLER_143_1808 ();
 FILLCELL_X32 FILLER_143_1840 ();
 FILLCELL_X32 FILLER_143_1872 ();
 FILLCELL_X32 FILLER_143_1904 ();
 FILLCELL_X32 FILLER_143_1936 ();
 FILLCELL_X32 FILLER_143_1968 ();
 FILLCELL_X32 FILLER_143_2000 ();
 FILLCELL_X32 FILLER_143_2032 ();
 FILLCELL_X32 FILLER_143_2064 ();
 FILLCELL_X32 FILLER_143_2096 ();
 FILLCELL_X32 FILLER_143_2128 ();
 FILLCELL_X32 FILLER_143_2160 ();
 FILLCELL_X32 FILLER_143_2192 ();
 FILLCELL_X32 FILLER_143_2224 ();
 FILLCELL_X32 FILLER_143_2256 ();
 FILLCELL_X32 FILLER_143_2288 ();
 FILLCELL_X32 FILLER_143_2320 ();
 FILLCELL_X32 FILLER_143_2352 ();
 FILLCELL_X32 FILLER_143_2384 ();
 FILLCELL_X32 FILLER_143_2416 ();
 FILLCELL_X32 FILLER_143_2448 ();
 FILLCELL_X32 FILLER_143_2480 ();
 FILLCELL_X8 FILLER_143_2512 ();
 FILLCELL_X4 FILLER_143_2520 ();
 FILLCELL_X2 FILLER_143_2524 ();
 FILLCELL_X32 FILLER_143_2527 ();
 FILLCELL_X32 FILLER_143_2559 ();
 FILLCELL_X32 FILLER_143_2591 ();
 FILLCELL_X32 FILLER_143_2623 ();
 FILLCELL_X32 FILLER_143_2655 ();
 FILLCELL_X32 FILLER_143_2687 ();
 FILLCELL_X32 FILLER_143_2719 ();
 FILLCELL_X32 FILLER_143_2751 ();
 FILLCELL_X32 FILLER_143_2783 ();
 FILLCELL_X32 FILLER_143_2815 ();
 FILLCELL_X32 FILLER_143_2847 ();
 FILLCELL_X32 FILLER_143_2879 ();
 FILLCELL_X32 FILLER_143_2911 ();
 FILLCELL_X32 FILLER_143_2943 ();
 FILLCELL_X32 FILLER_143_2975 ();
 FILLCELL_X32 FILLER_143_3007 ();
 FILLCELL_X32 FILLER_143_3039 ();
 FILLCELL_X32 FILLER_143_3071 ();
 FILLCELL_X32 FILLER_143_3103 ();
 FILLCELL_X32 FILLER_143_3135 ();
 FILLCELL_X32 FILLER_143_3167 ();
 FILLCELL_X32 FILLER_143_3199 ();
 FILLCELL_X32 FILLER_143_3231 ();
 FILLCELL_X32 FILLER_143_3263 ();
 FILLCELL_X32 FILLER_143_3295 ();
 FILLCELL_X32 FILLER_143_3327 ();
 FILLCELL_X32 FILLER_143_3359 ();
 FILLCELL_X32 FILLER_143_3391 ();
 FILLCELL_X32 FILLER_143_3423 ();
 FILLCELL_X32 FILLER_143_3455 ();
 FILLCELL_X32 FILLER_143_3487 ();
 FILLCELL_X32 FILLER_143_3519 ();
 FILLCELL_X32 FILLER_143_3551 ();
 FILLCELL_X32 FILLER_143_3583 ();
 FILLCELL_X32 FILLER_143_3615 ();
 FILLCELL_X32 FILLER_143_3647 ();
 FILLCELL_X32 FILLER_143_3679 ();
 FILLCELL_X16 FILLER_143_3711 ();
 FILLCELL_X8 FILLER_143_3727 ();
 FILLCELL_X2 FILLER_143_3735 ();
 FILLCELL_X1 FILLER_143_3737 ();
 FILLCELL_X32 FILLER_144_1 ();
 FILLCELL_X32 FILLER_144_33 ();
 FILLCELL_X32 FILLER_144_65 ();
 FILLCELL_X32 FILLER_144_97 ();
 FILLCELL_X32 FILLER_144_129 ();
 FILLCELL_X32 FILLER_144_161 ();
 FILLCELL_X32 FILLER_144_193 ();
 FILLCELL_X32 FILLER_144_225 ();
 FILLCELL_X32 FILLER_144_257 ();
 FILLCELL_X32 FILLER_144_289 ();
 FILLCELL_X32 FILLER_144_321 ();
 FILLCELL_X32 FILLER_144_353 ();
 FILLCELL_X32 FILLER_144_385 ();
 FILLCELL_X32 FILLER_144_417 ();
 FILLCELL_X32 FILLER_144_449 ();
 FILLCELL_X32 FILLER_144_481 ();
 FILLCELL_X32 FILLER_144_513 ();
 FILLCELL_X32 FILLER_144_545 ();
 FILLCELL_X32 FILLER_144_577 ();
 FILLCELL_X16 FILLER_144_609 ();
 FILLCELL_X4 FILLER_144_625 ();
 FILLCELL_X2 FILLER_144_629 ();
 FILLCELL_X32 FILLER_144_632 ();
 FILLCELL_X32 FILLER_144_664 ();
 FILLCELL_X32 FILLER_144_696 ();
 FILLCELL_X32 FILLER_144_728 ();
 FILLCELL_X32 FILLER_144_760 ();
 FILLCELL_X32 FILLER_144_792 ();
 FILLCELL_X32 FILLER_144_824 ();
 FILLCELL_X32 FILLER_144_856 ();
 FILLCELL_X32 FILLER_144_888 ();
 FILLCELL_X32 FILLER_144_920 ();
 FILLCELL_X32 FILLER_144_952 ();
 FILLCELL_X32 FILLER_144_984 ();
 FILLCELL_X32 FILLER_144_1016 ();
 FILLCELL_X32 FILLER_144_1048 ();
 FILLCELL_X32 FILLER_144_1080 ();
 FILLCELL_X32 FILLER_144_1112 ();
 FILLCELL_X32 FILLER_144_1144 ();
 FILLCELL_X32 FILLER_144_1176 ();
 FILLCELL_X32 FILLER_144_1208 ();
 FILLCELL_X32 FILLER_144_1240 ();
 FILLCELL_X32 FILLER_144_1272 ();
 FILLCELL_X32 FILLER_144_1304 ();
 FILLCELL_X32 FILLER_144_1336 ();
 FILLCELL_X32 FILLER_144_1368 ();
 FILLCELL_X32 FILLER_144_1400 ();
 FILLCELL_X32 FILLER_144_1432 ();
 FILLCELL_X32 FILLER_144_1464 ();
 FILLCELL_X32 FILLER_144_1496 ();
 FILLCELL_X32 FILLER_144_1528 ();
 FILLCELL_X32 FILLER_144_1560 ();
 FILLCELL_X32 FILLER_144_1592 ();
 FILLCELL_X32 FILLER_144_1624 ();
 FILLCELL_X32 FILLER_144_1656 ();
 FILLCELL_X32 FILLER_144_1688 ();
 FILLCELL_X32 FILLER_144_1720 ();
 FILLCELL_X32 FILLER_144_1752 ();
 FILLCELL_X32 FILLER_144_1784 ();
 FILLCELL_X32 FILLER_144_1816 ();
 FILLCELL_X32 FILLER_144_1848 ();
 FILLCELL_X8 FILLER_144_1880 ();
 FILLCELL_X4 FILLER_144_1888 ();
 FILLCELL_X2 FILLER_144_1892 ();
 FILLCELL_X32 FILLER_144_1895 ();
 FILLCELL_X32 FILLER_144_1927 ();
 FILLCELL_X32 FILLER_144_1959 ();
 FILLCELL_X32 FILLER_144_1991 ();
 FILLCELL_X32 FILLER_144_2023 ();
 FILLCELL_X32 FILLER_144_2055 ();
 FILLCELL_X32 FILLER_144_2087 ();
 FILLCELL_X32 FILLER_144_2119 ();
 FILLCELL_X32 FILLER_144_2151 ();
 FILLCELL_X32 FILLER_144_2183 ();
 FILLCELL_X32 FILLER_144_2215 ();
 FILLCELL_X32 FILLER_144_2247 ();
 FILLCELL_X32 FILLER_144_2279 ();
 FILLCELL_X32 FILLER_144_2311 ();
 FILLCELL_X32 FILLER_144_2343 ();
 FILLCELL_X32 FILLER_144_2375 ();
 FILLCELL_X32 FILLER_144_2407 ();
 FILLCELL_X32 FILLER_144_2439 ();
 FILLCELL_X32 FILLER_144_2471 ();
 FILLCELL_X32 FILLER_144_2503 ();
 FILLCELL_X32 FILLER_144_2535 ();
 FILLCELL_X32 FILLER_144_2567 ();
 FILLCELL_X32 FILLER_144_2599 ();
 FILLCELL_X32 FILLER_144_2631 ();
 FILLCELL_X32 FILLER_144_2663 ();
 FILLCELL_X32 FILLER_144_2695 ();
 FILLCELL_X32 FILLER_144_2727 ();
 FILLCELL_X32 FILLER_144_2759 ();
 FILLCELL_X32 FILLER_144_2791 ();
 FILLCELL_X32 FILLER_144_2823 ();
 FILLCELL_X32 FILLER_144_2855 ();
 FILLCELL_X32 FILLER_144_2887 ();
 FILLCELL_X32 FILLER_144_2919 ();
 FILLCELL_X32 FILLER_144_2951 ();
 FILLCELL_X32 FILLER_144_2983 ();
 FILLCELL_X32 FILLER_144_3015 ();
 FILLCELL_X32 FILLER_144_3047 ();
 FILLCELL_X32 FILLER_144_3079 ();
 FILLCELL_X32 FILLER_144_3111 ();
 FILLCELL_X8 FILLER_144_3143 ();
 FILLCELL_X4 FILLER_144_3151 ();
 FILLCELL_X2 FILLER_144_3155 ();
 FILLCELL_X32 FILLER_144_3158 ();
 FILLCELL_X32 FILLER_144_3190 ();
 FILLCELL_X32 FILLER_144_3222 ();
 FILLCELL_X32 FILLER_144_3254 ();
 FILLCELL_X32 FILLER_144_3286 ();
 FILLCELL_X32 FILLER_144_3318 ();
 FILLCELL_X32 FILLER_144_3350 ();
 FILLCELL_X32 FILLER_144_3382 ();
 FILLCELL_X32 FILLER_144_3414 ();
 FILLCELL_X32 FILLER_144_3446 ();
 FILLCELL_X32 FILLER_144_3478 ();
 FILLCELL_X32 FILLER_144_3510 ();
 FILLCELL_X32 FILLER_144_3542 ();
 FILLCELL_X32 FILLER_144_3574 ();
 FILLCELL_X32 FILLER_144_3606 ();
 FILLCELL_X32 FILLER_144_3638 ();
 FILLCELL_X32 FILLER_144_3670 ();
 FILLCELL_X32 FILLER_144_3702 ();
 FILLCELL_X4 FILLER_144_3734 ();
 FILLCELL_X32 FILLER_145_1 ();
 FILLCELL_X32 FILLER_145_33 ();
 FILLCELL_X32 FILLER_145_65 ();
 FILLCELL_X32 FILLER_145_97 ();
 FILLCELL_X32 FILLER_145_129 ();
 FILLCELL_X32 FILLER_145_161 ();
 FILLCELL_X32 FILLER_145_193 ();
 FILLCELL_X32 FILLER_145_225 ();
 FILLCELL_X32 FILLER_145_257 ();
 FILLCELL_X32 FILLER_145_289 ();
 FILLCELL_X32 FILLER_145_321 ();
 FILLCELL_X32 FILLER_145_353 ();
 FILLCELL_X32 FILLER_145_385 ();
 FILLCELL_X32 FILLER_145_417 ();
 FILLCELL_X32 FILLER_145_449 ();
 FILLCELL_X32 FILLER_145_481 ();
 FILLCELL_X32 FILLER_145_513 ();
 FILLCELL_X32 FILLER_145_545 ();
 FILLCELL_X32 FILLER_145_577 ();
 FILLCELL_X32 FILLER_145_609 ();
 FILLCELL_X32 FILLER_145_641 ();
 FILLCELL_X32 FILLER_145_673 ();
 FILLCELL_X32 FILLER_145_705 ();
 FILLCELL_X32 FILLER_145_737 ();
 FILLCELL_X32 FILLER_145_769 ();
 FILLCELL_X32 FILLER_145_801 ();
 FILLCELL_X32 FILLER_145_833 ();
 FILLCELL_X32 FILLER_145_865 ();
 FILLCELL_X32 FILLER_145_897 ();
 FILLCELL_X32 FILLER_145_929 ();
 FILLCELL_X32 FILLER_145_961 ();
 FILLCELL_X32 FILLER_145_993 ();
 FILLCELL_X32 FILLER_145_1025 ();
 FILLCELL_X32 FILLER_145_1057 ();
 FILLCELL_X32 FILLER_145_1089 ();
 FILLCELL_X32 FILLER_145_1121 ();
 FILLCELL_X32 FILLER_145_1153 ();
 FILLCELL_X32 FILLER_145_1185 ();
 FILLCELL_X32 FILLER_145_1217 ();
 FILLCELL_X8 FILLER_145_1249 ();
 FILLCELL_X4 FILLER_145_1257 ();
 FILLCELL_X2 FILLER_145_1261 ();
 FILLCELL_X32 FILLER_145_1264 ();
 FILLCELL_X32 FILLER_145_1296 ();
 FILLCELL_X32 FILLER_145_1328 ();
 FILLCELL_X32 FILLER_145_1360 ();
 FILLCELL_X32 FILLER_145_1392 ();
 FILLCELL_X32 FILLER_145_1424 ();
 FILLCELL_X32 FILLER_145_1456 ();
 FILLCELL_X32 FILLER_145_1488 ();
 FILLCELL_X32 FILLER_145_1520 ();
 FILLCELL_X32 FILLER_145_1552 ();
 FILLCELL_X32 FILLER_145_1584 ();
 FILLCELL_X32 FILLER_145_1616 ();
 FILLCELL_X32 FILLER_145_1648 ();
 FILLCELL_X32 FILLER_145_1680 ();
 FILLCELL_X32 FILLER_145_1712 ();
 FILLCELL_X32 FILLER_145_1744 ();
 FILLCELL_X32 FILLER_145_1776 ();
 FILLCELL_X32 FILLER_145_1808 ();
 FILLCELL_X32 FILLER_145_1840 ();
 FILLCELL_X32 FILLER_145_1872 ();
 FILLCELL_X32 FILLER_145_1904 ();
 FILLCELL_X32 FILLER_145_1936 ();
 FILLCELL_X32 FILLER_145_1968 ();
 FILLCELL_X32 FILLER_145_2000 ();
 FILLCELL_X32 FILLER_145_2032 ();
 FILLCELL_X32 FILLER_145_2064 ();
 FILLCELL_X32 FILLER_145_2096 ();
 FILLCELL_X32 FILLER_145_2128 ();
 FILLCELL_X32 FILLER_145_2160 ();
 FILLCELL_X32 FILLER_145_2192 ();
 FILLCELL_X32 FILLER_145_2224 ();
 FILLCELL_X32 FILLER_145_2256 ();
 FILLCELL_X32 FILLER_145_2288 ();
 FILLCELL_X32 FILLER_145_2320 ();
 FILLCELL_X32 FILLER_145_2352 ();
 FILLCELL_X32 FILLER_145_2384 ();
 FILLCELL_X32 FILLER_145_2416 ();
 FILLCELL_X32 FILLER_145_2448 ();
 FILLCELL_X32 FILLER_145_2480 ();
 FILLCELL_X8 FILLER_145_2512 ();
 FILLCELL_X4 FILLER_145_2520 ();
 FILLCELL_X2 FILLER_145_2524 ();
 FILLCELL_X32 FILLER_145_2527 ();
 FILLCELL_X32 FILLER_145_2559 ();
 FILLCELL_X32 FILLER_145_2591 ();
 FILLCELL_X32 FILLER_145_2623 ();
 FILLCELL_X32 FILLER_145_2655 ();
 FILLCELL_X32 FILLER_145_2687 ();
 FILLCELL_X32 FILLER_145_2719 ();
 FILLCELL_X32 FILLER_145_2751 ();
 FILLCELL_X32 FILLER_145_2783 ();
 FILLCELL_X32 FILLER_145_2815 ();
 FILLCELL_X32 FILLER_145_2847 ();
 FILLCELL_X32 FILLER_145_2879 ();
 FILLCELL_X32 FILLER_145_2911 ();
 FILLCELL_X32 FILLER_145_2943 ();
 FILLCELL_X32 FILLER_145_2975 ();
 FILLCELL_X32 FILLER_145_3007 ();
 FILLCELL_X32 FILLER_145_3039 ();
 FILLCELL_X32 FILLER_145_3071 ();
 FILLCELL_X32 FILLER_145_3103 ();
 FILLCELL_X32 FILLER_145_3135 ();
 FILLCELL_X32 FILLER_145_3167 ();
 FILLCELL_X32 FILLER_145_3199 ();
 FILLCELL_X32 FILLER_145_3231 ();
 FILLCELL_X32 FILLER_145_3263 ();
 FILLCELL_X32 FILLER_145_3295 ();
 FILLCELL_X32 FILLER_145_3327 ();
 FILLCELL_X32 FILLER_145_3359 ();
 FILLCELL_X32 FILLER_145_3391 ();
 FILLCELL_X32 FILLER_145_3423 ();
 FILLCELL_X32 FILLER_145_3455 ();
 FILLCELL_X32 FILLER_145_3487 ();
 FILLCELL_X32 FILLER_145_3519 ();
 FILLCELL_X32 FILLER_145_3551 ();
 FILLCELL_X32 FILLER_145_3583 ();
 FILLCELL_X32 FILLER_145_3615 ();
 FILLCELL_X32 FILLER_145_3647 ();
 FILLCELL_X32 FILLER_145_3679 ();
 FILLCELL_X16 FILLER_145_3711 ();
 FILLCELL_X8 FILLER_145_3727 ();
 FILLCELL_X2 FILLER_145_3735 ();
 FILLCELL_X1 FILLER_145_3737 ();
 FILLCELL_X32 FILLER_146_1 ();
 FILLCELL_X32 FILLER_146_33 ();
 FILLCELL_X32 FILLER_146_65 ();
 FILLCELL_X32 FILLER_146_97 ();
 FILLCELL_X32 FILLER_146_129 ();
 FILLCELL_X32 FILLER_146_161 ();
 FILLCELL_X32 FILLER_146_193 ();
 FILLCELL_X32 FILLER_146_225 ();
 FILLCELL_X32 FILLER_146_257 ();
 FILLCELL_X32 FILLER_146_289 ();
 FILLCELL_X32 FILLER_146_321 ();
 FILLCELL_X32 FILLER_146_353 ();
 FILLCELL_X32 FILLER_146_385 ();
 FILLCELL_X32 FILLER_146_417 ();
 FILLCELL_X32 FILLER_146_449 ();
 FILLCELL_X32 FILLER_146_481 ();
 FILLCELL_X32 FILLER_146_513 ();
 FILLCELL_X32 FILLER_146_545 ();
 FILLCELL_X32 FILLER_146_577 ();
 FILLCELL_X16 FILLER_146_609 ();
 FILLCELL_X4 FILLER_146_625 ();
 FILLCELL_X2 FILLER_146_629 ();
 FILLCELL_X32 FILLER_146_632 ();
 FILLCELL_X32 FILLER_146_664 ();
 FILLCELL_X32 FILLER_146_696 ();
 FILLCELL_X32 FILLER_146_728 ();
 FILLCELL_X32 FILLER_146_760 ();
 FILLCELL_X32 FILLER_146_792 ();
 FILLCELL_X32 FILLER_146_824 ();
 FILLCELL_X32 FILLER_146_856 ();
 FILLCELL_X32 FILLER_146_888 ();
 FILLCELL_X32 FILLER_146_920 ();
 FILLCELL_X32 FILLER_146_952 ();
 FILLCELL_X32 FILLER_146_984 ();
 FILLCELL_X32 FILLER_146_1016 ();
 FILLCELL_X32 FILLER_146_1048 ();
 FILLCELL_X32 FILLER_146_1080 ();
 FILLCELL_X32 FILLER_146_1112 ();
 FILLCELL_X32 FILLER_146_1144 ();
 FILLCELL_X32 FILLER_146_1176 ();
 FILLCELL_X32 FILLER_146_1208 ();
 FILLCELL_X32 FILLER_146_1240 ();
 FILLCELL_X32 FILLER_146_1272 ();
 FILLCELL_X32 FILLER_146_1304 ();
 FILLCELL_X32 FILLER_146_1336 ();
 FILLCELL_X32 FILLER_146_1368 ();
 FILLCELL_X32 FILLER_146_1400 ();
 FILLCELL_X32 FILLER_146_1432 ();
 FILLCELL_X32 FILLER_146_1464 ();
 FILLCELL_X32 FILLER_146_1496 ();
 FILLCELL_X32 FILLER_146_1528 ();
 FILLCELL_X32 FILLER_146_1560 ();
 FILLCELL_X32 FILLER_146_1592 ();
 FILLCELL_X32 FILLER_146_1624 ();
 FILLCELL_X32 FILLER_146_1656 ();
 FILLCELL_X32 FILLER_146_1688 ();
 FILLCELL_X32 FILLER_146_1720 ();
 FILLCELL_X32 FILLER_146_1752 ();
 FILLCELL_X32 FILLER_146_1784 ();
 FILLCELL_X32 FILLER_146_1816 ();
 FILLCELL_X32 FILLER_146_1848 ();
 FILLCELL_X8 FILLER_146_1880 ();
 FILLCELL_X4 FILLER_146_1888 ();
 FILLCELL_X2 FILLER_146_1892 ();
 FILLCELL_X32 FILLER_146_1895 ();
 FILLCELL_X32 FILLER_146_1927 ();
 FILLCELL_X32 FILLER_146_1959 ();
 FILLCELL_X32 FILLER_146_1991 ();
 FILLCELL_X32 FILLER_146_2023 ();
 FILLCELL_X32 FILLER_146_2055 ();
 FILLCELL_X32 FILLER_146_2087 ();
 FILLCELL_X32 FILLER_146_2119 ();
 FILLCELL_X32 FILLER_146_2151 ();
 FILLCELL_X32 FILLER_146_2183 ();
 FILLCELL_X32 FILLER_146_2215 ();
 FILLCELL_X32 FILLER_146_2247 ();
 FILLCELL_X32 FILLER_146_2279 ();
 FILLCELL_X32 FILLER_146_2311 ();
 FILLCELL_X32 FILLER_146_2343 ();
 FILLCELL_X32 FILLER_146_2375 ();
 FILLCELL_X32 FILLER_146_2407 ();
 FILLCELL_X32 FILLER_146_2439 ();
 FILLCELL_X32 FILLER_146_2471 ();
 FILLCELL_X32 FILLER_146_2503 ();
 FILLCELL_X32 FILLER_146_2535 ();
 FILLCELL_X32 FILLER_146_2567 ();
 FILLCELL_X32 FILLER_146_2599 ();
 FILLCELL_X32 FILLER_146_2631 ();
 FILLCELL_X32 FILLER_146_2663 ();
 FILLCELL_X32 FILLER_146_2695 ();
 FILLCELL_X32 FILLER_146_2727 ();
 FILLCELL_X32 FILLER_146_2759 ();
 FILLCELL_X32 FILLER_146_2791 ();
 FILLCELL_X32 FILLER_146_2823 ();
 FILLCELL_X32 FILLER_146_2855 ();
 FILLCELL_X32 FILLER_146_2887 ();
 FILLCELL_X32 FILLER_146_2919 ();
 FILLCELL_X32 FILLER_146_2951 ();
 FILLCELL_X32 FILLER_146_2983 ();
 FILLCELL_X32 FILLER_146_3015 ();
 FILLCELL_X32 FILLER_146_3047 ();
 FILLCELL_X32 FILLER_146_3079 ();
 FILLCELL_X32 FILLER_146_3111 ();
 FILLCELL_X8 FILLER_146_3143 ();
 FILLCELL_X4 FILLER_146_3151 ();
 FILLCELL_X2 FILLER_146_3155 ();
 FILLCELL_X32 FILLER_146_3158 ();
 FILLCELL_X32 FILLER_146_3190 ();
 FILLCELL_X32 FILLER_146_3222 ();
 FILLCELL_X32 FILLER_146_3254 ();
 FILLCELL_X32 FILLER_146_3286 ();
 FILLCELL_X32 FILLER_146_3318 ();
 FILLCELL_X32 FILLER_146_3350 ();
 FILLCELL_X32 FILLER_146_3382 ();
 FILLCELL_X32 FILLER_146_3414 ();
 FILLCELL_X32 FILLER_146_3446 ();
 FILLCELL_X32 FILLER_146_3478 ();
 FILLCELL_X32 FILLER_146_3510 ();
 FILLCELL_X32 FILLER_146_3542 ();
 FILLCELL_X32 FILLER_146_3574 ();
 FILLCELL_X32 FILLER_146_3606 ();
 FILLCELL_X32 FILLER_146_3638 ();
 FILLCELL_X32 FILLER_146_3670 ();
 FILLCELL_X32 FILLER_146_3702 ();
 FILLCELL_X4 FILLER_146_3734 ();
 FILLCELL_X32 FILLER_147_1 ();
 FILLCELL_X32 FILLER_147_33 ();
 FILLCELL_X32 FILLER_147_65 ();
 FILLCELL_X32 FILLER_147_97 ();
 FILLCELL_X32 FILLER_147_129 ();
 FILLCELL_X32 FILLER_147_161 ();
 FILLCELL_X32 FILLER_147_193 ();
 FILLCELL_X32 FILLER_147_225 ();
 FILLCELL_X32 FILLER_147_257 ();
 FILLCELL_X32 FILLER_147_289 ();
 FILLCELL_X32 FILLER_147_321 ();
 FILLCELL_X32 FILLER_147_353 ();
 FILLCELL_X32 FILLER_147_385 ();
 FILLCELL_X32 FILLER_147_417 ();
 FILLCELL_X32 FILLER_147_449 ();
 FILLCELL_X32 FILLER_147_481 ();
 FILLCELL_X32 FILLER_147_513 ();
 FILLCELL_X32 FILLER_147_545 ();
 FILLCELL_X32 FILLER_147_577 ();
 FILLCELL_X32 FILLER_147_609 ();
 FILLCELL_X32 FILLER_147_641 ();
 FILLCELL_X32 FILLER_147_673 ();
 FILLCELL_X32 FILLER_147_705 ();
 FILLCELL_X32 FILLER_147_737 ();
 FILLCELL_X32 FILLER_147_769 ();
 FILLCELL_X32 FILLER_147_801 ();
 FILLCELL_X32 FILLER_147_833 ();
 FILLCELL_X32 FILLER_147_865 ();
 FILLCELL_X32 FILLER_147_897 ();
 FILLCELL_X32 FILLER_147_929 ();
 FILLCELL_X32 FILLER_147_961 ();
 FILLCELL_X32 FILLER_147_993 ();
 FILLCELL_X32 FILLER_147_1025 ();
 FILLCELL_X32 FILLER_147_1057 ();
 FILLCELL_X32 FILLER_147_1089 ();
 FILLCELL_X32 FILLER_147_1121 ();
 FILLCELL_X32 FILLER_147_1153 ();
 FILLCELL_X32 FILLER_147_1185 ();
 FILLCELL_X32 FILLER_147_1217 ();
 FILLCELL_X8 FILLER_147_1249 ();
 FILLCELL_X4 FILLER_147_1257 ();
 FILLCELL_X2 FILLER_147_1261 ();
 FILLCELL_X32 FILLER_147_1264 ();
 FILLCELL_X32 FILLER_147_1296 ();
 FILLCELL_X32 FILLER_147_1328 ();
 FILLCELL_X32 FILLER_147_1360 ();
 FILLCELL_X32 FILLER_147_1392 ();
 FILLCELL_X32 FILLER_147_1424 ();
 FILLCELL_X32 FILLER_147_1456 ();
 FILLCELL_X32 FILLER_147_1488 ();
 FILLCELL_X32 FILLER_147_1520 ();
 FILLCELL_X32 FILLER_147_1552 ();
 FILLCELL_X32 FILLER_147_1584 ();
 FILLCELL_X32 FILLER_147_1616 ();
 FILLCELL_X32 FILLER_147_1648 ();
 FILLCELL_X32 FILLER_147_1680 ();
 FILLCELL_X32 FILLER_147_1712 ();
 FILLCELL_X32 FILLER_147_1744 ();
 FILLCELL_X32 FILLER_147_1776 ();
 FILLCELL_X32 FILLER_147_1808 ();
 FILLCELL_X32 FILLER_147_1840 ();
 FILLCELL_X32 FILLER_147_1872 ();
 FILLCELL_X32 FILLER_147_1904 ();
 FILLCELL_X32 FILLER_147_1936 ();
 FILLCELL_X32 FILLER_147_1968 ();
 FILLCELL_X32 FILLER_147_2000 ();
 FILLCELL_X32 FILLER_147_2032 ();
 FILLCELL_X32 FILLER_147_2064 ();
 FILLCELL_X32 FILLER_147_2096 ();
 FILLCELL_X32 FILLER_147_2128 ();
 FILLCELL_X32 FILLER_147_2160 ();
 FILLCELL_X32 FILLER_147_2192 ();
 FILLCELL_X32 FILLER_147_2224 ();
 FILLCELL_X32 FILLER_147_2256 ();
 FILLCELL_X32 FILLER_147_2288 ();
 FILLCELL_X32 FILLER_147_2320 ();
 FILLCELL_X32 FILLER_147_2352 ();
 FILLCELL_X32 FILLER_147_2384 ();
 FILLCELL_X32 FILLER_147_2416 ();
 FILLCELL_X32 FILLER_147_2448 ();
 FILLCELL_X32 FILLER_147_2480 ();
 FILLCELL_X8 FILLER_147_2512 ();
 FILLCELL_X4 FILLER_147_2520 ();
 FILLCELL_X2 FILLER_147_2524 ();
 FILLCELL_X32 FILLER_147_2527 ();
 FILLCELL_X32 FILLER_147_2559 ();
 FILLCELL_X32 FILLER_147_2591 ();
 FILLCELL_X32 FILLER_147_2623 ();
 FILLCELL_X32 FILLER_147_2655 ();
 FILLCELL_X32 FILLER_147_2687 ();
 FILLCELL_X32 FILLER_147_2719 ();
 FILLCELL_X32 FILLER_147_2751 ();
 FILLCELL_X32 FILLER_147_2783 ();
 FILLCELL_X32 FILLER_147_2815 ();
 FILLCELL_X32 FILLER_147_2847 ();
 FILLCELL_X32 FILLER_147_2879 ();
 FILLCELL_X32 FILLER_147_2911 ();
 FILLCELL_X32 FILLER_147_2943 ();
 FILLCELL_X32 FILLER_147_2975 ();
 FILLCELL_X32 FILLER_147_3007 ();
 FILLCELL_X32 FILLER_147_3039 ();
 FILLCELL_X32 FILLER_147_3071 ();
 FILLCELL_X32 FILLER_147_3103 ();
 FILLCELL_X32 FILLER_147_3135 ();
 FILLCELL_X32 FILLER_147_3167 ();
 FILLCELL_X32 FILLER_147_3199 ();
 FILLCELL_X32 FILLER_147_3231 ();
 FILLCELL_X32 FILLER_147_3263 ();
 FILLCELL_X32 FILLER_147_3295 ();
 FILLCELL_X32 FILLER_147_3327 ();
 FILLCELL_X32 FILLER_147_3359 ();
 FILLCELL_X32 FILLER_147_3391 ();
 FILLCELL_X32 FILLER_147_3423 ();
 FILLCELL_X32 FILLER_147_3455 ();
 FILLCELL_X32 FILLER_147_3487 ();
 FILLCELL_X32 FILLER_147_3519 ();
 FILLCELL_X32 FILLER_147_3551 ();
 FILLCELL_X32 FILLER_147_3583 ();
 FILLCELL_X32 FILLER_147_3615 ();
 FILLCELL_X32 FILLER_147_3647 ();
 FILLCELL_X32 FILLER_147_3679 ();
 FILLCELL_X16 FILLER_147_3711 ();
 FILLCELL_X8 FILLER_147_3727 ();
 FILLCELL_X2 FILLER_147_3735 ();
 FILLCELL_X1 FILLER_147_3737 ();
 FILLCELL_X32 FILLER_148_1 ();
 FILLCELL_X32 FILLER_148_33 ();
 FILLCELL_X32 FILLER_148_65 ();
 FILLCELL_X32 FILLER_148_97 ();
 FILLCELL_X32 FILLER_148_129 ();
 FILLCELL_X32 FILLER_148_161 ();
 FILLCELL_X32 FILLER_148_193 ();
 FILLCELL_X32 FILLER_148_225 ();
 FILLCELL_X32 FILLER_148_257 ();
 FILLCELL_X32 FILLER_148_289 ();
 FILLCELL_X32 FILLER_148_321 ();
 FILLCELL_X32 FILLER_148_353 ();
 FILLCELL_X32 FILLER_148_385 ();
 FILLCELL_X32 FILLER_148_417 ();
 FILLCELL_X32 FILLER_148_449 ();
 FILLCELL_X32 FILLER_148_481 ();
 FILLCELL_X32 FILLER_148_513 ();
 FILLCELL_X32 FILLER_148_545 ();
 FILLCELL_X32 FILLER_148_577 ();
 FILLCELL_X16 FILLER_148_609 ();
 FILLCELL_X4 FILLER_148_625 ();
 FILLCELL_X2 FILLER_148_629 ();
 FILLCELL_X32 FILLER_148_632 ();
 FILLCELL_X32 FILLER_148_664 ();
 FILLCELL_X32 FILLER_148_696 ();
 FILLCELL_X32 FILLER_148_728 ();
 FILLCELL_X32 FILLER_148_760 ();
 FILLCELL_X32 FILLER_148_792 ();
 FILLCELL_X32 FILLER_148_824 ();
 FILLCELL_X32 FILLER_148_856 ();
 FILLCELL_X32 FILLER_148_888 ();
 FILLCELL_X32 FILLER_148_920 ();
 FILLCELL_X32 FILLER_148_952 ();
 FILLCELL_X32 FILLER_148_984 ();
 FILLCELL_X32 FILLER_148_1016 ();
 FILLCELL_X32 FILLER_148_1048 ();
 FILLCELL_X32 FILLER_148_1080 ();
 FILLCELL_X32 FILLER_148_1112 ();
 FILLCELL_X32 FILLER_148_1144 ();
 FILLCELL_X32 FILLER_148_1176 ();
 FILLCELL_X32 FILLER_148_1208 ();
 FILLCELL_X32 FILLER_148_1240 ();
 FILLCELL_X32 FILLER_148_1272 ();
 FILLCELL_X32 FILLER_148_1304 ();
 FILLCELL_X32 FILLER_148_1336 ();
 FILLCELL_X32 FILLER_148_1368 ();
 FILLCELL_X32 FILLER_148_1400 ();
 FILLCELL_X32 FILLER_148_1432 ();
 FILLCELL_X32 FILLER_148_1464 ();
 FILLCELL_X32 FILLER_148_1496 ();
 FILLCELL_X32 FILLER_148_1528 ();
 FILLCELL_X32 FILLER_148_1560 ();
 FILLCELL_X32 FILLER_148_1592 ();
 FILLCELL_X32 FILLER_148_1624 ();
 FILLCELL_X32 FILLER_148_1656 ();
 FILLCELL_X32 FILLER_148_1688 ();
 FILLCELL_X32 FILLER_148_1720 ();
 FILLCELL_X32 FILLER_148_1752 ();
 FILLCELL_X32 FILLER_148_1784 ();
 FILLCELL_X32 FILLER_148_1816 ();
 FILLCELL_X32 FILLER_148_1848 ();
 FILLCELL_X8 FILLER_148_1880 ();
 FILLCELL_X4 FILLER_148_1888 ();
 FILLCELL_X2 FILLER_148_1892 ();
 FILLCELL_X32 FILLER_148_1895 ();
 FILLCELL_X32 FILLER_148_1927 ();
 FILLCELL_X32 FILLER_148_1959 ();
 FILLCELL_X32 FILLER_148_1991 ();
 FILLCELL_X32 FILLER_148_2023 ();
 FILLCELL_X32 FILLER_148_2055 ();
 FILLCELL_X32 FILLER_148_2087 ();
 FILLCELL_X32 FILLER_148_2119 ();
 FILLCELL_X32 FILLER_148_2151 ();
 FILLCELL_X32 FILLER_148_2183 ();
 FILLCELL_X32 FILLER_148_2215 ();
 FILLCELL_X32 FILLER_148_2247 ();
 FILLCELL_X32 FILLER_148_2279 ();
 FILLCELL_X32 FILLER_148_2311 ();
 FILLCELL_X32 FILLER_148_2343 ();
 FILLCELL_X32 FILLER_148_2375 ();
 FILLCELL_X32 FILLER_148_2407 ();
 FILLCELL_X32 FILLER_148_2439 ();
 FILLCELL_X32 FILLER_148_2471 ();
 FILLCELL_X32 FILLER_148_2503 ();
 FILLCELL_X32 FILLER_148_2535 ();
 FILLCELL_X32 FILLER_148_2567 ();
 FILLCELL_X32 FILLER_148_2599 ();
 FILLCELL_X32 FILLER_148_2631 ();
 FILLCELL_X32 FILLER_148_2663 ();
 FILLCELL_X32 FILLER_148_2695 ();
 FILLCELL_X32 FILLER_148_2727 ();
 FILLCELL_X32 FILLER_148_2759 ();
 FILLCELL_X32 FILLER_148_2791 ();
 FILLCELL_X32 FILLER_148_2823 ();
 FILLCELL_X32 FILLER_148_2855 ();
 FILLCELL_X32 FILLER_148_2887 ();
 FILLCELL_X32 FILLER_148_2919 ();
 FILLCELL_X32 FILLER_148_2951 ();
 FILLCELL_X32 FILLER_148_2983 ();
 FILLCELL_X32 FILLER_148_3015 ();
 FILLCELL_X32 FILLER_148_3047 ();
 FILLCELL_X32 FILLER_148_3079 ();
 FILLCELL_X32 FILLER_148_3111 ();
 FILLCELL_X8 FILLER_148_3143 ();
 FILLCELL_X4 FILLER_148_3151 ();
 FILLCELL_X2 FILLER_148_3155 ();
 FILLCELL_X32 FILLER_148_3158 ();
 FILLCELL_X32 FILLER_148_3190 ();
 FILLCELL_X32 FILLER_148_3222 ();
 FILLCELL_X32 FILLER_148_3254 ();
 FILLCELL_X32 FILLER_148_3286 ();
 FILLCELL_X32 FILLER_148_3318 ();
 FILLCELL_X32 FILLER_148_3350 ();
 FILLCELL_X32 FILLER_148_3382 ();
 FILLCELL_X32 FILLER_148_3414 ();
 FILLCELL_X32 FILLER_148_3446 ();
 FILLCELL_X32 FILLER_148_3478 ();
 FILLCELL_X32 FILLER_148_3510 ();
 FILLCELL_X32 FILLER_148_3542 ();
 FILLCELL_X32 FILLER_148_3574 ();
 FILLCELL_X32 FILLER_148_3606 ();
 FILLCELL_X32 FILLER_148_3638 ();
 FILLCELL_X32 FILLER_148_3670 ();
 FILLCELL_X32 FILLER_148_3702 ();
 FILLCELL_X4 FILLER_148_3734 ();
 FILLCELL_X32 FILLER_149_1 ();
 FILLCELL_X32 FILLER_149_33 ();
 FILLCELL_X32 FILLER_149_65 ();
 FILLCELL_X32 FILLER_149_97 ();
 FILLCELL_X32 FILLER_149_129 ();
 FILLCELL_X32 FILLER_149_161 ();
 FILLCELL_X32 FILLER_149_193 ();
 FILLCELL_X32 FILLER_149_225 ();
 FILLCELL_X32 FILLER_149_257 ();
 FILLCELL_X32 FILLER_149_289 ();
 FILLCELL_X32 FILLER_149_321 ();
 FILLCELL_X32 FILLER_149_353 ();
 FILLCELL_X32 FILLER_149_385 ();
 FILLCELL_X32 FILLER_149_417 ();
 FILLCELL_X32 FILLER_149_449 ();
 FILLCELL_X32 FILLER_149_481 ();
 FILLCELL_X32 FILLER_149_513 ();
 FILLCELL_X32 FILLER_149_545 ();
 FILLCELL_X32 FILLER_149_577 ();
 FILLCELL_X32 FILLER_149_609 ();
 FILLCELL_X32 FILLER_149_641 ();
 FILLCELL_X32 FILLER_149_673 ();
 FILLCELL_X32 FILLER_149_705 ();
 FILLCELL_X32 FILLER_149_737 ();
 FILLCELL_X32 FILLER_149_769 ();
 FILLCELL_X32 FILLER_149_801 ();
 FILLCELL_X32 FILLER_149_833 ();
 FILLCELL_X32 FILLER_149_865 ();
 FILLCELL_X32 FILLER_149_897 ();
 FILLCELL_X32 FILLER_149_929 ();
 FILLCELL_X32 FILLER_149_961 ();
 FILLCELL_X32 FILLER_149_993 ();
 FILLCELL_X32 FILLER_149_1025 ();
 FILLCELL_X32 FILLER_149_1057 ();
 FILLCELL_X32 FILLER_149_1089 ();
 FILLCELL_X32 FILLER_149_1121 ();
 FILLCELL_X32 FILLER_149_1153 ();
 FILLCELL_X32 FILLER_149_1185 ();
 FILLCELL_X32 FILLER_149_1217 ();
 FILLCELL_X8 FILLER_149_1249 ();
 FILLCELL_X4 FILLER_149_1257 ();
 FILLCELL_X2 FILLER_149_1261 ();
 FILLCELL_X32 FILLER_149_1264 ();
 FILLCELL_X32 FILLER_149_1296 ();
 FILLCELL_X32 FILLER_149_1328 ();
 FILLCELL_X32 FILLER_149_1360 ();
 FILLCELL_X32 FILLER_149_1392 ();
 FILLCELL_X32 FILLER_149_1424 ();
 FILLCELL_X32 FILLER_149_1456 ();
 FILLCELL_X32 FILLER_149_1488 ();
 FILLCELL_X32 FILLER_149_1520 ();
 FILLCELL_X32 FILLER_149_1552 ();
 FILLCELL_X32 FILLER_149_1584 ();
 FILLCELL_X32 FILLER_149_1616 ();
 FILLCELL_X32 FILLER_149_1648 ();
 FILLCELL_X32 FILLER_149_1680 ();
 FILLCELL_X32 FILLER_149_1712 ();
 FILLCELL_X32 FILLER_149_1744 ();
 FILLCELL_X32 FILLER_149_1776 ();
 FILLCELL_X32 FILLER_149_1808 ();
 FILLCELL_X32 FILLER_149_1840 ();
 FILLCELL_X32 FILLER_149_1872 ();
 FILLCELL_X32 FILLER_149_1904 ();
 FILLCELL_X32 FILLER_149_1936 ();
 FILLCELL_X32 FILLER_149_1968 ();
 FILLCELL_X32 FILLER_149_2000 ();
 FILLCELL_X32 FILLER_149_2032 ();
 FILLCELL_X32 FILLER_149_2064 ();
 FILLCELL_X32 FILLER_149_2096 ();
 FILLCELL_X32 FILLER_149_2128 ();
 FILLCELL_X32 FILLER_149_2160 ();
 FILLCELL_X32 FILLER_149_2192 ();
 FILLCELL_X32 FILLER_149_2224 ();
 FILLCELL_X32 FILLER_149_2256 ();
 FILLCELL_X32 FILLER_149_2288 ();
 FILLCELL_X32 FILLER_149_2320 ();
 FILLCELL_X32 FILLER_149_2352 ();
 FILLCELL_X32 FILLER_149_2384 ();
 FILLCELL_X32 FILLER_149_2416 ();
 FILLCELL_X32 FILLER_149_2448 ();
 FILLCELL_X32 FILLER_149_2480 ();
 FILLCELL_X8 FILLER_149_2512 ();
 FILLCELL_X4 FILLER_149_2520 ();
 FILLCELL_X2 FILLER_149_2524 ();
 FILLCELL_X32 FILLER_149_2527 ();
 FILLCELL_X32 FILLER_149_2559 ();
 FILLCELL_X32 FILLER_149_2591 ();
 FILLCELL_X32 FILLER_149_2623 ();
 FILLCELL_X32 FILLER_149_2655 ();
 FILLCELL_X32 FILLER_149_2687 ();
 FILLCELL_X32 FILLER_149_2719 ();
 FILLCELL_X32 FILLER_149_2751 ();
 FILLCELL_X32 FILLER_149_2783 ();
 FILLCELL_X32 FILLER_149_2815 ();
 FILLCELL_X32 FILLER_149_2847 ();
 FILLCELL_X32 FILLER_149_2879 ();
 FILLCELL_X32 FILLER_149_2911 ();
 FILLCELL_X32 FILLER_149_2943 ();
 FILLCELL_X32 FILLER_149_2975 ();
 FILLCELL_X32 FILLER_149_3007 ();
 FILLCELL_X32 FILLER_149_3039 ();
 FILLCELL_X32 FILLER_149_3071 ();
 FILLCELL_X32 FILLER_149_3103 ();
 FILLCELL_X32 FILLER_149_3135 ();
 FILLCELL_X32 FILLER_149_3167 ();
 FILLCELL_X32 FILLER_149_3199 ();
 FILLCELL_X32 FILLER_149_3231 ();
 FILLCELL_X32 FILLER_149_3263 ();
 FILLCELL_X32 FILLER_149_3295 ();
 FILLCELL_X32 FILLER_149_3327 ();
 FILLCELL_X32 FILLER_149_3359 ();
 FILLCELL_X32 FILLER_149_3391 ();
 FILLCELL_X32 FILLER_149_3423 ();
 FILLCELL_X32 FILLER_149_3455 ();
 FILLCELL_X32 FILLER_149_3487 ();
 FILLCELL_X32 FILLER_149_3519 ();
 FILLCELL_X32 FILLER_149_3551 ();
 FILLCELL_X32 FILLER_149_3583 ();
 FILLCELL_X32 FILLER_149_3615 ();
 FILLCELL_X32 FILLER_149_3647 ();
 FILLCELL_X32 FILLER_149_3679 ();
 FILLCELL_X16 FILLER_149_3711 ();
 FILLCELL_X8 FILLER_149_3727 ();
 FILLCELL_X2 FILLER_149_3735 ();
 FILLCELL_X1 FILLER_149_3737 ();
 FILLCELL_X32 FILLER_150_1 ();
 FILLCELL_X32 FILLER_150_33 ();
 FILLCELL_X32 FILLER_150_65 ();
 FILLCELL_X32 FILLER_150_97 ();
 FILLCELL_X32 FILLER_150_129 ();
 FILLCELL_X32 FILLER_150_161 ();
 FILLCELL_X32 FILLER_150_193 ();
 FILLCELL_X32 FILLER_150_225 ();
 FILLCELL_X32 FILLER_150_257 ();
 FILLCELL_X32 FILLER_150_289 ();
 FILLCELL_X32 FILLER_150_321 ();
 FILLCELL_X32 FILLER_150_353 ();
 FILLCELL_X32 FILLER_150_385 ();
 FILLCELL_X32 FILLER_150_417 ();
 FILLCELL_X32 FILLER_150_449 ();
 FILLCELL_X32 FILLER_150_481 ();
 FILLCELL_X32 FILLER_150_513 ();
 FILLCELL_X32 FILLER_150_545 ();
 FILLCELL_X32 FILLER_150_577 ();
 FILLCELL_X16 FILLER_150_609 ();
 FILLCELL_X4 FILLER_150_625 ();
 FILLCELL_X2 FILLER_150_629 ();
 FILLCELL_X32 FILLER_150_632 ();
 FILLCELL_X32 FILLER_150_664 ();
 FILLCELL_X32 FILLER_150_696 ();
 FILLCELL_X32 FILLER_150_728 ();
 FILLCELL_X32 FILLER_150_760 ();
 FILLCELL_X32 FILLER_150_792 ();
 FILLCELL_X32 FILLER_150_824 ();
 FILLCELL_X32 FILLER_150_856 ();
 FILLCELL_X32 FILLER_150_888 ();
 FILLCELL_X32 FILLER_150_920 ();
 FILLCELL_X32 FILLER_150_952 ();
 FILLCELL_X32 FILLER_150_984 ();
 FILLCELL_X32 FILLER_150_1016 ();
 FILLCELL_X32 FILLER_150_1048 ();
 FILLCELL_X32 FILLER_150_1080 ();
 FILLCELL_X32 FILLER_150_1112 ();
 FILLCELL_X32 FILLER_150_1144 ();
 FILLCELL_X32 FILLER_150_1176 ();
 FILLCELL_X32 FILLER_150_1208 ();
 FILLCELL_X32 FILLER_150_1240 ();
 FILLCELL_X32 FILLER_150_1272 ();
 FILLCELL_X32 FILLER_150_1304 ();
 FILLCELL_X32 FILLER_150_1336 ();
 FILLCELL_X32 FILLER_150_1368 ();
 FILLCELL_X32 FILLER_150_1400 ();
 FILLCELL_X32 FILLER_150_1432 ();
 FILLCELL_X32 FILLER_150_1464 ();
 FILLCELL_X32 FILLER_150_1496 ();
 FILLCELL_X32 FILLER_150_1528 ();
 FILLCELL_X32 FILLER_150_1560 ();
 FILLCELL_X32 FILLER_150_1592 ();
 FILLCELL_X32 FILLER_150_1624 ();
 FILLCELL_X32 FILLER_150_1656 ();
 FILLCELL_X32 FILLER_150_1688 ();
 FILLCELL_X32 FILLER_150_1720 ();
 FILLCELL_X32 FILLER_150_1752 ();
 FILLCELL_X32 FILLER_150_1784 ();
 FILLCELL_X32 FILLER_150_1816 ();
 FILLCELL_X32 FILLER_150_1848 ();
 FILLCELL_X8 FILLER_150_1880 ();
 FILLCELL_X4 FILLER_150_1888 ();
 FILLCELL_X2 FILLER_150_1892 ();
 FILLCELL_X32 FILLER_150_1895 ();
 FILLCELL_X32 FILLER_150_1927 ();
 FILLCELL_X32 FILLER_150_1959 ();
 FILLCELL_X32 FILLER_150_1991 ();
 FILLCELL_X32 FILLER_150_2023 ();
 FILLCELL_X32 FILLER_150_2055 ();
 FILLCELL_X32 FILLER_150_2087 ();
 FILLCELL_X32 FILLER_150_2119 ();
 FILLCELL_X32 FILLER_150_2151 ();
 FILLCELL_X32 FILLER_150_2183 ();
 FILLCELL_X32 FILLER_150_2215 ();
 FILLCELL_X32 FILLER_150_2247 ();
 FILLCELL_X32 FILLER_150_2279 ();
 FILLCELL_X32 FILLER_150_2311 ();
 FILLCELL_X32 FILLER_150_2343 ();
 FILLCELL_X32 FILLER_150_2375 ();
 FILLCELL_X32 FILLER_150_2407 ();
 FILLCELL_X32 FILLER_150_2439 ();
 FILLCELL_X32 FILLER_150_2471 ();
 FILLCELL_X32 FILLER_150_2503 ();
 FILLCELL_X32 FILLER_150_2535 ();
 FILLCELL_X32 FILLER_150_2567 ();
 FILLCELL_X32 FILLER_150_2599 ();
 FILLCELL_X32 FILLER_150_2631 ();
 FILLCELL_X32 FILLER_150_2663 ();
 FILLCELL_X32 FILLER_150_2695 ();
 FILLCELL_X32 FILLER_150_2727 ();
 FILLCELL_X32 FILLER_150_2759 ();
 FILLCELL_X32 FILLER_150_2791 ();
 FILLCELL_X32 FILLER_150_2823 ();
 FILLCELL_X32 FILLER_150_2855 ();
 FILLCELL_X32 FILLER_150_2887 ();
 FILLCELL_X32 FILLER_150_2919 ();
 FILLCELL_X32 FILLER_150_2951 ();
 FILLCELL_X32 FILLER_150_2983 ();
 FILLCELL_X32 FILLER_150_3015 ();
 FILLCELL_X32 FILLER_150_3047 ();
 FILLCELL_X32 FILLER_150_3079 ();
 FILLCELL_X32 FILLER_150_3111 ();
 FILLCELL_X8 FILLER_150_3143 ();
 FILLCELL_X4 FILLER_150_3151 ();
 FILLCELL_X2 FILLER_150_3155 ();
 FILLCELL_X32 FILLER_150_3158 ();
 FILLCELL_X32 FILLER_150_3190 ();
 FILLCELL_X32 FILLER_150_3222 ();
 FILLCELL_X32 FILLER_150_3254 ();
 FILLCELL_X32 FILLER_150_3286 ();
 FILLCELL_X32 FILLER_150_3318 ();
 FILLCELL_X32 FILLER_150_3350 ();
 FILLCELL_X32 FILLER_150_3382 ();
 FILLCELL_X32 FILLER_150_3414 ();
 FILLCELL_X32 FILLER_150_3446 ();
 FILLCELL_X32 FILLER_150_3478 ();
 FILLCELL_X32 FILLER_150_3510 ();
 FILLCELL_X32 FILLER_150_3542 ();
 FILLCELL_X32 FILLER_150_3574 ();
 FILLCELL_X32 FILLER_150_3606 ();
 FILLCELL_X32 FILLER_150_3638 ();
 FILLCELL_X32 FILLER_150_3670 ();
 FILLCELL_X32 FILLER_150_3702 ();
 FILLCELL_X4 FILLER_150_3734 ();
 FILLCELL_X32 FILLER_151_1 ();
 FILLCELL_X32 FILLER_151_33 ();
 FILLCELL_X32 FILLER_151_65 ();
 FILLCELL_X32 FILLER_151_97 ();
 FILLCELL_X32 FILLER_151_129 ();
 FILLCELL_X32 FILLER_151_161 ();
 FILLCELL_X32 FILLER_151_193 ();
 FILLCELL_X32 FILLER_151_225 ();
 FILLCELL_X32 FILLER_151_257 ();
 FILLCELL_X32 FILLER_151_289 ();
 FILLCELL_X32 FILLER_151_321 ();
 FILLCELL_X32 FILLER_151_353 ();
 FILLCELL_X32 FILLER_151_385 ();
 FILLCELL_X32 FILLER_151_417 ();
 FILLCELL_X32 FILLER_151_449 ();
 FILLCELL_X32 FILLER_151_481 ();
 FILLCELL_X32 FILLER_151_513 ();
 FILLCELL_X32 FILLER_151_545 ();
 FILLCELL_X32 FILLER_151_577 ();
 FILLCELL_X32 FILLER_151_609 ();
 FILLCELL_X32 FILLER_151_641 ();
 FILLCELL_X32 FILLER_151_673 ();
 FILLCELL_X32 FILLER_151_705 ();
 FILLCELL_X32 FILLER_151_737 ();
 FILLCELL_X32 FILLER_151_769 ();
 FILLCELL_X32 FILLER_151_801 ();
 FILLCELL_X32 FILLER_151_833 ();
 FILLCELL_X32 FILLER_151_865 ();
 FILLCELL_X32 FILLER_151_897 ();
 FILLCELL_X32 FILLER_151_929 ();
 FILLCELL_X32 FILLER_151_961 ();
 FILLCELL_X32 FILLER_151_993 ();
 FILLCELL_X32 FILLER_151_1025 ();
 FILLCELL_X32 FILLER_151_1057 ();
 FILLCELL_X32 FILLER_151_1089 ();
 FILLCELL_X32 FILLER_151_1121 ();
 FILLCELL_X32 FILLER_151_1153 ();
 FILLCELL_X32 FILLER_151_1185 ();
 FILLCELL_X32 FILLER_151_1217 ();
 FILLCELL_X8 FILLER_151_1249 ();
 FILLCELL_X4 FILLER_151_1257 ();
 FILLCELL_X2 FILLER_151_1261 ();
 FILLCELL_X32 FILLER_151_1264 ();
 FILLCELL_X32 FILLER_151_1296 ();
 FILLCELL_X32 FILLER_151_1328 ();
 FILLCELL_X32 FILLER_151_1360 ();
 FILLCELL_X32 FILLER_151_1392 ();
 FILLCELL_X32 FILLER_151_1424 ();
 FILLCELL_X32 FILLER_151_1456 ();
 FILLCELL_X32 FILLER_151_1488 ();
 FILLCELL_X32 FILLER_151_1520 ();
 FILLCELL_X32 FILLER_151_1552 ();
 FILLCELL_X32 FILLER_151_1584 ();
 FILLCELL_X32 FILLER_151_1616 ();
 FILLCELL_X32 FILLER_151_1648 ();
 FILLCELL_X32 FILLER_151_1680 ();
 FILLCELL_X32 FILLER_151_1712 ();
 FILLCELL_X32 FILLER_151_1744 ();
 FILLCELL_X32 FILLER_151_1776 ();
 FILLCELL_X32 FILLER_151_1808 ();
 FILLCELL_X32 FILLER_151_1840 ();
 FILLCELL_X32 FILLER_151_1872 ();
 FILLCELL_X32 FILLER_151_1904 ();
 FILLCELL_X32 FILLER_151_1936 ();
 FILLCELL_X32 FILLER_151_1968 ();
 FILLCELL_X32 FILLER_151_2000 ();
 FILLCELL_X32 FILLER_151_2032 ();
 FILLCELL_X32 FILLER_151_2064 ();
 FILLCELL_X32 FILLER_151_2096 ();
 FILLCELL_X32 FILLER_151_2128 ();
 FILLCELL_X32 FILLER_151_2160 ();
 FILLCELL_X32 FILLER_151_2192 ();
 FILLCELL_X32 FILLER_151_2224 ();
 FILLCELL_X32 FILLER_151_2256 ();
 FILLCELL_X32 FILLER_151_2288 ();
 FILLCELL_X32 FILLER_151_2320 ();
 FILLCELL_X32 FILLER_151_2352 ();
 FILLCELL_X32 FILLER_151_2384 ();
 FILLCELL_X32 FILLER_151_2416 ();
 FILLCELL_X32 FILLER_151_2448 ();
 FILLCELL_X32 FILLER_151_2480 ();
 FILLCELL_X8 FILLER_151_2512 ();
 FILLCELL_X4 FILLER_151_2520 ();
 FILLCELL_X2 FILLER_151_2524 ();
 FILLCELL_X32 FILLER_151_2527 ();
 FILLCELL_X32 FILLER_151_2559 ();
 FILLCELL_X32 FILLER_151_2591 ();
 FILLCELL_X32 FILLER_151_2623 ();
 FILLCELL_X32 FILLER_151_2655 ();
 FILLCELL_X32 FILLER_151_2687 ();
 FILLCELL_X32 FILLER_151_2719 ();
 FILLCELL_X32 FILLER_151_2751 ();
 FILLCELL_X32 FILLER_151_2783 ();
 FILLCELL_X32 FILLER_151_2815 ();
 FILLCELL_X32 FILLER_151_2847 ();
 FILLCELL_X32 FILLER_151_2879 ();
 FILLCELL_X32 FILLER_151_2911 ();
 FILLCELL_X32 FILLER_151_2943 ();
 FILLCELL_X32 FILLER_151_2975 ();
 FILLCELL_X32 FILLER_151_3007 ();
 FILLCELL_X32 FILLER_151_3039 ();
 FILLCELL_X32 FILLER_151_3071 ();
 FILLCELL_X32 FILLER_151_3103 ();
 FILLCELL_X32 FILLER_151_3135 ();
 FILLCELL_X32 FILLER_151_3167 ();
 FILLCELL_X32 FILLER_151_3199 ();
 FILLCELL_X32 FILLER_151_3231 ();
 FILLCELL_X32 FILLER_151_3263 ();
 FILLCELL_X32 FILLER_151_3295 ();
 FILLCELL_X32 FILLER_151_3327 ();
 FILLCELL_X32 FILLER_151_3359 ();
 FILLCELL_X32 FILLER_151_3391 ();
 FILLCELL_X32 FILLER_151_3423 ();
 FILLCELL_X32 FILLER_151_3455 ();
 FILLCELL_X32 FILLER_151_3487 ();
 FILLCELL_X32 FILLER_151_3519 ();
 FILLCELL_X32 FILLER_151_3551 ();
 FILLCELL_X32 FILLER_151_3583 ();
 FILLCELL_X32 FILLER_151_3615 ();
 FILLCELL_X32 FILLER_151_3647 ();
 FILLCELL_X32 FILLER_151_3679 ();
 FILLCELL_X16 FILLER_151_3711 ();
 FILLCELL_X8 FILLER_151_3727 ();
 FILLCELL_X2 FILLER_151_3735 ();
 FILLCELL_X1 FILLER_151_3737 ();
 FILLCELL_X32 FILLER_152_1 ();
 FILLCELL_X32 FILLER_152_33 ();
 FILLCELL_X32 FILLER_152_65 ();
 FILLCELL_X32 FILLER_152_97 ();
 FILLCELL_X32 FILLER_152_129 ();
 FILLCELL_X32 FILLER_152_161 ();
 FILLCELL_X32 FILLER_152_193 ();
 FILLCELL_X32 FILLER_152_225 ();
 FILLCELL_X32 FILLER_152_257 ();
 FILLCELL_X32 FILLER_152_289 ();
 FILLCELL_X32 FILLER_152_321 ();
 FILLCELL_X32 FILLER_152_353 ();
 FILLCELL_X32 FILLER_152_385 ();
 FILLCELL_X32 FILLER_152_417 ();
 FILLCELL_X32 FILLER_152_449 ();
 FILLCELL_X32 FILLER_152_481 ();
 FILLCELL_X32 FILLER_152_513 ();
 FILLCELL_X32 FILLER_152_545 ();
 FILLCELL_X32 FILLER_152_577 ();
 FILLCELL_X16 FILLER_152_609 ();
 FILLCELL_X4 FILLER_152_625 ();
 FILLCELL_X2 FILLER_152_629 ();
 FILLCELL_X32 FILLER_152_632 ();
 FILLCELL_X32 FILLER_152_664 ();
 FILLCELL_X32 FILLER_152_696 ();
 FILLCELL_X32 FILLER_152_728 ();
 FILLCELL_X32 FILLER_152_760 ();
 FILLCELL_X32 FILLER_152_792 ();
 FILLCELL_X32 FILLER_152_824 ();
 FILLCELL_X32 FILLER_152_856 ();
 FILLCELL_X32 FILLER_152_888 ();
 FILLCELL_X32 FILLER_152_920 ();
 FILLCELL_X32 FILLER_152_952 ();
 FILLCELL_X32 FILLER_152_984 ();
 FILLCELL_X32 FILLER_152_1016 ();
 FILLCELL_X32 FILLER_152_1048 ();
 FILLCELL_X32 FILLER_152_1080 ();
 FILLCELL_X32 FILLER_152_1112 ();
 FILLCELL_X32 FILLER_152_1144 ();
 FILLCELL_X32 FILLER_152_1176 ();
 FILLCELL_X32 FILLER_152_1208 ();
 FILLCELL_X32 FILLER_152_1240 ();
 FILLCELL_X32 FILLER_152_1272 ();
 FILLCELL_X32 FILLER_152_1304 ();
 FILLCELL_X32 FILLER_152_1336 ();
 FILLCELL_X32 FILLER_152_1368 ();
 FILLCELL_X32 FILLER_152_1400 ();
 FILLCELL_X32 FILLER_152_1432 ();
 FILLCELL_X32 FILLER_152_1464 ();
 FILLCELL_X32 FILLER_152_1496 ();
 FILLCELL_X32 FILLER_152_1528 ();
 FILLCELL_X32 FILLER_152_1560 ();
 FILLCELL_X32 FILLER_152_1592 ();
 FILLCELL_X32 FILLER_152_1624 ();
 FILLCELL_X32 FILLER_152_1656 ();
 FILLCELL_X32 FILLER_152_1688 ();
 FILLCELL_X32 FILLER_152_1720 ();
 FILLCELL_X32 FILLER_152_1752 ();
 FILLCELL_X32 FILLER_152_1784 ();
 FILLCELL_X32 FILLER_152_1816 ();
 FILLCELL_X32 FILLER_152_1848 ();
 FILLCELL_X8 FILLER_152_1880 ();
 FILLCELL_X4 FILLER_152_1888 ();
 FILLCELL_X2 FILLER_152_1892 ();
 FILLCELL_X32 FILLER_152_1895 ();
 FILLCELL_X32 FILLER_152_1927 ();
 FILLCELL_X32 FILLER_152_1959 ();
 FILLCELL_X32 FILLER_152_1991 ();
 FILLCELL_X32 FILLER_152_2023 ();
 FILLCELL_X32 FILLER_152_2055 ();
 FILLCELL_X32 FILLER_152_2087 ();
 FILLCELL_X32 FILLER_152_2119 ();
 FILLCELL_X32 FILLER_152_2151 ();
 FILLCELL_X32 FILLER_152_2183 ();
 FILLCELL_X32 FILLER_152_2215 ();
 FILLCELL_X32 FILLER_152_2247 ();
 FILLCELL_X32 FILLER_152_2279 ();
 FILLCELL_X32 FILLER_152_2311 ();
 FILLCELL_X32 FILLER_152_2343 ();
 FILLCELL_X32 FILLER_152_2375 ();
 FILLCELL_X32 FILLER_152_2407 ();
 FILLCELL_X32 FILLER_152_2439 ();
 FILLCELL_X32 FILLER_152_2471 ();
 FILLCELL_X32 FILLER_152_2503 ();
 FILLCELL_X32 FILLER_152_2535 ();
 FILLCELL_X32 FILLER_152_2567 ();
 FILLCELL_X32 FILLER_152_2599 ();
 FILLCELL_X32 FILLER_152_2631 ();
 FILLCELL_X32 FILLER_152_2663 ();
 FILLCELL_X32 FILLER_152_2695 ();
 FILLCELL_X32 FILLER_152_2727 ();
 FILLCELL_X32 FILLER_152_2759 ();
 FILLCELL_X32 FILLER_152_2791 ();
 FILLCELL_X32 FILLER_152_2823 ();
 FILLCELL_X32 FILLER_152_2855 ();
 FILLCELL_X32 FILLER_152_2887 ();
 FILLCELL_X32 FILLER_152_2919 ();
 FILLCELL_X32 FILLER_152_2951 ();
 FILLCELL_X32 FILLER_152_2983 ();
 FILLCELL_X32 FILLER_152_3015 ();
 FILLCELL_X32 FILLER_152_3047 ();
 FILLCELL_X32 FILLER_152_3079 ();
 FILLCELL_X32 FILLER_152_3111 ();
 FILLCELL_X8 FILLER_152_3143 ();
 FILLCELL_X4 FILLER_152_3151 ();
 FILLCELL_X2 FILLER_152_3155 ();
 FILLCELL_X32 FILLER_152_3158 ();
 FILLCELL_X32 FILLER_152_3190 ();
 FILLCELL_X32 FILLER_152_3222 ();
 FILLCELL_X32 FILLER_152_3254 ();
 FILLCELL_X32 FILLER_152_3286 ();
 FILLCELL_X32 FILLER_152_3318 ();
 FILLCELL_X32 FILLER_152_3350 ();
 FILLCELL_X32 FILLER_152_3382 ();
 FILLCELL_X32 FILLER_152_3414 ();
 FILLCELL_X32 FILLER_152_3446 ();
 FILLCELL_X32 FILLER_152_3478 ();
 FILLCELL_X32 FILLER_152_3510 ();
 FILLCELL_X32 FILLER_152_3542 ();
 FILLCELL_X32 FILLER_152_3574 ();
 FILLCELL_X32 FILLER_152_3606 ();
 FILLCELL_X32 FILLER_152_3638 ();
 FILLCELL_X32 FILLER_152_3670 ();
 FILLCELL_X32 FILLER_152_3702 ();
 FILLCELL_X4 FILLER_152_3734 ();
 FILLCELL_X32 FILLER_153_1 ();
 FILLCELL_X32 FILLER_153_33 ();
 FILLCELL_X32 FILLER_153_65 ();
 FILLCELL_X32 FILLER_153_97 ();
 FILLCELL_X32 FILLER_153_129 ();
 FILLCELL_X32 FILLER_153_161 ();
 FILLCELL_X32 FILLER_153_193 ();
 FILLCELL_X32 FILLER_153_225 ();
 FILLCELL_X32 FILLER_153_257 ();
 FILLCELL_X32 FILLER_153_289 ();
 FILLCELL_X32 FILLER_153_321 ();
 FILLCELL_X32 FILLER_153_353 ();
 FILLCELL_X32 FILLER_153_385 ();
 FILLCELL_X32 FILLER_153_417 ();
 FILLCELL_X32 FILLER_153_449 ();
 FILLCELL_X32 FILLER_153_481 ();
 FILLCELL_X32 FILLER_153_513 ();
 FILLCELL_X32 FILLER_153_545 ();
 FILLCELL_X32 FILLER_153_577 ();
 FILLCELL_X32 FILLER_153_609 ();
 FILLCELL_X32 FILLER_153_641 ();
 FILLCELL_X32 FILLER_153_673 ();
 FILLCELL_X32 FILLER_153_705 ();
 FILLCELL_X32 FILLER_153_737 ();
 FILLCELL_X32 FILLER_153_769 ();
 FILLCELL_X32 FILLER_153_801 ();
 FILLCELL_X32 FILLER_153_833 ();
 FILLCELL_X32 FILLER_153_865 ();
 FILLCELL_X32 FILLER_153_897 ();
 FILLCELL_X32 FILLER_153_929 ();
 FILLCELL_X32 FILLER_153_961 ();
 FILLCELL_X32 FILLER_153_993 ();
 FILLCELL_X32 FILLER_153_1025 ();
 FILLCELL_X32 FILLER_153_1057 ();
 FILLCELL_X32 FILLER_153_1089 ();
 FILLCELL_X32 FILLER_153_1121 ();
 FILLCELL_X32 FILLER_153_1153 ();
 FILLCELL_X32 FILLER_153_1185 ();
 FILLCELL_X32 FILLER_153_1217 ();
 FILLCELL_X8 FILLER_153_1249 ();
 FILLCELL_X4 FILLER_153_1257 ();
 FILLCELL_X2 FILLER_153_1261 ();
 FILLCELL_X32 FILLER_153_1264 ();
 FILLCELL_X32 FILLER_153_1296 ();
 FILLCELL_X32 FILLER_153_1328 ();
 FILLCELL_X32 FILLER_153_1360 ();
 FILLCELL_X32 FILLER_153_1392 ();
 FILLCELL_X32 FILLER_153_1424 ();
 FILLCELL_X32 FILLER_153_1456 ();
 FILLCELL_X32 FILLER_153_1488 ();
 FILLCELL_X32 FILLER_153_1520 ();
 FILLCELL_X32 FILLER_153_1552 ();
 FILLCELL_X32 FILLER_153_1584 ();
 FILLCELL_X32 FILLER_153_1616 ();
 FILLCELL_X32 FILLER_153_1648 ();
 FILLCELL_X32 FILLER_153_1680 ();
 FILLCELL_X32 FILLER_153_1712 ();
 FILLCELL_X32 FILLER_153_1744 ();
 FILLCELL_X32 FILLER_153_1776 ();
 FILLCELL_X32 FILLER_153_1808 ();
 FILLCELL_X32 FILLER_153_1840 ();
 FILLCELL_X32 FILLER_153_1872 ();
 FILLCELL_X32 FILLER_153_1904 ();
 FILLCELL_X32 FILLER_153_1936 ();
 FILLCELL_X32 FILLER_153_1968 ();
 FILLCELL_X32 FILLER_153_2000 ();
 FILLCELL_X32 FILLER_153_2032 ();
 FILLCELL_X32 FILLER_153_2064 ();
 FILLCELL_X32 FILLER_153_2096 ();
 FILLCELL_X32 FILLER_153_2128 ();
 FILLCELL_X32 FILLER_153_2160 ();
 FILLCELL_X32 FILLER_153_2192 ();
 FILLCELL_X32 FILLER_153_2224 ();
 FILLCELL_X32 FILLER_153_2256 ();
 FILLCELL_X32 FILLER_153_2288 ();
 FILLCELL_X32 FILLER_153_2320 ();
 FILLCELL_X32 FILLER_153_2352 ();
 FILLCELL_X32 FILLER_153_2384 ();
 FILLCELL_X32 FILLER_153_2416 ();
 FILLCELL_X32 FILLER_153_2448 ();
 FILLCELL_X32 FILLER_153_2480 ();
 FILLCELL_X8 FILLER_153_2512 ();
 FILLCELL_X4 FILLER_153_2520 ();
 FILLCELL_X2 FILLER_153_2524 ();
 FILLCELL_X32 FILLER_153_2527 ();
 FILLCELL_X32 FILLER_153_2559 ();
 FILLCELL_X32 FILLER_153_2591 ();
 FILLCELL_X32 FILLER_153_2623 ();
 FILLCELL_X32 FILLER_153_2655 ();
 FILLCELL_X32 FILLER_153_2687 ();
 FILLCELL_X32 FILLER_153_2719 ();
 FILLCELL_X32 FILLER_153_2751 ();
 FILLCELL_X32 FILLER_153_2783 ();
 FILLCELL_X32 FILLER_153_2815 ();
 FILLCELL_X32 FILLER_153_2847 ();
 FILLCELL_X32 FILLER_153_2879 ();
 FILLCELL_X32 FILLER_153_2911 ();
 FILLCELL_X32 FILLER_153_2943 ();
 FILLCELL_X32 FILLER_153_2975 ();
 FILLCELL_X32 FILLER_153_3007 ();
 FILLCELL_X32 FILLER_153_3039 ();
 FILLCELL_X32 FILLER_153_3071 ();
 FILLCELL_X32 FILLER_153_3103 ();
 FILLCELL_X32 FILLER_153_3135 ();
 FILLCELL_X32 FILLER_153_3167 ();
 FILLCELL_X32 FILLER_153_3199 ();
 FILLCELL_X32 FILLER_153_3231 ();
 FILLCELL_X32 FILLER_153_3263 ();
 FILLCELL_X32 FILLER_153_3295 ();
 FILLCELL_X32 FILLER_153_3327 ();
 FILLCELL_X32 FILLER_153_3359 ();
 FILLCELL_X32 FILLER_153_3391 ();
 FILLCELL_X32 FILLER_153_3423 ();
 FILLCELL_X32 FILLER_153_3455 ();
 FILLCELL_X32 FILLER_153_3487 ();
 FILLCELL_X32 FILLER_153_3519 ();
 FILLCELL_X32 FILLER_153_3551 ();
 FILLCELL_X32 FILLER_153_3583 ();
 FILLCELL_X32 FILLER_153_3615 ();
 FILLCELL_X32 FILLER_153_3647 ();
 FILLCELL_X32 FILLER_153_3679 ();
 FILLCELL_X16 FILLER_153_3711 ();
 FILLCELL_X8 FILLER_153_3727 ();
 FILLCELL_X2 FILLER_153_3735 ();
 FILLCELL_X1 FILLER_153_3737 ();
 FILLCELL_X32 FILLER_154_1 ();
 FILLCELL_X32 FILLER_154_33 ();
 FILLCELL_X32 FILLER_154_65 ();
 FILLCELL_X32 FILLER_154_97 ();
 FILLCELL_X32 FILLER_154_129 ();
 FILLCELL_X32 FILLER_154_161 ();
 FILLCELL_X32 FILLER_154_193 ();
 FILLCELL_X32 FILLER_154_225 ();
 FILLCELL_X32 FILLER_154_257 ();
 FILLCELL_X32 FILLER_154_289 ();
 FILLCELL_X32 FILLER_154_321 ();
 FILLCELL_X32 FILLER_154_353 ();
 FILLCELL_X32 FILLER_154_385 ();
 FILLCELL_X32 FILLER_154_417 ();
 FILLCELL_X32 FILLER_154_449 ();
 FILLCELL_X32 FILLER_154_481 ();
 FILLCELL_X32 FILLER_154_513 ();
 FILLCELL_X32 FILLER_154_545 ();
 FILLCELL_X32 FILLER_154_577 ();
 FILLCELL_X16 FILLER_154_609 ();
 FILLCELL_X4 FILLER_154_625 ();
 FILLCELL_X2 FILLER_154_629 ();
 FILLCELL_X32 FILLER_154_632 ();
 FILLCELL_X32 FILLER_154_664 ();
 FILLCELL_X32 FILLER_154_696 ();
 FILLCELL_X32 FILLER_154_728 ();
 FILLCELL_X32 FILLER_154_760 ();
 FILLCELL_X32 FILLER_154_792 ();
 FILLCELL_X32 FILLER_154_824 ();
 FILLCELL_X32 FILLER_154_856 ();
 FILLCELL_X32 FILLER_154_888 ();
 FILLCELL_X32 FILLER_154_920 ();
 FILLCELL_X32 FILLER_154_952 ();
 FILLCELL_X32 FILLER_154_984 ();
 FILLCELL_X32 FILLER_154_1016 ();
 FILLCELL_X32 FILLER_154_1048 ();
 FILLCELL_X32 FILLER_154_1080 ();
 FILLCELL_X32 FILLER_154_1112 ();
 FILLCELL_X32 FILLER_154_1144 ();
 FILLCELL_X32 FILLER_154_1176 ();
 FILLCELL_X32 FILLER_154_1208 ();
 FILLCELL_X32 FILLER_154_1240 ();
 FILLCELL_X32 FILLER_154_1272 ();
 FILLCELL_X32 FILLER_154_1304 ();
 FILLCELL_X32 FILLER_154_1336 ();
 FILLCELL_X32 FILLER_154_1368 ();
 FILLCELL_X32 FILLER_154_1400 ();
 FILLCELL_X32 FILLER_154_1432 ();
 FILLCELL_X32 FILLER_154_1464 ();
 FILLCELL_X32 FILLER_154_1496 ();
 FILLCELL_X32 FILLER_154_1528 ();
 FILLCELL_X32 FILLER_154_1560 ();
 FILLCELL_X32 FILLER_154_1592 ();
 FILLCELL_X32 FILLER_154_1624 ();
 FILLCELL_X32 FILLER_154_1656 ();
 FILLCELL_X32 FILLER_154_1688 ();
 FILLCELL_X32 FILLER_154_1720 ();
 FILLCELL_X32 FILLER_154_1752 ();
 FILLCELL_X32 FILLER_154_1784 ();
 FILLCELL_X32 FILLER_154_1816 ();
 FILLCELL_X32 FILLER_154_1848 ();
 FILLCELL_X8 FILLER_154_1880 ();
 FILLCELL_X4 FILLER_154_1888 ();
 FILLCELL_X2 FILLER_154_1892 ();
 FILLCELL_X32 FILLER_154_1895 ();
 FILLCELL_X32 FILLER_154_1927 ();
 FILLCELL_X32 FILLER_154_1959 ();
 FILLCELL_X32 FILLER_154_1991 ();
 FILLCELL_X32 FILLER_154_2023 ();
 FILLCELL_X32 FILLER_154_2055 ();
 FILLCELL_X32 FILLER_154_2087 ();
 FILLCELL_X32 FILLER_154_2119 ();
 FILLCELL_X32 FILLER_154_2151 ();
 FILLCELL_X32 FILLER_154_2183 ();
 FILLCELL_X32 FILLER_154_2215 ();
 FILLCELL_X32 FILLER_154_2247 ();
 FILLCELL_X32 FILLER_154_2279 ();
 FILLCELL_X32 FILLER_154_2311 ();
 FILLCELL_X32 FILLER_154_2343 ();
 FILLCELL_X32 FILLER_154_2375 ();
 FILLCELL_X32 FILLER_154_2407 ();
 FILLCELL_X32 FILLER_154_2439 ();
 FILLCELL_X32 FILLER_154_2471 ();
 FILLCELL_X32 FILLER_154_2503 ();
 FILLCELL_X32 FILLER_154_2535 ();
 FILLCELL_X32 FILLER_154_2567 ();
 FILLCELL_X32 FILLER_154_2599 ();
 FILLCELL_X32 FILLER_154_2631 ();
 FILLCELL_X32 FILLER_154_2663 ();
 FILLCELL_X32 FILLER_154_2695 ();
 FILLCELL_X32 FILLER_154_2727 ();
 FILLCELL_X32 FILLER_154_2759 ();
 FILLCELL_X32 FILLER_154_2791 ();
 FILLCELL_X32 FILLER_154_2823 ();
 FILLCELL_X32 FILLER_154_2855 ();
 FILLCELL_X32 FILLER_154_2887 ();
 FILLCELL_X32 FILLER_154_2919 ();
 FILLCELL_X32 FILLER_154_2951 ();
 FILLCELL_X32 FILLER_154_2983 ();
 FILLCELL_X32 FILLER_154_3015 ();
 FILLCELL_X32 FILLER_154_3047 ();
 FILLCELL_X32 FILLER_154_3079 ();
 FILLCELL_X32 FILLER_154_3111 ();
 FILLCELL_X8 FILLER_154_3143 ();
 FILLCELL_X4 FILLER_154_3151 ();
 FILLCELL_X2 FILLER_154_3155 ();
 FILLCELL_X32 FILLER_154_3158 ();
 FILLCELL_X32 FILLER_154_3190 ();
 FILLCELL_X32 FILLER_154_3222 ();
 FILLCELL_X32 FILLER_154_3254 ();
 FILLCELL_X32 FILLER_154_3286 ();
 FILLCELL_X32 FILLER_154_3318 ();
 FILLCELL_X32 FILLER_154_3350 ();
 FILLCELL_X32 FILLER_154_3382 ();
 FILLCELL_X32 FILLER_154_3414 ();
 FILLCELL_X32 FILLER_154_3446 ();
 FILLCELL_X32 FILLER_154_3478 ();
 FILLCELL_X32 FILLER_154_3510 ();
 FILLCELL_X32 FILLER_154_3542 ();
 FILLCELL_X32 FILLER_154_3574 ();
 FILLCELL_X32 FILLER_154_3606 ();
 FILLCELL_X32 FILLER_154_3638 ();
 FILLCELL_X32 FILLER_154_3670 ();
 FILLCELL_X32 FILLER_154_3702 ();
 FILLCELL_X4 FILLER_154_3734 ();
 FILLCELL_X32 FILLER_155_1 ();
 FILLCELL_X32 FILLER_155_33 ();
 FILLCELL_X32 FILLER_155_65 ();
 FILLCELL_X32 FILLER_155_97 ();
 FILLCELL_X32 FILLER_155_129 ();
 FILLCELL_X32 FILLER_155_161 ();
 FILLCELL_X32 FILLER_155_193 ();
 FILLCELL_X32 FILLER_155_225 ();
 FILLCELL_X32 FILLER_155_257 ();
 FILLCELL_X32 FILLER_155_289 ();
 FILLCELL_X32 FILLER_155_321 ();
 FILLCELL_X32 FILLER_155_353 ();
 FILLCELL_X32 FILLER_155_385 ();
 FILLCELL_X32 FILLER_155_417 ();
 FILLCELL_X32 FILLER_155_449 ();
 FILLCELL_X32 FILLER_155_481 ();
 FILLCELL_X32 FILLER_155_513 ();
 FILLCELL_X32 FILLER_155_545 ();
 FILLCELL_X32 FILLER_155_577 ();
 FILLCELL_X32 FILLER_155_609 ();
 FILLCELL_X32 FILLER_155_641 ();
 FILLCELL_X32 FILLER_155_673 ();
 FILLCELL_X32 FILLER_155_705 ();
 FILLCELL_X32 FILLER_155_737 ();
 FILLCELL_X32 FILLER_155_769 ();
 FILLCELL_X32 FILLER_155_801 ();
 FILLCELL_X32 FILLER_155_833 ();
 FILLCELL_X32 FILLER_155_865 ();
 FILLCELL_X32 FILLER_155_897 ();
 FILLCELL_X32 FILLER_155_929 ();
 FILLCELL_X32 FILLER_155_961 ();
 FILLCELL_X32 FILLER_155_993 ();
 FILLCELL_X32 FILLER_155_1025 ();
 FILLCELL_X32 FILLER_155_1057 ();
 FILLCELL_X32 FILLER_155_1089 ();
 FILLCELL_X32 FILLER_155_1121 ();
 FILLCELL_X32 FILLER_155_1153 ();
 FILLCELL_X32 FILLER_155_1185 ();
 FILLCELL_X32 FILLER_155_1217 ();
 FILLCELL_X8 FILLER_155_1249 ();
 FILLCELL_X4 FILLER_155_1257 ();
 FILLCELL_X2 FILLER_155_1261 ();
 FILLCELL_X32 FILLER_155_1264 ();
 FILLCELL_X32 FILLER_155_1296 ();
 FILLCELL_X32 FILLER_155_1328 ();
 FILLCELL_X32 FILLER_155_1360 ();
 FILLCELL_X32 FILLER_155_1392 ();
 FILLCELL_X32 FILLER_155_1424 ();
 FILLCELL_X32 FILLER_155_1456 ();
 FILLCELL_X32 FILLER_155_1488 ();
 FILLCELL_X32 FILLER_155_1520 ();
 FILLCELL_X32 FILLER_155_1552 ();
 FILLCELL_X32 FILLER_155_1584 ();
 FILLCELL_X32 FILLER_155_1616 ();
 FILLCELL_X32 FILLER_155_1648 ();
 FILLCELL_X32 FILLER_155_1680 ();
 FILLCELL_X32 FILLER_155_1712 ();
 FILLCELL_X32 FILLER_155_1744 ();
 FILLCELL_X32 FILLER_155_1776 ();
 FILLCELL_X32 FILLER_155_1808 ();
 FILLCELL_X32 FILLER_155_1840 ();
 FILLCELL_X32 FILLER_155_1872 ();
 FILLCELL_X32 FILLER_155_1904 ();
 FILLCELL_X32 FILLER_155_1936 ();
 FILLCELL_X32 FILLER_155_1968 ();
 FILLCELL_X32 FILLER_155_2000 ();
 FILLCELL_X32 FILLER_155_2032 ();
 FILLCELL_X32 FILLER_155_2064 ();
 FILLCELL_X32 FILLER_155_2096 ();
 FILLCELL_X32 FILLER_155_2128 ();
 FILLCELL_X32 FILLER_155_2160 ();
 FILLCELL_X32 FILLER_155_2192 ();
 FILLCELL_X32 FILLER_155_2224 ();
 FILLCELL_X32 FILLER_155_2256 ();
 FILLCELL_X32 FILLER_155_2288 ();
 FILLCELL_X32 FILLER_155_2320 ();
 FILLCELL_X32 FILLER_155_2352 ();
 FILLCELL_X32 FILLER_155_2384 ();
 FILLCELL_X32 FILLER_155_2416 ();
 FILLCELL_X32 FILLER_155_2448 ();
 FILLCELL_X32 FILLER_155_2480 ();
 FILLCELL_X8 FILLER_155_2512 ();
 FILLCELL_X4 FILLER_155_2520 ();
 FILLCELL_X2 FILLER_155_2524 ();
 FILLCELL_X32 FILLER_155_2527 ();
 FILLCELL_X32 FILLER_155_2559 ();
 FILLCELL_X32 FILLER_155_2591 ();
 FILLCELL_X32 FILLER_155_2623 ();
 FILLCELL_X32 FILLER_155_2655 ();
 FILLCELL_X32 FILLER_155_2687 ();
 FILLCELL_X32 FILLER_155_2719 ();
 FILLCELL_X32 FILLER_155_2751 ();
 FILLCELL_X32 FILLER_155_2783 ();
 FILLCELL_X32 FILLER_155_2815 ();
 FILLCELL_X32 FILLER_155_2847 ();
 FILLCELL_X32 FILLER_155_2879 ();
 FILLCELL_X32 FILLER_155_2911 ();
 FILLCELL_X32 FILLER_155_2943 ();
 FILLCELL_X32 FILLER_155_2975 ();
 FILLCELL_X32 FILLER_155_3007 ();
 FILLCELL_X32 FILLER_155_3039 ();
 FILLCELL_X32 FILLER_155_3071 ();
 FILLCELL_X32 FILLER_155_3103 ();
 FILLCELL_X32 FILLER_155_3135 ();
 FILLCELL_X32 FILLER_155_3167 ();
 FILLCELL_X32 FILLER_155_3199 ();
 FILLCELL_X32 FILLER_155_3231 ();
 FILLCELL_X32 FILLER_155_3263 ();
 FILLCELL_X32 FILLER_155_3295 ();
 FILLCELL_X32 FILLER_155_3327 ();
 FILLCELL_X32 FILLER_155_3359 ();
 FILLCELL_X32 FILLER_155_3391 ();
 FILLCELL_X32 FILLER_155_3423 ();
 FILLCELL_X32 FILLER_155_3455 ();
 FILLCELL_X32 FILLER_155_3487 ();
 FILLCELL_X32 FILLER_155_3519 ();
 FILLCELL_X32 FILLER_155_3551 ();
 FILLCELL_X32 FILLER_155_3583 ();
 FILLCELL_X32 FILLER_155_3615 ();
 FILLCELL_X32 FILLER_155_3647 ();
 FILLCELL_X32 FILLER_155_3679 ();
 FILLCELL_X16 FILLER_155_3711 ();
 FILLCELL_X8 FILLER_155_3727 ();
 FILLCELL_X2 FILLER_155_3735 ();
 FILLCELL_X1 FILLER_155_3737 ();
 FILLCELL_X32 FILLER_156_1 ();
 FILLCELL_X32 FILLER_156_33 ();
 FILLCELL_X32 FILLER_156_65 ();
 FILLCELL_X32 FILLER_156_97 ();
 FILLCELL_X32 FILLER_156_129 ();
 FILLCELL_X32 FILLER_156_161 ();
 FILLCELL_X32 FILLER_156_193 ();
 FILLCELL_X32 FILLER_156_225 ();
 FILLCELL_X32 FILLER_156_257 ();
 FILLCELL_X32 FILLER_156_289 ();
 FILLCELL_X32 FILLER_156_321 ();
 FILLCELL_X32 FILLER_156_353 ();
 FILLCELL_X32 FILLER_156_385 ();
 FILLCELL_X32 FILLER_156_417 ();
 FILLCELL_X32 FILLER_156_449 ();
 FILLCELL_X32 FILLER_156_481 ();
 FILLCELL_X32 FILLER_156_513 ();
 FILLCELL_X32 FILLER_156_545 ();
 FILLCELL_X32 FILLER_156_577 ();
 FILLCELL_X16 FILLER_156_609 ();
 FILLCELL_X4 FILLER_156_625 ();
 FILLCELL_X2 FILLER_156_629 ();
 FILLCELL_X32 FILLER_156_632 ();
 FILLCELL_X32 FILLER_156_664 ();
 FILLCELL_X32 FILLER_156_696 ();
 FILLCELL_X32 FILLER_156_728 ();
 FILLCELL_X32 FILLER_156_760 ();
 FILLCELL_X32 FILLER_156_792 ();
 FILLCELL_X32 FILLER_156_824 ();
 FILLCELL_X32 FILLER_156_856 ();
 FILLCELL_X32 FILLER_156_888 ();
 FILLCELL_X32 FILLER_156_920 ();
 FILLCELL_X32 FILLER_156_952 ();
 FILLCELL_X32 FILLER_156_984 ();
 FILLCELL_X32 FILLER_156_1016 ();
 FILLCELL_X32 FILLER_156_1048 ();
 FILLCELL_X32 FILLER_156_1080 ();
 FILLCELL_X32 FILLER_156_1112 ();
 FILLCELL_X32 FILLER_156_1144 ();
 FILLCELL_X32 FILLER_156_1176 ();
 FILLCELL_X32 FILLER_156_1208 ();
 FILLCELL_X32 FILLER_156_1240 ();
 FILLCELL_X32 FILLER_156_1272 ();
 FILLCELL_X32 FILLER_156_1304 ();
 FILLCELL_X32 FILLER_156_1336 ();
 FILLCELL_X32 FILLER_156_1368 ();
 FILLCELL_X32 FILLER_156_1400 ();
 FILLCELL_X32 FILLER_156_1432 ();
 FILLCELL_X32 FILLER_156_1464 ();
 FILLCELL_X32 FILLER_156_1496 ();
 FILLCELL_X32 FILLER_156_1528 ();
 FILLCELL_X32 FILLER_156_1560 ();
 FILLCELL_X32 FILLER_156_1592 ();
 FILLCELL_X32 FILLER_156_1624 ();
 FILLCELL_X32 FILLER_156_1656 ();
 FILLCELL_X32 FILLER_156_1688 ();
 FILLCELL_X32 FILLER_156_1720 ();
 FILLCELL_X32 FILLER_156_1752 ();
 FILLCELL_X32 FILLER_156_1784 ();
 FILLCELL_X32 FILLER_156_1816 ();
 FILLCELL_X32 FILLER_156_1848 ();
 FILLCELL_X8 FILLER_156_1880 ();
 FILLCELL_X4 FILLER_156_1888 ();
 FILLCELL_X2 FILLER_156_1892 ();
 FILLCELL_X32 FILLER_156_1895 ();
 FILLCELL_X32 FILLER_156_1927 ();
 FILLCELL_X32 FILLER_156_1959 ();
 FILLCELL_X32 FILLER_156_1991 ();
 FILLCELL_X32 FILLER_156_2023 ();
 FILLCELL_X32 FILLER_156_2055 ();
 FILLCELL_X32 FILLER_156_2087 ();
 FILLCELL_X32 FILLER_156_2119 ();
 FILLCELL_X32 FILLER_156_2151 ();
 FILLCELL_X32 FILLER_156_2183 ();
 FILLCELL_X32 FILLER_156_2215 ();
 FILLCELL_X32 FILLER_156_2247 ();
 FILLCELL_X32 FILLER_156_2279 ();
 FILLCELL_X32 FILLER_156_2311 ();
 FILLCELL_X32 FILLER_156_2343 ();
 FILLCELL_X32 FILLER_156_2375 ();
 FILLCELL_X32 FILLER_156_2407 ();
 FILLCELL_X32 FILLER_156_2439 ();
 FILLCELL_X32 FILLER_156_2471 ();
 FILLCELL_X32 FILLER_156_2503 ();
 FILLCELL_X32 FILLER_156_2535 ();
 FILLCELL_X32 FILLER_156_2567 ();
 FILLCELL_X32 FILLER_156_2599 ();
 FILLCELL_X32 FILLER_156_2631 ();
 FILLCELL_X32 FILLER_156_2663 ();
 FILLCELL_X32 FILLER_156_2695 ();
 FILLCELL_X32 FILLER_156_2727 ();
 FILLCELL_X32 FILLER_156_2759 ();
 FILLCELL_X32 FILLER_156_2791 ();
 FILLCELL_X32 FILLER_156_2823 ();
 FILLCELL_X32 FILLER_156_2855 ();
 FILLCELL_X32 FILLER_156_2887 ();
 FILLCELL_X32 FILLER_156_2919 ();
 FILLCELL_X32 FILLER_156_2951 ();
 FILLCELL_X32 FILLER_156_2983 ();
 FILLCELL_X32 FILLER_156_3015 ();
 FILLCELL_X32 FILLER_156_3047 ();
 FILLCELL_X32 FILLER_156_3079 ();
 FILLCELL_X32 FILLER_156_3111 ();
 FILLCELL_X8 FILLER_156_3143 ();
 FILLCELL_X4 FILLER_156_3151 ();
 FILLCELL_X2 FILLER_156_3155 ();
 FILLCELL_X32 FILLER_156_3158 ();
 FILLCELL_X32 FILLER_156_3190 ();
 FILLCELL_X32 FILLER_156_3222 ();
 FILLCELL_X32 FILLER_156_3254 ();
 FILLCELL_X32 FILLER_156_3286 ();
 FILLCELL_X32 FILLER_156_3318 ();
 FILLCELL_X32 FILLER_156_3350 ();
 FILLCELL_X32 FILLER_156_3382 ();
 FILLCELL_X32 FILLER_156_3414 ();
 FILLCELL_X32 FILLER_156_3446 ();
 FILLCELL_X32 FILLER_156_3478 ();
 FILLCELL_X32 FILLER_156_3510 ();
 FILLCELL_X32 FILLER_156_3542 ();
 FILLCELL_X32 FILLER_156_3574 ();
 FILLCELL_X32 FILLER_156_3606 ();
 FILLCELL_X32 FILLER_156_3638 ();
 FILLCELL_X32 FILLER_156_3670 ();
 FILLCELL_X32 FILLER_156_3702 ();
 FILLCELL_X4 FILLER_156_3734 ();
 FILLCELL_X32 FILLER_157_1 ();
 FILLCELL_X32 FILLER_157_33 ();
 FILLCELL_X32 FILLER_157_65 ();
 FILLCELL_X32 FILLER_157_97 ();
 FILLCELL_X32 FILLER_157_129 ();
 FILLCELL_X32 FILLER_157_161 ();
 FILLCELL_X32 FILLER_157_193 ();
 FILLCELL_X32 FILLER_157_225 ();
 FILLCELL_X32 FILLER_157_257 ();
 FILLCELL_X32 FILLER_157_289 ();
 FILLCELL_X32 FILLER_157_321 ();
 FILLCELL_X32 FILLER_157_353 ();
 FILLCELL_X32 FILLER_157_385 ();
 FILLCELL_X32 FILLER_157_417 ();
 FILLCELL_X32 FILLER_157_449 ();
 FILLCELL_X32 FILLER_157_481 ();
 FILLCELL_X32 FILLER_157_513 ();
 FILLCELL_X32 FILLER_157_545 ();
 FILLCELL_X32 FILLER_157_577 ();
 FILLCELL_X32 FILLER_157_609 ();
 FILLCELL_X32 FILLER_157_641 ();
 FILLCELL_X32 FILLER_157_673 ();
 FILLCELL_X32 FILLER_157_705 ();
 FILLCELL_X32 FILLER_157_737 ();
 FILLCELL_X32 FILLER_157_769 ();
 FILLCELL_X32 FILLER_157_801 ();
 FILLCELL_X32 FILLER_157_833 ();
 FILLCELL_X32 FILLER_157_865 ();
 FILLCELL_X32 FILLER_157_897 ();
 FILLCELL_X32 FILLER_157_929 ();
 FILLCELL_X32 FILLER_157_961 ();
 FILLCELL_X32 FILLER_157_993 ();
 FILLCELL_X32 FILLER_157_1025 ();
 FILLCELL_X32 FILLER_157_1057 ();
 FILLCELL_X32 FILLER_157_1089 ();
 FILLCELL_X32 FILLER_157_1121 ();
 FILLCELL_X32 FILLER_157_1153 ();
 FILLCELL_X32 FILLER_157_1185 ();
 FILLCELL_X32 FILLER_157_1217 ();
 FILLCELL_X8 FILLER_157_1249 ();
 FILLCELL_X4 FILLER_157_1257 ();
 FILLCELL_X2 FILLER_157_1261 ();
 FILLCELL_X32 FILLER_157_1264 ();
 FILLCELL_X32 FILLER_157_1296 ();
 FILLCELL_X32 FILLER_157_1328 ();
 FILLCELL_X32 FILLER_157_1360 ();
 FILLCELL_X32 FILLER_157_1392 ();
 FILLCELL_X32 FILLER_157_1424 ();
 FILLCELL_X32 FILLER_157_1456 ();
 FILLCELL_X32 FILLER_157_1488 ();
 FILLCELL_X32 FILLER_157_1520 ();
 FILLCELL_X32 FILLER_157_1552 ();
 FILLCELL_X32 FILLER_157_1584 ();
 FILLCELL_X32 FILLER_157_1616 ();
 FILLCELL_X32 FILLER_157_1648 ();
 FILLCELL_X32 FILLER_157_1680 ();
 FILLCELL_X32 FILLER_157_1712 ();
 FILLCELL_X32 FILLER_157_1744 ();
 FILLCELL_X32 FILLER_157_1776 ();
 FILLCELL_X32 FILLER_157_1808 ();
 FILLCELL_X32 FILLER_157_1840 ();
 FILLCELL_X32 FILLER_157_1872 ();
 FILLCELL_X32 FILLER_157_1904 ();
 FILLCELL_X32 FILLER_157_1936 ();
 FILLCELL_X32 FILLER_157_1968 ();
 FILLCELL_X32 FILLER_157_2000 ();
 FILLCELL_X32 FILLER_157_2032 ();
 FILLCELL_X32 FILLER_157_2064 ();
 FILLCELL_X32 FILLER_157_2096 ();
 FILLCELL_X32 FILLER_157_2128 ();
 FILLCELL_X32 FILLER_157_2160 ();
 FILLCELL_X32 FILLER_157_2192 ();
 FILLCELL_X32 FILLER_157_2224 ();
 FILLCELL_X32 FILLER_157_2256 ();
 FILLCELL_X32 FILLER_157_2288 ();
 FILLCELL_X32 FILLER_157_2320 ();
 FILLCELL_X32 FILLER_157_2352 ();
 FILLCELL_X32 FILLER_157_2384 ();
 FILLCELL_X32 FILLER_157_2416 ();
 FILLCELL_X32 FILLER_157_2448 ();
 FILLCELL_X32 FILLER_157_2480 ();
 FILLCELL_X8 FILLER_157_2512 ();
 FILLCELL_X4 FILLER_157_2520 ();
 FILLCELL_X2 FILLER_157_2524 ();
 FILLCELL_X32 FILLER_157_2527 ();
 FILLCELL_X32 FILLER_157_2559 ();
 FILLCELL_X32 FILLER_157_2591 ();
 FILLCELL_X32 FILLER_157_2623 ();
 FILLCELL_X32 FILLER_157_2655 ();
 FILLCELL_X32 FILLER_157_2687 ();
 FILLCELL_X32 FILLER_157_2719 ();
 FILLCELL_X32 FILLER_157_2751 ();
 FILLCELL_X32 FILLER_157_2783 ();
 FILLCELL_X32 FILLER_157_2815 ();
 FILLCELL_X32 FILLER_157_2847 ();
 FILLCELL_X32 FILLER_157_2879 ();
 FILLCELL_X32 FILLER_157_2911 ();
 FILLCELL_X32 FILLER_157_2943 ();
 FILLCELL_X32 FILLER_157_2975 ();
 FILLCELL_X32 FILLER_157_3007 ();
 FILLCELL_X32 FILLER_157_3039 ();
 FILLCELL_X32 FILLER_157_3071 ();
 FILLCELL_X32 FILLER_157_3103 ();
 FILLCELL_X32 FILLER_157_3135 ();
 FILLCELL_X32 FILLER_157_3167 ();
 FILLCELL_X32 FILLER_157_3199 ();
 FILLCELL_X32 FILLER_157_3231 ();
 FILLCELL_X32 FILLER_157_3263 ();
 FILLCELL_X32 FILLER_157_3295 ();
 FILLCELL_X32 FILLER_157_3327 ();
 FILLCELL_X32 FILLER_157_3359 ();
 FILLCELL_X32 FILLER_157_3391 ();
 FILLCELL_X32 FILLER_157_3423 ();
 FILLCELL_X32 FILLER_157_3455 ();
 FILLCELL_X32 FILLER_157_3487 ();
 FILLCELL_X32 FILLER_157_3519 ();
 FILLCELL_X32 FILLER_157_3551 ();
 FILLCELL_X32 FILLER_157_3583 ();
 FILLCELL_X32 FILLER_157_3615 ();
 FILLCELL_X32 FILLER_157_3647 ();
 FILLCELL_X32 FILLER_157_3679 ();
 FILLCELL_X16 FILLER_157_3711 ();
 FILLCELL_X8 FILLER_157_3727 ();
 FILLCELL_X2 FILLER_157_3735 ();
 FILLCELL_X1 FILLER_157_3737 ();
 FILLCELL_X32 FILLER_158_1 ();
 FILLCELL_X32 FILLER_158_33 ();
 FILLCELL_X32 FILLER_158_65 ();
 FILLCELL_X32 FILLER_158_97 ();
 FILLCELL_X32 FILLER_158_129 ();
 FILLCELL_X32 FILLER_158_161 ();
 FILLCELL_X32 FILLER_158_193 ();
 FILLCELL_X32 FILLER_158_225 ();
 FILLCELL_X32 FILLER_158_257 ();
 FILLCELL_X32 FILLER_158_289 ();
 FILLCELL_X32 FILLER_158_321 ();
 FILLCELL_X32 FILLER_158_353 ();
 FILLCELL_X32 FILLER_158_385 ();
 FILLCELL_X32 FILLER_158_417 ();
 FILLCELL_X32 FILLER_158_449 ();
 FILLCELL_X32 FILLER_158_481 ();
 FILLCELL_X32 FILLER_158_513 ();
 FILLCELL_X32 FILLER_158_545 ();
 FILLCELL_X32 FILLER_158_577 ();
 FILLCELL_X16 FILLER_158_609 ();
 FILLCELL_X4 FILLER_158_625 ();
 FILLCELL_X2 FILLER_158_629 ();
 FILLCELL_X32 FILLER_158_632 ();
 FILLCELL_X32 FILLER_158_664 ();
 FILLCELL_X32 FILLER_158_696 ();
 FILLCELL_X32 FILLER_158_728 ();
 FILLCELL_X32 FILLER_158_760 ();
 FILLCELL_X32 FILLER_158_792 ();
 FILLCELL_X32 FILLER_158_824 ();
 FILLCELL_X32 FILLER_158_856 ();
 FILLCELL_X32 FILLER_158_888 ();
 FILLCELL_X32 FILLER_158_920 ();
 FILLCELL_X32 FILLER_158_952 ();
 FILLCELL_X32 FILLER_158_984 ();
 FILLCELL_X32 FILLER_158_1016 ();
 FILLCELL_X32 FILLER_158_1048 ();
 FILLCELL_X32 FILLER_158_1080 ();
 FILLCELL_X32 FILLER_158_1112 ();
 FILLCELL_X32 FILLER_158_1144 ();
 FILLCELL_X32 FILLER_158_1176 ();
 FILLCELL_X32 FILLER_158_1208 ();
 FILLCELL_X32 FILLER_158_1240 ();
 FILLCELL_X32 FILLER_158_1272 ();
 FILLCELL_X32 FILLER_158_1304 ();
 FILLCELL_X32 FILLER_158_1336 ();
 FILLCELL_X32 FILLER_158_1368 ();
 FILLCELL_X32 FILLER_158_1400 ();
 FILLCELL_X32 FILLER_158_1432 ();
 FILLCELL_X32 FILLER_158_1464 ();
 FILLCELL_X32 FILLER_158_1496 ();
 FILLCELL_X32 FILLER_158_1528 ();
 FILLCELL_X32 FILLER_158_1560 ();
 FILLCELL_X32 FILLER_158_1592 ();
 FILLCELL_X32 FILLER_158_1624 ();
 FILLCELL_X32 FILLER_158_1656 ();
 FILLCELL_X32 FILLER_158_1688 ();
 FILLCELL_X32 FILLER_158_1720 ();
 FILLCELL_X32 FILLER_158_1752 ();
 FILLCELL_X32 FILLER_158_1784 ();
 FILLCELL_X32 FILLER_158_1816 ();
 FILLCELL_X32 FILLER_158_1848 ();
 FILLCELL_X8 FILLER_158_1880 ();
 FILLCELL_X4 FILLER_158_1888 ();
 FILLCELL_X2 FILLER_158_1892 ();
 FILLCELL_X32 FILLER_158_1895 ();
 FILLCELL_X32 FILLER_158_1927 ();
 FILLCELL_X32 FILLER_158_1959 ();
 FILLCELL_X32 FILLER_158_1991 ();
 FILLCELL_X32 FILLER_158_2023 ();
 FILLCELL_X32 FILLER_158_2055 ();
 FILLCELL_X32 FILLER_158_2087 ();
 FILLCELL_X32 FILLER_158_2119 ();
 FILLCELL_X32 FILLER_158_2151 ();
 FILLCELL_X32 FILLER_158_2183 ();
 FILLCELL_X32 FILLER_158_2215 ();
 FILLCELL_X32 FILLER_158_2247 ();
 FILLCELL_X32 FILLER_158_2279 ();
 FILLCELL_X32 FILLER_158_2311 ();
 FILLCELL_X32 FILLER_158_2343 ();
 FILLCELL_X32 FILLER_158_2375 ();
 FILLCELL_X32 FILLER_158_2407 ();
 FILLCELL_X32 FILLER_158_2439 ();
 FILLCELL_X32 FILLER_158_2471 ();
 FILLCELL_X32 FILLER_158_2503 ();
 FILLCELL_X32 FILLER_158_2535 ();
 FILLCELL_X32 FILLER_158_2567 ();
 FILLCELL_X32 FILLER_158_2599 ();
 FILLCELL_X32 FILLER_158_2631 ();
 FILLCELL_X32 FILLER_158_2663 ();
 FILLCELL_X32 FILLER_158_2695 ();
 FILLCELL_X32 FILLER_158_2727 ();
 FILLCELL_X32 FILLER_158_2759 ();
 FILLCELL_X32 FILLER_158_2791 ();
 FILLCELL_X32 FILLER_158_2823 ();
 FILLCELL_X32 FILLER_158_2855 ();
 FILLCELL_X32 FILLER_158_2887 ();
 FILLCELL_X32 FILLER_158_2919 ();
 FILLCELL_X32 FILLER_158_2951 ();
 FILLCELL_X32 FILLER_158_2983 ();
 FILLCELL_X32 FILLER_158_3015 ();
 FILLCELL_X32 FILLER_158_3047 ();
 FILLCELL_X32 FILLER_158_3079 ();
 FILLCELL_X32 FILLER_158_3111 ();
 FILLCELL_X8 FILLER_158_3143 ();
 FILLCELL_X4 FILLER_158_3151 ();
 FILLCELL_X2 FILLER_158_3155 ();
 FILLCELL_X32 FILLER_158_3158 ();
 FILLCELL_X32 FILLER_158_3190 ();
 FILLCELL_X32 FILLER_158_3222 ();
 FILLCELL_X32 FILLER_158_3254 ();
 FILLCELL_X32 FILLER_158_3286 ();
 FILLCELL_X32 FILLER_158_3318 ();
 FILLCELL_X32 FILLER_158_3350 ();
 FILLCELL_X32 FILLER_158_3382 ();
 FILLCELL_X32 FILLER_158_3414 ();
 FILLCELL_X32 FILLER_158_3446 ();
 FILLCELL_X32 FILLER_158_3478 ();
 FILLCELL_X32 FILLER_158_3510 ();
 FILLCELL_X32 FILLER_158_3542 ();
 FILLCELL_X32 FILLER_158_3574 ();
 FILLCELL_X32 FILLER_158_3606 ();
 FILLCELL_X32 FILLER_158_3638 ();
 FILLCELL_X32 FILLER_158_3670 ();
 FILLCELL_X32 FILLER_158_3702 ();
 FILLCELL_X4 FILLER_158_3734 ();
 FILLCELL_X32 FILLER_159_1 ();
 FILLCELL_X32 FILLER_159_33 ();
 FILLCELL_X32 FILLER_159_65 ();
 FILLCELL_X32 FILLER_159_97 ();
 FILLCELL_X32 FILLER_159_129 ();
 FILLCELL_X32 FILLER_159_161 ();
 FILLCELL_X32 FILLER_159_193 ();
 FILLCELL_X32 FILLER_159_225 ();
 FILLCELL_X32 FILLER_159_257 ();
 FILLCELL_X32 FILLER_159_289 ();
 FILLCELL_X32 FILLER_159_321 ();
 FILLCELL_X32 FILLER_159_353 ();
 FILLCELL_X32 FILLER_159_385 ();
 FILLCELL_X32 FILLER_159_417 ();
 FILLCELL_X32 FILLER_159_449 ();
 FILLCELL_X32 FILLER_159_481 ();
 FILLCELL_X32 FILLER_159_513 ();
 FILLCELL_X32 FILLER_159_545 ();
 FILLCELL_X32 FILLER_159_577 ();
 FILLCELL_X32 FILLER_159_609 ();
 FILLCELL_X32 FILLER_159_641 ();
 FILLCELL_X32 FILLER_159_673 ();
 FILLCELL_X32 FILLER_159_705 ();
 FILLCELL_X32 FILLER_159_737 ();
 FILLCELL_X32 FILLER_159_769 ();
 FILLCELL_X32 FILLER_159_801 ();
 FILLCELL_X32 FILLER_159_833 ();
 FILLCELL_X32 FILLER_159_865 ();
 FILLCELL_X32 FILLER_159_897 ();
 FILLCELL_X32 FILLER_159_929 ();
 FILLCELL_X32 FILLER_159_961 ();
 FILLCELL_X32 FILLER_159_993 ();
 FILLCELL_X32 FILLER_159_1025 ();
 FILLCELL_X32 FILLER_159_1057 ();
 FILLCELL_X32 FILLER_159_1089 ();
 FILLCELL_X32 FILLER_159_1121 ();
 FILLCELL_X32 FILLER_159_1153 ();
 FILLCELL_X32 FILLER_159_1185 ();
 FILLCELL_X32 FILLER_159_1217 ();
 FILLCELL_X8 FILLER_159_1249 ();
 FILLCELL_X4 FILLER_159_1257 ();
 FILLCELL_X2 FILLER_159_1261 ();
 FILLCELL_X32 FILLER_159_1264 ();
 FILLCELL_X32 FILLER_159_1296 ();
 FILLCELL_X32 FILLER_159_1328 ();
 FILLCELL_X32 FILLER_159_1360 ();
 FILLCELL_X32 FILLER_159_1392 ();
 FILLCELL_X32 FILLER_159_1424 ();
 FILLCELL_X32 FILLER_159_1456 ();
 FILLCELL_X32 FILLER_159_1488 ();
 FILLCELL_X32 FILLER_159_1520 ();
 FILLCELL_X32 FILLER_159_1552 ();
 FILLCELL_X32 FILLER_159_1584 ();
 FILLCELL_X32 FILLER_159_1616 ();
 FILLCELL_X32 FILLER_159_1648 ();
 FILLCELL_X32 FILLER_159_1680 ();
 FILLCELL_X32 FILLER_159_1712 ();
 FILLCELL_X32 FILLER_159_1744 ();
 FILLCELL_X32 FILLER_159_1776 ();
 FILLCELL_X32 FILLER_159_1808 ();
 FILLCELL_X32 FILLER_159_1840 ();
 FILLCELL_X32 FILLER_159_1872 ();
 FILLCELL_X32 FILLER_159_1904 ();
 FILLCELL_X32 FILLER_159_1936 ();
 FILLCELL_X32 FILLER_159_1968 ();
 FILLCELL_X32 FILLER_159_2000 ();
 FILLCELL_X32 FILLER_159_2032 ();
 FILLCELL_X32 FILLER_159_2064 ();
 FILLCELL_X32 FILLER_159_2096 ();
 FILLCELL_X32 FILLER_159_2128 ();
 FILLCELL_X32 FILLER_159_2160 ();
 FILLCELL_X32 FILLER_159_2192 ();
 FILLCELL_X32 FILLER_159_2224 ();
 FILLCELL_X32 FILLER_159_2256 ();
 FILLCELL_X32 FILLER_159_2288 ();
 FILLCELL_X32 FILLER_159_2320 ();
 FILLCELL_X32 FILLER_159_2352 ();
 FILLCELL_X32 FILLER_159_2384 ();
 FILLCELL_X32 FILLER_159_2416 ();
 FILLCELL_X32 FILLER_159_2448 ();
 FILLCELL_X32 FILLER_159_2480 ();
 FILLCELL_X8 FILLER_159_2512 ();
 FILLCELL_X4 FILLER_159_2520 ();
 FILLCELL_X2 FILLER_159_2524 ();
 FILLCELL_X32 FILLER_159_2527 ();
 FILLCELL_X32 FILLER_159_2559 ();
 FILLCELL_X32 FILLER_159_2591 ();
 FILLCELL_X32 FILLER_159_2623 ();
 FILLCELL_X32 FILLER_159_2655 ();
 FILLCELL_X32 FILLER_159_2687 ();
 FILLCELL_X32 FILLER_159_2719 ();
 FILLCELL_X32 FILLER_159_2751 ();
 FILLCELL_X32 FILLER_159_2783 ();
 FILLCELL_X32 FILLER_159_2815 ();
 FILLCELL_X32 FILLER_159_2847 ();
 FILLCELL_X32 FILLER_159_2879 ();
 FILLCELL_X32 FILLER_159_2911 ();
 FILLCELL_X32 FILLER_159_2943 ();
 FILLCELL_X32 FILLER_159_2975 ();
 FILLCELL_X32 FILLER_159_3007 ();
 FILLCELL_X32 FILLER_159_3039 ();
 FILLCELL_X32 FILLER_159_3071 ();
 FILLCELL_X32 FILLER_159_3103 ();
 FILLCELL_X32 FILLER_159_3135 ();
 FILLCELL_X32 FILLER_159_3167 ();
 FILLCELL_X32 FILLER_159_3199 ();
 FILLCELL_X32 FILLER_159_3231 ();
 FILLCELL_X32 FILLER_159_3263 ();
 FILLCELL_X32 FILLER_159_3295 ();
 FILLCELL_X32 FILLER_159_3327 ();
 FILLCELL_X32 FILLER_159_3359 ();
 FILLCELL_X32 FILLER_159_3391 ();
 FILLCELL_X32 FILLER_159_3423 ();
 FILLCELL_X32 FILLER_159_3455 ();
 FILLCELL_X32 FILLER_159_3487 ();
 FILLCELL_X32 FILLER_159_3519 ();
 FILLCELL_X32 FILLER_159_3551 ();
 FILLCELL_X32 FILLER_159_3583 ();
 FILLCELL_X32 FILLER_159_3615 ();
 FILLCELL_X32 FILLER_159_3647 ();
 FILLCELL_X32 FILLER_159_3679 ();
 FILLCELL_X16 FILLER_159_3711 ();
 FILLCELL_X8 FILLER_159_3727 ();
 FILLCELL_X2 FILLER_159_3735 ();
 FILLCELL_X1 FILLER_159_3737 ();
 FILLCELL_X32 FILLER_160_1 ();
 FILLCELL_X32 FILLER_160_33 ();
 FILLCELL_X32 FILLER_160_65 ();
 FILLCELL_X32 FILLER_160_97 ();
 FILLCELL_X32 FILLER_160_129 ();
 FILLCELL_X32 FILLER_160_161 ();
 FILLCELL_X32 FILLER_160_193 ();
 FILLCELL_X32 FILLER_160_225 ();
 FILLCELL_X32 FILLER_160_257 ();
 FILLCELL_X32 FILLER_160_289 ();
 FILLCELL_X32 FILLER_160_321 ();
 FILLCELL_X32 FILLER_160_353 ();
 FILLCELL_X32 FILLER_160_385 ();
 FILLCELL_X32 FILLER_160_417 ();
 FILLCELL_X32 FILLER_160_449 ();
 FILLCELL_X32 FILLER_160_481 ();
 FILLCELL_X32 FILLER_160_513 ();
 FILLCELL_X32 FILLER_160_545 ();
 FILLCELL_X32 FILLER_160_577 ();
 FILLCELL_X16 FILLER_160_609 ();
 FILLCELL_X4 FILLER_160_625 ();
 FILLCELL_X2 FILLER_160_629 ();
 FILLCELL_X32 FILLER_160_632 ();
 FILLCELL_X32 FILLER_160_664 ();
 FILLCELL_X32 FILLER_160_696 ();
 FILLCELL_X32 FILLER_160_728 ();
 FILLCELL_X32 FILLER_160_760 ();
 FILLCELL_X32 FILLER_160_792 ();
 FILLCELL_X32 FILLER_160_824 ();
 FILLCELL_X32 FILLER_160_856 ();
 FILLCELL_X32 FILLER_160_888 ();
 FILLCELL_X32 FILLER_160_920 ();
 FILLCELL_X32 FILLER_160_952 ();
 FILLCELL_X32 FILLER_160_984 ();
 FILLCELL_X32 FILLER_160_1016 ();
 FILLCELL_X32 FILLER_160_1048 ();
 FILLCELL_X32 FILLER_160_1080 ();
 FILLCELL_X32 FILLER_160_1112 ();
 FILLCELL_X32 FILLER_160_1144 ();
 FILLCELL_X32 FILLER_160_1176 ();
 FILLCELL_X32 FILLER_160_1208 ();
 FILLCELL_X32 FILLER_160_1240 ();
 FILLCELL_X32 FILLER_160_1272 ();
 FILLCELL_X32 FILLER_160_1304 ();
 FILLCELL_X32 FILLER_160_1336 ();
 FILLCELL_X32 FILLER_160_1368 ();
 FILLCELL_X32 FILLER_160_1400 ();
 FILLCELL_X32 FILLER_160_1432 ();
 FILLCELL_X32 FILLER_160_1464 ();
 FILLCELL_X32 FILLER_160_1496 ();
 FILLCELL_X32 FILLER_160_1528 ();
 FILLCELL_X32 FILLER_160_1560 ();
 FILLCELL_X32 FILLER_160_1592 ();
 FILLCELL_X32 FILLER_160_1624 ();
 FILLCELL_X32 FILLER_160_1656 ();
 FILLCELL_X32 FILLER_160_1688 ();
 FILLCELL_X32 FILLER_160_1720 ();
 FILLCELL_X32 FILLER_160_1752 ();
 FILLCELL_X32 FILLER_160_1784 ();
 FILLCELL_X32 FILLER_160_1816 ();
 FILLCELL_X32 FILLER_160_1848 ();
 FILLCELL_X8 FILLER_160_1880 ();
 FILLCELL_X4 FILLER_160_1888 ();
 FILLCELL_X2 FILLER_160_1892 ();
 FILLCELL_X32 FILLER_160_1895 ();
 FILLCELL_X32 FILLER_160_1927 ();
 FILLCELL_X32 FILLER_160_1959 ();
 FILLCELL_X32 FILLER_160_1991 ();
 FILLCELL_X32 FILLER_160_2023 ();
 FILLCELL_X32 FILLER_160_2055 ();
 FILLCELL_X32 FILLER_160_2087 ();
 FILLCELL_X32 FILLER_160_2119 ();
 FILLCELL_X32 FILLER_160_2151 ();
 FILLCELL_X32 FILLER_160_2183 ();
 FILLCELL_X32 FILLER_160_2215 ();
 FILLCELL_X32 FILLER_160_2247 ();
 FILLCELL_X32 FILLER_160_2279 ();
 FILLCELL_X32 FILLER_160_2311 ();
 FILLCELL_X32 FILLER_160_2343 ();
 FILLCELL_X32 FILLER_160_2375 ();
 FILLCELL_X32 FILLER_160_2407 ();
 FILLCELL_X32 FILLER_160_2439 ();
 FILLCELL_X32 FILLER_160_2471 ();
 FILLCELL_X32 FILLER_160_2503 ();
 FILLCELL_X32 FILLER_160_2535 ();
 FILLCELL_X32 FILLER_160_2567 ();
 FILLCELL_X32 FILLER_160_2599 ();
 FILLCELL_X32 FILLER_160_2631 ();
 FILLCELL_X32 FILLER_160_2663 ();
 FILLCELL_X32 FILLER_160_2695 ();
 FILLCELL_X32 FILLER_160_2727 ();
 FILLCELL_X32 FILLER_160_2759 ();
 FILLCELL_X32 FILLER_160_2791 ();
 FILLCELL_X32 FILLER_160_2823 ();
 FILLCELL_X32 FILLER_160_2855 ();
 FILLCELL_X32 FILLER_160_2887 ();
 FILLCELL_X32 FILLER_160_2919 ();
 FILLCELL_X32 FILLER_160_2951 ();
 FILLCELL_X32 FILLER_160_2983 ();
 FILLCELL_X32 FILLER_160_3015 ();
 FILLCELL_X32 FILLER_160_3047 ();
 FILLCELL_X32 FILLER_160_3079 ();
 FILLCELL_X32 FILLER_160_3111 ();
 FILLCELL_X8 FILLER_160_3143 ();
 FILLCELL_X4 FILLER_160_3151 ();
 FILLCELL_X2 FILLER_160_3155 ();
 FILLCELL_X32 FILLER_160_3158 ();
 FILLCELL_X32 FILLER_160_3190 ();
 FILLCELL_X32 FILLER_160_3222 ();
 FILLCELL_X32 FILLER_160_3254 ();
 FILLCELL_X32 FILLER_160_3286 ();
 FILLCELL_X32 FILLER_160_3318 ();
 FILLCELL_X32 FILLER_160_3350 ();
 FILLCELL_X32 FILLER_160_3382 ();
 FILLCELL_X32 FILLER_160_3414 ();
 FILLCELL_X32 FILLER_160_3446 ();
 FILLCELL_X32 FILLER_160_3478 ();
 FILLCELL_X32 FILLER_160_3510 ();
 FILLCELL_X32 FILLER_160_3542 ();
 FILLCELL_X32 FILLER_160_3574 ();
 FILLCELL_X32 FILLER_160_3606 ();
 FILLCELL_X32 FILLER_160_3638 ();
 FILLCELL_X32 FILLER_160_3670 ();
 FILLCELL_X32 FILLER_160_3702 ();
 FILLCELL_X4 FILLER_160_3734 ();
 FILLCELL_X32 FILLER_161_1 ();
 FILLCELL_X32 FILLER_161_33 ();
 FILLCELL_X32 FILLER_161_65 ();
 FILLCELL_X32 FILLER_161_97 ();
 FILLCELL_X32 FILLER_161_129 ();
 FILLCELL_X32 FILLER_161_161 ();
 FILLCELL_X32 FILLER_161_193 ();
 FILLCELL_X32 FILLER_161_225 ();
 FILLCELL_X32 FILLER_161_257 ();
 FILLCELL_X32 FILLER_161_289 ();
 FILLCELL_X32 FILLER_161_321 ();
 FILLCELL_X32 FILLER_161_353 ();
 FILLCELL_X32 FILLER_161_385 ();
 FILLCELL_X32 FILLER_161_417 ();
 FILLCELL_X32 FILLER_161_449 ();
 FILLCELL_X32 FILLER_161_481 ();
 FILLCELL_X32 FILLER_161_513 ();
 FILLCELL_X32 FILLER_161_545 ();
 FILLCELL_X32 FILLER_161_577 ();
 FILLCELL_X32 FILLER_161_609 ();
 FILLCELL_X32 FILLER_161_641 ();
 FILLCELL_X32 FILLER_161_673 ();
 FILLCELL_X32 FILLER_161_705 ();
 FILLCELL_X32 FILLER_161_737 ();
 FILLCELL_X32 FILLER_161_769 ();
 FILLCELL_X32 FILLER_161_801 ();
 FILLCELL_X32 FILLER_161_833 ();
 FILLCELL_X32 FILLER_161_865 ();
 FILLCELL_X32 FILLER_161_897 ();
 FILLCELL_X32 FILLER_161_929 ();
 FILLCELL_X32 FILLER_161_961 ();
 FILLCELL_X32 FILLER_161_993 ();
 FILLCELL_X32 FILLER_161_1025 ();
 FILLCELL_X32 FILLER_161_1057 ();
 FILLCELL_X32 FILLER_161_1089 ();
 FILLCELL_X32 FILLER_161_1121 ();
 FILLCELL_X32 FILLER_161_1153 ();
 FILLCELL_X32 FILLER_161_1185 ();
 FILLCELL_X32 FILLER_161_1217 ();
 FILLCELL_X8 FILLER_161_1249 ();
 FILLCELL_X4 FILLER_161_1257 ();
 FILLCELL_X2 FILLER_161_1261 ();
 FILLCELL_X32 FILLER_161_1264 ();
 FILLCELL_X32 FILLER_161_1296 ();
 FILLCELL_X32 FILLER_161_1328 ();
 FILLCELL_X32 FILLER_161_1360 ();
 FILLCELL_X32 FILLER_161_1392 ();
 FILLCELL_X32 FILLER_161_1424 ();
 FILLCELL_X32 FILLER_161_1456 ();
 FILLCELL_X32 FILLER_161_1488 ();
 FILLCELL_X32 FILLER_161_1520 ();
 FILLCELL_X32 FILLER_161_1552 ();
 FILLCELL_X32 FILLER_161_1584 ();
 FILLCELL_X32 FILLER_161_1616 ();
 FILLCELL_X32 FILLER_161_1648 ();
 FILLCELL_X32 FILLER_161_1680 ();
 FILLCELL_X32 FILLER_161_1712 ();
 FILLCELL_X32 FILLER_161_1744 ();
 FILLCELL_X32 FILLER_161_1776 ();
 FILLCELL_X32 FILLER_161_1808 ();
 FILLCELL_X32 FILLER_161_1840 ();
 FILLCELL_X32 FILLER_161_1872 ();
 FILLCELL_X32 FILLER_161_1904 ();
 FILLCELL_X32 FILLER_161_1936 ();
 FILLCELL_X32 FILLER_161_1968 ();
 FILLCELL_X32 FILLER_161_2000 ();
 FILLCELL_X32 FILLER_161_2032 ();
 FILLCELL_X32 FILLER_161_2064 ();
 FILLCELL_X32 FILLER_161_2096 ();
 FILLCELL_X32 FILLER_161_2128 ();
 FILLCELL_X32 FILLER_161_2160 ();
 FILLCELL_X32 FILLER_161_2192 ();
 FILLCELL_X32 FILLER_161_2224 ();
 FILLCELL_X32 FILLER_161_2256 ();
 FILLCELL_X32 FILLER_161_2288 ();
 FILLCELL_X32 FILLER_161_2320 ();
 FILLCELL_X32 FILLER_161_2352 ();
 FILLCELL_X32 FILLER_161_2384 ();
 FILLCELL_X32 FILLER_161_2416 ();
 FILLCELL_X32 FILLER_161_2448 ();
 FILLCELL_X32 FILLER_161_2480 ();
 FILLCELL_X8 FILLER_161_2512 ();
 FILLCELL_X4 FILLER_161_2520 ();
 FILLCELL_X2 FILLER_161_2524 ();
 FILLCELL_X32 FILLER_161_2527 ();
 FILLCELL_X32 FILLER_161_2559 ();
 FILLCELL_X32 FILLER_161_2591 ();
 FILLCELL_X32 FILLER_161_2623 ();
 FILLCELL_X32 FILLER_161_2655 ();
 FILLCELL_X32 FILLER_161_2687 ();
 FILLCELL_X32 FILLER_161_2719 ();
 FILLCELL_X32 FILLER_161_2751 ();
 FILLCELL_X32 FILLER_161_2783 ();
 FILLCELL_X32 FILLER_161_2815 ();
 FILLCELL_X32 FILLER_161_2847 ();
 FILLCELL_X32 FILLER_161_2879 ();
 FILLCELL_X32 FILLER_161_2911 ();
 FILLCELL_X32 FILLER_161_2943 ();
 FILLCELL_X32 FILLER_161_2975 ();
 FILLCELL_X32 FILLER_161_3007 ();
 FILLCELL_X32 FILLER_161_3039 ();
 FILLCELL_X32 FILLER_161_3071 ();
 FILLCELL_X32 FILLER_161_3103 ();
 FILLCELL_X32 FILLER_161_3135 ();
 FILLCELL_X32 FILLER_161_3167 ();
 FILLCELL_X32 FILLER_161_3199 ();
 FILLCELL_X32 FILLER_161_3231 ();
 FILLCELL_X32 FILLER_161_3263 ();
 FILLCELL_X32 FILLER_161_3295 ();
 FILLCELL_X32 FILLER_161_3327 ();
 FILLCELL_X32 FILLER_161_3359 ();
 FILLCELL_X32 FILLER_161_3391 ();
 FILLCELL_X32 FILLER_161_3423 ();
 FILLCELL_X32 FILLER_161_3455 ();
 FILLCELL_X32 FILLER_161_3487 ();
 FILLCELL_X32 FILLER_161_3519 ();
 FILLCELL_X32 FILLER_161_3551 ();
 FILLCELL_X32 FILLER_161_3583 ();
 FILLCELL_X32 FILLER_161_3615 ();
 FILLCELL_X32 FILLER_161_3647 ();
 FILLCELL_X32 FILLER_161_3679 ();
 FILLCELL_X16 FILLER_161_3711 ();
 FILLCELL_X8 FILLER_161_3727 ();
 FILLCELL_X2 FILLER_161_3735 ();
 FILLCELL_X1 FILLER_161_3737 ();
 FILLCELL_X32 FILLER_162_1 ();
 FILLCELL_X32 FILLER_162_33 ();
 FILLCELL_X32 FILLER_162_65 ();
 FILLCELL_X32 FILLER_162_97 ();
 FILLCELL_X32 FILLER_162_129 ();
 FILLCELL_X32 FILLER_162_161 ();
 FILLCELL_X32 FILLER_162_193 ();
 FILLCELL_X32 FILLER_162_225 ();
 FILLCELL_X32 FILLER_162_257 ();
 FILLCELL_X32 FILLER_162_289 ();
 FILLCELL_X32 FILLER_162_321 ();
 FILLCELL_X32 FILLER_162_353 ();
 FILLCELL_X32 FILLER_162_385 ();
 FILLCELL_X32 FILLER_162_417 ();
 FILLCELL_X32 FILLER_162_449 ();
 FILLCELL_X32 FILLER_162_481 ();
 FILLCELL_X32 FILLER_162_513 ();
 FILLCELL_X32 FILLER_162_545 ();
 FILLCELL_X32 FILLER_162_577 ();
 FILLCELL_X16 FILLER_162_609 ();
 FILLCELL_X4 FILLER_162_625 ();
 FILLCELL_X2 FILLER_162_629 ();
 FILLCELL_X32 FILLER_162_632 ();
 FILLCELL_X32 FILLER_162_664 ();
 FILLCELL_X32 FILLER_162_696 ();
 FILLCELL_X32 FILLER_162_728 ();
 FILLCELL_X32 FILLER_162_760 ();
 FILLCELL_X32 FILLER_162_792 ();
 FILLCELL_X32 FILLER_162_824 ();
 FILLCELL_X32 FILLER_162_856 ();
 FILLCELL_X32 FILLER_162_888 ();
 FILLCELL_X32 FILLER_162_920 ();
 FILLCELL_X32 FILLER_162_952 ();
 FILLCELL_X32 FILLER_162_984 ();
 FILLCELL_X32 FILLER_162_1016 ();
 FILLCELL_X32 FILLER_162_1048 ();
 FILLCELL_X32 FILLER_162_1080 ();
 FILLCELL_X32 FILLER_162_1112 ();
 FILLCELL_X32 FILLER_162_1144 ();
 FILLCELL_X32 FILLER_162_1176 ();
 FILLCELL_X32 FILLER_162_1208 ();
 FILLCELL_X32 FILLER_162_1240 ();
 FILLCELL_X32 FILLER_162_1272 ();
 FILLCELL_X32 FILLER_162_1304 ();
 FILLCELL_X32 FILLER_162_1336 ();
 FILLCELL_X32 FILLER_162_1368 ();
 FILLCELL_X32 FILLER_162_1400 ();
 FILLCELL_X32 FILLER_162_1432 ();
 FILLCELL_X32 FILLER_162_1464 ();
 FILLCELL_X32 FILLER_162_1496 ();
 FILLCELL_X32 FILLER_162_1528 ();
 FILLCELL_X32 FILLER_162_1560 ();
 FILLCELL_X32 FILLER_162_1592 ();
 FILLCELL_X32 FILLER_162_1624 ();
 FILLCELL_X32 FILLER_162_1656 ();
 FILLCELL_X32 FILLER_162_1688 ();
 FILLCELL_X32 FILLER_162_1720 ();
 FILLCELL_X32 FILLER_162_1752 ();
 FILLCELL_X32 FILLER_162_1784 ();
 FILLCELL_X32 FILLER_162_1816 ();
 FILLCELL_X32 FILLER_162_1848 ();
 FILLCELL_X8 FILLER_162_1880 ();
 FILLCELL_X4 FILLER_162_1888 ();
 FILLCELL_X2 FILLER_162_1892 ();
 FILLCELL_X32 FILLER_162_1895 ();
 FILLCELL_X32 FILLER_162_1927 ();
 FILLCELL_X32 FILLER_162_1959 ();
 FILLCELL_X32 FILLER_162_1991 ();
 FILLCELL_X32 FILLER_162_2023 ();
 FILLCELL_X32 FILLER_162_2055 ();
 FILLCELL_X32 FILLER_162_2087 ();
 FILLCELL_X32 FILLER_162_2119 ();
 FILLCELL_X32 FILLER_162_2151 ();
 FILLCELL_X32 FILLER_162_2183 ();
 FILLCELL_X32 FILLER_162_2215 ();
 FILLCELL_X32 FILLER_162_2247 ();
 FILLCELL_X32 FILLER_162_2279 ();
 FILLCELL_X32 FILLER_162_2311 ();
 FILLCELL_X32 FILLER_162_2343 ();
 FILLCELL_X32 FILLER_162_2375 ();
 FILLCELL_X32 FILLER_162_2407 ();
 FILLCELL_X32 FILLER_162_2439 ();
 FILLCELL_X32 FILLER_162_2471 ();
 FILLCELL_X32 FILLER_162_2503 ();
 FILLCELL_X32 FILLER_162_2535 ();
 FILLCELL_X32 FILLER_162_2567 ();
 FILLCELL_X32 FILLER_162_2599 ();
 FILLCELL_X32 FILLER_162_2631 ();
 FILLCELL_X32 FILLER_162_2663 ();
 FILLCELL_X32 FILLER_162_2695 ();
 FILLCELL_X32 FILLER_162_2727 ();
 FILLCELL_X32 FILLER_162_2759 ();
 FILLCELL_X32 FILLER_162_2791 ();
 FILLCELL_X32 FILLER_162_2823 ();
 FILLCELL_X32 FILLER_162_2855 ();
 FILLCELL_X32 FILLER_162_2887 ();
 FILLCELL_X32 FILLER_162_2919 ();
 FILLCELL_X32 FILLER_162_2951 ();
 FILLCELL_X32 FILLER_162_2983 ();
 FILLCELL_X32 FILLER_162_3015 ();
 FILLCELL_X32 FILLER_162_3047 ();
 FILLCELL_X32 FILLER_162_3079 ();
 FILLCELL_X32 FILLER_162_3111 ();
 FILLCELL_X8 FILLER_162_3143 ();
 FILLCELL_X4 FILLER_162_3151 ();
 FILLCELL_X2 FILLER_162_3155 ();
 FILLCELL_X32 FILLER_162_3158 ();
 FILLCELL_X32 FILLER_162_3190 ();
 FILLCELL_X32 FILLER_162_3222 ();
 FILLCELL_X32 FILLER_162_3254 ();
 FILLCELL_X32 FILLER_162_3286 ();
 FILLCELL_X32 FILLER_162_3318 ();
 FILLCELL_X32 FILLER_162_3350 ();
 FILLCELL_X32 FILLER_162_3382 ();
 FILLCELL_X32 FILLER_162_3414 ();
 FILLCELL_X32 FILLER_162_3446 ();
 FILLCELL_X32 FILLER_162_3478 ();
 FILLCELL_X32 FILLER_162_3510 ();
 FILLCELL_X32 FILLER_162_3542 ();
 FILLCELL_X32 FILLER_162_3574 ();
 FILLCELL_X32 FILLER_162_3606 ();
 FILLCELL_X32 FILLER_162_3638 ();
 FILLCELL_X32 FILLER_162_3670 ();
 FILLCELL_X32 FILLER_162_3702 ();
 FILLCELL_X4 FILLER_162_3734 ();
 FILLCELL_X32 FILLER_163_1 ();
 FILLCELL_X32 FILLER_163_33 ();
 FILLCELL_X32 FILLER_163_65 ();
 FILLCELL_X32 FILLER_163_97 ();
 FILLCELL_X32 FILLER_163_129 ();
 FILLCELL_X32 FILLER_163_161 ();
 FILLCELL_X32 FILLER_163_193 ();
 FILLCELL_X32 FILLER_163_225 ();
 FILLCELL_X32 FILLER_163_257 ();
 FILLCELL_X32 FILLER_163_289 ();
 FILLCELL_X32 FILLER_163_321 ();
 FILLCELL_X32 FILLER_163_353 ();
 FILLCELL_X32 FILLER_163_385 ();
 FILLCELL_X32 FILLER_163_417 ();
 FILLCELL_X32 FILLER_163_449 ();
 FILLCELL_X32 FILLER_163_481 ();
 FILLCELL_X32 FILLER_163_513 ();
 FILLCELL_X32 FILLER_163_545 ();
 FILLCELL_X32 FILLER_163_577 ();
 FILLCELL_X32 FILLER_163_609 ();
 FILLCELL_X32 FILLER_163_641 ();
 FILLCELL_X32 FILLER_163_673 ();
 FILLCELL_X32 FILLER_163_705 ();
 FILLCELL_X32 FILLER_163_737 ();
 FILLCELL_X32 FILLER_163_769 ();
 FILLCELL_X32 FILLER_163_801 ();
 FILLCELL_X32 FILLER_163_833 ();
 FILLCELL_X32 FILLER_163_865 ();
 FILLCELL_X32 FILLER_163_897 ();
 FILLCELL_X32 FILLER_163_929 ();
 FILLCELL_X32 FILLER_163_961 ();
 FILLCELL_X32 FILLER_163_993 ();
 FILLCELL_X32 FILLER_163_1025 ();
 FILLCELL_X32 FILLER_163_1057 ();
 FILLCELL_X32 FILLER_163_1089 ();
 FILLCELL_X32 FILLER_163_1121 ();
 FILLCELL_X32 FILLER_163_1153 ();
 FILLCELL_X32 FILLER_163_1185 ();
 FILLCELL_X32 FILLER_163_1217 ();
 FILLCELL_X8 FILLER_163_1249 ();
 FILLCELL_X4 FILLER_163_1257 ();
 FILLCELL_X2 FILLER_163_1261 ();
 FILLCELL_X32 FILLER_163_1264 ();
 FILLCELL_X32 FILLER_163_1296 ();
 FILLCELL_X32 FILLER_163_1328 ();
 FILLCELL_X32 FILLER_163_1360 ();
 FILLCELL_X32 FILLER_163_1392 ();
 FILLCELL_X32 FILLER_163_1424 ();
 FILLCELL_X32 FILLER_163_1456 ();
 FILLCELL_X32 FILLER_163_1488 ();
 FILLCELL_X32 FILLER_163_1520 ();
 FILLCELL_X32 FILLER_163_1552 ();
 FILLCELL_X32 FILLER_163_1584 ();
 FILLCELL_X32 FILLER_163_1616 ();
 FILLCELL_X32 FILLER_163_1648 ();
 FILLCELL_X32 FILLER_163_1680 ();
 FILLCELL_X32 FILLER_163_1712 ();
 FILLCELL_X32 FILLER_163_1744 ();
 FILLCELL_X32 FILLER_163_1776 ();
 FILLCELL_X32 FILLER_163_1808 ();
 FILLCELL_X32 FILLER_163_1840 ();
 FILLCELL_X32 FILLER_163_1872 ();
 FILLCELL_X32 FILLER_163_1904 ();
 FILLCELL_X32 FILLER_163_1936 ();
 FILLCELL_X32 FILLER_163_1968 ();
 FILLCELL_X32 FILLER_163_2000 ();
 FILLCELL_X32 FILLER_163_2032 ();
 FILLCELL_X32 FILLER_163_2064 ();
 FILLCELL_X32 FILLER_163_2096 ();
 FILLCELL_X32 FILLER_163_2128 ();
 FILLCELL_X32 FILLER_163_2160 ();
 FILLCELL_X32 FILLER_163_2192 ();
 FILLCELL_X32 FILLER_163_2224 ();
 FILLCELL_X32 FILLER_163_2256 ();
 FILLCELL_X32 FILLER_163_2288 ();
 FILLCELL_X32 FILLER_163_2320 ();
 FILLCELL_X32 FILLER_163_2352 ();
 FILLCELL_X32 FILLER_163_2384 ();
 FILLCELL_X32 FILLER_163_2416 ();
 FILLCELL_X32 FILLER_163_2448 ();
 FILLCELL_X32 FILLER_163_2480 ();
 FILLCELL_X8 FILLER_163_2512 ();
 FILLCELL_X4 FILLER_163_2520 ();
 FILLCELL_X2 FILLER_163_2524 ();
 FILLCELL_X32 FILLER_163_2527 ();
 FILLCELL_X32 FILLER_163_2559 ();
 FILLCELL_X32 FILLER_163_2591 ();
 FILLCELL_X32 FILLER_163_2623 ();
 FILLCELL_X32 FILLER_163_2655 ();
 FILLCELL_X32 FILLER_163_2687 ();
 FILLCELL_X32 FILLER_163_2719 ();
 FILLCELL_X32 FILLER_163_2751 ();
 FILLCELL_X32 FILLER_163_2783 ();
 FILLCELL_X32 FILLER_163_2815 ();
 FILLCELL_X32 FILLER_163_2847 ();
 FILLCELL_X32 FILLER_163_2879 ();
 FILLCELL_X32 FILLER_163_2911 ();
 FILLCELL_X32 FILLER_163_2943 ();
 FILLCELL_X32 FILLER_163_2975 ();
 FILLCELL_X32 FILLER_163_3007 ();
 FILLCELL_X32 FILLER_163_3039 ();
 FILLCELL_X32 FILLER_163_3071 ();
 FILLCELL_X32 FILLER_163_3103 ();
 FILLCELL_X32 FILLER_163_3135 ();
 FILLCELL_X32 FILLER_163_3167 ();
 FILLCELL_X32 FILLER_163_3199 ();
 FILLCELL_X32 FILLER_163_3231 ();
 FILLCELL_X32 FILLER_163_3263 ();
 FILLCELL_X32 FILLER_163_3295 ();
 FILLCELL_X32 FILLER_163_3327 ();
 FILLCELL_X32 FILLER_163_3359 ();
 FILLCELL_X32 FILLER_163_3391 ();
 FILLCELL_X32 FILLER_163_3423 ();
 FILLCELL_X32 FILLER_163_3455 ();
 FILLCELL_X32 FILLER_163_3487 ();
 FILLCELL_X32 FILLER_163_3519 ();
 FILLCELL_X32 FILLER_163_3551 ();
 FILLCELL_X32 FILLER_163_3583 ();
 FILLCELL_X32 FILLER_163_3615 ();
 FILLCELL_X32 FILLER_163_3647 ();
 FILLCELL_X32 FILLER_163_3679 ();
 FILLCELL_X16 FILLER_163_3711 ();
 FILLCELL_X8 FILLER_163_3727 ();
 FILLCELL_X2 FILLER_163_3735 ();
 FILLCELL_X1 FILLER_163_3737 ();
 FILLCELL_X32 FILLER_164_1 ();
 FILLCELL_X32 FILLER_164_33 ();
 FILLCELL_X32 FILLER_164_65 ();
 FILLCELL_X32 FILLER_164_97 ();
 FILLCELL_X32 FILLER_164_129 ();
 FILLCELL_X32 FILLER_164_161 ();
 FILLCELL_X32 FILLER_164_193 ();
 FILLCELL_X32 FILLER_164_225 ();
 FILLCELL_X32 FILLER_164_257 ();
 FILLCELL_X32 FILLER_164_289 ();
 FILLCELL_X32 FILLER_164_321 ();
 FILLCELL_X32 FILLER_164_353 ();
 FILLCELL_X32 FILLER_164_385 ();
 FILLCELL_X32 FILLER_164_417 ();
 FILLCELL_X32 FILLER_164_449 ();
 FILLCELL_X32 FILLER_164_481 ();
 FILLCELL_X32 FILLER_164_513 ();
 FILLCELL_X32 FILLER_164_545 ();
 FILLCELL_X32 FILLER_164_577 ();
 FILLCELL_X16 FILLER_164_609 ();
 FILLCELL_X4 FILLER_164_625 ();
 FILLCELL_X2 FILLER_164_629 ();
 FILLCELL_X32 FILLER_164_632 ();
 FILLCELL_X32 FILLER_164_664 ();
 FILLCELL_X32 FILLER_164_696 ();
 FILLCELL_X32 FILLER_164_728 ();
 FILLCELL_X32 FILLER_164_760 ();
 FILLCELL_X32 FILLER_164_792 ();
 FILLCELL_X32 FILLER_164_824 ();
 FILLCELL_X32 FILLER_164_856 ();
 FILLCELL_X32 FILLER_164_888 ();
 FILLCELL_X32 FILLER_164_920 ();
 FILLCELL_X32 FILLER_164_952 ();
 FILLCELL_X32 FILLER_164_984 ();
 FILLCELL_X32 FILLER_164_1016 ();
 FILLCELL_X32 FILLER_164_1048 ();
 FILLCELL_X32 FILLER_164_1080 ();
 FILLCELL_X32 FILLER_164_1112 ();
 FILLCELL_X32 FILLER_164_1144 ();
 FILLCELL_X32 FILLER_164_1176 ();
 FILLCELL_X32 FILLER_164_1208 ();
 FILLCELL_X32 FILLER_164_1240 ();
 FILLCELL_X32 FILLER_164_1272 ();
 FILLCELL_X32 FILLER_164_1304 ();
 FILLCELL_X32 FILLER_164_1336 ();
 FILLCELL_X32 FILLER_164_1368 ();
 FILLCELL_X32 FILLER_164_1400 ();
 FILLCELL_X32 FILLER_164_1432 ();
 FILLCELL_X32 FILLER_164_1464 ();
 FILLCELL_X32 FILLER_164_1496 ();
 FILLCELL_X32 FILLER_164_1528 ();
 FILLCELL_X32 FILLER_164_1560 ();
 FILLCELL_X32 FILLER_164_1592 ();
 FILLCELL_X32 FILLER_164_1624 ();
 FILLCELL_X32 FILLER_164_1656 ();
 FILLCELL_X32 FILLER_164_1688 ();
 FILLCELL_X32 FILLER_164_1720 ();
 FILLCELL_X32 FILLER_164_1752 ();
 FILLCELL_X32 FILLER_164_1784 ();
 FILLCELL_X32 FILLER_164_1816 ();
 FILLCELL_X32 FILLER_164_1848 ();
 FILLCELL_X8 FILLER_164_1880 ();
 FILLCELL_X4 FILLER_164_1888 ();
 FILLCELL_X2 FILLER_164_1892 ();
 FILLCELL_X16 FILLER_164_1895 ();
 FILLCELL_X4 FILLER_164_1911 ();
 FILLCELL_X1 FILLER_164_1915 ();
 FILLCELL_X32 FILLER_164_1921 ();
 FILLCELL_X32 FILLER_164_1953 ();
 FILLCELL_X32 FILLER_164_1985 ();
 FILLCELL_X32 FILLER_164_2017 ();
 FILLCELL_X32 FILLER_164_2049 ();
 FILLCELL_X32 FILLER_164_2081 ();
 FILLCELL_X32 FILLER_164_2113 ();
 FILLCELL_X32 FILLER_164_2145 ();
 FILLCELL_X32 FILLER_164_2177 ();
 FILLCELL_X32 FILLER_164_2209 ();
 FILLCELL_X32 FILLER_164_2241 ();
 FILLCELL_X32 FILLER_164_2273 ();
 FILLCELL_X32 FILLER_164_2305 ();
 FILLCELL_X32 FILLER_164_2337 ();
 FILLCELL_X32 FILLER_164_2369 ();
 FILLCELL_X32 FILLER_164_2401 ();
 FILLCELL_X32 FILLER_164_2433 ();
 FILLCELL_X32 FILLER_164_2465 ();
 FILLCELL_X32 FILLER_164_2497 ();
 FILLCELL_X32 FILLER_164_2529 ();
 FILLCELL_X32 FILLER_164_2561 ();
 FILLCELL_X32 FILLER_164_2593 ();
 FILLCELL_X32 FILLER_164_2625 ();
 FILLCELL_X32 FILLER_164_2657 ();
 FILLCELL_X32 FILLER_164_2689 ();
 FILLCELL_X32 FILLER_164_2721 ();
 FILLCELL_X32 FILLER_164_2753 ();
 FILLCELL_X32 FILLER_164_2785 ();
 FILLCELL_X32 FILLER_164_2817 ();
 FILLCELL_X32 FILLER_164_2849 ();
 FILLCELL_X32 FILLER_164_2881 ();
 FILLCELL_X32 FILLER_164_2913 ();
 FILLCELL_X32 FILLER_164_2945 ();
 FILLCELL_X32 FILLER_164_2977 ();
 FILLCELL_X32 FILLER_164_3009 ();
 FILLCELL_X32 FILLER_164_3041 ();
 FILLCELL_X32 FILLER_164_3073 ();
 FILLCELL_X32 FILLER_164_3105 ();
 FILLCELL_X16 FILLER_164_3137 ();
 FILLCELL_X4 FILLER_164_3153 ();
 FILLCELL_X32 FILLER_164_3158 ();
 FILLCELL_X32 FILLER_164_3190 ();
 FILLCELL_X32 FILLER_164_3222 ();
 FILLCELL_X32 FILLER_164_3254 ();
 FILLCELL_X32 FILLER_164_3286 ();
 FILLCELL_X32 FILLER_164_3318 ();
 FILLCELL_X32 FILLER_164_3350 ();
 FILLCELL_X32 FILLER_164_3382 ();
 FILLCELL_X32 FILLER_164_3414 ();
 FILLCELL_X32 FILLER_164_3446 ();
 FILLCELL_X32 FILLER_164_3478 ();
 FILLCELL_X32 FILLER_164_3510 ();
 FILLCELL_X32 FILLER_164_3542 ();
 FILLCELL_X32 FILLER_164_3574 ();
 FILLCELL_X32 FILLER_164_3606 ();
 FILLCELL_X32 FILLER_164_3638 ();
 FILLCELL_X32 FILLER_164_3670 ();
 FILLCELL_X32 FILLER_164_3702 ();
 FILLCELL_X4 FILLER_164_3734 ();
 FILLCELL_X32 FILLER_165_1 ();
 FILLCELL_X32 FILLER_165_33 ();
 FILLCELL_X32 FILLER_165_65 ();
 FILLCELL_X32 FILLER_165_97 ();
 FILLCELL_X32 FILLER_165_129 ();
 FILLCELL_X32 FILLER_165_161 ();
 FILLCELL_X32 FILLER_165_193 ();
 FILLCELL_X32 FILLER_165_225 ();
 FILLCELL_X32 FILLER_165_257 ();
 FILLCELL_X32 FILLER_165_289 ();
 FILLCELL_X32 FILLER_165_321 ();
 FILLCELL_X32 FILLER_165_353 ();
 FILLCELL_X32 FILLER_165_385 ();
 FILLCELL_X32 FILLER_165_417 ();
 FILLCELL_X32 FILLER_165_449 ();
 FILLCELL_X32 FILLER_165_481 ();
 FILLCELL_X32 FILLER_165_513 ();
 FILLCELL_X32 FILLER_165_545 ();
 FILLCELL_X32 FILLER_165_577 ();
 FILLCELL_X32 FILLER_165_609 ();
 FILLCELL_X32 FILLER_165_641 ();
 FILLCELL_X32 FILLER_165_673 ();
 FILLCELL_X32 FILLER_165_705 ();
 FILLCELL_X32 FILLER_165_737 ();
 FILLCELL_X32 FILLER_165_769 ();
 FILLCELL_X32 FILLER_165_801 ();
 FILLCELL_X32 FILLER_165_833 ();
 FILLCELL_X32 FILLER_165_865 ();
 FILLCELL_X32 FILLER_165_897 ();
 FILLCELL_X32 FILLER_165_929 ();
 FILLCELL_X32 FILLER_165_961 ();
 FILLCELL_X32 FILLER_165_993 ();
 FILLCELL_X32 FILLER_165_1025 ();
 FILLCELL_X32 FILLER_165_1057 ();
 FILLCELL_X32 FILLER_165_1089 ();
 FILLCELL_X32 FILLER_165_1121 ();
 FILLCELL_X32 FILLER_165_1153 ();
 FILLCELL_X32 FILLER_165_1185 ();
 FILLCELL_X32 FILLER_165_1217 ();
 FILLCELL_X8 FILLER_165_1249 ();
 FILLCELL_X4 FILLER_165_1257 ();
 FILLCELL_X2 FILLER_165_1261 ();
 FILLCELL_X32 FILLER_165_1264 ();
 FILLCELL_X32 FILLER_165_1296 ();
 FILLCELL_X32 FILLER_165_1328 ();
 FILLCELL_X32 FILLER_165_1360 ();
 FILLCELL_X32 FILLER_165_1392 ();
 FILLCELL_X32 FILLER_165_1424 ();
 FILLCELL_X32 FILLER_165_1456 ();
 FILLCELL_X32 FILLER_165_1488 ();
 FILLCELL_X32 FILLER_165_1520 ();
 FILLCELL_X32 FILLER_165_1552 ();
 FILLCELL_X32 FILLER_165_1584 ();
 FILLCELL_X32 FILLER_165_1616 ();
 FILLCELL_X32 FILLER_165_1648 ();
 FILLCELL_X32 FILLER_165_1680 ();
 FILLCELL_X32 FILLER_165_1712 ();
 FILLCELL_X32 FILLER_165_1744 ();
 FILLCELL_X32 FILLER_165_1776 ();
 FILLCELL_X32 FILLER_165_1808 ();
 FILLCELL_X32 FILLER_165_1840 ();
 FILLCELL_X32 FILLER_165_1872 ();
 FILLCELL_X32 FILLER_165_1904 ();
 FILLCELL_X32 FILLER_165_1936 ();
 FILLCELL_X32 FILLER_165_1968 ();
 FILLCELL_X32 FILLER_165_2000 ();
 FILLCELL_X32 FILLER_165_2032 ();
 FILLCELL_X32 FILLER_165_2064 ();
 FILLCELL_X32 FILLER_165_2096 ();
 FILLCELL_X32 FILLER_165_2128 ();
 FILLCELL_X32 FILLER_165_2160 ();
 FILLCELL_X32 FILLER_165_2192 ();
 FILLCELL_X32 FILLER_165_2224 ();
 FILLCELL_X32 FILLER_165_2256 ();
 FILLCELL_X32 FILLER_165_2288 ();
 FILLCELL_X32 FILLER_165_2320 ();
 FILLCELL_X32 FILLER_165_2352 ();
 FILLCELL_X32 FILLER_165_2384 ();
 FILLCELL_X32 FILLER_165_2416 ();
 FILLCELL_X32 FILLER_165_2448 ();
 FILLCELL_X32 FILLER_165_2480 ();
 FILLCELL_X8 FILLER_165_2512 ();
 FILLCELL_X4 FILLER_165_2520 ();
 FILLCELL_X2 FILLER_165_2524 ();
 FILLCELL_X32 FILLER_165_2527 ();
 FILLCELL_X32 FILLER_165_2559 ();
 FILLCELL_X32 FILLER_165_2591 ();
 FILLCELL_X32 FILLER_165_2623 ();
 FILLCELL_X32 FILLER_165_2655 ();
 FILLCELL_X32 FILLER_165_2687 ();
 FILLCELL_X32 FILLER_165_2719 ();
 FILLCELL_X32 FILLER_165_2751 ();
 FILLCELL_X32 FILLER_165_2783 ();
 FILLCELL_X32 FILLER_165_2815 ();
 FILLCELL_X32 FILLER_165_2847 ();
 FILLCELL_X32 FILLER_165_2879 ();
 FILLCELL_X32 FILLER_165_2911 ();
 FILLCELL_X32 FILLER_165_2943 ();
 FILLCELL_X32 FILLER_165_2975 ();
 FILLCELL_X32 FILLER_165_3007 ();
 FILLCELL_X32 FILLER_165_3039 ();
 FILLCELL_X32 FILLER_165_3071 ();
 FILLCELL_X32 FILLER_165_3103 ();
 FILLCELL_X32 FILLER_165_3135 ();
 FILLCELL_X32 FILLER_165_3167 ();
 FILLCELL_X32 FILLER_165_3199 ();
 FILLCELL_X32 FILLER_165_3231 ();
 FILLCELL_X32 FILLER_165_3263 ();
 FILLCELL_X32 FILLER_165_3295 ();
 FILLCELL_X32 FILLER_165_3327 ();
 FILLCELL_X32 FILLER_165_3359 ();
 FILLCELL_X32 FILLER_165_3391 ();
 FILLCELL_X32 FILLER_165_3423 ();
 FILLCELL_X32 FILLER_165_3455 ();
 FILLCELL_X32 FILLER_165_3487 ();
 FILLCELL_X32 FILLER_165_3519 ();
 FILLCELL_X32 FILLER_165_3551 ();
 FILLCELL_X32 FILLER_165_3583 ();
 FILLCELL_X32 FILLER_165_3615 ();
 FILLCELL_X32 FILLER_165_3647 ();
 FILLCELL_X32 FILLER_165_3679 ();
 FILLCELL_X16 FILLER_165_3711 ();
 FILLCELL_X8 FILLER_165_3727 ();
 FILLCELL_X2 FILLER_165_3735 ();
 FILLCELL_X1 FILLER_165_3737 ();
 FILLCELL_X32 FILLER_166_1 ();
 FILLCELL_X32 FILLER_166_33 ();
 FILLCELL_X32 FILLER_166_65 ();
 FILLCELL_X32 FILLER_166_97 ();
 FILLCELL_X32 FILLER_166_129 ();
 FILLCELL_X32 FILLER_166_161 ();
 FILLCELL_X32 FILLER_166_193 ();
 FILLCELL_X32 FILLER_166_225 ();
 FILLCELL_X32 FILLER_166_257 ();
 FILLCELL_X32 FILLER_166_289 ();
 FILLCELL_X32 FILLER_166_321 ();
 FILLCELL_X32 FILLER_166_353 ();
 FILLCELL_X32 FILLER_166_385 ();
 FILLCELL_X32 FILLER_166_417 ();
 FILLCELL_X32 FILLER_166_449 ();
 FILLCELL_X32 FILLER_166_481 ();
 FILLCELL_X32 FILLER_166_513 ();
 FILLCELL_X32 FILLER_166_545 ();
 FILLCELL_X32 FILLER_166_577 ();
 FILLCELL_X16 FILLER_166_609 ();
 FILLCELL_X4 FILLER_166_625 ();
 FILLCELL_X2 FILLER_166_629 ();
 FILLCELL_X32 FILLER_166_632 ();
 FILLCELL_X32 FILLER_166_664 ();
 FILLCELL_X32 FILLER_166_696 ();
 FILLCELL_X32 FILLER_166_728 ();
 FILLCELL_X32 FILLER_166_760 ();
 FILLCELL_X32 FILLER_166_792 ();
 FILLCELL_X32 FILLER_166_824 ();
 FILLCELL_X32 FILLER_166_856 ();
 FILLCELL_X32 FILLER_166_888 ();
 FILLCELL_X32 FILLER_166_920 ();
 FILLCELL_X32 FILLER_166_952 ();
 FILLCELL_X32 FILLER_166_984 ();
 FILLCELL_X32 FILLER_166_1016 ();
 FILLCELL_X32 FILLER_166_1048 ();
 FILLCELL_X32 FILLER_166_1080 ();
 FILLCELL_X32 FILLER_166_1112 ();
 FILLCELL_X32 FILLER_166_1144 ();
 FILLCELL_X32 FILLER_166_1176 ();
 FILLCELL_X32 FILLER_166_1208 ();
 FILLCELL_X32 FILLER_166_1240 ();
 FILLCELL_X32 FILLER_166_1272 ();
 FILLCELL_X32 FILLER_166_1304 ();
 FILLCELL_X32 FILLER_166_1336 ();
 FILLCELL_X32 FILLER_166_1368 ();
 FILLCELL_X32 FILLER_166_1400 ();
 FILLCELL_X32 FILLER_166_1432 ();
 FILLCELL_X32 FILLER_166_1464 ();
 FILLCELL_X32 FILLER_166_1496 ();
 FILLCELL_X32 FILLER_166_1528 ();
 FILLCELL_X32 FILLER_166_1560 ();
 FILLCELL_X32 FILLER_166_1592 ();
 FILLCELL_X32 FILLER_166_1624 ();
 FILLCELL_X32 FILLER_166_1656 ();
 FILLCELL_X32 FILLER_166_1688 ();
 FILLCELL_X32 FILLER_166_1720 ();
 FILLCELL_X32 FILLER_166_1752 ();
 FILLCELL_X32 FILLER_166_1784 ();
 FILLCELL_X32 FILLER_166_1816 ();
 FILLCELL_X32 FILLER_166_1848 ();
 FILLCELL_X8 FILLER_166_1880 ();
 FILLCELL_X4 FILLER_166_1888 ();
 FILLCELL_X2 FILLER_166_1892 ();
 FILLCELL_X32 FILLER_166_1895 ();
 FILLCELL_X32 FILLER_166_1927 ();
 FILLCELL_X32 FILLER_166_1959 ();
 FILLCELL_X32 FILLER_166_1991 ();
 FILLCELL_X32 FILLER_166_2023 ();
 FILLCELL_X32 FILLER_166_2055 ();
 FILLCELL_X32 FILLER_166_2087 ();
 FILLCELL_X32 FILLER_166_2119 ();
 FILLCELL_X32 FILLER_166_2151 ();
 FILLCELL_X32 FILLER_166_2183 ();
 FILLCELL_X32 FILLER_166_2215 ();
 FILLCELL_X32 FILLER_166_2247 ();
 FILLCELL_X32 FILLER_166_2279 ();
 FILLCELL_X32 FILLER_166_2311 ();
 FILLCELL_X32 FILLER_166_2343 ();
 FILLCELL_X32 FILLER_166_2375 ();
 FILLCELL_X32 FILLER_166_2407 ();
 FILLCELL_X32 FILLER_166_2439 ();
 FILLCELL_X32 FILLER_166_2471 ();
 FILLCELL_X32 FILLER_166_2503 ();
 FILLCELL_X32 FILLER_166_2535 ();
 FILLCELL_X32 FILLER_166_2567 ();
 FILLCELL_X32 FILLER_166_2599 ();
 FILLCELL_X32 FILLER_166_2631 ();
 FILLCELL_X32 FILLER_166_2663 ();
 FILLCELL_X32 FILLER_166_2695 ();
 FILLCELL_X32 FILLER_166_2727 ();
 FILLCELL_X32 FILLER_166_2759 ();
 FILLCELL_X32 FILLER_166_2791 ();
 FILLCELL_X32 FILLER_166_2823 ();
 FILLCELL_X32 FILLER_166_2855 ();
 FILLCELL_X32 FILLER_166_2887 ();
 FILLCELL_X32 FILLER_166_2919 ();
 FILLCELL_X32 FILLER_166_2951 ();
 FILLCELL_X32 FILLER_166_2983 ();
 FILLCELL_X32 FILLER_166_3015 ();
 FILLCELL_X32 FILLER_166_3047 ();
 FILLCELL_X32 FILLER_166_3079 ();
 FILLCELL_X32 FILLER_166_3111 ();
 FILLCELL_X8 FILLER_166_3143 ();
 FILLCELL_X4 FILLER_166_3151 ();
 FILLCELL_X2 FILLER_166_3155 ();
 FILLCELL_X32 FILLER_166_3158 ();
 FILLCELL_X32 FILLER_166_3190 ();
 FILLCELL_X32 FILLER_166_3222 ();
 FILLCELL_X32 FILLER_166_3254 ();
 FILLCELL_X32 FILLER_166_3286 ();
 FILLCELL_X32 FILLER_166_3318 ();
 FILLCELL_X32 FILLER_166_3350 ();
 FILLCELL_X32 FILLER_166_3382 ();
 FILLCELL_X32 FILLER_166_3414 ();
 FILLCELL_X32 FILLER_166_3446 ();
 FILLCELL_X32 FILLER_166_3478 ();
 FILLCELL_X32 FILLER_166_3510 ();
 FILLCELL_X32 FILLER_166_3542 ();
 FILLCELL_X32 FILLER_166_3574 ();
 FILLCELL_X32 FILLER_166_3606 ();
 FILLCELL_X32 FILLER_166_3638 ();
 FILLCELL_X32 FILLER_166_3670 ();
 FILLCELL_X32 FILLER_166_3702 ();
 FILLCELL_X4 FILLER_166_3734 ();
 FILLCELL_X32 FILLER_167_1 ();
 FILLCELL_X32 FILLER_167_33 ();
 FILLCELL_X32 FILLER_167_65 ();
 FILLCELL_X32 FILLER_167_97 ();
 FILLCELL_X32 FILLER_167_129 ();
 FILLCELL_X32 FILLER_167_161 ();
 FILLCELL_X32 FILLER_167_193 ();
 FILLCELL_X32 FILLER_167_225 ();
 FILLCELL_X32 FILLER_167_257 ();
 FILLCELL_X32 FILLER_167_289 ();
 FILLCELL_X32 FILLER_167_321 ();
 FILLCELL_X32 FILLER_167_353 ();
 FILLCELL_X32 FILLER_167_385 ();
 FILLCELL_X32 FILLER_167_417 ();
 FILLCELL_X32 FILLER_167_449 ();
 FILLCELL_X32 FILLER_167_481 ();
 FILLCELL_X32 FILLER_167_513 ();
 FILLCELL_X32 FILLER_167_545 ();
 FILLCELL_X32 FILLER_167_577 ();
 FILLCELL_X32 FILLER_167_609 ();
 FILLCELL_X32 FILLER_167_641 ();
 FILLCELL_X32 FILLER_167_673 ();
 FILLCELL_X32 FILLER_167_705 ();
 FILLCELL_X32 FILLER_167_737 ();
 FILLCELL_X32 FILLER_167_769 ();
 FILLCELL_X32 FILLER_167_801 ();
 FILLCELL_X32 FILLER_167_833 ();
 FILLCELL_X32 FILLER_167_865 ();
 FILLCELL_X32 FILLER_167_897 ();
 FILLCELL_X32 FILLER_167_929 ();
 FILLCELL_X32 FILLER_167_961 ();
 FILLCELL_X32 FILLER_167_993 ();
 FILLCELL_X32 FILLER_167_1025 ();
 FILLCELL_X32 FILLER_167_1057 ();
 FILLCELL_X32 FILLER_167_1089 ();
 FILLCELL_X32 FILLER_167_1121 ();
 FILLCELL_X32 FILLER_167_1153 ();
 FILLCELL_X32 FILLER_167_1185 ();
 FILLCELL_X32 FILLER_167_1217 ();
 FILLCELL_X8 FILLER_167_1249 ();
 FILLCELL_X4 FILLER_167_1257 ();
 FILLCELL_X2 FILLER_167_1261 ();
 FILLCELL_X32 FILLER_167_1264 ();
 FILLCELL_X32 FILLER_167_1296 ();
 FILLCELL_X32 FILLER_167_1328 ();
 FILLCELL_X32 FILLER_167_1360 ();
 FILLCELL_X32 FILLER_167_1392 ();
 FILLCELL_X32 FILLER_167_1424 ();
 FILLCELL_X32 FILLER_167_1456 ();
 FILLCELL_X32 FILLER_167_1488 ();
 FILLCELL_X32 FILLER_167_1520 ();
 FILLCELL_X32 FILLER_167_1552 ();
 FILLCELL_X32 FILLER_167_1584 ();
 FILLCELL_X32 FILLER_167_1616 ();
 FILLCELL_X32 FILLER_167_1648 ();
 FILLCELL_X32 FILLER_167_1680 ();
 FILLCELL_X32 FILLER_167_1712 ();
 FILLCELL_X32 FILLER_167_1744 ();
 FILLCELL_X32 FILLER_167_1776 ();
 FILLCELL_X32 FILLER_167_1808 ();
 FILLCELL_X32 FILLER_167_1840 ();
 FILLCELL_X32 FILLER_167_1872 ();
 FILLCELL_X32 FILLER_167_1904 ();
 FILLCELL_X32 FILLER_167_1936 ();
 FILLCELL_X32 FILLER_167_1968 ();
 FILLCELL_X32 FILLER_167_2000 ();
 FILLCELL_X32 FILLER_167_2032 ();
 FILLCELL_X32 FILLER_167_2064 ();
 FILLCELL_X32 FILLER_167_2096 ();
 FILLCELL_X32 FILLER_167_2128 ();
 FILLCELL_X32 FILLER_167_2160 ();
 FILLCELL_X32 FILLER_167_2192 ();
 FILLCELL_X32 FILLER_167_2224 ();
 FILLCELL_X32 FILLER_167_2256 ();
 FILLCELL_X32 FILLER_167_2288 ();
 FILLCELL_X32 FILLER_167_2320 ();
 FILLCELL_X32 FILLER_167_2352 ();
 FILLCELL_X32 FILLER_167_2384 ();
 FILLCELL_X32 FILLER_167_2416 ();
 FILLCELL_X32 FILLER_167_2448 ();
 FILLCELL_X32 FILLER_167_2480 ();
 FILLCELL_X8 FILLER_167_2512 ();
 FILLCELL_X4 FILLER_167_2520 ();
 FILLCELL_X2 FILLER_167_2524 ();
 FILLCELL_X32 FILLER_167_2527 ();
 FILLCELL_X32 FILLER_167_2559 ();
 FILLCELL_X32 FILLER_167_2591 ();
 FILLCELL_X32 FILLER_167_2623 ();
 FILLCELL_X32 FILLER_167_2655 ();
 FILLCELL_X32 FILLER_167_2687 ();
 FILLCELL_X32 FILLER_167_2719 ();
 FILLCELL_X32 FILLER_167_2751 ();
 FILLCELL_X32 FILLER_167_2783 ();
 FILLCELL_X32 FILLER_167_2815 ();
 FILLCELL_X32 FILLER_167_2847 ();
 FILLCELL_X32 FILLER_167_2879 ();
 FILLCELL_X32 FILLER_167_2911 ();
 FILLCELL_X32 FILLER_167_2943 ();
 FILLCELL_X32 FILLER_167_2975 ();
 FILLCELL_X32 FILLER_167_3007 ();
 FILLCELL_X32 FILLER_167_3039 ();
 FILLCELL_X32 FILLER_167_3071 ();
 FILLCELL_X32 FILLER_167_3103 ();
 FILLCELL_X32 FILLER_167_3135 ();
 FILLCELL_X32 FILLER_167_3167 ();
 FILLCELL_X32 FILLER_167_3199 ();
 FILLCELL_X32 FILLER_167_3231 ();
 FILLCELL_X32 FILLER_167_3263 ();
 FILLCELL_X32 FILLER_167_3295 ();
 FILLCELL_X32 FILLER_167_3327 ();
 FILLCELL_X32 FILLER_167_3359 ();
 FILLCELL_X32 FILLER_167_3391 ();
 FILLCELL_X32 FILLER_167_3423 ();
 FILLCELL_X32 FILLER_167_3455 ();
 FILLCELL_X32 FILLER_167_3487 ();
 FILLCELL_X32 FILLER_167_3519 ();
 FILLCELL_X32 FILLER_167_3551 ();
 FILLCELL_X32 FILLER_167_3583 ();
 FILLCELL_X32 FILLER_167_3615 ();
 FILLCELL_X32 FILLER_167_3647 ();
 FILLCELL_X32 FILLER_167_3679 ();
 FILLCELL_X16 FILLER_167_3711 ();
 FILLCELL_X8 FILLER_167_3727 ();
 FILLCELL_X2 FILLER_167_3735 ();
 FILLCELL_X1 FILLER_167_3737 ();
 FILLCELL_X32 FILLER_168_1 ();
 FILLCELL_X32 FILLER_168_33 ();
 FILLCELL_X32 FILLER_168_65 ();
 FILLCELL_X32 FILLER_168_97 ();
 FILLCELL_X32 FILLER_168_129 ();
 FILLCELL_X32 FILLER_168_161 ();
 FILLCELL_X32 FILLER_168_193 ();
 FILLCELL_X32 FILLER_168_225 ();
 FILLCELL_X32 FILLER_168_257 ();
 FILLCELL_X32 FILLER_168_289 ();
 FILLCELL_X32 FILLER_168_321 ();
 FILLCELL_X32 FILLER_168_353 ();
 FILLCELL_X32 FILLER_168_385 ();
 FILLCELL_X32 FILLER_168_417 ();
 FILLCELL_X32 FILLER_168_449 ();
 FILLCELL_X32 FILLER_168_481 ();
 FILLCELL_X32 FILLER_168_513 ();
 FILLCELL_X32 FILLER_168_545 ();
 FILLCELL_X32 FILLER_168_577 ();
 FILLCELL_X16 FILLER_168_609 ();
 FILLCELL_X4 FILLER_168_625 ();
 FILLCELL_X2 FILLER_168_629 ();
 FILLCELL_X32 FILLER_168_632 ();
 FILLCELL_X32 FILLER_168_664 ();
 FILLCELL_X32 FILLER_168_696 ();
 FILLCELL_X32 FILLER_168_728 ();
 FILLCELL_X32 FILLER_168_760 ();
 FILLCELL_X32 FILLER_168_792 ();
 FILLCELL_X32 FILLER_168_824 ();
 FILLCELL_X32 FILLER_168_856 ();
 FILLCELL_X32 FILLER_168_888 ();
 FILLCELL_X32 FILLER_168_920 ();
 FILLCELL_X32 FILLER_168_952 ();
 FILLCELL_X32 FILLER_168_984 ();
 FILLCELL_X32 FILLER_168_1016 ();
 FILLCELL_X32 FILLER_168_1048 ();
 FILLCELL_X32 FILLER_168_1080 ();
 FILLCELL_X32 FILLER_168_1112 ();
 FILLCELL_X32 FILLER_168_1144 ();
 FILLCELL_X32 FILLER_168_1176 ();
 FILLCELL_X32 FILLER_168_1208 ();
 FILLCELL_X32 FILLER_168_1240 ();
 FILLCELL_X32 FILLER_168_1272 ();
 FILLCELL_X32 FILLER_168_1304 ();
 FILLCELL_X32 FILLER_168_1336 ();
 FILLCELL_X32 FILLER_168_1368 ();
 FILLCELL_X32 FILLER_168_1400 ();
 FILLCELL_X32 FILLER_168_1432 ();
 FILLCELL_X32 FILLER_168_1464 ();
 FILLCELL_X32 FILLER_168_1496 ();
 FILLCELL_X32 FILLER_168_1528 ();
 FILLCELL_X32 FILLER_168_1560 ();
 FILLCELL_X32 FILLER_168_1592 ();
 FILLCELL_X32 FILLER_168_1624 ();
 FILLCELL_X32 FILLER_168_1656 ();
 FILLCELL_X32 FILLER_168_1688 ();
 FILLCELL_X32 FILLER_168_1720 ();
 FILLCELL_X32 FILLER_168_1752 ();
 FILLCELL_X32 FILLER_168_1784 ();
 FILLCELL_X32 FILLER_168_1816 ();
 FILLCELL_X32 FILLER_168_1848 ();
 FILLCELL_X8 FILLER_168_1880 ();
 FILLCELL_X4 FILLER_168_1888 ();
 FILLCELL_X2 FILLER_168_1892 ();
 FILLCELL_X32 FILLER_168_1895 ();
 FILLCELL_X32 FILLER_168_1927 ();
 FILLCELL_X32 FILLER_168_1959 ();
 FILLCELL_X32 FILLER_168_1991 ();
 FILLCELL_X32 FILLER_168_2023 ();
 FILLCELL_X32 FILLER_168_2055 ();
 FILLCELL_X32 FILLER_168_2087 ();
 FILLCELL_X32 FILLER_168_2119 ();
 FILLCELL_X32 FILLER_168_2151 ();
 FILLCELL_X32 FILLER_168_2183 ();
 FILLCELL_X32 FILLER_168_2215 ();
 FILLCELL_X32 FILLER_168_2247 ();
 FILLCELL_X32 FILLER_168_2279 ();
 FILLCELL_X32 FILLER_168_2311 ();
 FILLCELL_X32 FILLER_168_2343 ();
 FILLCELL_X32 FILLER_168_2375 ();
 FILLCELL_X32 FILLER_168_2407 ();
 FILLCELL_X32 FILLER_168_2439 ();
 FILLCELL_X32 FILLER_168_2471 ();
 FILLCELL_X32 FILLER_168_2503 ();
 FILLCELL_X32 FILLER_168_2535 ();
 FILLCELL_X32 FILLER_168_2567 ();
 FILLCELL_X32 FILLER_168_2599 ();
 FILLCELL_X32 FILLER_168_2631 ();
 FILLCELL_X32 FILLER_168_2663 ();
 FILLCELL_X32 FILLER_168_2695 ();
 FILLCELL_X32 FILLER_168_2727 ();
 FILLCELL_X32 FILLER_168_2759 ();
 FILLCELL_X32 FILLER_168_2791 ();
 FILLCELL_X32 FILLER_168_2823 ();
 FILLCELL_X32 FILLER_168_2855 ();
 FILLCELL_X32 FILLER_168_2887 ();
 FILLCELL_X32 FILLER_168_2919 ();
 FILLCELL_X32 FILLER_168_2951 ();
 FILLCELL_X32 FILLER_168_2983 ();
 FILLCELL_X32 FILLER_168_3015 ();
 FILLCELL_X32 FILLER_168_3047 ();
 FILLCELL_X32 FILLER_168_3079 ();
 FILLCELL_X32 FILLER_168_3111 ();
 FILLCELL_X8 FILLER_168_3143 ();
 FILLCELL_X4 FILLER_168_3151 ();
 FILLCELL_X2 FILLER_168_3155 ();
 FILLCELL_X32 FILLER_168_3158 ();
 FILLCELL_X32 FILLER_168_3190 ();
 FILLCELL_X32 FILLER_168_3222 ();
 FILLCELL_X32 FILLER_168_3254 ();
 FILLCELL_X32 FILLER_168_3286 ();
 FILLCELL_X32 FILLER_168_3318 ();
 FILLCELL_X32 FILLER_168_3350 ();
 FILLCELL_X32 FILLER_168_3382 ();
 FILLCELL_X32 FILLER_168_3414 ();
 FILLCELL_X32 FILLER_168_3446 ();
 FILLCELL_X32 FILLER_168_3478 ();
 FILLCELL_X32 FILLER_168_3510 ();
 FILLCELL_X32 FILLER_168_3542 ();
 FILLCELL_X32 FILLER_168_3574 ();
 FILLCELL_X32 FILLER_168_3606 ();
 FILLCELL_X32 FILLER_168_3638 ();
 FILLCELL_X32 FILLER_168_3670 ();
 FILLCELL_X32 FILLER_168_3702 ();
 FILLCELL_X4 FILLER_168_3734 ();
 FILLCELL_X32 FILLER_169_1 ();
 FILLCELL_X32 FILLER_169_33 ();
 FILLCELL_X32 FILLER_169_65 ();
 FILLCELL_X32 FILLER_169_97 ();
 FILLCELL_X32 FILLER_169_129 ();
 FILLCELL_X32 FILLER_169_161 ();
 FILLCELL_X32 FILLER_169_193 ();
 FILLCELL_X32 FILLER_169_225 ();
 FILLCELL_X32 FILLER_169_257 ();
 FILLCELL_X32 FILLER_169_289 ();
 FILLCELL_X32 FILLER_169_321 ();
 FILLCELL_X32 FILLER_169_353 ();
 FILLCELL_X32 FILLER_169_385 ();
 FILLCELL_X32 FILLER_169_417 ();
 FILLCELL_X32 FILLER_169_449 ();
 FILLCELL_X32 FILLER_169_481 ();
 FILLCELL_X32 FILLER_169_513 ();
 FILLCELL_X32 FILLER_169_545 ();
 FILLCELL_X32 FILLER_169_577 ();
 FILLCELL_X32 FILLER_169_609 ();
 FILLCELL_X32 FILLER_169_641 ();
 FILLCELL_X32 FILLER_169_673 ();
 FILLCELL_X32 FILLER_169_705 ();
 FILLCELL_X32 FILLER_169_737 ();
 FILLCELL_X32 FILLER_169_769 ();
 FILLCELL_X32 FILLER_169_801 ();
 FILLCELL_X32 FILLER_169_833 ();
 FILLCELL_X32 FILLER_169_865 ();
 FILLCELL_X32 FILLER_169_897 ();
 FILLCELL_X32 FILLER_169_929 ();
 FILLCELL_X32 FILLER_169_961 ();
 FILLCELL_X32 FILLER_169_993 ();
 FILLCELL_X32 FILLER_169_1025 ();
 FILLCELL_X32 FILLER_169_1057 ();
 FILLCELL_X32 FILLER_169_1089 ();
 FILLCELL_X32 FILLER_169_1121 ();
 FILLCELL_X32 FILLER_169_1153 ();
 FILLCELL_X32 FILLER_169_1185 ();
 FILLCELL_X32 FILLER_169_1217 ();
 FILLCELL_X8 FILLER_169_1249 ();
 FILLCELL_X4 FILLER_169_1257 ();
 FILLCELL_X2 FILLER_169_1261 ();
 FILLCELL_X32 FILLER_169_1264 ();
 FILLCELL_X32 FILLER_169_1296 ();
 FILLCELL_X32 FILLER_169_1328 ();
 FILLCELL_X32 FILLER_169_1360 ();
 FILLCELL_X32 FILLER_169_1392 ();
 FILLCELL_X32 FILLER_169_1424 ();
 FILLCELL_X32 FILLER_169_1456 ();
 FILLCELL_X32 FILLER_169_1488 ();
 FILLCELL_X32 FILLER_169_1520 ();
 FILLCELL_X32 FILLER_169_1552 ();
 FILLCELL_X32 FILLER_169_1584 ();
 FILLCELL_X32 FILLER_169_1616 ();
 FILLCELL_X32 FILLER_169_1648 ();
 FILLCELL_X32 FILLER_169_1680 ();
 FILLCELL_X32 FILLER_169_1712 ();
 FILLCELL_X32 FILLER_169_1744 ();
 FILLCELL_X32 FILLER_169_1776 ();
 FILLCELL_X32 FILLER_169_1808 ();
 FILLCELL_X32 FILLER_169_1840 ();
 FILLCELL_X32 FILLER_169_1872 ();
 FILLCELL_X32 FILLER_169_1904 ();
 FILLCELL_X32 FILLER_169_1936 ();
 FILLCELL_X32 FILLER_169_1968 ();
 FILLCELL_X32 FILLER_169_2000 ();
 FILLCELL_X32 FILLER_169_2032 ();
 FILLCELL_X32 FILLER_169_2064 ();
 FILLCELL_X32 FILLER_169_2096 ();
 FILLCELL_X32 FILLER_169_2128 ();
 FILLCELL_X32 FILLER_169_2160 ();
 FILLCELL_X32 FILLER_169_2192 ();
 FILLCELL_X32 FILLER_169_2224 ();
 FILLCELL_X32 FILLER_169_2256 ();
 FILLCELL_X32 FILLER_169_2288 ();
 FILLCELL_X32 FILLER_169_2320 ();
 FILLCELL_X32 FILLER_169_2352 ();
 FILLCELL_X32 FILLER_169_2384 ();
 FILLCELL_X32 FILLER_169_2416 ();
 FILLCELL_X32 FILLER_169_2448 ();
 FILLCELL_X32 FILLER_169_2480 ();
 FILLCELL_X8 FILLER_169_2512 ();
 FILLCELL_X4 FILLER_169_2520 ();
 FILLCELL_X2 FILLER_169_2524 ();
 FILLCELL_X32 FILLER_169_2527 ();
 FILLCELL_X32 FILLER_169_2559 ();
 FILLCELL_X32 FILLER_169_2591 ();
 FILLCELL_X32 FILLER_169_2623 ();
 FILLCELL_X32 FILLER_169_2655 ();
 FILLCELL_X32 FILLER_169_2687 ();
 FILLCELL_X32 FILLER_169_2719 ();
 FILLCELL_X32 FILLER_169_2751 ();
 FILLCELL_X32 FILLER_169_2783 ();
 FILLCELL_X32 FILLER_169_2815 ();
 FILLCELL_X32 FILLER_169_2847 ();
 FILLCELL_X32 FILLER_169_2879 ();
 FILLCELL_X32 FILLER_169_2911 ();
 FILLCELL_X32 FILLER_169_2943 ();
 FILLCELL_X32 FILLER_169_2975 ();
 FILLCELL_X32 FILLER_169_3007 ();
 FILLCELL_X32 FILLER_169_3039 ();
 FILLCELL_X32 FILLER_169_3071 ();
 FILLCELL_X32 FILLER_169_3103 ();
 FILLCELL_X32 FILLER_169_3135 ();
 FILLCELL_X32 FILLER_169_3167 ();
 FILLCELL_X32 FILLER_169_3199 ();
 FILLCELL_X32 FILLER_169_3231 ();
 FILLCELL_X32 FILLER_169_3263 ();
 FILLCELL_X32 FILLER_169_3295 ();
 FILLCELL_X32 FILLER_169_3327 ();
 FILLCELL_X32 FILLER_169_3359 ();
 FILLCELL_X32 FILLER_169_3391 ();
 FILLCELL_X32 FILLER_169_3423 ();
 FILLCELL_X32 FILLER_169_3455 ();
 FILLCELL_X32 FILLER_169_3487 ();
 FILLCELL_X32 FILLER_169_3519 ();
 FILLCELL_X32 FILLER_169_3551 ();
 FILLCELL_X32 FILLER_169_3583 ();
 FILLCELL_X32 FILLER_169_3615 ();
 FILLCELL_X32 FILLER_169_3647 ();
 FILLCELL_X32 FILLER_169_3679 ();
 FILLCELL_X16 FILLER_169_3711 ();
 FILLCELL_X8 FILLER_169_3727 ();
 FILLCELL_X2 FILLER_169_3735 ();
 FILLCELL_X1 FILLER_169_3737 ();
 FILLCELL_X32 FILLER_170_1 ();
 FILLCELL_X32 FILLER_170_33 ();
 FILLCELL_X32 FILLER_170_65 ();
 FILLCELL_X32 FILLER_170_97 ();
 FILLCELL_X32 FILLER_170_129 ();
 FILLCELL_X32 FILLER_170_161 ();
 FILLCELL_X32 FILLER_170_193 ();
 FILLCELL_X32 FILLER_170_225 ();
 FILLCELL_X32 FILLER_170_257 ();
 FILLCELL_X32 FILLER_170_289 ();
 FILLCELL_X32 FILLER_170_321 ();
 FILLCELL_X32 FILLER_170_353 ();
 FILLCELL_X32 FILLER_170_385 ();
 FILLCELL_X32 FILLER_170_417 ();
 FILLCELL_X32 FILLER_170_449 ();
 FILLCELL_X32 FILLER_170_481 ();
 FILLCELL_X32 FILLER_170_513 ();
 FILLCELL_X32 FILLER_170_545 ();
 FILLCELL_X32 FILLER_170_577 ();
 FILLCELL_X16 FILLER_170_609 ();
 FILLCELL_X4 FILLER_170_625 ();
 FILLCELL_X2 FILLER_170_629 ();
 FILLCELL_X32 FILLER_170_632 ();
 FILLCELL_X32 FILLER_170_664 ();
 FILLCELL_X32 FILLER_170_696 ();
 FILLCELL_X32 FILLER_170_728 ();
 FILLCELL_X32 FILLER_170_760 ();
 FILLCELL_X32 FILLER_170_792 ();
 FILLCELL_X32 FILLER_170_824 ();
 FILLCELL_X32 FILLER_170_856 ();
 FILLCELL_X32 FILLER_170_888 ();
 FILLCELL_X32 FILLER_170_920 ();
 FILLCELL_X32 FILLER_170_952 ();
 FILLCELL_X32 FILLER_170_984 ();
 FILLCELL_X32 FILLER_170_1016 ();
 FILLCELL_X32 FILLER_170_1048 ();
 FILLCELL_X32 FILLER_170_1080 ();
 FILLCELL_X32 FILLER_170_1112 ();
 FILLCELL_X32 FILLER_170_1144 ();
 FILLCELL_X32 FILLER_170_1176 ();
 FILLCELL_X32 FILLER_170_1208 ();
 FILLCELL_X32 FILLER_170_1240 ();
 FILLCELL_X32 FILLER_170_1272 ();
 FILLCELL_X32 FILLER_170_1304 ();
 FILLCELL_X32 FILLER_170_1336 ();
 FILLCELL_X32 FILLER_170_1368 ();
 FILLCELL_X32 FILLER_170_1400 ();
 FILLCELL_X32 FILLER_170_1432 ();
 FILLCELL_X32 FILLER_170_1464 ();
 FILLCELL_X32 FILLER_170_1496 ();
 FILLCELL_X32 FILLER_170_1528 ();
 FILLCELL_X32 FILLER_170_1560 ();
 FILLCELL_X32 FILLER_170_1592 ();
 FILLCELL_X32 FILLER_170_1624 ();
 FILLCELL_X32 FILLER_170_1656 ();
 FILLCELL_X32 FILLER_170_1688 ();
 FILLCELL_X32 FILLER_170_1720 ();
 FILLCELL_X32 FILLER_170_1752 ();
 FILLCELL_X32 FILLER_170_1784 ();
 FILLCELL_X32 FILLER_170_1816 ();
 FILLCELL_X32 FILLER_170_1848 ();
 FILLCELL_X8 FILLER_170_1880 ();
 FILLCELL_X4 FILLER_170_1888 ();
 FILLCELL_X2 FILLER_170_1892 ();
 FILLCELL_X32 FILLER_170_1895 ();
 FILLCELL_X32 FILLER_170_1927 ();
 FILLCELL_X32 FILLER_170_1959 ();
 FILLCELL_X32 FILLER_170_1991 ();
 FILLCELL_X32 FILLER_170_2023 ();
 FILLCELL_X32 FILLER_170_2055 ();
 FILLCELL_X32 FILLER_170_2087 ();
 FILLCELL_X32 FILLER_170_2119 ();
 FILLCELL_X32 FILLER_170_2151 ();
 FILLCELL_X32 FILLER_170_2183 ();
 FILLCELL_X32 FILLER_170_2215 ();
 FILLCELL_X32 FILLER_170_2247 ();
 FILLCELL_X32 FILLER_170_2279 ();
 FILLCELL_X32 FILLER_170_2311 ();
 FILLCELL_X32 FILLER_170_2343 ();
 FILLCELL_X32 FILLER_170_2375 ();
 FILLCELL_X32 FILLER_170_2407 ();
 FILLCELL_X32 FILLER_170_2439 ();
 FILLCELL_X32 FILLER_170_2471 ();
 FILLCELL_X32 FILLER_170_2503 ();
 FILLCELL_X32 FILLER_170_2535 ();
 FILLCELL_X32 FILLER_170_2567 ();
 FILLCELL_X32 FILLER_170_2599 ();
 FILLCELL_X32 FILLER_170_2631 ();
 FILLCELL_X32 FILLER_170_2663 ();
 FILLCELL_X32 FILLER_170_2695 ();
 FILLCELL_X32 FILLER_170_2727 ();
 FILLCELL_X32 FILLER_170_2759 ();
 FILLCELL_X32 FILLER_170_2791 ();
 FILLCELL_X32 FILLER_170_2823 ();
 FILLCELL_X32 FILLER_170_2855 ();
 FILLCELL_X32 FILLER_170_2887 ();
 FILLCELL_X32 FILLER_170_2919 ();
 FILLCELL_X32 FILLER_170_2951 ();
 FILLCELL_X32 FILLER_170_2983 ();
 FILLCELL_X32 FILLER_170_3015 ();
 FILLCELL_X32 FILLER_170_3047 ();
 FILLCELL_X32 FILLER_170_3079 ();
 FILLCELL_X32 FILLER_170_3111 ();
 FILLCELL_X8 FILLER_170_3143 ();
 FILLCELL_X4 FILLER_170_3151 ();
 FILLCELL_X2 FILLER_170_3155 ();
 FILLCELL_X32 FILLER_170_3158 ();
 FILLCELL_X32 FILLER_170_3190 ();
 FILLCELL_X32 FILLER_170_3222 ();
 FILLCELL_X32 FILLER_170_3254 ();
 FILLCELL_X32 FILLER_170_3286 ();
 FILLCELL_X32 FILLER_170_3318 ();
 FILLCELL_X32 FILLER_170_3350 ();
 FILLCELL_X32 FILLER_170_3382 ();
 FILLCELL_X32 FILLER_170_3414 ();
 FILLCELL_X32 FILLER_170_3446 ();
 FILLCELL_X32 FILLER_170_3478 ();
 FILLCELL_X32 FILLER_170_3510 ();
 FILLCELL_X32 FILLER_170_3542 ();
 FILLCELL_X32 FILLER_170_3574 ();
 FILLCELL_X32 FILLER_170_3606 ();
 FILLCELL_X32 FILLER_170_3638 ();
 FILLCELL_X32 FILLER_170_3670 ();
 FILLCELL_X32 FILLER_170_3702 ();
 FILLCELL_X4 FILLER_170_3734 ();
 FILLCELL_X32 FILLER_171_1 ();
 FILLCELL_X32 FILLER_171_33 ();
 FILLCELL_X32 FILLER_171_65 ();
 FILLCELL_X32 FILLER_171_97 ();
 FILLCELL_X32 FILLER_171_129 ();
 FILLCELL_X32 FILLER_171_161 ();
 FILLCELL_X32 FILLER_171_193 ();
 FILLCELL_X32 FILLER_171_225 ();
 FILLCELL_X32 FILLER_171_257 ();
 FILLCELL_X32 FILLER_171_289 ();
 FILLCELL_X32 FILLER_171_321 ();
 FILLCELL_X32 FILLER_171_353 ();
 FILLCELL_X32 FILLER_171_385 ();
 FILLCELL_X32 FILLER_171_417 ();
 FILLCELL_X32 FILLER_171_449 ();
 FILLCELL_X32 FILLER_171_481 ();
 FILLCELL_X32 FILLER_171_513 ();
 FILLCELL_X32 FILLER_171_545 ();
 FILLCELL_X32 FILLER_171_577 ();
 FILLCELL_X32 FILLER_171_609 ();
 FILLCELL_X32 FILLER_171_641 ();
 FILLCELL_X32 FILLER_171_673 ();
 FILLCELL_X32 FILLER_171_705 ();
 FILLCELL_X32 FILLER_171_737 ();
 FILLCELL_X32 FILLER_171_769 ();
 FILLCELL_X32 FILLER_171_801 ();
 FILLCELL_X32 FILLER_171_833 ();
 FILLCELL_X32 FILLER_171_865 ();
 FILLCELL_X32 FILLER_171_897 ();
 FILLCELL_X32 FILLER_171_929 ();
 FILLCELL_X32 FILLER_171_961 ();
 FILLCELL_X32 FILLER_171_993 ();
 FILLCELL_X32 FILLER_171_1025 ();
 FILLCELL_X32 FILLER_171_1057 ();
 FILLCELL_X32 FILLER_171_1089 ();
 FILLCELL_X32 FILLER_171_1121 ();
 FILLCELL_X32 FILLER_171_1153 ();
 FILLCELL_X32 FILLER_171_1185 ();
 FILLCELL_X32 FILLER_171_1217 ();
 FILLCELL_X8 FILLER_171_1249 ();
 FILLCELL_X4 FILLER_171_1257 ();
 FILLCELL_X2 FILLER_171_1261 ();
 FILLCELL_X32 FILLER_171_1264 ();
 FILLCELL_X32 FILLER_171_1296 ();
 FILLCELL_X32 FILLER_171_1328 ();
 FILLCELL_X32 FILLER_171_1360 ();
 FILLCELL_X32 FILLER_171_1392 ();
 FILLCELL_X32 FILLER_171_1424 ();
 FILLCELL_X32 FILLER_171_1456 ();
 FILLCELL_X32 FILLER_171_1488 ();
 FILLCELL_X32 FILLER_171_1520 ();
 FILLCELL_X32 FILLER_171_1552 ();
 FILLCELL_X32 FILLER_171_1584 ();
 FILLCELL_X32 FILLER_171_1616 ();
 FILLCELL_X32 FILLER_171_1648 ();
 FILLCELL_X32 FILLER_171_1680 ();
 FILLCELL_X32 FILLER_171_1712 ();
 FILLCELL_X32 FILLER_171_1744 ();
 FILLCELL_X32 FILLER_171_1776 ();
 FILLCELL_X32 FILLER_171_1808 ();
 FILLCELL_X32 FILLER_171_1840 ();
 FILLCELL_X32 FILLER_171_1872 ();
 FILLCELL_X32 FILLER_171_1904 ();
 FILLCELL_X32 FILLER_171_1936 ();
 FILLCELL_X32 FILLER_171_1968 ();
 FILLCELL_X32 FILLER_171_2000 ();
 FILLCELL_X32 FILLER_171_2032 ();
 FILLCELL_X32 FILLER_171_2064 ();
 FILLCELL_X32 FILLER_171_2096 ();
 FILLCELL_X32 FILLER_171_2128 ();
 FILLCELL_X32 FILLER_171_2160 ();
 FILLCELL_X32 FILLER_171_2192 ();
 FILLCELL_X32 FILLER_171_2224 ();
 FILLCELL_X32 FILLER_171_2256 ();
 FILLCELL_X32 FILLER_171_2288 ();
 FILLCELL_X32 FILLER_171_2320 ();
 FILLCELL_X32 FILLER_171_2352 ();
 FILLCELL_X32 FILLER_171_2384 ();
 FILLCELL_X32 FILLER_171_2416 ();
 FILLCELL_X32 FILLER_171_2448 ();
 FILLCELL_X32 FILLER_171_2480 ();
 FILLCELL_X8 FILLER_171_2512 ();
 FILLCELL_X4 FILLER_171_2520 ();
 FILLCELL_X2 FILLER_171_2524 ();
 FILLCELL_X32 FILLER_171_2527 ();
 FILLCELL_X32 FILLER_171_2559 ();
 FILLCELL_X32 FILLER_171_2591 ();
 FILLCELL_X32 FILLER_171_2623 ();
 FILLCELL_X32 FILLER_171_2655 ();
 FILLCELL_X32 FILLER_171_2687 ();
 FILLCELL_X32 FILLER_171_2719 ();
 FILLCELL_X32 FILLER_171_2751 ();
 FILLCELL_X32 FILLER_171_2783 ();
 FILLCELL_X32 FILLER_171_2815 ();
 FILLCELL_X32 FILLER_171_2847 ();
 FILLCELL_X32 FILLER_171_2879 ();
 FILLCELL_X32 FILLER_171_2911 ();
 FILLCELL_X32 FILLER_171_2943 ();
 FILLCELL_X32 FILLER_171_2975 ();
 FILLCELL_X32 FILLER_171_3007 ();
 FILLCELL_X32 FILLER_171_3039 ();
 FILLCELL_X32 FILLER_171_3071 ();
 FILLCELL_X32 FILLER_171_3103 ();
 FILLCELL_X32 FILLER_171_3135 ();
 FILLCELL_X32 FILLER_171_3167 ();
 FILLCELL_X32 FILLER_171_3199 ();
 FILLCELL_X32 FILLER_171_3231 ();
 FILLCELL_X32 FILLER_171_3263 ();
 FILLCELL_X32 FILLER_171_3295 ();
 FILLCELL_X32 FILLER_171_3327 ();
 FILLCELL_X32 FILLER_171_3359 ();
 FILLCELL_X32 FILLER_171_3391 ();
 FILLCELL_X32 FILLER_171_3423 ();
 FILLCELL_X32 FILLER_171_3455 ();
 FILLCELL_X32 FILLER_171_3487 ();
 FILLCELL_X32 FILLER_171_3519 ();
 FILLCELL_X32 FILLER_171_3551 ();
 FILLCELL_X32 FILLER_171_3583 ();
 FILLCELL_X32 FILLER_171_3615 ();
 FILLCELL_X32 FILLER_171_3647 ();
 FILLCELL_X32 FILLER_171_3679 ();
 FILLCELL_X16 FILLER_171_3711 ();
 FILLCELL_X8 FILLER_171_3727 ();
 FILLCELL_X2 FILLER_171_3735 ();
 FILLCELL_X1 FILLER_171_3737 ();
 FILLCELL_X32 FILLER_172_1 ();
 FILLCELL_X32 FILLER_172_33 ();
 FILLCELL_X32 FILLER_172_65 ();
 FILLCELL_X32 FILLER_172_97 ();
 FILLCELL_X32 FILLER_172_129 ();
 FILLCELL_X32 FILLER_172_161 ();
 FILLCELL_X32 FILLER_172_193 ();
 FILLCELL_X32 FILLER_172_225 ();
 FILLCELL_X32 FILLER_172_257 ();
 FILLCELL_X32 FILLER_172_289 ();
 FILLCELL_X32 FILLER_172_321 ();
 FILLCELL_X32 FILLER_172_353 ();
 FILLCELL_X32 FILLER_172_385 ();
 FILLCELL_X32 FILLER_172_417 ();
 FILLCELL_X32 FILLER_172_449 ();
 FILLCELL_X32 FILLER_172_481 ();
 FILLCELL_X32 FILLER_172_513 ();
 FILLCELL_X32 FILLER_172_545 ();
 FILLCELL_X32 FILLER_172_577 ();
 FILLCELL_X16 FILLER_172_609 ();
 FILLCELL_X4 FILLER_172_625 ();
 FILLCELL_X2 FILLER_172_629 ();
 FILLCELL_X32 FILLER_172_632 ();
 FILLCELL_X32 FILLER_172_664 ();
 FILLCELL_X32 FILLER_172_696 ();
 FILLCELL_X32 FILLER_172_728 ();
 FILLCELL_X32 FILLER_172_760 ();
 FILLCELL_X32 FILLER_172_792 ();
 FILLCELL_X32 FILLER_172_824 ();
 FILLCELL_X32 FILLER_172_856 ();
 FILLCELL_X32 FILLER_172_888 ();
 FILLCELL_X32 FILLER_172_920 ();
 FILLCELL_X32 FILLER_172_952 ();
 FILLCELL_X32 FILLER_172_984 ();
 FILLCELL_X32 FILLER_172_1016 ();
 FILLCELL_X32 FILLER_172_1048 ();
 FILLCELL_X32 FILLER_172_1080 ();
 FILLCELL_X32 FILLER_172_1112 ();
 FILLCELL_X32 FILLER_172_1144 ();
 FILLCELL_X32 FILLER_172_1176 ();
 FILLCELL_X32 FILLER_172_1208 ();
 FILLCELL_X32 FILLER_172_1240 ();
 FILLCELL_X32 FILLER_172_1272 ();
 FILLCELL_X32 FILLER_172_1304 ();
 FILLCELL_X32 FILLER_172_1336 ();
 FILLCELL_X32 FILLER_172_1368 ();
 FILLCELL_X32 FILLER_172_1400 ();
 FILLCELL_X32 FILLER_172_1432 ();
 FILLCELL_X32 FILLER_172_1464 ();
 FILLCELL_X32 FILLER_172_1496 ();
 FILLCELL_X32 FILLER_172_1528 ();
 FILLCELL_X32 FILLER_172_1560 ();
 FILLCELL_X32 FILLER_172_1592 ();
 FILLCELL_X32 FILLER_172_1624 ();
 FILLCELL_X32 FILLER_172_1656 ();
 FILLCELL_X32 FILLER_172_1688 ();
 FILLCELL_X32 FILLER_172_1720 ();
 FILLCELL_X32 FILLER_172_1752 ();
 FILLCELL_X32 FILLER_172_1784 ();
 FILLCELL_X32 FILLER_172_1816 ();
 FILLCELL_X32 FILLER_172_1848 ();
 FILLCELL_X8 FILLER_172_1880 ();
 FILLCELL_X4 FILLER_172_1888 ();
 FILLCELL_X2 FILLER_172_1892 ();
 FILLCELL_X32 FILLER_172_1895 ();
 FILLCELL_X32 FILLER_172_1927 ();
 FILLCELL_X32 FILLER_172_1959 ();
 FILLCELL_X32 FILLER_172_1991 ();
 FILLCELL_X32 FILLER_172_2023 ();
 FILLCELL_X32 FILLER_172_2055 ();
 FILLCELL_X32 FILLER_172_2087 ();
 FILLCELL_X32 FILLER_172_2119 ();
 FILLCELL_X32 FILLER_172_2151 ();
 FILLCELL_X32 FILLER_172_2183 ();
 FILLCELL_X32 FILLER_172_2215 ();
 FILLCELL_X32 FILLER_172_2247 ();
 FILLCELL_X32 FILLER_172_2279 ();
 FILLCELL_X32 FILLER_172_2311 ();
 FILLCELL_X32 FILLER_172_2343 ();
 FILLCELL_X32 FILLER_172_2375 ();
 FILLCELL_X32 FILLER_172_2407 ();
 FILLCELL_X32 FILLER_172_2439 ();
 FILLCELL_X32 FILLER_172_2471 ();
 FILLCELL_X32 FILLER_172_2503 ();
 FILLCELL_X32 FILLER_172_2535 ();
 FILLCELL_X32 FILLER_172_2567 ();
 FILLCELL_X32 FILLER_172_2599 ();
 FILLCELL_X32 FILLER_172_2631 ();
 FILLCELL_X32 FILLER_172_2663 ();
 FILLCELL_X32 FILLER_172_2695 ();
 FILLCELL_X32 FILLER_172_2727 ();
 FILLCELL_X32 FILLER_172_2759 ();
 FILLCELL_X32 FILLER_172_2791 ();
 FILLCELL_X32 FILLER_172_2823 ();
 FILLCELL_X32 FILLER_172_2855 ();
 FILLCELL_X32 FILLER_172_2887 ();
 FILLCELL_X32 FILLER_172_2919 ();
 FILLCELL_X32 FILLER_172_2951 ();
 FILLCELL_X32 FILLER_172_2983 ();
 FILLCELL_X32 FILLER_172_3015 ();
 FILLCELL_X32 FILLER_172_3047 ();
 FILLCELL_X32 FILLER_172_3079 ();
 FILLCELL_X32 FILLER_172_3111 ();
 FILLCELL_X8 FILLER_172_3143 ();
 FILLCELL_X4 FILLER_172_3151 ();
 FILLCELL_X2 FILLER_172_3155 ();
 FILLCELL_X32 FILLER_172_3158 ();
 FILLCELL_X32 FILLER_172_3190 ();
 FILLCELL_X32 FILLER_172_3222 ();
 FILLCELL_X32 FILLER_172_3254 ();
 FILLCELL_X32 FILLER_172_3286 ();
 FILLCELL_X32 FILLER_172_3318 ();
 FILLCELL_X32 FILLER_172_3350 ();
 FILLCELL_X32 FILLER_172_3382 ();
 FILLCELL_X32 FILLER_172_3414 ();
 FILLCELL_X32 FILLER_172_3446 ();
 FILLCELL_X32 FILLER_172_3478 ();
 FILLCELL_X32 FILLER_172_3510 ();
 FILLCELL_X32 FILLER_172_3542 ();
 FILLCELL_X32 FILLER_172_3574 ();
 FILLCELL_X32 FILLER_172_3606 ();
 FILLCELL_X32 FILLER_172_3638 ();
 FILLCELL_X32 FILLER_172_3670 ();
 FILLCELL_X32 FILLER_172_3702 ();
 FILLCELL_X4 FILLER_172_3734 ();
 FILLCELL_X32 FILLER_173_1 ();
 FILLCELL_X32 FILLER_173_33 ();
 FILLCELL_X32 FILLER_173_65 ();
 FILLCELL_X32 FILLER_173_97 ();
 FILLCELL_X32 FILLER_173_129 ();
 FILLCELL_X32 FILLER_173_161 ();
 FILLCELL_X32 FILLER_173_193 ();
 FILLCELL_X32 FILLER_173_225 ();
 FILLCELL_X32 FILLER_173_257 ();
 FILLCELL_X32 FILLER_173_289 ();
 FILLCELL_X32 FILLER_173_321 ();
 FILLCELL_X32 FILLER_173_353 ();
 FILLCELL_X32 FILLER_173_385 ();
 FILLCELL_X32 FILLER_173_417 ();
 FILLCELL_X32 FILLER_173_449 ();
 FILLCELL_X32 FILLER_173_481 ();
 FILLCELL_X32 FILLER_173_513 ();
 FILLCELL_X32 FILLER_173_545 ();
 FILLCELL_X32 FILLER_173_577 ();
 FILLCELL_X32 FILLER_173_609 ();
 FILLCELL_X32 FILLER_173_641 ();
 FILLCELL_X32 FILLER_173_673 ();
 FILLCELL_X32 FILLER_173_705 ();
 FILLCELL_X32 FILLER_173_737 ();
 FILLCELL_X32 FILLER_173_769 ();
 FILLCELL_X32 FILLER_173_801 ();
 FILLCELL_X32 FILLER_173_833 ();
 FILLCELL_X32 FILLER_173_865 ();
 FILLCELL_X32 FILLER_173_897 ();
 FILLCELL_X32 FILLER_173_929 ();
 FILLCELL_X32 FILLER_173_961 ();
 FILLCELL_X32 FILLER_173_993 ();
 FILLCELL_X32 FILLER_173_1025 ();
 FILLCELL_X32 FILLER_173_1057 ();
 FILLCELL_X32 FILLER_173_1089 ();
 FILLCELL_X32 FILLER_173_1121 ();
 FILLCELL_X32 FILLER_173_1153 ();
 FILLCELL_X32 FILLER_173_1185 ();
 FILLCELL_X32 FILLER_173_1217 ();
 FILLCELL_X8 FILLER_173_1249 ();
 FILLCELL_X4 FILLER_173_1257 ();
 FILLCELL_X2 FILLER_173_1261 ();
 FILLCELL_X32 FILLER_173_1264 ();
 FILLCELL_X32 FILLER_173_1296 ();
 FILLCELL_X32 FILLER_173_1328 ();
 FILLCELL_X32 FILLER_173_1360 ();
 FILLCELL_X32 FILLER_173_1392 ();
 FILLCELL_X32 FILLER_173_1424 ();
 FILLCELL_X32 FILLER_173_1456 ();
 FILLCELL_X32 FILLER_173_1488 ();
 FILLCELL_X32 FILLER_173_1520 ();
 FILLCELL_X32 FILLER_173_1552 ();
 FILLCELL_X32 FILLER_173_1584 ();
 FILLCELL_X32 FILLER_173_1616 ();
 FILLCELL_X32 FILLER_173_1648 ();
 FILLCELL_X32 FILLER_173_1680 ();
 FILLCELL_X32 FILLER_173_1712 ();
 FILLCELL_X32 FILLER_173_1744 ();
 FILLCELL_X32 FILLER_173_1776 ();
 FILLCELL_X32 FILLER_173_1808 ();
 FILLCELL_X32 FILLER_173_1840 ();
 FILLCELL_X32 FILLER_173_1872 ();
 FILLCELL_X32 FILLER_173_1904 ();
 FILLCELL_X32 FILLER_173_1936 ();
 FILLCELL_X32 FILLER_173_1968 ();
 FILLCELL_X32 FILLER_173_2000 ();
 FILLCELL_X32 FILLER_173_2032 ();
 FILLCELL_X32 FILLER_173_2064 ();
 FILLCELL_X32 FILLER_173_2096 ();
 FILLCELL_X32 FILLER_173_2128 ();
 FILLCELL_X32 FILLER_173_2160 ();
 FILLCELL_X32 FILLER_173_2192 ();
 FILLCELL_X32 FILLER_173_2224 ();
 FILLCELL_X32 FILLER_173_2256 ();
 FILLCELL_X32 FILLER_173_2288 ();
 FILLCELL_X32 FILLER_173_2320 ();
 FILLCELL_X32 FILLER_173_2352 ();
 FILLCELL_X32 FILLER_173_2384 ();
 FILLCELL_X32 FILLER_173_2416 ();
 FILLCELL_X32 FILLER_173_2448 ();
 FILLCELL_X32 FILLER_173_2480 ();
 FILLCELL_X8 FILLER_173_2512 ();
 FILLCELL_X4 FILLER_173_2520 ();
 FILLCELL_X2 FILLER_173_2524 ();
 FILLCELL_X32 FILLER_173_2527 ();
 FILLCELL_X32 FILLER_173_2559 ();
 FILLCELL_X32 FILLER_173_2591 ();
 FILLCELL_X32 FILLER_173_2623 ();
 FILLCELL_X32 FILLER_173_2655 ();
 FILLCELL_X32 FILLER_173_2687 ();
 FILLCELL_X32 FILLER_173_2719 ();
 FILLCELL_X32 FILLER_173_2751 ();
 FILLCELL_X32 FILLER_173_2783 ();
 FILLCELL_X32 FILLER_173_2815 ();
 FILLCELL_X32 FILLER_173_2847 ();
 FILLCELL_X32 FILLER_173_2879 ();
 FILLCELL_X32 FILLER_173_2911 ();
 FILLCELL_X32 FILLER_173_2943 ();
 FILLCELL_X32 FILLER_173_2975 ();
 FILLCELL_X32 FILLER_173_3007 ();
 FILLCELL_X32 FILLER_173_3039 ();
 FILLCELL_X32 FILLER_173_3071 ();
 FILLCELL_X32 FILLER_173_3103 ();
 FILLCELL_X32 FILLER_173_3135 ();
 FILLCELL_X32 FILLER_173_3167 ();
 FILLCELL_X32 FILLER_173_3199 ();
 FILLCELL_X32 FILLER_173_3231 ();
 FILLCELL_X32 FILLER_173_3263 ();
 FILLCELL_X32 FILLER_173_3295 ();
 FILLCELL_X32 FILLER_173_3327 ();
 FILLCELL_X32 FILLER_173_3359 ();
 FILLCELL_X32 FILLER_173_3391 ();
 FILLCELL_X32 FILLER_173_3423 ();
 FILLCELL_X32 FILLER_173_3455 ();
 FILLCELL_X32 FILLER_173_3487 ();
 FILLCELL_X32 FILLER_173_3519 ();
 FILLCELL_X32 FILLER_173_3551 ();
 FILLCELL_X32 FILLER_173_3583 ();
 FILLCELL_X32 FILLER_173_3615 ();
 FILLCELL_X32 FILLER_173_3647 ();
 FILLCELL_X32 FILLER_173_3679 ();
 FILLCELL_X16 FILLER_173_3711 ();
 FILLCELL_X8 FILLER_173_3727 ();
 FILLCELL_X2 FILLER_173_3735 ();
 FILLCELL_X1 FILLER_173_3737 ();
 FILLCELL_X32 FILLER_174_1 ();
 FILLCELL_X32 FILLER_174_33 ();
 FILLCELL_X32 FILLER_174_65 ();
 FILLCELL_X32 FILLER_174_97 ();
 FILLCELL_X32 FILLER_174_129 ();
 FILLCELL_X32 FILLER_174_161 ();
 FILLCELL_X32 FILLER_174_193 ();
 FILLCELL_X32 FILLER_174_225 ();
 FILLCELL_X32 FILLER_174_257 ();
 FILLCELL_X32 FILLER_174_289 ();
 FILLCELL_X32 FILLER_174_321 ();
 FILLCELL_X32 FILLER_174_353 ();
 FILLCELL_X32 FILLER_174_385 ();
 FILLCELL_X32 FILLER_174_417 ();
 FILLCELL_X32 FILLER_174_449 ();
 FILLCELL_X32 FILLER_174_481 ();
 FILLCELL_X32 FILLER_174_513 ();
 FILLCELL_X32 FILLER_174_545 ();
 FILLCELL_X32 FILLER_174_577 ();
 FILLCELL_X16 FILLER_174_609 ();
 FILLCELL_X4 FILLER_174_625 ();
 FILLCELL_X2 FILLER_174_629 ();
 FILLCELL_X32 FILLER_174_632 ();
 FILLCELL_X32 FILLER_174_664 ();
 FILLCELL_X32 FILLER_174_696 ();
 FILLCELL_X32 FILLER_174_728 ();
 FILLCELL_X32 FILLER_174_760 ();
 FILLCELL_X32 FILLER_174_792 ();
 FILLCELL_X32 FILLER_174_824 ();
 FILLCELL_X32 FILLER_174_856 ();
 FILLCELL_X32 FILLER_174_888 ();
 FILLCELL_X32 FILLER_174_920 ();
 FILLCELL_X32 FILLER_174_952 ();
 FILLCELL_X32 FILLER_174_984 ();
 FILLCELL_X32 FILLER_174_1016 ();
 FILLCELL_X32 FILLER_174_1048 ();
 FILLCELL_X32 FILLER_174_1080 ();
 FILLCELL_X32 FILLER_174_1112 ();
 FILLCELL_X32 FILLER_174_1144 ();
 FILLCELL_X32 FILLER_174_1176 ();
 FILLCELL_X32 FILLER_174_1208 ();
 FILLCELL_X32 FILLER_174_1240 ();
 FILLCELL_X32 FILLER_174_1272 ();
 FILLCELL_X32 FILLER_174_1304 ();
 FILLCELL_X32 FILLER_174_1336 ();
 FILLCELL_X32 FILLER_174_1368 ();
 FILLCELL_X32 FILLER_174_1400 ();
 FILLCELL_X32 FILLER_174_1432 ();
 FILLCELL_X32 FILLER_174_1464 ();
 FILLCELL_X32 FILLER_174_1496 ();
 FILLCELL_X32 FILLER_174_1528 ();
 FILLCELL_X32 FILLER_174_1560 ();
 FILLCELL_X32 FILLER_174_1592 ();
 FILLCELL_X32 FILLER_174_1624 ();
 FILLCELL_X32 FILLER_174_1656 ();
 FILLCELL_X32 FILLER_174_1688 ();
 FILLCELL_X32 FILLER_174_1720 ();
 FILLCELL_X32 FILLER_174_1752 ();
 FILLCELL_X32 FILLER_174_1784 ();
 FILLCELL_X32 FILLER_174_1816 ();
 FILLCELL_X32 FILLER_174_1848 ();
 FILLCELL_X8 FILLER_174_1880 ();
 FILLCELL_X4 FILLER_174_1888 ();
 FILLCELL_X2 FILLER_174_1892 ();
 FILLCELL_X32 FILLER_174_1895 ();
 FILLCELL_X32 FILLER_174_1927 ();
 FILLCELL_X32 FILLER_174_1959 ();
 FILLCELL_X32 FILLER_174_1991 ();
 FILLCELL_X32 FILLER_174_2023 ();
 FILLCELL_X32 FILLER_174_2055 ();
 FILLCELL_X32 FILLER_174_2087 ();
 FILLCELL_X32 FILLER_174_2119 ();
 FILLCELL_X32 FILLER_174_2151 ();
 FILLCELL_X32 FILLER_174_2183 ();
 FILLCELL_X32 FILLER_174_2215 ();
 FILLCELL_X32 FILLER_174_2247 ();
 FILLCELL_X32 FILLER_174_2279 ();
 FILLCELL_X32 FILLER_174_2311 ();
 FILLCELL_X32 FILLER_174_2343 ();
 FILLCELL_X32 FILLER_174_2375 ();
 FILLCELL_X32 FILLER_174_2407 ();
 FILLCELL_X32 FILLER_174_2439 ();
 FILLCELL_X32 FILLER_174_2471 ();
 FILLCELL_X32 FILLER_174_2503 ();
 FILLCELL_X32 FILLER_174_2535 ();
 FILLCELL_X32 FILLER_174_2567 ();
 FILLCELL_X32 FILLER_174_2599 ();
 FILLCELL_X32 FILLER_174_2631 ();
 FILLCELL_X32 FILLER_174_2663 ();
 FILLCELL_X32 FILLER_174_2695 ();
 FILLCELL_X32 FILLER_174_2727 ();
 FILLCELL_X32 FILLER_174_2759 ();
 FILLCELL_X32 FILLER_174_2791 ();
 FILLCELL_X32 FILLER_174_2823 ();
 FILLCELL_X32 FILLER_174_2855 ();
 FILLCELL_X32 FILLER_174_2887 ();
 FILLCELL_X32 FILLER_174_2919 ();
 FILLCELL_X32 FILLER_174_2951 ();
 FILLCELL_X32 FILLER_174_2983 ();
 FILLCELL_X32 FILLER_174_3015 ();
 FILLCELL_X32 FILLER_174_3047 ();
 FILLCELL_X32 FILLER_174_3079 ();
 FILLCELL_X32 FILLER_174_3111 ();
 FILLCELL_X8 FILLER_174_3143 ();
 FILLCELL_X4 FILLER_174_3151 ();
 FILLCELL_X2 FILLER_174_3155 ();
 FILLCELL_X32 FILLER_174_3158 ();
 FILLCELL_X32 FILLER_174_3190 ();
 FILLCELL_X32 FILLER_174_3222 ();
 FILLCELL_X32 FILLER_174_3254 ();
 FILLCELL_X32 FILLER_174_3286 ();
 FILLCELL_X32 FILLER_174_3318 ();
 FILLCELL_X32 FILLER_174_3350 ();
 FILLCELL_X32 FILLER_174_3382 ();
 FILLCELL_X32 FILLER_174_3414 ();
 FILLCELL_X32 FILLER_174_3446 ();
 FILLCELL_X32 FILLER_174_3478 ();
 FILLCELL_X32 FILLER_174_3510 ();
 FILLCELL_X32 FILLER_174_3542 ();
 FILLCELL_X32 FILLER_174_3574 ();
 FILLCELL_X32 FILLER_174_3606 ();
 FILLCELL_X32 FILLER_174_3638 ();
 FILLCELL_X32 FILLER_174_3670 ();
 FILLCELL_X32 FILLER_174_3702 ();
 FILLCELL_X4 FILLER_174_3734 ();
 FILLCELL_X32 FILLER_175_1 ();
 FILLCELL_X32 FILLER_175_33 ();
 FILLCELL_X32 FILLER_175_65 ();
 FILLCELL_X32 FILLER_175_97 ();
 FILLCELL_X32 FILLER_175_129 ();
 FILLCELL_X32 FILLER_175_161 ();
 FILLCELL_X32 FILLER_175_193 ();
 FILLCELL_X32 FILLER_175_225 ();
 FILLCELL_X32 FILLER_175_257 ();
 FILLCELL_X32 FILLER_175_289 ();
 FILLCELL_X32 FILLER_175_321 ();
 FILLCELL_X32 FILLER_175_353 ();
 FILLCELL_X32 FILLER_175_385 ();
 FILLCELL_X32 FILLER_175_417 ();
 FILLCELL_X32 FILLER_175_449 ();
 FILLCELL_X32 FILLER_175_481 ();
 FILLCELL_X32 FILLER_175_513 ();
 FILLCELL_X32 FILLER_175_545 ();
 FILLCELL_X32 FILLER_175_577 ();
 FILLCELL_X32 FILLER_175_609 ();
 FILLCELL_X32 FILLER_175_641 ();
 FILLCELL_X32 FILLER_175_673 ();
 FILLCELL_X32 FILLER_175_705 ();
 FILLCELL_X32 FILLER_175_737 ();
 FILLCELL_X32 FILLER_175_769 ();
 FILLCELL_X32 FILLER_175_801 ();
 FILLCELL_X32 FILLER_175_833 ();
 FILLCELL_X32 FILLER_175_865 ();
 FILLCELL_X32 FILLER_175_897 ();
 FILLCELL_X32 FILLER_175_929 ();
 FILLCELL_X32 FILLER_175_961 ();
 FILLCELL_X32 FILLER_175_993 ();
 FILLCELL_X32 FILLER_175_1025 ();
 FILLCELL_X32 FILLER_175_1057 ();
 FILLCELL_X32 FILLER_175_1089 ();
 FILLCELL_X32 FILLER_175_1121 ();
 FILLCELL_X32 FILLER_175_1153 ();
 FILLCELL_X32 FILLER_175_1185 ();
 FILLCELL_X32 FILLER_175_1217 ();
 FILLCELL_X8 FILLER_175_1249 ();
 FILLCELL_X4 FILLER_175_1257 ();
 FILLCELL_X2 FILLER_175_1261 ();
 FILLCELL_X32 FILLER_175_1264 ();
 FILLCELL_X32 FILLER_175_1296 ();
 FILLCELL_X32 FILLER_175_1328 ();
 FILLCELL_X32 FILLER_175_1360 ();
 FILLCELL_X32 FILLER_175_1392 ();
 FILLCELL_X32 FILLER_175_1424 ();
 FILLCELL_X32 FILLER_175_1456 ();
 FILLCELL_X32 FILLER_175_1488 ();
 FILLCELL_X32 FILLER_175_1520 ();
 FILLCELL_X32 FILLER_175_1552 ();
 FILLCELL_X32 FILLER_175_1584 ();
 FILLCELL_X32 FILLER_175_1616 ();
 FILLCELL_X32 FILLER_175_1648 ();
 FILLCELL_X32 FILLER_175_1680 ();
 FILLCELL_X32 FILLER_175_1712 ();
 FILLCELL_X32 FILLER_175_1744 ();
 FILLCELL_X32 FILLER_175_1776 ();
 FILLCELL_X32 FILLER_175_1808 ();
 FILLCELL_X32 FILLER_175_1840 ();
 FILLCELL_X32 FILLER_175_1872 ();
 FILLCELL_X32 FILLER_175_1904 ();
 FILLCELL_X32 FILLER_175_1936 ();
 FILLCELL_X32 FILLER_175_1968 ();
 FILLCELL_X32 FILLER_175_2000 ();
 FILLCELL_X32 FILLER_175_2032 ();
 FILLCELL_X32 FILLER_175_2064 ();
 FILLCELL_X32 FILLER_175_2096 ();
 FILLCELL_X32 FILLER_175_2128 ();
 FILLCELL_X32 FILLER_175_2160 ();
 FILLCELL_X32 FILLER_175_2192 ();
 FILLCELL_X32 FILLER_175_2224 ();
 FILLCELL_X32 FILLER_175_2256 ();
 FILLCELL_X32 FILLER_175_2288 ();
 FILLCELL_X32 FILLER_175_2320 ();
 FILLCELL_X32 FILLER_175_2352 ();
 FILLCELL_X32 FILLER_175_2384 ();
 FILLCELL_X32 FILLER_175_2416 ();
 FILLCELL_X32 FILLER_175_2448 ();
 FILLCELL_X32 FILLER_175_2480 ();
 FILLCELL_X8 FILLER_175_2512 ();
 FILLCELL_X4 FILLER_175_2520 ();
 FILLCELL_X2 FILLER_175_2524 ();
 FILLCELL_X32 FILLER_175_2527 ();
 FILLCELL_X32 FILLER_175_2559 ();
 FILLCELL_X32 FILLER_175_2591 ();
 FILLCELL_X32 FILLER_175_2623 ();
 FILLCELL_X32 FILLER_175_2655 ();
 FILLCELL_X32 FILLER_175_2687 ();
 FILLCELL_X32 FILLER_175_2719 ();
 FILLCELL_X32 FILLER_175_2751 ();
 FILLCELL_X32 FILLER_175_2783 ();
 FILLCELL_X32 FILLER_175_2815 ();
 FILLCELL_X32 FILLER_175_2847 ();
 FILLCELL_X32 FILLER_175_2879 ();
 FILLCELL_X32 FILLER_175_2911 ();
 FILLCELL_X32 FILLER_175_2943 ();
 FILLCELL_X32 FILLER_175_2975 ();
 FILLCELL_X32 FILLER_175_3007 ();
 FILLCELL_X32 FILLER_175_3039 ();
 FILLCELL_X32 FILLER_175_3071 ();
 FILLCELL_X32 FILLER_175_3103 ();
 FILLCELL_X32 FILLER_175_3135 ();
 FILLCELL_X32 FILLER_175_3167 ();
 FILLCELL_X32 FILLER_175_3199 ();
 FILLCELL_X32 FILLER_175_3231 ();
 FILLCELL_X32 FILLER_175_3263 ();
 FILLCELL_X32 FILLER_175_3295 ();
 FILLCELL_X32 FILLER_175_3327 ();
 FILLCELL_X32 FILLER_175_3359 ();
 FILLCELL_X32 FILLER_175_3391 ();
 FILLCELL_X32 FILLER_175_3423 ();
 FILLCELL_X32 FILLER_175_3455 ();
 FILLCELL_X32 FILLER_175_3487 ();
 FILLCELL_X32 FILLER_175_3519 ();
 FILLCELL_X32 FILLER_175_3551 ();
 FILLCELL_X32 FILLER_175_3583 ();
 FILLCELL_X32 FILLER_175_3615 ();
 FILLCELL_X32 FILLER_175_3647 ();
 FILLCELL_X32 FILLER_175_3679 ();
 FILLCELL_X16 FILLER_175_3711 ();
 FILLCELL_X8 FILLER_175_3727 ();
 FILLCELL_X2 FILLER_175_3735 ();
 FILLCELL_X1 FILLER_175_3737 ();
 FILLCELL_X32 FILLER_176_1 ();
 FILLCELL_X32 FILLER_176_33 ();
 FILLCELL_X32 FILLER_176_65 ();
 FILLCELL_X32 FILLER_176_97 ();
 FILLCELL_X32 FILLER_176_129 ();
 FILLCELL_X32 FILLER_176_161 ();
 FILLCELL_X32 FILLER_176_193 ();
 FILLCELL_X32 FILLER_176_225 ();
 FILLCELL_X32 FILLER_176_257 ();
 FILLCELL_X32 FILLER_176_289 ();
 FILLCELL_X32 FILLER_176_321 ();
 FILLCELL_X32 FILLER_176_353 ();
 FILLCELL_X32 FILLER_176_385 ();
 FILLCELL_X32 FILLER_176_417 ();
 FILLCELL_X32 FILLER_176_449 ();
 FILLCELL_X32 FILLER_176_481 ();
 FILLCELL_X32 FILLER_176_513 ();
 FILLCELL_X32 FILLER_176_545 ();
 FILLCELL_X32 FILLER_176_577 ();
 FILLCELL_X16 FILLER_176_609 ();
 FILLCELL_X4 FILLER_176_625 ();
 FILLCELL_X2 FILLER_176_629 ();
 FILLCELL_X32 FILLER_176_632 ();
 FILLCELL_X32 FILLER_176_664 ();
 FILLCELL_X32 FILLER_176_696 ();
 FILLCELL_X32 FILLER_176_728 ();
 FILLCELL_X32 FILLER_176_760 ();
 FILLCELL_X32 FILLER_176_792 ();
 FILLCELL_X32 FILLER_176_824 ();
 FILLCELL_X32 FILLER_176_856 ();
 FILLCELL_X32 FILLER_176_888 ();
 FILLCELL_X32 FILLER_176_920 ();
 FILLCELL_X32 FILLER_176_952 ();
 FILLCELL_X32 FILLER_176_984 ();
 FILLCELL_X32 FILLER_176_1016 ();
 FILLCELL_X32 FILLER_176_1048 ();
 FILLCELL_X32 FILLER_176_1080 ();
 FILLCELL_X32 FILLER_176_1112 ();
 FILLCELL_X32 FILLER_176_1144 ();
 FILLCELL_X32 FILLER_176_1176 ();
 FILLCELL_X32 FILLER_176_1208 ();
 FILLCELL_X32 FILLER_176_1240 ();
 FILLCELL_X32 FILLER_176_1272 ();
 FILLCELL_X32 FILLER_176_1304 ();
 FILLCELL_X32 FILLER_176_1336 ();
 FILLCELL_X32 FILLER_176_1368 ();
 FILLCELL_X32 FILLER_176_1400 ();
 FILLCELL_X32 FILLER_176_1432 ();
 FILLCELL_X32 FILLER_176_1464 ();
 FILLCELL_X32 FILLER_176_1496 ();
 FILLCELL_X32 FILLER_176_1528 ();
 FILLCELL_X32 FILLER_176_1560 ();
 FILLCELL_X32 FILLER_176_1592 ();
 FILLCELL_X32 FILLER_176_1624 ();
 FILLCELL_X32 FILLER_176_1656 ();
 FILLCELL_X32 FILLER_176_1688 ();
 FILLCELL_X32 FILLER_176_1720 ();
 FILLCELL_X32 FILLER_176_1752 ();
 FILLCELL_X32 FILLER_176_1784 ();
 FILLCELL_X32 FILLER_176_1816 ();
 FILLCELL_X32 FILLER_176_1848 ();
 FILLCELL_X8 FILLER_176_1880 ();
 FILLCELL_X4 FILLER_176_1888 ();
 FILLCELL_X2 FILLER_176_1892 ();
 FILLCELL_X32 FILLER_176_1895 ();
 FILLCELL_X32 FILLER_176_1927 ();
 FILLCELL_X32 FILLER_176_1959 ();
 FILLCELL_X32 FILLER_176_1991 ();
 FILLCELL_X32 FILLER_176_2023 ();
 FILLCELL_X32 FILLER_176_2055 ();
 FILLCELL_X32 FILLER_176_2087 ();
 FILLCELL_X32 FILLER_176_2119 ();
 FILLCELL_X32 FILLER_176_2151 ();
 FILLCELL_X32 FILLER_176_2183 ();
 FILLCELL_X32 FILLER_176_2215 ();
 FILLCELL_X32 FILLER_176_2247 ();
 FILLCELL_X32 FILLER_176_2279 ();
 FILLCELL_X32 FILLER_176_2311 ();
 FILLCELL_X32 FILLER_176_2343 ();
 FILLCELL_X32 FILLER_176_2375 ();
 FILLCELL_X32 FILLER_176_2407 ();
 FILLCELL_X32 FILLER_176_2439 ();
 FILLCELL_X32 FILLER_176_2471 ();
 FILLCELL_X32 FILLER_176_2503 ();
 FILLCELL_X32 FILLER_176_2535 ();
 FILLCELL_X32 FILLER_176_2567 ();
 FILLCELL_X32 FILLER_176_2599 ();
 FILLCELL_X32 FILLER_176_2631 ();
 FILLCELL_X32 FILLER_176_2663 ();
 FILLCELL_X32 FILLER_176_2695 ();
 FILLCELL_X32 FILLER_176_2727 ();
 FILLCELL_X32 FILLER_176_2759 ();
 FILLCELL_X32 FILLER_176_2791 ();
 FILLCELL_X32 FILLER_176_2823 ();
 FILLCELL_X32 FILLER_176_2855 ();
 FILLCELL_X32 FILLER_176_2887 ();
 FILLCELL_X32 FILLER_176_2919 ();
 FILLCELL_X32 FILLER_176_2951 ();
 FILLCELL_X32 FILLER_176_2983 ();
 FILLCELL_X32 FILLER_176_3015 ();
 FILLCELL_X32 FILLER_176_3047 ();
 FILLCELL_X32 FILLER_176_3079 ();
 FILLCELL_X32 FILLER_176_3111 ();
 FILLCELL_X8 FILLER_176_3143 ();
 FILLCELL_X4 FILLER_176_3151 ();
 FILLCELL_X2 FILLER_176_3155 ();
 FILLCELL_X32 FILLER_176_3158 ();
 FILLCELL_X32 FILLER_176_3190 ();
 FILLCELL_X32 FILLER_176_3222 ();
 FILLCELL_X32 FILLER_176_3254 ();
 FILLCELL_X32 FILLER_176_3286 ();
 FILLCELL_X32 FILLER_176_3318 ();
 FILLCELL_X32 FILLER_176_3350 ();
 FILLCELL_X32 FILLER_176_3382 ();
 FILLCELL_X32 FILLER_176_3414 ();
 FILLCELL_X32 FILLER_176_3446 ();
 FILLCELL_X32 FILLER_176_3478 ();
 FILLCELL_X32 FILLER_176_3510 ();
 FILLCELL_X32 FILLER_176_3542 ();
 FILLCELL_X32 FILLER_176_3574 ();
 FILLCELL_X32 FILLER_176_3606 ();
 FILLCELL_X32 FILLER_176_3638 ();
 FILLCELL_X32 FILLER_176_3670 ();
 FILLCELL_X32 FILLER_176_3702 ();
 FILLCELL_X4 FILLER_176_3734 ();
 FILLCELL_X32 FILLER_177_1 ();
 FILLCELL_X32 FILLER_177_33 ();
 FILLCELL_X32 FILLER_177_65 ();
 FILLCELL_X32 FILLER_177_97 ();
 FILLCELL_X32 FILLER_177_129 ();
 FILLCELL_X32 FILLER_177_161 ();
 FILLCELL_X32 FILLER_177_193 ();
 FILLCELL_X32 FILLER_177_225 ();
 FILLCELL_X32 FILLER_177_257 ();
 FILLCELL_X32 FILLER_177_289 ();
 FILLCELL_X32 FILLER_177_321 ();
 FILLCELL_X32 FILLER_177_353 ();
 FILLCELL_X32 FILLER_177_385 ();
 FILLCELL_X32 FILLER_177_417 ();
 FILLCELL_X32 FILLER_177_449 ();
 FILLCELL_X32 FILLER_177_481 ();
 FILLCELL_X32 FILLER_177_513 ();
 FILLCELL_X32 FILLER_177_545 ();
 FILLCELL_X32 FILLER_177_577 ();
 FILLCELL_X32 FILLER_177_609 ();
 FILLCELL_X32 FILLER_177_641 ();
 FILLCELL_X32 FILLER_177_673 ();
 FILLCELL_X32 FILLER_177_705 ();
 FILLCELL_X32 FILLER_177_737 ();
 FILLCELL_X32 FILLER_177_769 ();
 FILLCELL_X32 FILLER_177_801 ();
 FILLCELL_X32 FILLER_177_833 ();
 FILLCELL_X32 FILLER_177_865 ();
 FILLCELL_X32 FILLER_177_897 ();
 FILLCELL_X32 FILLER_177_929 ();
 FILLCELL_X32 FILLER_177_961 ();
 FILLCELL_X32 FILLER_177_993 ();
 FILLCELL_X32 FILLER_177_1025 ();
 FILLCELL_X32 FILLER_177_1057 ();
 FILLCELL_X32 FILLER_177_1089 ();
 FILLCELL_X32 FILLER_177_1121 ();
 FILLCELL_X32 FILLER_177_1153 ();
 FILLCELL_X32 FILLER_177_1185 ();
 FILLCELL_X32 FILLER_177_1217 ();
 FILLCELL_X8 FILLER_177_1249 ();
 FILLCELL_X4 FILLER_177_1257 ();
 FILLCELL_X2 FILLER_177_1261 ();
 FILLCELL_X32 FILLER_177_1264 ();
 FILLCELL_X32 FILLER_177_1296 ();
 FILLCELL_X32 FILLER_177_1328 ();
 FILLCELL_X32 FILLER_177_1360 ();
 FILLCELL_X32 FILLER_177_1392 ();
 FILLCELL_X32 FILLER_177_1424 ();
 FILLCELL_X32 FILLER_177_1456 ();
 FILLCELL_X32 FILLER_177_1488 ();
 FILLCELL_X32 FILLER_177_1520 ();
 FILLCELL_X32 FILLER_177_1552 ();
 FILLCELL_X32 FILLER_177_1584 ();
 FILLCELL_X32 FILLER_177_1616 ();
 FILLCELL_X32 FILLER_177_1648 ();
 FILLCELL_X32 FILLER_177_1680 ();
 FILLCELL_X32 FILLER_177_1712 ();
 FILLCELL_X32 FILLER_177_1744 ();
 FILLCELL_X32 FILLER_177_1776 ();
 FILLCELL_X32 FILLER_177_1808 ();
 FILLCELL_X32 FILLER_177_1840 ();
 FILLCELL_X32 FILLER_177_1872 ();
 FILLCELL_X32 FILLER_177_1904 ();
 FILLCELL_X32 FILLER_177_1936 ();
 FILLCELL_X32 FILLER_177_1968 ();
 FILLCELL_X32 FILLER_177_2000 ();
 FILLCELL_X32 FILLER_177_2032 ();
 FILLCELL_X32 FILLER_177_2064 ();
 FILLCELL_X32 FILLER_177_2096 ();
 FILLCELL_X32 FILLER_177_2128 ();
 FILLCELL_X32 FILLER_177_2160 ();
 FILLCELL_X32 FILLER_177_2192 ();
 FILLCELL_X32 FILLER_177_2224 ();
 FILLCELL_X32 FILLER_177_2256 ();
 FILLCELL_X32 FILLER_177_2288 ();
 FILLCELL_X32 FILLER_177_2320 ();
 FILLCELL_X32 FILLER_177_2352 ();
 FILLCELL_X32 FILLER_177_2384 ();
 FILLCELL_X32 FILLER_177_2416 ();
 FILLCELL_X32 FILLER_177_2448 ();
 FILLCELL_X32 FILLER_177_2480 ();
 FILLCELL_X8 FILLER_177_2512 ();
 FILLCELL_X4 FILLER_177_2520 ();
 FILLCELL_X2 FILLER_177_2524 ();
 FILLCELL_X32 FILLER_177_2527 ();
 FILLCELL_X32 FILLER_177_2559 ();
 FILLCELL_X32 FILLER_177_2591 ();
 FILLCELL_X32 FILLER_177_2623 ();
 FILLCELL_X32 FILLER_177_2655 ();
 FILLCELL_X32 FILLER_177_2687 ();
 FILLCELL_X32 FILLER_177_2719 ();
 FILLCELL_X32 FILLER_177_2751 ();
 FILLCELL_X32 FILLER_177_2783 ();
 FILLCELL_X32 FILLER_177_2815 ();
 FILLCELL_X32 FILLER_177_2847 ();
 FILLCELL_X32 FILLER_177_2879 ();
 FILLCELL_X32 FILLER_177_2911 ();
 FILLCELL_X32 FILLER_177_2943 ();
 FILLCELL_X32 FILLER_177_2975 ();
 FILLCELL_X32 FILLER_177_3007 ();
 FILLCELL_X32 FILLER_177_3039 ();
 FILLCELL_X32 FILLER_177_3071 ();
 FILLCELL_X32 FILLER_177_3103 ();
 FILLCELL_X32 FILLER_177_3135 ();
 FILLCELL_X32 FILLER_177_3167 ();
 FILLCELL_X32 FILLER_177_3199 ();
 FILLCELL_X32 FILLER_177_3231 ();
 FILLCELL_X32 FILLER_177_3263 ();
 FILLCELL_X32 FILLER_177_3295 ();
 FILLCELL_X32 FILLER_177_3327 ();
 FILLCELL_X32 FILLER_177_3359 ();
 FILLCELL_X32 FILLER_177_3391 ();
 FILLCELL_X32 FILLER_177_3423 ();
 FILLCELL_X32 FILLER_177_3455 ();
 FILLCELL_X32 FILLER_177_3487 ();
 FILLCELL_X32 FILLER_177_3519 ();
 FILLCELL_X32 FILLER_177_3551 ();
 FILLCELL_X32 FILLER_177_3583 ();
 FILLCELL_X32 FILLER_177_3615 ();
 FILLCELL_X32 FILLER_177_3647 ();
 FILLCELL_X32 FILLER_177_3679 ();
 FILLCELL_X16 FILLER_177_3711 ();
 FILLCELL_X8 FILLER_177_3727 ();
 FILLCELL_X2 FILLER_177_3735 ();
 FILLCELL_X1 FILLER_177_3737 ();
 FILLCELL_X32 FILLER_178_1 ();
 FILLCELL_X32 FILLER_178_33 ();
 FILLCELL_X32 FILLER_178_65 ();
 FILLCELL_X32 FILLER_178_97 ();
 FILLCELL_X32 FILLER_178_129 ();
 FILLCELL_X32 FILLER_178_161 ();
 FILLCELL_X32 FILLER_178_193 ();
 FILLCELL_X32 FILLER_178_225 ();
 FILLCELL_X32 FILLER_178_257 ();
 FILLCELL_X32 FILLER_178_289 ();
 FILLCELL_X32 FILLER_178_321 ();
 FILLCELL_X32 FILLER_178_353 ();
 FILLCELL_X32 FILLER_178_385 ();
 FILLCELL_X32 FILLER_178_417 ();
 FILLCELL_X32 FILLER_178_449 ();
 FILLCELL_X32 FILLER_178_481 ();
 FILLCELL_X32 FILLER_178_513 ();
 FILLCELL_X32 FILLER_178_545 ();
 FILLCELL_X32 FILLER_178_577 ();
 FILLCELL_X16 FILLER_178_609 ();
 FILLCELL_X4 FILLER_178_625 ();
 FILLCELL_X2 FILLER_178_629 ();
 FILLCELL_X32 FILLER_178_632 ();
 FILLCELL_X32 FILLER_178_664 ();
 FILLCELL_X32 FILLER_178_696 ();
 FILLCELL_X32 FILLER_178_728 ();
 FILLCELL_X32 FILLER_178_760 ();
 FILLCELL_X32 FILLER_178_792 ();
 FILLCELL_X32 FILLER_178_824 ();
 FILLCELL_X32 FILLER_178_856 ();
 FILLCELL_X32 FILLER_178_888 ();
 FILLCELL_X32 FILLER_178_920 ();
 FILLCELL_X32 FILLER_178_952 ();
 FILLCELL_X32 FILLER_178_984 ();
 FILLCELL_X32 FILLER_178_1016 ();
 FILLCELL_X32 FILLER_178_1048 ();
 FILLCELL_X32 FILLER_178_1080 ();
 FILLCELL_X32 FILLER_178_1112 ();
 FILLCELL_X32 FILLER_178_1144 ();
 FILLCELL_X32 FILLER_178_1176 ();
 FILLCELL_X32 FILLER_178_1208 ();
 FILLCELL_X32 FILLER_178_1240 ();
 FILLCELL_X32 FILLER_178_1272 ();
 FILLCELL_X32 FILLER_178_1304 ();
 FILLCELL_X32 FILLER_178_1336 ();
 FILLCELL_X32 FILLER_178_1368 ();
 FILLCELL_X32 FILLER_178_1400 ();
 FILLCELL_X32 FILLER_178_1432 ();
 FILLCELL_X32 FILLER_178_1464 ();
 FILLCELL_X32 FILLER_178_1496 ();
 FILLCELL_X32 FILLER_178_1528 ();
 FILLCELL_X32 FILLER_178_1560 ();
 FILLCELL_X32 FILLER_178_1592 ();
 FILLCELL_X32 FILLER_178_1624 ();
 FILLCELL_X32 FILLER_178_1656 ();
 FILLCELL_X32 FILLER_178_1688 ();
 FILLCELL_X32 FILLER_178_1720 ();
 FILLCELL_X32 FILLER_178_1752 ();
 FILLCELL_X32 FILLER_178_1784 ();
 FILLCELL_X32 FILLER_178_1816 ();
 FILLCELL_X32 FILLER_178_1848 ();
 FILLCELL_X8 FILLER_178_1880 ();
 FILLCELL_X4 FILLER_178_1888 ();
 FILLCELL_X2 FILLER_178_1892 ();
 FILLCELL_X32 FILLER_178_1895 ();
 FILLCELL_X32 FILLER_178_1927 ();
 FILLCELL_X32 FILLER_178_1959 ();
 FILLCELL_X32 FILLER_178_1991 ();
 FILLCELL_X32 FILLER_178_2023 ();
 FILLCELL_X32 FILLER_178_2055 ();
 FILLCELL_X32 FILLER_178_2087 ();
 FILLCELL_X32 FILLER_178_2119 ();
 FILLCELL_X32 FILLER_178_2151 ();
 FILLCELL_X32 FILLER_178_2183 ();
 FILLCELL_X32 FILLER_178_2215 ();
 FILLCELL_X32 FILLER_178_2247 ();
 FILLCELL_X32 FILLER_178_2279 ();
 FILLCELL_X32 FILLER_178_2311 ();
 FILLCELL_X32 FILLER_178_2343 ();
 FILLCELL_X32 FILLER_178_2375 ();
 FILLCELL_X32 FILLER_178_2407 ();
 FILLCELL_X32 FILLER_178_2439 ();
 FILLCELL_X32 FILLER_178_2471 ();
 FILLCELL_X32 FILLER_178_2503 ();
 FILLCELL_X32 FILLER_178_2535 ();
 FILLCELL_X32 FILLER_178_2567 ();
 FILLCELL_X32 FILLER_178_2599 ();
 FILLCELL_X32 FILLER_178_2631 ();
 FILLCELL_X32 FILLER_178_2663 ();
 FILLCELL_X32 FILLER_178_2695 ();
 FILLCELL_X32 FILLER_178_2727 ();
 FILLCELL_X32 FILLER_178_2759 ();
 FILLCELL_X32 FILLER_178_2791 ();
 FILLCELL_X32 FILLER_178_2823 ();
 FILLCELL_X32 FILLER_178_2855 ();
 FILLCELL_X32 FILLER_178_2887 ();
 FILLCELL_X32 FILLER_178_2919 ();
 FILLCELL_X32 FILLER_178_2951 ();
 FILLCELL_X32 FILLER_178_2983 ();
 FILLCELL_X32 FILLER_178_3015 ();
 FILLCELL_X32 FILLER_178_3047 ();
 FILLCELL_X32 FILLER_178_3079 ();
 FILLCELL_X32 FILLER_178_3111 ();
 FILLCELL_X8 FILLER_178_3143 ();
 FILLCELL_X4 FILLER_178_3151 ();
 FILLCELL_X2 FILLER_178_3155 ();
 FILLCELL_X32 FILLER_178_3158 ();
 FILLCELL_X32 FILLER_178_3190 ();
 FILLCELL_X32 FILLER_178_3222 ();
 FILLCELL_X32 FILLER_178_3254 ();
 FILLCELL_X32 FILLER_178_3286 ();
 FILLCELL_X32 FILLER_178_3318 ();
 FILLCELL_X32 FILLER_178_3350 ();
 FILLCELL_X32 FILLER_178_3382 ();
 FILLCELL_X32 FILLER_178_3414 ();
 FILLCELL_X32 FILLER_178_3446 ();
 FILLCELL_X32 FILLER_178_3478 ();
 FILLCELL_X32 FILLER_178_3510 ();
 FILLCELL_X32 FILLER_178_3542 ();
 FILLCELL_X32 FILLER_178_3574 ();
 FILLCELL_X32 FILLER_178_3606 ();
 FILLCELL_X32 FILLER_178_3638 ();
 FILLCELL_X32 FILLER_178_3670 ();
 FILLCELL_X32 FILLER_178_3702 ();
 FILLCELL_X4 FILLER_178_3734 ();
 FILLCELL_X32 FILLER_179_1 ();
 FILLCELL_X32 FILLER_179_33 ();
 FILLCELL_X32 FILLER_179_65 ();
 FILLCELL_X32 FILLER_179_97 ();
 FILLCELL_X32 FILLER_179_129 ();
 FILLCELL_X32 FILLER_179_161 ();
 FILLCELL_X32 FILLER_179_193 ();
 FILLCELL_X32 FILLER_179_225 ();
 FILLCELL_X32 FILLER_179_257 ();
 FILLCELL_X32 FILLER_179_289 ();
 FILLCELL_X32 FILLER_179_321 ();
 FILLCELL_X32 FILLER_179_353 ();
 FILLCELL_X32 FILLER_179_385 ();
 FILLCELL_X32 FILLER_179_417 ();
 FILLCELL_X32 FILLER_179_449 ();
 FILLCELL_X32 FILLER_179_481 ();
 FILLCELL_X32 FILLER_179_513 ();
 FILLCELL_X32 FILLER_179_545 ();
 FILLCELL_X32 FILLER_179_577 ();
 FILLCELL_X32 FILLER_179_609 ();
 FILLCELL_X32 FILLER_179_641 ();
 FILLCELL_X32 FILLER_179_673 ();
 FILLCELL_X32 FILLER_179_705 ();
 FILLCELL_X32 FILLER_179_737 ();
 FILLCELL_X32 FILLER_179_769 ();
 FILLCELL_X32 FILLER_179_801 ();
 FILLCELL_X32 FILLER_179_833 ();
 FILLCELL_X32 FILLER_179_865 ();
 FILLCELL_X32 FILLER_179_897 ();
 FILLCELL_X32 FILLER_179_929 ();
 FILLCELL_X32 FILLER_179_961 ();
 FILLCELL_X32 FILLER_179_993 ();
 FILLCELL_X32 FILLER_179_1025 ();
 FILLCELL_X32 FILLER_179_1057 ();
 FILLCELL_X32 FILLER_179_1089 ();
 FILLCELL_X32 FILLER_179_1121 ();
 FILLCELL_X32 FILLER_179_1153 ();
 FILLCELL_X32 FILLER_179_1185 ();
 FILLCELL_X32 FILLER_179_1217 ();
 FILLCELL_X8 FILLER_179_1249 ();
 FILLCELL_X4 FILLER_179_1257 ();
 FILLCELL_X2 FILLER_179_1261 ();
 FILLCELL_X32 FILLER_179_1264 ();
 FILLCELL_X32 FILLER_179_1296 ();
 FILLCELL_X32 FILLER_179_1328 ();
 FILLCELL_X32 FILLER_179_1360 ();
 FILLCELL_X32 FILLER_179_1392 ();
 FILLCELL_X32 FILLER_179_1424 ();
 FILLCELL_X32 FILLER_179_1456 ();
 FILLCELL_X32 FILLER_179_1488 ();
 FILLCELL_X32 FILLER_179_1520 ();
 FILLCELL_X32 FILLER_179_1552 ();
 FILLCELL_X32 FILLER_179_1584 ();
 FILLCELL_X32 FILLER_179_1616 ();
 FILLCELL_X32 FILLER_179_1648 ();
 FILLCELL_X32 FILLER_179_1680 ();
 FILLCELL_X32 FILLER_179_1712 ();
 FILLCELL_X32 FILLER_179_1744 ();
 FILLCELL_X32 FILLER_179_1776 ();
 FILLCELL_X32 FILLER_179_1808 ();
 FILLCELL_X32 FILLER_179_1840 ();
 FILLCELL_X32 FILLER_179_1872 ();
 FILLCELL_X32 FILLER_179_1904 ();
 FILLCELL_X32 FILLER_179_1936 ();
 FILLCELL_X32 FILLER_179_1968 ();
 FILLCELL_X32 FILLER_179_2000 ();
 FILLCELL_X32 FILLER_179_2032 ();
 FILLCELL_X32 FILLER_179_2064 ();
 FILLCELL_X32 FILLER_179_2096 ();
 FILLCELL_X32 FILLER_179_2128 ();
 FILLCELL_X32 FILLER_179_2160 ();
 FILLCELL_X32 FILLER_179_2192 ();
 FILLCELL_X32 FILLER_179_2224 ();
 FILLCELL_X32 FILLER_179_2256 ();
 FILLCELL_X32 FILLER_179_2288 ();
 FILLCELL_X32 FILLER_179_2320 ();
 FILLCELL_X32 FILLER_179_2352 ();
 FILLCELL_X32 FILLER_179_2384 ();
 FILLCELL_X32 FILLER_179_2416 ();
 FILLCELL_X32 FILLER_179_2448 ();
 FILLCELL_X32 FILLER_179_2480 ();
 FILLCELL_X8 FILLER_179_2512 ();
 FILLCELL_X4 FILLER_179_2520 ();
 FILLCELL_X2 FILLER_179_2524 ();
 FILLCELL_X32 FILLER_179_2527 ();
 FILLCELL_X32 FILLER_179_2559 ();
 FILLCELL_X32 FILLER_179_2591 ();
 FILLCELL_X32 FILLER_179_2623 ();
 FILLCELL_X32 FILLER_179_2655 ();
 FILLCELL_X32 FILLER_179_2687 ();
 FILLCELL_X32 FILLER_179_2719 ();
 FILLCELL_X32 FILLER_179_2751 ();
 FILLCELL_X32 FILLER_179_2783 ();
 FILLCELL_X32 FILLER_179_2815 ();
 FILLCELL_X32 FILLER_179_2847 ();
 FILLCELL_X32 FILLER_179_2879 ();
 FILLCELL_X32 FILLER_179_2911 ();
 FILLCELL_X32 FILLER_179_2943 ();
 FILLCELL_X32 FILLER_179_2975 ();
 FILLCELL_X32 FILLER_179_3007 ();
 FILLCELL_X32 FILLER_179_3039 ();
 FILLCELL_X32 FILLER_179_3071 ();
 FILLCELL_X32 FILLER_179_3103 ();
 FILLCELL_X32 FILLER_179_3135 ();
 FILLCELL_X32 FILLER_179_3167 ();
 FILLCELL_X32 FILLER_179_3199 ();
 FILLCELL_X32 FILLER_179_3231 ();
 FILLCELL_X32 FILLER_179_3263 ();
 FILLCELL_X32 FILLER_179_3295 ();
 FILLCELL_X32 FILLER_179_3327 ();
 FILLCELL_X32 FILLER_179_3359 ();
 FILLCELL_X32 FILLER_179_3391 ();
 FILLCELL_X32 FILLER_179_3423 ();
 FILLCELL_X32 FILLER_179_3455 ();
 FILLCELL_X32 FILLER_179_3487 ();
 FILLCELL_X32 FILLER_179_3519 ();
 FILLCELL_X32 FILLER_179_3551 ();
 FILLCELL_X32 FILLER_179_3583 ();
 FILLCELL_X32 FILLER_179_3615 ();
 FILLCELL_X32 FILLER_179_3647 ();
 FILLCELL_X32 FILLER_179_3679 ();
 FILLCELL_X16 FILLER_179_3711 ();
 FILLCELL_X8 FILLER_179_3727 ();
 FILLCELL_X2 FILLER_179_3735 ();
 FILLCELL_X1 FILLER_179_3737 ();
 FILLCELL_X32 FILLER_180_1 ();
 FILLCELL_X32 FILLER_180_33 ();
 FILLCELL_X32 FILLER_180_65 ();
 FILLCELL_X32 FILLER_180_97 ();
 FILLCELL_X32 FILLER_180_129 ();
 FILLCELL_X32 FILLER_180_161 ();
 FILLCELL_X32 FILLER_180_193 ();
 FILLCELL_X32 FILLER_180_225 ();
 FILLCELL_X32 FILLER_180_257 ();
 FILLCELL_X32 FILLER_180_289 ();
 FILLCELL_X32 FILLER_180_321 ();
 FILLCELL_X32 FILLER_180_353 ();
 FILLCELL_X32 FILLER_180_385 ();
 FILLCELL_X32 FILLER_180_417 ();
 FILLCELL_X32 FILLER_180_449 ();
 FILLCELL_X32 FILLER_180_481 ();
 FILLCELL_X32 FILLER_180_513 ();
 FILLCELL_X32 FILLER_180_545 ();
 FILLCELL_X32 FILLER_180_577 ();
 FILLCELL_X16 FILLER_180_609 ();
 FILLCELL_X4 FILLER_180_625 ();
 FILLCELL_X2 FILLER_180_629 ();
 FILLCELL_X32 FILLER_180_632 ();
 FILLCELL_X32 FILLER_180_664 ();
 FILLCELL_X32 FILLER_180_696 ();
 FILLCELL_X32 FILLER_180_728 ();
 FILLCELL_X32 FILLER_180_760 ();
 FILLCELL_X32 FILLER_180_792 ();
 FILLCELL_X32 FILLER_180_824 ();
 FILLCELL_X32 FILLER_180_856 ();
 FILLCELL_X32 FILLER_180_888 ();
 FILLCELL_X32 FILLER_180_920 ();
 FILLCELL_X32 FILLER_180_952 ();
 FILLCELL_X32 FILLER_180_984 ();
 FILLCELL_X32 FILLER_180_1016 ();
 FILLCELL_X32 FILLER_180_1048 ();
 FILLCELL_X32 FILLER_180_1080 ();
 FILLCELL_X32 FILLER_180_1112 ();
 FILLCELL_X32 FILLER_180_1144 ();
 FILLCELL_X32 FILLER_180_1176 ();
 FILLCELL_X32 FILLER_180_1208 ();
 FILLCELL_X32 FILLER_180_1240 ();
 FILLCELL_X32 FILLER_180_1272 ();
 FILLCELL_X32 FILLER_180_1304 ();
 FILLCELL_X32 FILLER_180_1336 ();
 FILLCELL_X32 FILLER_180_1368 ();
 FILLCELL_X32 FILLER_180_1400 ();
 FILLCELL_X32 FILLER_180_1432 ();
 FILLCELL_X32 FILLER_180_1464 ();
 FILLCELL_X32 FILLER_180_1496 ();
 FILLCELL_X32 FILLER_180_1528 ();
 FILLCELL_X32 FILLER_180_1560 ();
 FILLCELL_X32 FILLER_180_1592 ();
 FILLCELL_X32 FILLER_180_1624 ();
 FILLCELL_X32 FILLER_180_1656 ();
 FILLCELL_X32 FILLER_180_1688 ();
 FILLCELL_X32 FILLER_180_1720 ();
 FILLCELL_X32 FILLER_180_1752 ();
 FILLCELL_X32 FILLER_180_1784 ();
 FILLCELL_X32 FILLER_180_1816 ();
 FILLCELL_X32 FILLER_180_1848 ();
 FILLCELL_X8 FILLER_180_1880 ();
 FILLCELL_X4 FILLER_180_1888 ();
 FILLCELL_X2 FILLER_180_1892 ();
 FILLCELL_X32 FILLER_180_1895 ();
 FILLCELL_X32 FILLER_180_1927 ();
 FILLCELL_X32 FILLER_180_1959 ();
 FILLCELL_X32 FILLER_180_1991 ();
 FILLCELL_X32 FILLER_180_2023 ();
 FILLCELL_X32 FILLER_180_2055 ();
 FILLCELL_X32 FILLER_180_2087 ();
 FILLCELL_X32 FILLER_180_2119 ();
 FILLCELL_X32 FILLER_180_2151 ();
 FILLCELL_X32 FILLER_180_2183 ();
 FILLCELL_X32 FILLER_180_2215 ();
 FILLCELL_X32 FILLER_180_2247 ();
 FILLCELL_X32 FILLER_180_2279 ();
 FILLCELL_X32 FILLER_180_2311 ();
 FILLCELL_X32 FILLER_180_2343 ();
 FILLCELL_X32 FILLER_180_2375 ();
 FILLCELL_X32 FILLER_180_2407 ();
 FILLCELL_X32 FILLER_180_2439 ();
 FILLCELL_X32 FILLER_180_2471 ();
 FILLCELL_X32 FILLER_180_2503 ();
 FILLCELL_X32 FILLER_180_2535 ();
 FILLCELL_X32 FILLER_180_2567 ();
 FILLCELL_X32 FILLER_180_2599 ();
 FILLCELL_X32 FILLER_180_2631 ();
 FILLCELL_X32 FILLER_180_2663 ();
 FILLCELL_X32 FILLER_180_2695 ();
 FILLCELL_X32 FILLER_180_2727 ();
 FILLCELL_X32 FILLER_180_2759 ();
 FILLCELL_X32 FILLER_180_2791 ();
 FILLCELL_X32 FILLER_180_2823 ();
 FILLCELL_X32 FILLER_180_2855 ();
 FILLCELL_X32 FILLER_180_2887 ();
 FILLCELL_X32 FILLER_180_2919 ();
 FILLCELL_X32 FILLER_180_2951 ();
 FILLCELL_X32 FILLER_180_2983 ();
 FILLCELL_X32 FILLER_180_3015 ();
 FILLCELL_X32 FILLER_180_3047 ();
 FILLCELL_X32 FILLER_180_3079 ();
 FILLCELL_X32 FILLER_180_3111 ();
 FILLCELL_X8 FILLER_180_3143 ();
 FILLCELL_X4 FILLER_180_3151 ();
 FILLCELL_X2 FILLER_180_3155 ();
 FILLCELL_X32 FILLER_180_3158 ();
 FILLCELL_X32 FILLER_180_3190 ();
 FILLCELL_X32 FILLER_180_3222 ();
 FILLCELL_X32 FILLER_180_3254 ();
 FILLCELL_X32 FILLER_180_3286 ();
 FILLCELL_X32 FILLER_180_3318 ();
 FILLCELL_X32 FILLER_180_3350 ();
 FILLCELL_X32 FILLER_180_3382 ();
 FILLCELL_X32 FILLER_180_3414 ();
 FILLCELL_X32 FILLER_180_3446 ();
 FILLCELL_X32 FILLER_180_3478 ();
 FILLCELL_X32 FILLER_180_3510 ();
 FILLCELL_X32 FILLER_180_3542 ();
 FILLCELL_X32 FILLER_180_3574 ();
 FILLCELL_X32 FILLER_180_3606 ();
 FILLCELL_X32 FILLER_180_3638 ();
 FILLCELL_X32 FILLER_180_3670 ();
 FILLCELL_X32 FILLER_180_3702 ();
 FILLCELL_X4 FILLER_180_3734 ();
 FILLCELL_X32 FILLER_181_1 ();
 FILLCELL_X32 FILLER_181_33 ();
 FILLCELL_X32 FILLER_181_65 ();
 FILLCELL_X32 FILLER_181_97 ();
 FILLCELL_X32 FILLER_181_129 ();
 FILLCELL_X32 FILLER_181_161 ();
 FILLCELL_X32 FILLER_181_193 ();
 FILLCELL_X32 FILLER_181_225 ();
 FILLCELL_X32 FILLER_181_257 ();
 FILLCELL_X32 FILLER_181_289 ();
 FILLCELL_X32 FILLER_181_321 ();
 FILLCELL_X32 FILLER_181_353 ();
 FILLCELL_X32 FILLER_181_385 ();
 FILLCELL_X32 FILLER_181_417 ();
 FILLCELL_X32 FILLER_181_449 ();
 FILLCELL_X32 FILLER_181_481 ();
 FILLCELL_X32 FILLER_181_513 ();
 FILLCELL_X32 FILLER_181_545 ();
 FILLCELL_X32 FILLER_181_577 ();
 FILLCELL_X32 FILLER_181_609 ();
 FILLCELL_X32 FILLER_181_641 ();
 FILLCELL_X32 FILLER_181_673 ();
 FILLCELL_X32 FILLER_181_705 ();
 FILLCELL_X32 FILLER_181_737 ();
 FILLCELL_X32 FILLER_181_769 ();
 FILLCELL_X32 FILLER_181_801 ();
 FILLCELL_X32 FILLER_181_833 ();
 FILLCELL_X32 FILLER_181_865 ();
 FILLCELL_X32 FILLER_181_897 ();
 FILLCELL_X32 FILLER_181_929 ();
 FILLCELL_X32 FILLER_181_961 ();
 FILLCELL_X32 FILLER_181_993 ();
 FILLCELL_X32 FILLER_181_1025 ();
 FILLCELL_X32 FILLER_181_1057 ();
 FILLCELL_X32 FILLER_181_1089 ();
 FILLCELL_X32 FILLER_181_1121 ();
 FILLCELL_X32 FILLER_181_1153 ();
 FILLCELL_X32 FILLER_181_1185 ();
 FILLCELL_X32 FILLER_181_1217 ();
 FILLCELL_X8 FILLER_181_1249 ();
 FILLCELL_X4 FILLER_181_1257 ();
 FILLCELL_X2 FILLER_181_1261 ();
 FILLCELL_X32 FILLER_181_1264 ();
 FILLCELL_X32 FILLER_181_1296 ();
 FILLCELL_X32 FILLER_181_1328 ();
 FILLCELL_X32 FILLER_181_1360 ();
 FILLCELL_X32 FILLER_181_1392 ();
 FILLCELL_X32 FILLER_181_1424 ();
 FILLCELL_X32 FILLER_181_1456 ();
 FILLCELL_X32 FILLER_181_1488 ();
 FILLCELL_X32 FILLER_181_1520 ();
 FILLCELL_X32 FILLER_181_1552 ();
 FILLCELL_X32 FILLER_181_1584 ();
 FILLCELL_X32 FILLER_181_1616 ();
 FILLCELL_X32 FILLER_181_1648 ();
 FILLCELL_X32 FILLER_181_1680 ();
 FILLCELL_X32 FILLER_181_1712 ();
 FILLCELL_X32 FILLER_181_1744 ();
 FILLCELL_X32 FILLER_181_1776 ();
 FILLCELL_X32 FILLER_181_1808 ();
 FILLCELL_X32 FILLER_181_1840 ();
 FILLCELL_X32 FILLER_181_1872 ();
 FILLCELL_X32 FILLER_181_1904 ();
 FILLCELL_X32 FILLER_181_1936 ();
 FILLCELL_X32 FILLER_181_1968 ();
 FILLCELL_X32 FILLER_181_2000 ();
 FILLCELL_X32 FILLER_181_2032 ();
 FILLCELL_X32 FILLER_181_2064 ();
 FILLCELL_X32 FILLER_181_2096 ();
 FILLCELL_X32 FILLER_181_2128 ();
 FILLCELL_X32 FILLER_181_2160 ();
 FILLCELL_X32 FILLER_181_2192 ();
 FILLCELL_X32 FILLER_181_2224 ();
 FILLCELL_X32 FILLER_181_2256 ();
 FILLCELL_X32 FILLER_181_2288 ();
 FILLCELL_X32 FILLER_181_2320 ();
 FILLCELL_X32 FILLER_181_2352 ();
 FILLCELL_X32 FILLER_181_2384 ();
 FILLCELL_X32 FILLER_181_2416 ();
 FILLCELL_X32 FILLER_181_2448 ();
 FILLCELL_X32 FILLER_181_2480 ();
 FILLCELL_X8 FILLER_181_2512 ();
 FILLCELL_X4 FILLER_181_2520 ();
 FILLCELL_X2 FILLER_181_2524 ();
 FILLCELL_X32 FILLER_181_2527 ();
 FILLCELL_X32 FILLER_181_2559 ();
 FILLCELL_X32 FILLER_181_2591 ();
 FILLCELL_X32 FILLER_181_2623 ();
 FILLCELL_X32 FILLER_181_2655 ();
 FILLCELL_X32 FILLER_181_2687 ();
 FILLCELL_X32 FILLER_181_2719 ();
 FILLCELL_X32 FILLER_181_2751 ();
 FILLCELL_X32 FILLER_181_2783 ();
 FILLCELL_X32 FILLER_181_2815 ();
 FILLCELL_X32 FILLER_181_2847 ();
 FILLCELL_X32 FILLER_181_2879 ();
 FILLCELL_X32 FILLER_181_2911 ();
 FILLCELL_X32 FILLER_181_2943 ();
 FILLCELL_X32 FILLER_181_2975 ();
 FILLCELL_X32 FILLER_181_3007 ();
 FILLCELL_X32 FILLER_181_3039 ();
 FILLCELL_X32 FILLER_181_3071 ();
 FILLCELL_X32 FILLER_181_3103 ();
 FILLCELL_X32 FILLER_181_3135 ();
 FILLCELL_X32 FILLER_181_3167 ();
 FILLCELL_X32 FILLER_181_3199 ();
 FILLCELL_X32 FILLER_181_3231 ();
 FILLCELL_X32 FILLER_181_3263 ();
 FILLCELL_X32 FILLER_181_3295 ();
 FILLCELL_X32 FILLER_181_3327 ();
 FILLCELL_X32 FILLER_181_3359 ();
 FILLCELL_X32 FILLER_181_3391 ();
 FILLCELL_X32 FILLER_181_3423 ();
 FILLCELL_X32 FILLER_181_3455 ();
 FILLCELL_X32 FILLER_181_3487 ();
 FILLCELL_X32 FILLER_181_3519 ();
 FILLCELL_X32 FILLER_181_3551 ();
 FILLCELL_X32 FILLER_181_3583 ();
 FILLCELL_X32 FILLER_181_3615 ();
 FILLCELL_X32 FILLER_181_3647 ();
 FILLCELL_X32 FILLER_181_3679 ();
 FILLCELL_X16 FILLER_181_3711 ();
 FILLCELL_X8 FILLER_181_3727 ();
 FILLCELL_X2 FILLER_181_3735 ();
 FILLCELL_X1 FILLER_181_3737 ();
 FILLCELL_X32 FILLER_182_1 ();
 FILLCELL_X32 FILLER_182_33 ();
 FILLCELL_X32 FILLER_182_65 ();
 FILLCELL_X32 FILLER_182_97 ();
 FILLCELL_X32 FILLER_182_129 ();
 FILLCELL_X32 FILLER_182_161 ();
 FILLCELL_X32 FILLER_182_193 ();
 FILLCELL_X32 FILLER_182_225 ();
 FILLCELL_X32 FILLER_182_257 ();
 FILLCELL_X32 FILLER_182_289 ();
 FILLCELL_X32 FILLER_182_321 ();
 FILLCELL_X32 FILLER_182_353 ();
 FILLCELL_X32 FILLER_182_385 ();
 FILLCELL_X32 FILLER_182_417 ();
 FILLCELL_X32 FILLER_182_449 ();
 FILLCELL_X32 FILLER_182_481 ();
 FILLCELL_X32 FILLER_182_513 ();
 FILLCELL_X32 FILLER_182_545 ();
 FILLCELL_X32 FILLER_182_577 ();
 FILLCELL_X16 FILLER_182_609 ();
 FILLCELL_X4 FILLER_182_625 ();
 FILLCELL_X2 FILLER_182_629 ();
 FILLCELL_X32 FILLER_182_632 ();
 FILLCELL_X32 FILLER_182_664 ();
 FILLCELL_X32 FILLER_182_696 ();
 FILLCELL_X32 FILLER_182_728 ();
 FILLCELL_X32 FILLER_182_760 ();
 FILLCELL_X32 FILLER_182_792 ();
 FILLCELL_X32 FILLER_182_824 ();
 FILLCELL_X32 FILLER_182_856 ();
 FILLCELL_X32 FILLER_182_888 ();
 FILLCELL_X32 FILLER_182_920 ();
 FILLCELL_X32 FILLER_182_952 ();
 FILLCELL_X32 FILLER_182_984 ();
 FILLCELL_X32 FILLER_182_1016 ();
 FILLCELL_X32 FILLER_182_1048 ();
 FILLCELL_X32 FILLER_182_1080 ();
 FILLCELL_X32 FILLER_182_1112 ();
 FILLCELL_X32 FILLER_182_1144 ();
 FILLCELL_X32 FILLER_182_1176 ();
 FILLCELL_X32 FILLER_182_1208 ();
 FILLCELL_X32 FILLER_182_1240 ();
 FILLCELL_X32 FILLER_182_1272 ();
 FILLCELL_X32 FILLER_182_1304 ();
 FILLCELL_X32 FILLER_182_1336 ();
 FILLCELL_X32 FILLER_182_1368 ();
 FILLCELL_X32 FILLER_182_1400 ();
 FILLCELL_X32 FILLER_182_1432 ();
 FILLCELL_X32 FILLER_182_1464 ();
 FILLCELL_X32 FILLER_182_1496 ();
 FILLCELL_X32 FILLER_182_1528 ();
 FILLCELL_X32 FILLER_182_1560 ();
 FILLCELL_X32 FILLER_182_1592 ();
 FILLCELL_X32 FILLER_182_1624 ();
 FILLCELL_X32 FILLER_182_1656 ();
 FILLCELL_X32 FILLER_182_1688 ();
 FILLCELL_X32 FILLER_182_1720 ();
 FILLCELL_X32 FILLER_182_1752 ();
 FILLCELL_X32 FILLER_182_1784 ();
 FILLCELL_X32 FILLER_182_1816 ();
 FILLCELL_X32 FILLER_182_1848 ();
 FILLCELL_X8 FILLER_182_1880 ();
 FILLCELL_X4 FILLER_182_1888 ();
 FILLCELL_X2 FILLER_182_1892 ();
 FILLCELL_X32 FILLER_182_1895 ();
 FILLCELL_X32 FILLER_182_1927 ();
 FILLCELL_X32 FILLER_182_1959 ();
 FILLCELL_X32 FILLER_182_1991 ();
 FILLCELL_X32 FILLER_182_2023 ();
 FILLCELL_X32 FILLER_182_2055 ();
 FILLCELL_X32 FILLER_182_2087 ();
 FILLCELL_X32 FILLER_182_2119 ();
 FILLCELL_X32 FILLER_182_2151 ();
 FILLCELL_X32 FILLER_182_2183 ();
 FILLCELL_X32 FILLER_182_2215 ();
 FILLCELL_X32 FILLER_182_2247 ();
 FILLCELL_X32 FILLER_182_2279 ();
 FILLCELL_X32 FILLER_182_2311 ();
 FILLCELL_X32 FILLER_182_2343 ();
 FILLCELL_X32 FILLER_182_2375 ();
 FILLCELL_X32 FILLER_182_2407 ();
 FILLCELL_X32 FILLER_182_2439 ();
 FILLCELL_X32 FILLER_182_2471 ();
 FILLCELL_X32 FILLER_182_2503 ();
 FILLCELL_X32 FILLER_182_2535 ();
 FILLCELL_X32 FILLER_182_2567 ();
 FILLCELL_X32 FILLER_182_2599 ();
 FILLCELL_X32 FILLER_182_2631 ();
 FILLCELL_X32 FILLER_182_2663 ();
 FILLCELL_X32 FILLER_182_2695 ();
 FILLCELL_X32 FILLER_182_2727 ();
 FILLCELL_X32 FILLER_182_2759 ();
 FILLCELL_X32 FILLER_182_2791 ();
 FILLCELL_X32 FILLER_182_2823 ();
 FILLCELL_X32 FILLER_182_2855 ();
 FILLCELL_X32 FILLER_182_2887 ();
 FILLCELL_X32 FILLER_182_2919 ();
 FILLCELL_X32 FILLER_182_2951 ();
 FILLCELL_X32 FILLER_182_2983 ();
 FILLCELL_X32 FILLER_182_3015 ();
 FILLCELL_X32 FILLER_182_3047 ();
 FILLCELL_X32 FILLER_182_3079 ();
 FILLCELL_X32 FILLER_182_3111 ();
 FILLCELL_X8 FILLER_182_3143 ();
 FILLCELL_X4 FILLER_182_3151 ();
 FILLCELL_X2 FILLER_182_3155 ();
 FILLCELL_X32 FILLER_182_3158 ();
 FILLCELL_X32 FILLER_182_3190 ();
 FILLCELL_X32 FILLER_182_3222 ();
 FILLCELL_X32 FILLER_182_3254 ();
 FILLCELL_X32 FILLER_182_3286 ();
 FILLCELL_X32 FILLER_182_3318 ();
 FILLCELL_X32 FILLER_182_3350 ();
 FILLCELL_X32 FILLER_182_3382 ();
 FILLCELL_X32 FILLER_182_3414 ();
 FILLCELL_X32 FILLER_182_3446 ();
 FILLCELL_X32 FILLER_182_3478 ();
 FILLCELL_X32 FILLER_182_3510 ();
 FILLCELL_X32 FILLER_182_3542 ();
 FILLCELL_X32 FILLER_182_3574 ();
 FILLCELL_X32 FILLER_182_3606 ();
 FILLCELL_X32 FILLER_182_3638 ();
 FILLCELL_X32 FILLER_182_3670 ();
 FILLCELL_X32 FILLER_182_3702 ();
 FILLCELL_X4 FILLER_182_3734 ();
 FILLCELL_X32 FILLER_183_1 ();
 FILLCELL_X32 FILLER_183_33 ();
 FILLCELL_X32 FILLER_183_65 ();
 FILLCELL_X32 FILLER_183_97 ();
 FILLCELL_X32 FILLER_183_129 ();
 FILLCELL_X32 FILLER_183_161 ();
 FILLCELL_X32 FILLER_183_193 ();
 FILLCELL_X32 FILLER_183_225 ();
 FILLCELL_X32 FILLER_183_257 ();
 FILLCELL_X32 FILLER_183_289 ();
 FILLCELL_X32 FILLER_183_321 ();
 FILLCELL_X32 FILLER_183_353 ();
 FILLCELL_X32 FILLER_183_385 ();
 FILLCELL_X32 FILLER_183_417 ();
 FILLCELL_X32 FILLER_183_449 ();
 FILLCELL_X32 FILLER_183_481 ();
 FILLCELL_X32 FILLER_183_513 ();
 FILLCELL_X32 FILLER_183_545 ();
 FILLCELL_X32 FILLER_183_577 ();
 FILLCELL_X32 FILLER_183_609 ();
 FILLCELL_X32 FILLER_183_641 ();
 FILLCELL_X32 FILLER_183_673 ();
 FILLCELL_X32 FILLER_183_705 ();
 FILLCELL_X32 FILLER_183_737 ();
 FILLCELL_X32 FILLER_183_769 ();
 FILLCELL_X32 FILLER_183_801 ();
 FILLCELL_X32 FILLER_183_833 ();
 FILLCELL_X32 FILLER_183_865 ();
 FILLCELL_X32 FILLER_183_897 ();
 FILLCELL_X32 FILLER_183_929 ();
 FILLCELL_X32 FILLER_183_961 ();
 FILLCELL_X32 FILLER_183_993 ();
 FILLCELL_X32 FILLER_183_1025 ();
 FILLCELL_X32 FILLER_183_1057 ();
 FILLCELL_X32 FILLER_183_1089 ();
 FILLCELL_X32 FILLER_183_1121 ();
 FILLCELL_X32 FILLER_183_1153 ();
 FILLCELL_X32 FILLER_183_1185 ();
 FILLCELL_X32 FILLER_183_1217 ();
 FILLCELL_X8 FILLER_183_1249 ();
 FILLCELL_X4 FILLER_183_1257 ();
 FILLCELL_X2 FILLER_183_1261 ();
 FILLCELL_X32 FILLER_183_1264 ();
 FILLCELL_X32 FILLER_183_1296 ();
 FILLCELL_X32 FILLER_183_1328 ();
 FILLCELL_X32 FILLER_183_1360 ();
 FILLCELL_X32 FILLER_183_1392 ();
 FILLCELL_X32 FILLER_183_1424 ();
 FILLCELL_X32 FILLER_183_1456 ();
 FILLCELL_X32 FILLER_183_1488 ();
 FILLCELL_X32 FILLER_183_1520 ();
 FILLCELL_X32 FILLER_183_1552 ();
 FILLCELL_X32 FILLER_183_1584 ();
 FILLCELL_X32 FILLER_183_1616 ();
 FILLCELL_X32 FILLER_183_1648 ();
 FILLCELL_X32 FILLER_183_1680 ();
 FILLCELL_X32 FILLER_183_1712 ();
 FILLCELL_X32 FILLER_183_1744 ();
 FILLCELL_X32 FILLER_183_1776 ();
 FILLCELL_X32 FILLER_183_1808 ();
 FILLCELL_X32 FILLER_183_1840 ();
 FILLCELL_X32 FILLER_183_1872 ();
 FILLCELL_X32 FILLER_183_1904 ();
 FILLCELL_X32 FILLER_183_1936 ();
 FILLCELL_X32 FILLER_183_1968 ();
 FILLCELL_X32 FILLER_183_2000 ();
 FILLCELL_X32 FILLER_183_2032 ();
 FILLCELL_X32 FILLER_183_2064 ();
 FILLCELL_X32 FILLER_183_2096 ();
 FILLCELL_X32 FILLER_183_2128 ();
 FILLCELL_X32 FILLER_183_2160 ();
 FILLCELL_X32 FILLER_183_2192 ();
 FILLCELL_X32 FILLER_183_2224 ();
 FILLCELL_X32 FILLER_183_2256 ();
 FILLCELL_X32 FILLER_183_2288 ();
 FILLCELL_X32 FILLER_183_2320 ();
 FILLCELL_X32 FILLER_183_2352 ();
 FILLCELL_X32 FILLER_183_2384 ();
 FILLCELL_X32 FILLER_183_2416 ();
 FILLCELL_X32 FILLER_183_2448 ();
 FILLCELL_X32 FILLER_183_2480 ();
 FILLCELL_X8 FILLER_183_2512 ();
 FILLCELL_X4 FILLER_183_2520 ();
 FILLCELL_X2 FILLER_183_2524 ();
 FILLCELL_X32 FILLER_183_2527 ();
 FILLCELL_X32 FILLER_183_2559 ();
 FILLCELL_X32 FILLER_183_2591 ();
 FILLCELL_X32 FILLER_183_2623 ();
 FILLCELL_X32 FILLER_183_2655 ();
 FILLCELL_X32 FILLER_183_2687 ();
 FILLCELL_X32 FILLER_183_2719 ();
 FILLCELL_X32 FILLER_183_2751 ();
 FILLCELL_X32 FILLER_183_2783 ();
 FILLCELL_X32 FILLER_183_2815 ();
 FILLCELL_X32 FILLER_183_2847 ();
 FILLCELL_X32 FILLER_183_2879 ();
 FILLCELL_X32 FILLER_183_2911 ();
 FILLCELL_X32 FILLER_183_2943 ();
 FILLCELL_X32 FILLER_183_2975 ();
 FILLCELL_X32 FILLER_183_3007 ();
 FILLCELL_X32 FILLER_183_3039 ();
 FILLCELL_X32 FILLER_183_3071 ();
 FILLCELL_X32 FILLER_183_3103 ();
 FILLCELL_X32 FILLER_183_3135 ();
 FILLCELL_X32 FILLER_183_3167 ();
 FILLCELL_X32 FILLER_183_3199 ();
 FILLCELL_X32 FILLER_183_3231 ();
 FILLCELL_X32 FILLER_183_3263 ();
 FILLCELL_X32 FILLER_183_3295 ();
 FILLCELL_X32 FILLER_183_3327 ();
 FILLCELL_X32 FILLER_183_3359 ();
 FILLCELL_X32 FILLER_183_3391 ();
 FILLCELL_X32 FILLER_183_3423 ();
 FILLCELL_X32 FILLER_183_3455 ();
 FILLCELL_X32 FILLER_183_3487 ();
 FILLCELL_X32 FILLER_183_3519 ();
 FILLCELL_X32 FILLER_183_3551 ();
 FILLCELL_X32 FILLER_183_3583 ();
 FILLCELL_X32 FILLER_183_3615 ();
 FILLCELL_X32 FILLER_183_3647 ();
 FILLCELL_X32 FILLER_183_3679 ();
 FILLCELL_X16 FILLER_183_3711 ();
 FILLCELL_X8 FILLER_183_3727 ();
 FILLCELL_X2 FILLER_183_3735 ();
 FILLCELL_X1 FILLER_183_3737 ();
 FILLCELL_X32 FILLER_184_1 ();
 FILLCELL_X32 FILLER_184_33 ();
 FILLCELL_X32 FILLER_184_65 ();
 FILLCELL_X32 FILLER_184_97 ();
 FILLCELL_X32 FILLER_184_129 ();
 FILLCELL_X32 FILLER_184_161 ();
 FILLCELL_X32 FILLER_184_193 ();
 FILLCELL_X32 FILLER_184_225 ();
 FILLCELL_X32 FILLER_184_257 ();
 FILLCELL_X32 FILLER_184_289 ();
 FILLCELL_X32 FILLER_184_321 ();
 FILLCELL_X32 FILLER_184_353 ();
 FILLCELL_X32 FILLER_184_385 ();
 FILLCELL_X32 FILLER_184_417 ();
 FILLCELL_X32 FILLER_184_449 ();
 FILLCELL_X32 FILLER_184_481 ();
 FILLCELL_X32 FILLER_184_513 ();
 FILLCELL_X32 FILLER_184_545 ();
 FILLCELL_X32 FILLER_184_577 ();
 FILLCELL_X16 FILLER_184_609 ();
 FILLCELL_X4 FILLER_184_625 ();
 FILLCELL_X2 FILLER_184_629 ();
 FILLCELL_X32 FILLER_184_632 ();
 FILLCELL_X32 FILLER_184_664 ();
 FILLCELL_X32 FILLER_184_696 ();
 FILLCELL_X32 FILLER_184_728 ();
 FILLCELL_X32 FILLER_184_760 ();
 FILLCELL_X32 FILLER_184_792 ();
 FILLCELL_X32 FILLER_184_824 ();
 FILLCELL_X32 FILLER_184_856 ();
 FILLCELL_X32 FILLER_184_888 ();
 FILLCELL_X32 FILLER_184_920 ();
 FILLCELL_X32 FILLER_184_952 ();
 FILLCELL_X32 FILLER_184_984 ();
 FILLCELL_X32 FILLER_184_1016 ();
 FILLCELL_X32 FILLER_184_1048 ();
 FILLCELL_X32 FILLER_184_1080 ();
 FILLCELL_X32 FILLER_184_1112 ();
 FILLCELL_X32 FILLER_184_1144 ();
 FILLCELL_X32 FILLER_184_1176 ();
 FILLCELL_X32 FILLER_184_1208 ();
 FILLCELL_X32 FILLER_184_1240 ();
 FILLCELL_X32 FILLER_184_1272 ();
 FILLCELL_X32 FILLER_184_1304 ();
 FILLCELL_X32 FILLER_184_1336 ();
 FILLCELL_X32 FILLER_184_1368 ();
 FILLCELL_X32 FILLER_184_1400 ();
 FILLCELL_X32 FILLER_184_1432 ();
 FILLCELL_X32 FILLER_184_1464 ();
 FILLCELL_X32 FILLER_184_1496 ();
 FILLCELL_X32 FILLER_184_1528 ();
 FILLCELL_X32 FILLER_184_1560 ();
 FILLCELL_X32 FILLER_184_1592 ();
 FILLCELL_X32 FILLER_184_1624 ();
 FILLCELL_X32 FILLER_184_1656 ();
 FILLCELL_X32 FILLER_184_1688 ();
 FILLCELL_X32 FILLER_184_1720 ();
 FILLCELL_X32 FILLER_184_1752 ();
 FILLCELL_X32 FILLER_184_1784 ();
 FILLCELL_X32 FILLER_184_1816 ();
 FILLCELL_X32 FILLER_184_1848 ();
 FILLCELL_X8 FILLER_184_1880 ();
 FILLCELL_X4 FILLER_184_1888 ();
 FILLCELL_X2 FILLER_184_1892 ();
 FILLCELL_X32 FILLER_184_1895 ();
 FILLCELL_X32 FILLER_184_1927 ();
 FILLCELL_X32 FILLER_184_1959 ();
 FILLCELL_X32 FILLER_184_1991 ();
 FILLCELL_X32 FILLER_184_2023 ();
 FILLCELL_X32 FILLER_184_2055 ();
 FILLCELL_X32 FILLER_184_2087 ();
 FILLCELL_X32 FILLER_184_2119 ();
 FILLCELL_X32 FILLER_184_2151 ();
 FILLCELL_X32 FILLER_184_2183 ();
 FILLCELL_X32 FILLER_184_2215 ();
 FILLCELL_X32 FILLER_184_2247 ();
 FILLCELL_X32 FILLER_184_2279 ();
 FILLCELL_X32 FILLER_184_2311 ();
 FILLCELL_X32 FILLER_184_2343 ();
 FILLCELL_X32 FILLER_184_2375 ();
 FILLCELL_X32 FILLER_184_2407 ();
 FILLCELL_X32 FILLER_184_2439 ();
 FILLCELL_X32 FILLER_184_2471 ();
 FILLCELL_X32 FILLER_184_2503 ();
 FILLCELL_X32 FILLER_184_2535 ();
 FILLCELL_X32 FILLER_184_2567 ();
 FILLCELL_X32 FILLER_184_2599 ();
 FILLCELL_X32 FILLER_184_2631 ();
 FILLCELL_X32 FILLER_184_2663 ();
 FILLCELL_X32 FILLER_184_2695 ();
 FILLCELL_X32 FILLER_184_2727 ();
 FILLCELL_X32 FILLER_184_2759 ();
 FILLCELL_X32 FILLER_184_2791 ();
 FILLCELL_X32 FILLER_184_2823 ();
 FILLCELL_X32 FILLER_184_2855 ();
 FILLCELL_X32 FILLER_184_2887 ();
 FILLCELL_X32 FILLER_184_2919 ();
 FILLCELL_X32 FILLER_184_2951 ();
 FILLCELL_X32 FILLER_184_2983 ();
 FILLCELL_X32 FILLER_184_3015 ();
 FILLCELL_X32 FILLER_184_3047 ();
 FILLCELL_X32 FILLER_184_3079 ();
 FILLCELL_X32 FILLER_184_3111 ();
 FILLCELL_X8 FILLER_184_3143 ();
 FILLCELL_X4 FILLER_184_3151 ();
 FILLCELL_X2 FILLER_184_3155 ();
 FILLCELL_X32 FILLER_184_3158 ();
 FILLCELL_X32 FILLER_184_3190 ();
 FILLCELL_X32 FILLER_184_3222 ();
 FILLCELL_X32 FILLER_184_3254 ();
 FILLCELL_X32 FILLER_184_3286 ();
 FILLCELL_X32 FILLER_184_3318 ();
 FILLCELL_X32 FILLER_184_3350 ();
 FILLCELL_X32 FILLER_184_3382 ();
 FILLCELL_X32 FILLER_184_3414 ();
 FILLCELL_X32 FILLER_184_3446 ();
 FILLCELL_X32 FILLER_184_3478 ();
 FILLCELL_X32 FILLER_184_3510 ();
 FILLCELL_X32 FILLER_184_3542 ();
 FILLCELL_X32 FILLER_184_3574 ();
 FILLCELL_X32 FILLER_184_3606 ();
 FILLCELL_X32 FILLER_184_3638 ();
 FILLCELL_X32 FILLER_184_3670 ();
 FILLCELL_X32 FILLER_184_3702 ();
 FILLCELL_X4 FILLER_184_3734 ();
 FILLCELL_X32 FILLER_185_1 ();
 FILLCELL_X32 FILLER_185_33 ();
 FILLCELL_X32 FILLER_185_65 ();
 FILLCELL_X32 FILLER_185_97 ();
 FILLCELL_X32 FILLER_185_129 ();
 FILLCELL_X32 FILLER_185_161 ();
 FILLCELL_X32 FILLER_185_193 ();
 FILLCELL_X32 FILLER_185_225 ();
 FILLCELL_X32 FILLER_185_257 ();
 FILLCELL_X32 FILLER_185_289 ();
 FILLCELL_X32 FILLER_185_321 ();
 FILLCELL_X32 FILLER_185_353 ();
 FILLCELL_X32 FILLER_185_385 ();
 FILLCELL_X32 FILLER_185_417 ();
 FILLCELL_X32 FILLER_185_449 ();
 FILLCELL_X32 FILLER_185_481 ();
 FILLCELL_X32 FILLER_185_513 ();
 FILLCELL_X32 FILLER_185_545 ();
 FILLCELL_X32 FILLER_185_577 ();
 FILLCELL_X32 FILLER_185_609 ();
 FILLCELL_X32 FILLER_185_641 ();
 FILLCELL_X32 FILLER_185_673 ();
 FILLCELL_X32 FILLER_185_705 ();
 FILLCELL_X32 FILLER_185_737 ();
 FILLCELL_X32 FILLER_185_769 ();
 FILLCELL_X32 FILLER_185_801 ();
 FILLCELL_X32 FILLER_185_833 ();
 FILLCELL_X32 FILLER_185_865 ();
 FILLCELL_X32 FILLER_185_897 ();
 FILLCELL_X32 FILLER_185_929 ();
 FILLCELL_X32 FILLER_185_961 ();
 FILLCELL_X32 FILLER_185_993 ();
 FILLCELL_X32 FILLER_185_1025 ();
 FILLCELL_X32 FILLER_185_1057 ();
 FILLCELL_X32 FILLER_185_1089 ();
 FILLCELL_X32 FILLER_185_1121 ();
 FILLCELL_X32 FILLER_185_1153 ();
 FILLCELL_X32 FILLER_185_1185 ();
 FILLCELL_X32 FILLER_185_1217 ();
 FILLCELL_X8 FILLER_185_1249 ();
 FILLCELL_X4 FILLER_185_1257 ();
 FILLCELL_X2 FILLER_185_1261 ();
 FILLCELL_X32 FILLER_185_1264 ();
 FILLCELL_X32 FILLER_185_1296 ();
 FILLCELL_X32 FILLER_185_1328 ();
 FILLCELL_X32 FILLER_185_1360 ();
 FILLCELL_X32 FILLER_185_1392 ();
 FILLCELL_X32 FILLER_185_1424 ();
 FILLCELL_X32 FILLER_185_1456 ();
 FILLCELL_X32 FILLER_185_1488 ();
 FILLCELL_X32 FILLER_185_1520 ();
 FILLCELL_X32 FILLER_185_1552 ();
 FILLCELL_X32 FILLER_185_1584 ();
 FILLCELL_X32 FILLER_185_1616 ();
 FILLCELL_X32 FILLER_185_1648 ();
 FILLCELL_X32 FILLER_185_1680 ();
 FILLCELL_X32 FILLER_185_1712 ();
 FILLCELL_X32 FILLER_185_1744 ();
 FILLCELL_X32 FILLER_185_1776 ();
 FILLCELL_X32 FILLER_185_1808 ();
 FILLCELL_X32 FILLER_185_1840 ();
 FILLCELL_X32 FILLER_185_1872 ();
 FILLCELL_X32 FILLER_185_1904 ();
 FILLCELL_X32 FILLER_185_1936 ();
 FILLCELL_X32 FILLER_185_1968 ();
 FILLCELL_X32 FILLER_185_2000 ();
 FILLCELL_X32 FILLER_185_2032 ();
 FILLCELL_X32 FILLER_185_2064 ();
 FILLCELL_X32 FILLER_185_2096 ();
 FILLCELL_X32 FILLER_185_2128 ();
 FILLCELL_X32 FILLER_185_2160 ();
 FILLCELL_X32 FILLER_185_2192 ();
 FILLCELL_X32 FILLER_185_2224 ();
 FILLCELL_X32 FILLER_185_2256 ();
 FILLCELL_X32 FILLER_185_2288 ();
 FILLCELL_X32 FILLER_185_2320 ();
 FILLCELL_X32 FILLER_185_2352 ();
 FILLCELL_X32 FILLER_185_2384 ();
 FILLCELL_X32 FILLER_185_2416 ();
 FILLCELL_X32 FILLER_185_2448 ();
 FILLCELL_X32 FILLER_185_2480 ();
 FILLCELL_X8 FILLER_185_2512 ();
 FILLCELL_X4 FILLER_185_2520 ();
 FILLCELL_X2 FILLER_185_2524 ();
 FILLCELL_X32 FILLER_185_2527 ();
 FILLCELL_X32 FILLER_185_2559 ();
 FILLCELL_X32 FILLER_185_2591 ();
 FILLCELL_X32 FILLER_185_2623 ();
 FILLCELL_X32 FILLER_185_2655 ();
 FILLCELL_X32 FILLER_185_2687 ();
 FILLCELL_X32 FILLER_185_2719 ();
 FILLCELL_X32 FILLER_185_2751 ();
 FILLCELL_X32 FILLER_185_2783 ();
 FILLCELL_X32 FILLER_185_2815 ();
 FILLCELL_X32 FILLER_185_2847 ();
 FILLCELL_X32 FILLER_185_2879 ();
 FILLCELL_X32 FILLER_185_2911 ();
 FILLCELL_X32 FILLER_185_2943 ();
 FILLCELL_X32 FILLER_185_2975 ();
 FILLCELL_X32 FILLER_185_3007 ();
 FILLCELL_X32 FILLER_185_3039 ();
 FILLCELL_X32 FILLER_185_3071 ();
 FILLCELL_X32 FILLER_185_3103 ();
 FILLCELL_X32 FILLER_185_3135 ();
 FILLCELL_X32 FILLER_185_3167 ();
 FILLCELL_X32 FILLER_185_3199 ();
 FILLCELL_X32 FILLER_185_3231 ();
 FILLCELL_X32 FILLER_185_3263 ();
 FILLCELL_X32 FILLER_185_3295 ();
 FILLCELL_X32 FILLER_185_3327 ();
 FILLCELL_X32 FILLER_185_3359 ();
 FILLCELL_X32 FILLER_185_3391 ();
 FILLCELL_X32 FILLER_185_3423 ();
 FILLCELL_X32 FILLER_185_3455 ();
 FILLCELL_X32 FILLER_185_3487 ();
 FILLCELL_X32 FILLER_185_3519 ();
 FILLCELL_X32 FILLER_185_3551 ();
 FILLCELL_X32 FILLER_185_3583 ();
 FILLCELL_X32 FILLER_185_3615 ();
 FILLCELL_X32 FILLER_185_3647 ();
 FILLCELL_X32 FILLER_185_3679 ();
 FILLCELL_X16 FILLER_185_3711 ();
 FILLCELL_X8 FILLER_185_3727 ();
 FILLCELL_X2 FILLER_185_3735 ();
 FILLCELL_X1 FILLER_185_3737 ();
 FILLCELL_X32 FILLER_186_1 ();
 FILLCELL_X32 FILLER_186_33 ();
 FILLCELL_X32 FILLER_186_65 ();
 FILLCELL_X32 FILLER_186_97 ();
 FILLCELL_X32 FILLER_186_129 ();
 FILLCELL_X32 FILLER_186_161 ();
 FILLCELL_X32 FILLER_186_193 ();
 FILLCELL_X32 FILLER_186_225 ();
 FILLCELL_X32 FILLER_186_257 ();
 FILLCELL_X32 FILLER_186_289 ();
 FILLCELL_X32 FILLER_186_321 ();
 FILLCELL_X32 FILLER_186_353 ();
 FILLCELL_X32 FILLER_186_385 ();
 FILLCELL_X32 FILLER_186_417 ();
 FILLCELL_X32 FILLER_186_449 ();
 FILLCELL_X32 FILLER_186_481 ();
 FILLCELL_X32 FILLER_186_513 ();
 FILLCELL_X32 FILLER_186_545 ();
 FILLCELL_X32 FILLER_186_577 ();
 FILLCELL_X16 FILLER_186_609 ();
 FILLCELL_X4 FILLER_186_625 ();
 FILLCELL_X2 FILLER_186_629 ();
 FILLCELL_X32 FILLER_186_632 ();
 FILLCELL_X32 FILLER_186_664 ();
 FILLCELL_X32 FILLER_186_696 ();
 FILLCELL_X32 FILLER_186_728 ();
 FILLCELL_X32 FILLER_186_760 ();
 FILLCELL_X32 FILLER_186_792 ();
 FILLCELL_X32 FILLER_186_824 ();
 FILLCELL_X32 FILLER_186_856 ();
 FILLCELL_X32 FILLER_186_888 ();
 FILLCELL_X32 FILLER_186_920 ();
 FILLCELL_X32 FILLER_186_952 ();
 FILLCELL_X32 FILLER_186_984 ();
 FILLCELL_X32 FILLER_186_1016 ();
 FILLCELL_X32 FILLER_186_1048 ();
 FILLCELL_X32 FILLER_186_1080 ();
 FILLCELL_X32 FILLER_186_1112 ();
 FILLCELL_X32 FILLER_186_1144 ();
 FILLCELL_X32 FILLER_186_1176 ();
 FILLCELL_X32 FILLER_186_1208 ();
 FILLCELL_X32 FILLER_186_1240 ();
 FILLCELL_X32 FILLER_186_1272 ();
 FILLCELL_X32 FILLER_186_1304 ();
 FILLCELL_X32 FILLER_186_1336 ();
 FILLCELL_X32 FILLER_186_1368 ();
 FILLCELL_X32 FILLER_186_1400 ();
 FILLCELL_X32 FILLER_186_1432 ();
 FILLCELL_X32 FILLER_186_1464 ();
 FILLCELL_X32 FILLER_186_1496 ();
 FILLCELL_X32 FILLER_186_1528 ();
 FILLCELL_X32 FILLER_186_1560 ();
 FILLCELL_X32 FILLER_186_1592 ();
 FILLCELL_X32 FILLER_186_1624 ();
 FILLCELL_X32 FILLER_186_1656 ();
 FILLCELL_X32 FILLER_186_1688 ();
 FILLCELL_X32 FILLER_186_1720 ();
 FILLCELL_X32 FILLER_186_1752 ();
 FILLCELL_X32 FILLER_186_1784 ();
 FILLCELL_X32 FILLER_186_1816 ();
 FILLCELL_X32 FILLER_186_1848 ();
 FILLCELL_X8 FILLER_186_1880 ();
 FILLCELL_X4 FILLER_186_1888 ();
 FILLCELL_X2 FILLER_186_1892 ();
 FILLCELL_X32 FILLER_186_1895 ();
 FILLCELL_X32 FILLER_186_1927 ();
 FILLCELL_X32 FILLER_186_1959 ();
 FILLCELL_X32 FILLER_186_1991 ();
 FILLCELL_X32 FILLER_186_2023 ();
 FILLCELL_X32 FILLER_186_2055 ();
 FILLCELL_X32 FILLER_186_2087 ();
 FILLCELL_X32 FILLER_186_2119 ();
 FILLCELL_X32 FILLER_186_2151 ();
 FILLCELL_X32 FILLER_186_2183 ();
 FILLCELL_X32 FILLER_186_2215 ();
 FILLCELL_X32 FILLER_186_2247 ();
 FILLCELL_X32 FILLER_186_2279 ();
 FILLCELL_X32 FILLER_186_2311 ();
 FILLCELL_X32 FILLER_186_2343 ();
 FILLCELL_X32 FILLER_186_2375 ();
 FILLCELL_X32 FILLER_186_2407 ();
 FILLCELL_X32 FILLER_186_2439 ();
 FILLCELL_X32 FILLER_186_2471 ();
 FILLCELL_X32 FILLER_186_2503 ();
 FILLCELL_X32 FILLER_186_2535 ();
 FILLCELL_X32 FILLER_186_2567 ();
 FILLCELL_X32 FILLER_186_2599 ();
 FILLCELL_X32 FILLER_186_2631 ();
 FILLCELL_X32 FILLER_186_2663 ();
 FILLCELL_X32 FILLER_186_2695 ();
 FILLCELL_X32 FILLER_186_2727 ();
 FILLCELL_X32 FILLER_186_2759 ();
 FILLCELL_X32 FILLER_186_2791 ();
 FILLCELL_X32 FILLER_186_2823 ();
 FILLCELL_X32 FILLER_186_2855 ();
 FILLCELL_X32 FILLER_186_2887 ();
 FILLCELL_X32 FILLER_186_2919 ();
 FILLCELL_X32 FILLER_186_2951 ();
 FILLCELL_X32 FILLER_186_2983 ();
 FILLCELL_X32 FILLER_186_3015 ();
 FILLCELL_X32 FILLER_186_3047 ();
 FILLCELL_X32 FILLER_186_3079 ();
 FILLCELL_X32 FILLER_186_3111 ();
 FILLCELL_X8 FILLER_186_3143 ();
 FILLCELL_X4 FILLER_186_3151 ();
 FILLCELL_X2 FILLER_186_3155 ();
 FILLCELL_X32 FILLER_186_3158 ();
 FILLCELL_X32 FILLER_186_3190 ();
 FILLCELL_X32 FILLER_186_3222 ();
 FILLCELL_X32 FILLER_186_3254 ();
 FILLCELL_X32 FILLER_186_3286 ();
 FILLCELL_X32 FILLER_186_3318 ();
 FILLCELL_X32 FILLER_186_3350 ();
 FILLCELL_X32 FILLER_186_3382 ();
 FILLCELL_X32 FILLER_186_3414 ();
 FILLCELL_X32 FILLER_186_3446 ();
 FILLCELL_X32 FILLER_186_3478 ();
 FILLCELL_X32 FILLER_186_3510 ();
 FILLCELL_X32 FILLER_186_3542 ();
 FILLCELL_X32 FILLER_186_3574 ();
 FILLCELL_X32 FILLER_186_3606 ();
 FILLCELL_X32 FILLER_186_3638 ();
 FILLCELL_X32 FILLER_186_3670 ();
 FILLCELL_X32 FILLER_186_3702 ();
 FILLCELL_X4 FILLER_186_3734 ();
 FILLCELL_X32 FILLER_187_1 ();
 FILLCELL_X32 FILLER_187_33 ();
 FILLCELL_X32 FILLER_187_65 ();
 FILLCELL_X32 FILLER_187_97 ();
 FILLCELL_X32 FILLER_187_129 ();
 FILLCELL_X32 FILLER_187_161 ();
 FILLCELL_X32 FILLER_187_193 ();
 FILLCELL_X32 FILLER_187_225 ();
 FILLCELL_X32 FILLER_187_257 ();
 FILLCELL_X32 FILLER_187_289 ();
 FILLCELL_X32 FILLER_187_321 ();
 FILLCELL_X32 FILLER_187_353 ();
 FILLCELL_X32 FILLER_187_385 ();
 FILLCELL_X32 FILLER_187_417 ();
 FILLCELL_X32 FILLER_187_449 ();
 FILLCELL_X32 FILLER_187_481 ();
 FILLCELL_X32 FILLER_187_513 ();
 FILLCELL_X32 FILLER_187_545 ();
 FILLCELL_X32 FILLER_187_577 ();
 FILLCELL_X32 FILLER_187_609 ();
 FILLCELL_X32 FILLER_187_641 ();
 FILLCELL_X32 FILLER_187_673 ();
 FILLCELL_X32 FILLER_187_705 ();
 FILLCELL_X32 FILLER_187_737 ();
 FILLCELL_X32 FILLER_187_769 ();
 FILLCELL_X32 FILLER_187_801 ();
 FILLCELL_X32 FILLER_187_833 ();
 FILLCELL_X32 FILLER_187_865 ();
 FILLCELL_X32 FILLER_187_897 ();
 FILLCELL_X32 FILLER_187_929 ();
 FILLCELL_X32 FILLER_187_961 ();
 FILLCELL_X32 FILLER_187_993 ();
 FILLCELL_X32 FILLER_187_1025 ();
 FILLCELL_X32 FILLER_187_1057 ();
 FILLCELL_X32 FILLER_187_1089 ();
 FILLCELL_X32 FILLER_187_1121 ();
 FILLCELL_X32 FILLER_187_1153 ();
 FILLCELL_X32 FILLER_187_1185 ();
 FILLCELL_X32 FILLER_187_1217 ();
 FILLCELL_X8 FILLER_187_1249 ();
 FILLCELL_X4 FILLER_187_1257 ();
 FILLCELL_X2 FILLER_187_1261 ();
 FILLCELL_X32 FILLER_187_1264 ();
 FILLCELL_X32 FILLER_187_1296 ();
 FILLCELL_X32 FILLER_187_1328 ();
 FILLCELL_X32 FILLER_187_1360 ();
 FILLCELL_X32 FILLER_187_1392 ();
 FILLCELL_X32 FILLER_187_1424 ();
 FILLCELL_X32 FILLER_187_1456 ();
 FILLCELL_X32 FILLER_187_1488 ();
 FILLCELL_X32 FILLER_187_1520 ();
 FILLCELL_X32 FILLER_187_1552 ();
 FILLCELL_X32 FILLER_187_1584 ();
 FILLCELL_X32 FILLER_187_1616 ();
 FILLCELL_X32 FILLER_187_1648 ();
 FILLCELL_X32 FILLER_187_1680 ();
 FILLCELL_X32 FILLER_187_1712 ();
 FILLCELL_X32 FILLER_187_1744 ();
 FILLCELL_X32 FILLER_187_1776 ();
 FILLCELL_X32 FILLER_187_1808 ();
 FILLCELL_X32 FILLER_187_1840 ();
 FILLCELL_X32 FILLER_187_1872 ();
 FILLCELL_X32 FILLER_187_1904 ();
 FILLCELL_X32 FILLER_187_1936 ();
 FILLCELL_X32 FILLER_187_1968 ();
 FILLCELL_X32 FILLER_187_2000 ();
 FILLCELL_X32 FILLER_187_2032 ();
 FILLCELL_X32 FILLER_187_2064 ();
 FILLCELL_X32 FILLER_187_2096 ();
 FILLCELL_X32 FILLER_187_2128 ();
 FILLCELL_X32 FILLER_187_2160 ();
 FILLCELL_X32 FILLER_187_2192 ();
 FILLCELL_X32 FILLER_187_2224 ();
 FILLCELL_X32 FILLER_187_2256 ();
 FILLCELL_X32 FILLER_187_2288 ();
 FILLCELL_X32 FILLER_187_2320 ();
 FILLCELL_X32 FILLER_187_2352 ();
 FILLCELL_X32 FILLER_187_2384 ();
 FILLCELL_X32 FILLER_187_2416 ();
 FILLCELL_X32 FILLER_187_2448 ();
 FILLCELL_X32 FILLER_187_2480 ();
 FILLCELL_X8 FILLER_187_2512 ();
 FILLCELL_X4 FILLER_187_2520 ();
 FILLCELL_X2 FILLER_187_2524 ();
 FILLCELL_X32 FILLER_187_2527 ();
 FILLCELL_X32 FILLER_187_2559 ();
 FILLCELL_X32 FILLER_187_2591 ();
 FILLCELL_X32 FILLER_187_2623 ();
 FILLCELL_X32 FILLER_187_2655 ();
 FILLCELL_X32 FILLER_187_2687 ();
 FILLCELL_X32 FILLER_187_2719 ();
 FILLCELL_X32 FILLER_187_2751 ();
 FILLCELL_X32 FILLER_187_2783 ();
 FILLCELL_X32 FILLER_187_2815 ();
 FILLCELL_X32 FILLER_187_2847 ();
 FILLCELL_X32 FILLER_187_2879 ();
 FILLCELL_X32 FILLER_187_2911 ();
 FILLCELL_X32 FILLER_187_2943 ();
 FILLCELL_X32 FILLER_187_2975 ();
 FILLCELL_X32 FILLER_187_3007 ();
 FILLCELL_X32 FILLER_187_3039 ();
 FILLCELL_X32 FILLER_187_3071 ();
 FILLCELL_X32 FILLER_187_3103 ();
 FILLCELL_X32 FILLER_187_3135 ();
 FILLCELL_X32 FILLER_187_3167 ();
 FILLCELL_X32 FILLER_187_3199 ();
 FILLCELL_X32 FILLER_187_3231 ();
 FILLCELL_X32 FILLER_187_3263 ();
 FILLCELL_X32 FILLER_187_3295 ();
 FILLCELL_X32 FILLER_187_3327 ();
 FILLCELL_X32 FILLER_187_3359 ();
 FILLCELL_X32 FILLER_187_3391 ();
 FILLCELL_X32 FILLER_187_3423 ();
 FILLCELL_X32 FILLER_187_3455 ();
 FILLCELL_X32 FILLER_187_3487 ();
 FILLCELL_X32 FILLER_187_3519 ();
 FILLCELL_X32 FILLER_187_3551 ();
 FILLCELL_X32 FILLER_187_3583 ();
 FILLCELL_X32 FILLER_187_3615 ();
 FILLCELL_X32 FILLER_187_3647 ();
 FILLCELL_X32 FILLER_187_3679 ();
 FILLCELL_X16 FILLER_187_3711 ();
 FILLCELL_X8 FILLER_187_3727 ();
 FILLCELL_X2 FILLER_187_3735 ();
 FILLCELL_X1 FILLER_187_3737 ();
 FILLCELL_X32 FILLER_188_1 ();
 FILLCELL_X32 FILLER_188_33 ();
 FILLCELL_X32 FILLER_188_65 ();
 FILLCELL_X32 FILLER_188_97 ();
 FILLCELL_X32 FILLER_188_129 ();
 FILLCELL_X32 FILLER_188_161 ();
 FILLCELL_X32 FILLER_188_193 ();
 FILLCELL_X32 FILLER_188_225 ();
 FILLCELL_X32 FILLER_188_257 ();
 FILLCELL_X32 FILLER_188_289 ();
 FILLCELL_X32 FILLER_188_321 ();
 FILLCELL_X32 FILLER_188_353 ();
 FILLCELL_X32 FILLER_188_385 ();
 FILLCELL_X32 FILLER_188_417 ();
 FILLCELL_X32 FILLER_188_449 ();
 FILLCELL_X32 FILLER_188_481 ();
 FILLCELL_X32 FILLER_188_513 ();
 FILLCELL_X32 FILLER_188_545 ();
 FILLCELL_X32 FILLER_188_577 ();
 FILLCELL_X16 FILLER_188_609 ();
 FILLCELL_X4 FILLER_188_625 ();
 FILLCELL_X2 FILLER_188_629 ();
 FILLCELL_X32 FILLER_188_632 ();
 FILLCELL_X32 FILLER_188_664 ();
 FILLCELL_X32 FILLER_188_696 ();
 FILLCELL_X32 FILLER_188_728 ();
 FILLCELL_X32 FILLER_188_760 ();
 FILLCELL_X32 FILLER_188_792 ();
 FILLCELL_X32 FILLER_188_824 ();
 FILLCELL_X32 FILLER_188_856 ();
 FILLCELL_X32 FILLER_188_888 ();
 FILLCELL_X32 FILLER_188_920 ();
 FILLCELL_X32 FILLER_188_952 ();
 FILLCELL_X32 FILLER_188_984 ();
 FILLCELL_X32 FILLER_188_1016 ();
 FILLCELL_X32 FILLER_188_1048 ();
 FILLCELL_X32 FILLER_188_1080 ();
 FILLCELL_X32 FILLER_188_1112 ();
 FILLCELL_X32 FILLER_188_1144 ();
 FILLCELL_X32 FILLER_188_1176 ();
 FILLCELL_X32 FILLER_188_1208 ();
 FILLCELL_X32 FILLER_188_1240 ();
 FILLCELL_X32 FILLER_188_1272 ();
 FILLCELL_X32 FILLER_188_1304 ();
 FILLCELL_X32 FILLER_188_1336 ();
 FILLCELL_X32 FILLER_188_1368 ();
 FILLCELL_X32 FILLER_188_1400 ();
 FILLCELL_X32 FILLER_188_1432 ();
 FILLCELL_X32 FILLER_188_1464 ();
 FILLCELL_X32 FILLER_188_1496 ();
 FILLCELL_X32 FILLER_188_1528 ();
 FILLCELL_X32 FILLER_188_1560 ();
 FILLCELL_X32 FILLER_188_1592 ();
 FILLCELL_X32 FILLER_188_1624 ();
 FILLCELL_X32 FILLER_188_1656 ();
 FILLCELL_X32 FILLER_188_1688 ();
 FILLCELL_X32 FILLER_188_1720 ();
 FILLCELL_X32 FILLER_188_1752 ();
 FILLCELL_X32 FILLER_188_1784 ();
 FILLCELL_X32 FILLER_188_1816 ();
 FILLCELL_X32 FILLER_188_1848 ();
 FILLCELL_X8 FILLER_188_1880 ();
 FILLCELL_X4 FILLER_188_1888 ();
 FILLCELL_X2 FILLER_188_1892 ();
 FILLCELL_X32 FILLER_188_1895 ();
 FILLCELL_X32 FILLER_188_1927 ();
 FILLCELL_X32 FILLER_188_1959 ();
 FILLCELL_X32 FILLER_188_1991 ();
 FILLCELL_X32 FILLER_188_2023 ();
 FILLCELL_X32 FILLER_188_2055 ();
 FILLCELL_X32 FILLER_188_2087 ();
 FILLCELL_X32 FILLER_188_2119 ();
 FILLCELL_X32 FILLER_188_2151 ();
 FILLCELL_X32 FILLER_188_2183 ();
 FILLCELL_X32 FILLER_188_2215 ();
 FILLCELL_X32 FILLER_188_2247 ();
 FILLCELL_X32 FILLER_188_2279 ();
 FILLCELL_X32 FILLER_188_2311 ();
 FILLCELL_X32 FILLER_188_2343 ();
 FILLCELL_X32 FILLER_188_2375 ();
 FILLCELL_X32 FILLER_188_2407 ();
 FILLCELL_X32 FILLER_188_2439 ();
 FILLCELL_X32 FILLER_188_2471 ();
 FILLCELL_X32 FILLER_188_2503 ();
 FILLCELL_X32 FILLER_188_2535 ();
 FILLCELL_X32 FILLER_188_2567 ();
 FILLCELL_X32 FILLER_188_2599 ();
 FILLCELL_X32 FILLER_188_2631 ();
 FILLCELL_X32 FILLER_188_2663 ();
 FILLCELL_X32 FILLER_188_2695 ();
 FILLCELL_X32 FILLER_188_2727 ();
 FILLCELL_X32 FILLER_188_2759 ();
 FILLCELL_X32 FILLER_188_2791 ();
 FILLCELL_X32 FILLER_188_2823 ();
 FILLCELL_X32 FILLER_188_2855 ();
 FILLCELL_X32 FILLER_188_2887 ();
 FILLCELL_X32 FILLER_188_2919 ();
 FILLCELL_X32 FILLER_188_2951 ();
 FILLCELL_X32 FILLER_188_2983 ();
 FILLCELL_X32 FILLER_188_3015 ();
 FILLCELL_X32 FILLER_188_3047 ();
 FILLCELL_X32 FILLER_188_3079 ();
 FILLCELL_X32 FILLER_188_3111 ();
 FILLCELL_X8 FILLER_188_3143 ();
 FILLCELL_X4 FILLER_188_3151 ();
 FILLCELL_X2 FILLER_188_3155 ();
 FILLCELL_X32 FILLER_188_3158 ();
 FILLCELL_X32 FILLER_188_3190 ();
 FILLCELL_X32 FILLER_188_3222 ();
 FILLCELL_X32 FILLER_188_3254 ();
 FILLCELL_X32 FILLER_188_3286 ();
 FILLCELL_X32 FILLER_188_3318 ();
 FILLCELL_X32 FILLER_188_3350 ();
 FILLCELL_X32 FILLER_188_3382 ();
 FILLCELL_X32 FILLER_188_3414 ();
 FILLCELL_X32 FILLER_188_3446 ();
 FILLCELL_X32 FILLER_188_3478 ();
 FILLCELL_X32 FILLER_188_3510 ();
 FILLCELL_X32 FILLER_188_3542 ();
 FILLCELL_X32 FILLER_188_3574 ();
 FILLCELL_X32 FILLER_188_3606 ();
 FILLCELL_X32 FILLER_188_3638 ();
 FILLCELL_X32 FILLER_188_3670 ();
 FILLCELL_X32 FILLER_188_3702 ();
 FILLCELL_X4 FILLER_188_3734 ();
 FILLCELL_X32 FILLER_189_1 ();
 FILLCELL_X32 FILLER_189_33 ();
 FILLCELL_X32 FILLER_189_65 ();
 FILLCELL_X32 FILLER_189_97 ();
 FILLCELL_X32 FILLER_189_129 ();
 FILLCELL_X32 FILLER_189_161 ();
 FILLCELL_X32 FILLER_189_193 ();
 FILLCELL_X32 FILLER_189_225 ();
 FILLCELL_X32 FILLER_189_257 ();
 FILLCELL_X32 FILLER_189_289 ();
 FILLCELL_X32 FILLER_189_321 ();
 FILLCELL_X32 FILLER_189_353 ();
 FILLCELL_X32 FILLER_189_385 ();
 FILLCELL_X32 FILLER_189_417 ();
 FILLCELL_X32 FILLER_189_449 ();
 FILLCELL_X32 FILLER_189_481 ();
 FILLCELL_X32 FILLER_189_513 ();
 FILLCELL_X32 FILLER_189_545 ();
 FILLCELL_X32 FILLER_189_577 ();
 FILLCELL_X32 FILLER_189_609 ();
 FILLCELL_X32 FILLER_189_641 ();
 FILLCELL_X32 FILLER_189_673 ();
 FILLCELL_X32 FILLER_189_705 ();
 FILLCELL_X32 FILLER_189_737 ();
 FILLCELL_X32 FILLER_189_769 ();
 FILLCELL_X32 FILLER_189_801 ();
 FILLCELL_X32 FILLER_189_833 ();
 FILLCELL_X32 FILLER_189_865 ();
 FILLCELL_X32 FILLER_189_897 ();
 FILLCELL_X32 FILLER_189_929 ();
 FILLCELL_X32 FILLER_189_961 ();
 FILLCELL_X32 FILLER_189_993 ();
 FILLCELL_X32 FILLER_189_1025 ();
 FILLCELL_X32 FILLER_189_1057 ();
 FILLCELL_X32 FILLER_189_1089 ();
 FILLCELL_X32 FILLER_189_1121 ();
 FILLCELL_X32 FILLER_189_1153 ();
 FILLCELL_X32 FILLER_189_1185 ();
 FILLCELL_X32 FILLER_189_1217 ();
 FILLCELL_X8 FILLER_189_1249 ();
 FILLCELL_X4 FILLER_189_1257 ();
 FILLCELL_X2 FILLER_189_1261 ();
 FILLCELL_X32 FILLER_189_1264 ();
 FILLCELL_X32 FILLER_189_1296 ();
 FILLCELL_X32 FILLER_189_1328 ();
 FILLCELL_X32 FILLER_189_1360 ();
 FILLCELL_X32 FILLER_189_1392 ();
 FILLCELL_X32 FILLER_189_1424 ();
 FILLCELL_X32 FILLER_189_1456 ();
 FILLCELL_X32 FILLER_189_1488 ();
 FILLCELL_X32 FILLER_189_1520 ();
 FILLCELL_X32 FILLER_189_1552 ();
 FILLCELL_X32 FILLER_189_1584 ();
 FILLCELL_X32 FILLER_189_1616 ();
 FILLCELL_X32 FILLER_189_1648 ();
 FILLCELL_X32 FILLER_189_1680 ();
 FILLCELL_X32 FILLER_189_1712 ();
 FILLCELL_X32 FILLER_189_1744 ();
 FILLCELL_X32 FILLER_189_1776 ();
 FILLCELL_X32 FILLER_189_1808 ();
 FILLCELL_X32 FILLER_189_1840 ();
 FILLCELL_X32 FILLER_189_1872 ();
 FILLCELL_X32 FILLER_189_1904 ();
 FILLCELL_X32 FILLER_189_1936 ();
 FILLCELL_X32 FILLER_189_1968 ();
 FILLCELL_X32 FILLER_189_2000 ();
 FILLCELL_X32 FILLER_189_2032 ();
 FILLCELL_X32 FILLER_189_2064 ();
 FILLCELL_X32 FILLER_189_2096 ();
 FILLCELL_X32 FILLER_189_2128 ();
 FILLCELL_X32 FILLER_189_2160 ();
 FILLCELL_X32 FILLER_189_2192 ();
 FILLCELL_X32 FILLER_189_2224 ();
 FILLCELL_X32 FILLER_189_2256 ();
 FILLCELL_X32 FILLER_189_2288 ();
 FILLCELL_X32 FILLER_189_2320 ();
 FILLCELL_X32 FILLER_189_2352 ();
 FILLCELL_X32 FILLER_189_2384 ();
 FILLCELL_X32 FILLER_189_2416 ();
 FILLCELL_X32 FILLER_189_2448 ();
 FILLCELL_X32 FILLER_189_2480 ();
 FILLCELL_X8 FILLER_189_2512 ();
 FILLCELL_X4 FILLER_189_2520 ();
 FILLCELL_X2 FILLER_189_2524 ();
 FILLCELL_X32 FILLER_189_2527 ();
 FILLCELL_X32 FILLER_189_2559 ();
 FILLCELL_X32 FILLER_189_2591 ();
 FILLCELL_X32 FILLER_189_2623 ();
 FILLCELL_X32 FILLER_189_2655 ();
 FILLCELL_X32 FILLER_189_2687 ();
 FILLCELL_X32 FILLER_189_2719 ();
 FILLCELL_X32 FILLER_189_2751 ();
 FILLCELL_X32 FILLER_189_2783 ();
 FILLCELL_X32 FILLER_189_2815 ();
 FILLCELL_X32 FILLER_189_2847 ();
 FILLCELL_X32 FILLER_189_2879 ();
 FILLCELL_X32 FILLER_189_2911 ();
 FILLCELL_X32 FILLER_189_2943 ();
 FILLCELL_X32 FILLER_189_2975 ();
 FILLCELL_X32 FILLER_189_3007 ();
 FILLCELL_X32 FILLER_189_3039 ();
 FILLCELL_X32 FILLER_189_3071 ();
 FILLCELL_X32 FILLER_189_3103 ();
 FILLCELL_X32 FILLER_189_3135 ();
 FILLCELL_X32 FILLER_189_3167 ();
 FILLCELL_X32 FILLER_189_3199 ();
 FILLCELL_X32 FILLER_189_3231 ();
 FILLCELL_X32 FILLER_189_3263 ();
 FILLCELL_X32 FILLER_189_3295 ();
 FILLCELL_X32 FILLER_189_3327 ();
 FILLCELL_X32 FILLER_189_3359 ();
 FILLCELL_X32 FILLER_189_3391 ();
 FILLCELL_X32 FILLER_189_3423 ();
 FILLCELL_X32 FILLER_189_3455 ();
 FILLCELL_X32 FILLER_189_3487 ();
 FILLCELL_X32 FILLER_189_3519 ();
 FILLCELL_X32 FILLER_189_3551 ();
 FILLCELL_X32 FILLER_189_3583 ();
 FILLCELL_X32 FILLER_189_3615 ();
 FILLCELL_X32 FILLER_189_3647 ();
 FILLCELL_X32 FILLER_189_3679 ();
 FILLCELL_X16 FILLER_189_3711 ();
 FILLCELL_X8 FILLER_189_3727 ();
 FILLCELL_X2 FILLER_189_3735 ();
 FILLCELL_X1 FILLER_189_3737 ();
 FILLCELL_X32 FILLER_190_1 ();
 FILLCELL_X32 FILLER_190_33 ();
 FILLCELL_X32 FILLER_190_65 ();
 FILLCELL_X32 FILLER_190_97 ();
 FILLCELL_X32 FILLER_190_129 ();
 FILLCELL_X32 FILLER_190_161 ();
 FILLCELL_X32 FILLER_190_193 ();
 FILLCELL_X32 FILLER_190_225 ();
 FILLCELL_X32 FILLER_190_257 ();
 FILLCELL_X32 FILLER_190_289 ();
 FILLCELL_X32 FILLER_190_321 ();
 FILLCELL_X32 FILLER_190_353 ();
 FILLCELL_X32 FILLER_190_385 ();
 FILLCELL_X32 FILLER_190_417 ();
 FILLCELL_X32 FILLER_190_449 ();
 FILLCELL_X32 FILLER_190_481 ();
 FILLCELL_X32 FILLER_190_513 ();
 FILLCELL_X32 FILLER_190_545 ();
 FILLCELL_X32 FILLER_190_577 ();
 FILLCELL_X16 FILLER_190_609 ();
 FILLCELL_X4 FILLER_190_625 ();
 FILLCELL_X2 FILLER_190_629 ();
 FILLCELL_X32 FILLER_190_632 ();
 FILLCELL_X32 FILLER_190_664 ();
 FILLCELL_X32 FILLER_190_696 ();
 FILLCELL_X32 FILLER_190_728 ();
 FILLCELL_X32 FILLER_190_760 ();
 FILLCELL_X32 FILLER_190_792 ();
 FILLCELL_X32 FILLER_190_824 ();
 FILLCELL_X32 FILLER_190_856 ();
 FILLCELL_X32 FILLER_190_888 ();
 FILLCELL_X32 FILLER_190_920 ();
 FILLCELL_X32 FILLER_190_952 ();
 FILLCELL_X32 FILLER_190_984 ();
 FILLCELL_X32 FILLER_190_1016 ();
 FILLCELL_X32 FILLER_190_1048 ();
 FILLCELL_X32 FILLER_190_1080 ();
 FILLCELL_X32 FILLER_190_1112 ();
 FILLCELL_X32 FILLER_190_1144 ();
 FILLCELL_X32 FILLER_190_1176 ();
 FILLCELL_X32 FILLER_190_1208 ();
 FILLCELL_X32 FILLER_190_1240 ();
 FILLCELL_X32 FILLER_190_1272 ();
 FILLCELL_X32 FILLER_190_1304 ();
 FILLCELL_X32 FILLER_190_1336 ();
 FILLCELL_X32 FILLER_190_1368 ();
 FILLCELL_X32 FILLER_190_1400 ();
 FILLCELL_X32 FILLER_190_1432 ();
 FILLCELL_X32 FILLER_190_1464 ();
 FILLCELL_X32 FILLER_190_1496 ();
 FILLCELL_X32 FILLER_190_1528 ();
 FILLCELL_X32 FILLER_190_1560 ();
 FILLCELL_X32 FILLER_190_1592 ();
 FILLCELL_X32 FILLER_190_1624 ();
 FILLCELL_X32 FILLER_190_1656 ();
 FILLCELL_X32 FILLER_190_1688 ();
 FILLCELL_X32 FILLER_190_1720 ();
 FILLCELL_X32 FILLER_190_1752 ();
 FILLCELL_X32 FILLER_190_1784 ();
 FILLCELL_X32 FILLER_190_1816 ();
 FILLCELL_X32 FILLER_190_1848 ();
 FILLCELL_X8 FILLER_190_1880 ();
 FILLCELL_X4 FILLER_190_1888 ();
 FILLCELL_X2 FILLER_190_1892 ();
 FILLCELL_X32 FILLER_190_1895 ();
 FILLCELL_X32 FILLER_190_1927 ();
 FILLCELL_X32 FILLER_190_1959 ();
 FILLCELL_X32 FILLER_190_1991 ();
 FILLCELL_X32 FILLER_190_2023 ();
 FILLCELL_X32 FILLER_190_2055 ();
 FILLCELL_X32 FILLER_190_2087 ();
 FILLCELL_X32 FILLER_190_2119 ();
 FILLCELL_X32 FILLER_190_2151 ();
 FILLCELL_X32 FILLER_190_2183 ();
 FILLCELL_X32 FILLER_190_2215 ();
 FILLCELL_X32 FILLER_190_2247 ();
 FILLCELL_X32 FILLER_190_2279 ();
 FILLCELL_X32 FILLER_190_2311 ();
 FILLCELL_X32 FILLER_190_2343 ();
 FILLCELL_X32 FILLER_190_2375 ();
 FILLCELL_X32 FILLER_190_2407 ();
 FILLCELL_X32 FILLER_190_2439 ();
 FILLCELL_X32 FILLER_190_2471 ();
 FILLCELL_X32 FILLER_190_2503 ();
 FILLCELL_X32 FILLER_190_2535 ();
 FILLCELL_X32 FILLER_190_2567 ();
 FILLCELL_X32 FILLER_190_2599 ();
 FILLCELL_X32 FILLER_190_2631 ();
 FILLCELL_X32 FILLER_190_2663 ();
 FILLCELL_X32 FILLER_190_2695 ();
 FILLCELL_X32 FILLER_190_2727 ();
 FILLCELL_X32 FILLER_190_2759 ();
 FILLCELL_X32 FILLER_190_2791 ();
 FILLCELL_X32 FILLER_190_2823 ();
 FILLCELL_X32 FILLER_190_2855 ();
 FILLCELL_X32 FILLER_190_2887 ();
 FILLCELL_X32 FILLER_190_2919 ();
 FILLCELL_X32 FILLER_190_2951 ();
 FILLCELL_X32 FILLER_190_2983 ();
 FILLCELL_X32 FILLER_190_3015 ();
 FILLCELL_X32 FILLER_190_3047 ();
 FILLCELL_X32 FILLER_190_3079 ();
 FILLCELL_X32 FILLER_190_3111 ();
 FILLCELL_X8 FILLER_190_3143 ();
 FILLCELL_X4 FILLER_190_3151 ();
 FILLCELL_X2 FILLER_190_3155 ();
 FILLCELL_X32 FILLER_190_3158 ();
 FILLCELL_X32 FILLER_190_3190 ();
 FILLCELL_X32 FILLER_190_3222 ();
 FILLCELL_X32 FILLER_190_3254 ();
 FILLCELL_X32 FILLER_190_3286 ();
 FILLCELL_X32 FILLER_190_3318 ();
 FILLCELL_X32 FILLER_190_3350 ();
 FILLCELL_X32 FILLER_190_3382 ();
 FILLCELL_X32 FILLER_190_3414 ();
 FILLCELL_X32 FILLER_190_3446 ();
 FILLCELL_X32 FILLER_190_3478 ();
 FILLCELL_X32 FILLER_190_3510 ();
 FILLCELL_X32 FILLER_190_3542 ();
 FILLCELL_X32 FILLER_190_3574 ();
 FILLCELL_X32 FILLER_190_3606 ();
 FILLCELL_X32 FILLER_190_3638 ();
 FILLCELL_X32 FILLER_190_3670 ();
 FILLCELL_X32 FILLER_190_3702 ();
 FILLCELL_X4 FILLER_190_3734 ();
 FILLCELL_X32 FILLER_191_1 ();
 FILLCELL_X32 FILLER_191_33 ();
 FILLCELL_X32 FILLER_191_65 ();
 FILLCELL_X32 FILLER_191_97 ();
 FILLCELL_X32 FILLER_191_129 ();
 FILLCELL_X32 FILLER_191_161 ();
 FILLCELL_X32 FILLER_191_193 ();
 FILLCELL_X32 FILLER_191_225 ();
 FILLCELL_X32 FILLER_191_257 ();
 FILLCELL_X32 FILLER_191_289 ();
 FILLCELL_X32 FILLER_191_321 ();
 FILLCELL_X32 FILLER_191_353 ();
 FILLCELL_X32 FILLER_191_385 ();
 FILLCELL_X32 FILLER_191_417 ();
 FILLCELL_X32 FILLER_191_449 ();
 FILLCELL_X32 FILLER_191_481 ();
 FILLCELL_X32 FILLER_191_513 ();
 FILLCELL_X32 FILLER_191_545 ();
 FILLCELL_X32 FILLER_191_577 ();
 FILLCELL_X32 FILLER_191_609 ();
 FILLCELL_X32 FILLER_191_641 ();
 FILLCELL_X32 FILLER_191_673 ();
 FILLCELL_X32 FILLER_191_705 ();
 FILLCELL_X32 FILLER_191_737 ();
 FILLCELL_X32 FILLER_191_769 ();
 FILLCELL_X32 FILLER_191_801 ();
 FILLCELL_X32 FILLER_191_833 ();
 FILLCELL_X32 FILLER_191_865 ();
 FILLCELL_X32 FILLER_191_897 ();
 FILLCELL_X32 FILLER_191_929 ();
 FILLCELL_X32 FILLER_191_961 ();
 FILLCELL_X32 FILLER_191_993 ();
 FILLCELL_X32 FILLER_191_1025 ();
 FILLCELL_X32 FILLER_191_1057 ();
 FILLCELL_X32 FILLER_191_1089 ();
 FILLCELL_X32 FILLER_191_1121 ();
 FILLCELL_X32 FILLER_191_1153 ();
 FILLCELL_X32 FILLER_191_1185 ();
 FILLCELL_X32 FILLER_191_1217 ();
 FILLCELL_X8 FILLER_191_1249 ();
 FILLCELL_X4 FILLER_191_1257 ();
 FILLCELL_X2 FILLER_191_1261 ();
 FILLCELL_X32 FILLER_191_1264 ();
 FILLCELL_X32 FILLER_191_1296 ();
 FILLCELL_X32 FILLER_191_1328 ();
 FILLCELL_X32 FILLER_191_1360 ();
 FILLCELL_X32 FILLER_191_1392 ();
 FILLCELL_X32 FILLER_191_1424 ();
 FILLCELL_X32 FILLER_191_1456 ();
 FILLCELL_X32 FILLER_191_1488 ();
 FILLCELL_X32 FILLER_191_1520 ();
 FILLCELL_X32 FILLER_191_1552 ();
 FILLCELL_X32 FILLER_191_1584 ();
 FILLCELL_X32 FILLER_191_1616 ();
 FILLCELL_X32 FILLER_191_1648 ();
 FILLCELL_X32 FILLER_191_1680 ();
 FILLCELL_X32 FILLER_191_1712 ();
 FILLCELL_X32 FILLER_191_1744 ();
 FILLCELL_X32 FILLER_191_1776 ();
 FILLCELL_X32 FILLER_191_1808 ();
 FILLCELL_X32 FILLER_191_1840 ();
 FILLCELL_X32 FILLER_191_1872 ();
 FILLCELL_X32 FILLER_191_1904 ();
 FILLCELL_X32 FILLER_191_1936 ();
 FILLCELL_X32 FILLER_191_1968 ();
 FILLCELL_X32 FILLER_191_2000 ();
 FILLCELL_X32 FILLER_191_2032 ();
 FILLCELL_X32 FILLER_191_2064 ();
 FILLCELL_X32 FILLER_191_2096 ();
 FILLCELL_X32 FILLER_191_2128 ();
 FILLCELL_X32 FILLER_191_2160 ();
 FILLCELL_X32 FILLER_191_2192 ();
 FILLCELL_X32 FILLER_191_2224 ();
 FILLCELL_X32 FILLER_191_2256 ();
 FILLCELL_X32 FILLER_191_2288 ();
 FILLCELL_X32 FILLER_191_2320 ();
 FILLCELL_X32 FILLER_191_2352 ();
 FILLCELL_X32 FILLER_191_2384 ();
 FILLCELL_X32 FILLER_191_2416 ();
 FILLCELL_X32 FILLER_191_2448 ();
 FILLCELL_X32 FILLER_191_2480 ();
 FILLCELL_X8 FILLER_191_2512 ();
 FILLCELL_X4 FILLER_191_2520 ();
 FILLCELL_X2 FILLER_191_2524 ();
 FILLCELL_X32 FILLER_191_2527 ();
 FILLCELL_X32 FILLER_191_2559 ();
 FILLCELL_X32 FILLER_191_2591 ();
 FILLCELL_X32 FILLER_191_2623 ();
 FILLCELL_X32 FILLER_191_2655 ();
 FILLCELL_X32 FILLER_191_2687 ();
 FILLCELL_X32 FILLER_191_2719 ();
 FILLCELL_X32 FILLER_191_2751 ();
 FILLCELL_X32 FILLER_191_2783 ();
 FILLCELL_X32 FILLER_191_2815 ();
 FILLCELL_X32 FILLER_191_2847 ();
 FILLCELL_X32 FILLER_191_2879 ();
 FILLCELL_X32 FILLER_191_2911 ();
 FILLCELL_X32 FILLER_191_2943 ();
 FILLCELL_X32 FILLER_191_2975 ();
 FILLCELL_X32 FILLER_191_3007 ();
 FILLCELL_X32 FILLER_191_3039 ();
 FILLCELL_X32 FILLER_191_3071 ();
 FILLCELL_X32 FILLER_191_3103 ();
 FILLCELL_X32 FILLER_191_3135 ();
 FILLCELL_X32 FILLER_191_3167 ();
 FILLCELL_X32 FILLER_191_3199 ();
 FILLCELL_X32 FILLER_191_3231 ();
 FILLCELL_X32 FILLER_191_3263 ();
 FILLCELL_X32 FILLER_191_3295 ();
 FILLCELL_X32 FILLER_191_3327 ();
 FILLCELL_X32 FILLER_191_3359 ();
 FILLCELL_X32 FILLER_191_3391 ();
 FILLCELL_X32 FILLER_191_3423 ();
 FILLCELL_X32 FILLER_191_3455 ();
 FILLCELL_X32 FILLER_191_3487 ();
 FILLCELL_X32 FILLER_191_3519 ();
 FILLCELL_X32 FILLER_191_3551 ();
 FILLCELL_X32 FILLER_191_3583 ();
 FILLCELL_X32 FILLER_191_3615 ();
 FILLCELL_X32 FILLER_191_3647 ();
 FILLCELL_X32 FILLER_191_3679 ();
 FILLCELL_X16 FILLER_191_3711 ();
 FILLCELL_X8 FILLER_191_3727 ();
 FILLCELL_X2 FILLER_191_3735 ();
 FILLCELL_X1 FILLER_191_3737 ();
 FILLCELL_X32 FILLER_192_1 ();
 FILLCELL_X32 FILLER_192_33 ();
 FILLCELL_X32 FILLER_192_65 ();
 FILLCELL_X32 FILLER_192_97 ();
 FILLCELL_X32 FILLER_192_129 ();
 FILLCELL_X32 FILLER_192_161 ();
 FILLCELL_X32 FILLER_192_193 ();
 FILLCELL_X32 FILLER_192_225 ();
 FILLCELL_X32 FILLER_192_257 ();
 FILLCELL_X32 FILLER_192_289 ();
 FILLCELL_X32 FILLER_192_321 ();
 FILLCELL_X32 FILLER_192_353 ();
 FILLCELL_X32 FILLER_192_385 ();
 FILLCELL_X32 FILLER_192_417 ();
 FILLCELL_X32 FILLER_192_449 ();
 FILLCELL_X32 FILLER_192_481 ();
 FILLCELL_X32 FILLER_192_513 ();
 FILLCELL_X32 FILLER_192_545 ();
 FILLCELL_X32 FILLER_192_577 ();
 FILLCELL_X16 FILLER_192_609 ();
 FILLCELL_X4 FILLER_192_625 ();
 FILLCELL_X2 FILLER_192_629 ();
 FILLCELL_X32 FILLER_192_632 ();
 FILLCELL_X32 FILLER_192_664 ();
 FILLCELL_X32 FILLER_192_696 ();
 FILLCELL_X32 FILLER_192_728 ();
 FILLCELL_X32 FILLER_192_760 ();
 FILLCELL_X32 FILLER_192_792 ();
 FILLCELL_X32 FILLER_192_824 ();
 FILLCELL_X32 FILLER_192_856 ();
 FILLCELL_X32 FILLER_192_888 ();
 FILLCELL_X32 FILLER_192_920 ();
 FILLCELL_X32 FILLER_192_952 ();
 FILLCELL_X32 FILLER_192_984 ();
 FILLCELL_X32 FILLER_192_1016 ();
 FILLCELL_X32 FILLER_192_1048 ();
 FILLCELL_X32 FILLER_192_1080 ();
 FILLCELL_X32 FILLER_192_1112 ();
 FILLCELL_X32 FILLER_192_1144 ();
 FILLCELL_X32 FILLER_192_1176 ();
 FILLCELL_X32 FILLER_192_1208 ();
 FILLCELL_X32 FILLER_192_1240 ();
 FILLCELL_X32 FILLER_192_1272 ();
 FILLCELL_X32 FILLER_192_1304 ();
 FILLCELL_X32 FILLER_192_1336 ();
 FILLCELL_X32 FILLER_192_1368 ();
 FILLCELL_X32 FILLER_192_1400 ();
 FILLCELL_X32 FILLER_192_1432 ();
 FILLCELL_X32 FILLER_192_1464 ();
 FILLCELL_X32 FILLER_192_1496 ();
 FILLCELL_X32 FILLER_192_1528 ();
 FILLCELL_X32 FILLER_192_1560 ();
 FILLCELL_X32 FILLER_192_1592 ();
 FILLCELL_X32 FILLER_192_1624 ();
 FILLCELL_X32 FILLER_192_1656 ();
 FILLCELL_X32 FILLER_192_1688 ();
 FILLCELL_X32 FILLER_192_1720 ();
 FILLCELL_X32 FILLER_192_1752 ();
 FILLCELL_X32 FILLER_192_1784 ();
 FILLCELL_X32 FILLER_192_1816 ();
 FILLCELL_X32 FILLER_192_1848 ();
 FILLCELL_X8 FILLER_192_1880 ();
 FILLCELL_X4 FILLER_192_1888 ();
 FILLCELL_X2 FILLER_192_1892 ();
 FILLCELL_X32 FILLER_192_1895 ();
 FILLCELL_X32 FILLER_192_1927 ();
 FILLCELL_X32 FILLER_192_1959 ();
 FILLCELL_X32 FILLER_192_1991 ();
 FILLCELL_X32 FILLER_192_2023 ();
 FILLCELL_X32 FILLER_192_2055 ();
 FILLCELL_X32 FILLER_192_2087 ();
 FILLCELL_X32 FILLER_192_2119 ();
 FILLCELL_X32 FILLER_192_2151 ();
 FILLCELL_X32 FILLER_192_2183 ();
 FILLCELL_X32 FILLER_192_2215 ();
 FILLCELL_X32 FILLER_192_2247 ();
 FILLCELL_X32 FILLER_192_2279 ();
 FILLCELL_X32 FILLER_192_2311 ();
 FILLCELL_X32 FILLER_192_2343 ();
 FILLCELL_X32 FILLER_192_2375 ();
 FILLCELL_X32 FILLER_192_2407 ();
 FILLCELL_X32 FILLER_192_2439 ();
 FILLCELL_X32 FILLER_192_2471 ();
 FILLCELL_X32 FILLER_192_2503 ();
 FILLCELL_X32 FILLER_192_2535 ();
 FILLCELL_X32 FILLER_192_2567 ();
 FILLCELL_X32 FILLER_192_2599 ();
 FILLCELL_X32 FILLER_192_2631 ();
 FILLCELL_X32 FILLER_192_2663 ();
 FILLCELL_X32 FILLER_192_2695 ();
 FILLCELL_X32 FILLER_192_2727 ();
 FILLCELL_X32 FILLER_192_2759 ();
 FILLCELL_X32 FILLER_192_2791 ();
 FILLCELL_X32 FILLER_192_2823 ();
 FILLCELL_X32 FILLER_192_2855 ();
 FILLCELL_X32 FILLER_192_2887 ();
 FILLCELL_X32 FILLER_192_2919 ();
 FILLCELL_X32 FILLER_192_2951 ();
 FILLCELL_X32 FILLER_192_2983 ();
 FILLCELL_X32 FILLER_192_3015 ();
 FILLCELL_X32 FILLER_192_3047 ();
 FILLCELL_X32 FILLER_192_3079 ();
 FILLCELL_X32 FILLER_192_3111 ();
 FILLCELL_X8 FILLER_192_3143 ();
 FILLCELL_X4 FILLER_192_3151 ();
 FILLCELL_X2 FILLER_192_3155 ();
 FILLCELL_X32 FILLER_192_3158 ();
 FILLCELL_X32 FILLER_192_3190 ();
 FILLCELL_X32 FILLER_192_3222 ();
 FILLCELL_X32 FILLER_192_3254 ();
 FILLCELL_X32 FILLER_192_3286 ();
 FILLCELL_X32 FILLER_192_3318 ();
 FILLCELL_X32 FILLER_192_3350 ();
 FILLCELL_X32 FILLER_192_3382 ();
 FILLCELL_X32 FILLER_192_3414 ();
 FILLCELL_X32 FILLER_192_3446 ();
 FILLCELL_X32 FILLER_192_3478 ();
 FILLCELL_X32 FILLER_192_3510 ();
 FILLCELL_X32 FILLER_192_3542 ();
 FILLCELL_X32 FILLER_192_3574 ();
 FILLCELL_X32 FILLER_192_3606 ();
 FILLCELL_X32 FILLER_192_3638 ();
 FILLCELL_X32 FILLER_192_3670 ();
 FILLCELL_X32 FILLER_192_3702 ();
 FILLCELL_X4 FILLER_192_3734 ();
 FILLCELL_X32 FILLER_193_1 ();
 FILLCELL_X32 FILLER_193_33 ();
 FILLCELL_X32 FILLER_193_65 ();
 FILLCELL_X32 FILLER_193_97 ();
 FILLCELL_X32 FILLER_193_129 ();
 FILLCELL_X32 FILLER_193_161 ();
 FILLCELL_X32 FILLER_193_193 ();
 FILLCELL_X32 FILLER_193_225 ();
 FILLCELL_X32 FILLER_193_257 ();
 FILLCELL_X32 FILLER_193_289 ();
 FILLCELL_X32 FILLER_193_321 ();
 FILLCELL_X32 FILLER_193_353 ();
 FILLCELL_X32 FILLER_193_385 ();
 FILLCELL_X32 FILLER_193_417 ();
 FILLCELL_X32 FILLER_193_449 ();
 FILLCELL_X32 FILLER_193_481 ();
 FILLCELL_X32 FILLER_193_513 ();
 FILLCELL_X32 FILLER_193_545 ();
 FILLCELL_X32 FILLER_193_577 ();
 FILLCELL_X32 FILLER_193_609 ();
 FILLCELL_X32 FILLER_193_641 ();
 FILLCELL_X32 FILLER_193_673 ();
 FILLCELL_X32 FILLER_193_705 ();
 FILLCELL_X32 FILLER_193_737 ();
 FILLCELL_X32 FILLER_193_769 ();
 FILLCELL_X32 FILLER_193_801 ();
 FILLCELL_X32 FILLER_193_833 ();
 FILLCELL_X32 FILLER_193_865 ();
 FILLCELL_X32 FILLER_193_897 ();
 FILLCELL_X32 FILLER_193_929 ();
 FILLCELL_X32 FILLER_193_961 ();
 FILLCELL_X32 FILLER_193_993 ();
 FILLCELL_X32 FILLER_193_1025 ();
 FILLCELL_X32 FILLER_193_1057 ();
 FILLCELL_X32 FILLER_193_1089 ();
 FILLCELL_X32 FILLER_193_1121 ();
 FILLCELL_X32 FILLER_193_1153 ();
 FILLCELL_X32 FILLER_193_1185 ();
 FILLCELL_X32 FILLER_193_1217 ();
 FILLCELL_X8 FILLER_193_1249 ();
 FILLCELL_X4 FILLER_193_1257 ();
 FILLCELL_X2 FILLER_193_1261 ();
 FILLCELL_X32 FILLER_193_1264 ();
 FILLCELL_X32 FILLER_193_1296 ();
 FILLCELL_X32 FILLER_193_1328 ();
 FILLCELL_X32 FILLER_193_1360 ();
 FILLCELL_X32 FILLER_193_1392 ();
 FILLCELL_X32 FILLER_193_1424 ();
 FILLCELL_X32 FILLER_193_1456 ();
 FILLCELL_X32 FILLER_193_1488 ();
 FILLCELL_X32 FILLER_193_1520 ();
 FILLCELL_X32 FILLER_193_1552 ();
 FILLCELL_X32 FILLER_193_1584 ();
 FILLCELL_X32 FILLER_193_1616 ();
 FILLCELL_X32 FILLER_193_1648 ();
 FILLCELL_X32 FILLER_193_1680 ();
 FILLCELL_X32 FILLER_193_1712 ();
 FILLCELL_X32 FILLER_193_1744 ();
 FILLCELL_X32 FILLER_193_1776 ();
 FILLCELL_X32 FILLER_193_1808 ();
 FILLCELL_X32 FILLER_193_1840 ();
 FILLCELL_X32 FILLER_193_1872 ();
 FILLCELL_X32 FILLER_193_1904 ();
 FILLCELL_X32 FILLER_193_1936 ();
 FILLCELL_X32 FILLER_193_1968 ();
 FILLCELL_X32 FILLER_193_2000 ();
 FILLCELL_X32 FILLER_193_2032 ();
 FILLCELL_X32 FILLER_193_2064 ();
 FILLCELL_X32 FILLER_193_2096 ();
 FILLCELL_X32 FILLER_193_2128 ();
 FILLCELL_X32 FILLER_193_2160 ();
 FILLCELL_X32 FILLER_193_2192 ();
 FILLCELL_X32 FILLER_193_2224 ();
 FILLCELL_X32 FILLER_193_2256 ();
 FILLCELL_X32 FILLER_193_2288 ();
 FILLCELL_X32 FILLER_193_2320 ();
 FILLCELL_X32 FILLER_193_2352 ();
 FILLCELL_X32 FILLER_193_2384 ();
 FILLCELL_X32 FILLER_193_2416 ();
 FILLCELL_X32 FILLER_193_2448 ();
 FILLCELL_X32 FILLER_193_2480 ();
 FILLCELL_X8 FILLER_193_2512 ();
 FILLCELL_X4 FILLER_193_2520 ();
 FILLCELL_X2 FILLER_193_2524 ();
 FILLCELL_X32 FILLER_193_2527 ();
 FILLCELL_X32 FILLER_193_2559 ();
 FILLCELL_X32 FILLER_193_2591 ();
 FILLCELL_X32 FILLER_193_2623 ();
 FILLCELL_X32 FILLER_193_2655 ();
 FILLCELL_X32 FILLER_193_2687 ();
 FILLCELL_X32 FILLER_193_2719 ();
 FILLCELL_X32 FILLER_193_2751 ();
 FILLCELL_X32 FILLER_193_2783 ();
 FILLCELL_X32 FILLER_193_2815 ();
 FILLCELL_X32 FILLER_193_2847 ();
 FILLCELL_X32 FILLER_193_2879 ();
 FILLCELL_X32 FILLER_193_2911 ();
 FILLCELL_X32 FILLER_193_2943 ();
 FILLCELL_X32 FILLER_193_2975 ();
 FILLCELL_X32 FILLER_193_3007 ();
 FILLCELL_X32 FILLER_193_3039 ();
 FILLCELL_X32 FILLER_193_3071 ();
 FILLCELL_X32 FILLER_193_3103 ();
 FILLCELL_X32 FILLER_193_3135 ();
 FILLCELL_X32 FILLER_193_3167 ();
 FILLCELL_X32 FILLER_193_3199 ();
 FILLCELL_X32 FILLER_193_3231 ();
 FILLCELL_X32 FILLER_193_3263 ();
 FILLCELL_X32 FILLER_193_3295 ();
 FILLCELL_X32 FILLER_193_3327 ();
 FILLCELL_X32 FILLER_193_3359 ();
 FILLCELL_X32 FILLER_193_3391 ();
 FILLCELL_X32 FILLER_193_3423 ();
 FILLCELL_X32 FILLER_193_3455 ();
 FILLCELL_X32 FILLER_193_3487 ();
 FILLCELL_X32 FILLER_193_3519 ();
 FILLCELL_X32 FILLER_193_3551 ();
 FILLCELL_X32 FILLER_193_3583 ();
 FILLCELL_X32 FILLER_193_3615 ();
 FILLCELL_X32 FILLER_193_3647 ();
 FILLCELL_X32 FILLER_193_3679 ();
 FILLCELL_X16 FILLER_193_3711 ();
 FILLCELL_X8 FILLER_193_3727 ();
 FILLCELL_X2 FILLER_193_3735 ();
 FILLCELL_X1 FILLER_193_3737 ();
 FILLCELL_X32 FILLER_194_1 ();
 FILLCELL_X32 FILLER_194_33 ();
 FILLCELL_X32 FILLER_194_65 ();
 FILLCELL_X32 FILLER_194_97 ();
 FILLCELL_X32 FILLER_194_129 ();
 FILLCELL_X32 FILLER_194_161 ();
 FILLCELL_X32 FILLER_194_193 ();
 FILLCELL_X32 FILLER_194_225 ();
 FILLCELL_X32 FILLER_194_257 ();
 FILLCELL_X32 FILLER_194_289 ();
 FILLCELL_X32 FILLER_194_321 ();
 FILLCELL_X32 FILLER_194_353 ();
 FILLCELL_X32 FILLER_194_385 ();
 FILLCELL_X32 FILLER_194_417 ();
 FILLCELL_X32 FILLER_194_449 ();
 FILLCELL_X32 FILLER_194_481 ();
 FILLCELL_X32 FILLER_194_513 ();
 FILLCELL_X32 FILLER_194_545 ();
 FILLCELL_X32 FILLER_194_577 ();
 FILLCELL_X16 FILLER_194_609 ();
 FILLCELL_X4 FILLER_194_625 ();
 FILLCELL_X2 FILLER_194_629 ();
 FILLCELL_X32 FILLER_194_632 ();
 FILLCELL_X32 FILLER_194_664 ();
 FILLCELL_X32 FILLER_194_696 ();
 FILLCELL_X32 FILLER_194_728 ();
 FILLCELL_X32 FILLER_194_760 ();
 FILLCELL_X32 FILLER_194_792 ();
 FILLCELL_X32 FILLER_194_824 ();
 FILLCELL_X32 FILLER_194_856 ();
 FILLCELL_X32 FILLER_194_888 ();
 FILLCELL_X32 FILLER_194_920 ();
 FILLCELL_X32 FILLER_194_952 ();
 FILLCELL_X32 FILLER_194_984 ();
 FILLCELL_X32 FILLER_194_1016 ();
 FILLCELL_X32 FILLER_194_1048 ();
 FILLCELL_X32 FILLER_194_1080 ();
 FILLCELL_X32 FILLER_194_1112 ();
 FILLCELL_X32 FILLER_194_1144 ();
 FILLCELL_X32 FILLER_194_1176 ();
 FILLCELL_X32 FILLER_194_1208 ();
 FILLCELL_X32 FILLER_194_1240 ();
 FILLCELL_X32 FILLER_194_1272 ();
 FILLCELL_X32 FILLER_194_1304 ();
 FILLCELL_X32 FILLER_194_1336 ();
 FILLCELL_X32 FILLER_194_1368 ();
 FILLCELL_X32 FILLER_194_1400 ();
 FILLCELL_X32 FILLER_194_1432 ();
 FILLCELL_X32 FILLER_194_1464 ();
 FILLCELL_X32 FILLER_194_1496 ();
 FILLCELL_X32 FILLER_194_1528 ();
 FILLCELL_X32 FILLER_194_1560 ();
 FILLCELL_X32 FILLER_194_1592 ();
 FILLCELL_X32 FILLER_194_1624 ();
 FILLCELL_X32 FILLER_194_1656 ();
 FILLCELL_X32 FILLER_194_1688 ();
 FILLCELL_X32 FILLER_194_1720 ();
 FILLCELL_X32 FILLER_194_1752 ();
 FILLCELL_X32 FILLER_194_1784 ();
 FILLCELL_X32 FILLER_194_1816 ();
 FILLCELL_X32 FILLER_194_1848 ();
 FILLCELL_X8 FILLER_194_1880 ();
 FILLCELL_X4 FILLER_194_1888 ();
 FILLCELL_X2 FILLER_194_1892 ();
 FILLCELL_X32 FILLER_194_1895 ();
 FILLCELL_X32 FILLER_194_1927 ();
 FILLCELL_X32 FILLER_194_1959 ();
 FILLCELL_X32 FILLER_194_1991 ();
 FILLCELL_X32 FILLER_194_2023 ();
 FILLCELL_X32 FILLER_194_2055 ();
 FILLCELL_X32 FILLER_194_2087 ();
 FILLCELL_X32 FILLER_194_2119 ();
 FILLCELL_X32 FILLER_194_2151 ();
 FILLCELL_X32 FILLER_194_2183 ();
 FILLCELL_X32 FILLER_194_2215 ();
 FILLCELL_X32 FILLER_194_2247 ();
 FILLCELL_X32 FILLER_194_2279 ();
 FILLCELL_X32 FILLER_194_2311 ();
 FILLCELL_X32 FILLER_194_2343 ();
 FILLCELL_X32 FILLER_194_2375 ();
 FILLCELL_X32 FILLER_194_2407 ();
 FILLCELL_X32 FILLER_194_2439 ();
 FILLCELL_X32 FILLER_194_2471 ();
 FILLCELL_X32 FILLER_194_2503 ();
 FILLCELL_X32 FILLER_194_2535 ();
 FILLCELL_X32 FILLER_194_2567 ();
 FILLCELL_X32 FILLER_194_2599 ();
 FILLCELL_X32 FILLER_194_2631 ();
 FILLCELL_X32 FILLER_194_2663 ();
 FILLCELL_X32 FILLER_194_2695 ();
 FILLCELL_X32 FILLER_194_2727 ();
 FILLCELL_X32 FILLER_194_2759 ();
 FILLCELL_X32 FILLER_194_2791 ();
 FILLCELL_X32 FILLER_194_2823 ();
 FILLCELL_X32 FILLER_194_2855 ();
 FILLCELL_X32 FILLER_194_2887 ();
 FILLCELL_X32 FILLER_194_2919 ();
 FILLCELL_X32 FILLER_194_2951 ();
 FILLCELL_X32 FILLER_194_2983 ();
 FILLCELL_X32 FILLER_194_3015 ();
 FILLCELL_X32 FILLER_194_3047 ();
 FILLCELL_X32 FILLER_194_3079 ();
 FILLCELL_X32 FILLER_194_3111 ();
 FILLCELL_X8 FILLER_194_3143 ();
 FILLCELL_X4 FILLER_194_3151 ();
 FILLCELL_X2 FILLER_194_3155 ();
 FILLCELL_X32 FILLER_194_3158 ();
 FILLCELL_X32 FILLER_194_3190 ();
 FILLCELL_X32 FILLER_194_3222 ();
 FILLCELL_X32 FILLER_194_3254 ();
 FILLCELL_X32 FILLER_194_3286 ();
 FILLCELL_X32 FILLER_194_3318 ();
 FILLCELL_X32 FILLER_194_3350 ();
 FILLCELL_X32 FILLER_194_3382 ();
 FILLCELL_X32 FILLER_194_3414 ();
 FILLCELL_X32 FILLER_194_3446 ();
 FILLCELL_X32 FILLER_194_3478 ();
 FILLCELL_X32 FILLER_194_3510 ();
 FILLCELL_X32 FILLER_194_3542 ();
 FILLCELL_X32 FILLER_194_3574 ();
 FILLCELL_X32 FILLER_194_3606 ();
 FILLCELL_X32 FILLER_194_3638 ();
 FILLCELL_X32 FILLER_194_3670 ();
 FILLCELL_X32 FILLER_194_3702 ();
 FILLCELL_X4 FILLER_194_3734 ();
 FILLCELL_X32 FILLER_195_1 ();
 FILLCELL_X32 FILLER_195_33 ();
 FILLCELL_X32 FILLER_195_65 ();
 FILLCELL_X32 FILLER_195_97 ();
 FILLCELL_X32 FILLER_195_129 ();
 FILLCELL_X32 FILLER_195_161 ();
 FILLCELL_X32 FILLER_195_193 ();
 FILLCELL_X32 FILLER_195_225 ();
 FILLCELL_X32 FILLER_195_257 ();
 FILLCELL_X32 FILLER_195_289 ();
 FILLCELL_X32 FILLER_195_321 ();
 FILLCELL_X32 FILLER_195_353 ();
 FILLCELL_X32 FILLER_195_385 ();
 FILLCELL_X32 FILLER_195_417 ();
 FILLCELL_X32 FILLER_195_449 ();
 FILLCELL_X32 FILLER_195_481 ();
 FILLCELL_X32 FILLER_195_513 ();
 FILLCELL_X32 FILLER_195_545 ();
 FILLCELL_X32 FILLER_195_577 ();
 FILLCELL_X32 FILLER_195_609 ();
 FILLCELL_X32 FILLER_195_641 ();
 FILLCELL_X32 FILLER_195_673 ();
 FILLCELL_X32 FILLER_195_705 ();
 FILLCELL_X32 FILLER_195_737 ();
 FILLCELL_X32 FILLER_195_769 ();
 FILLCELL_X32 FILLER_195_801 ();
 FILLCELL_X32 FILLER_195_833 ();
 FILLCELL_X32 FILLER_195_865 ();
 FILLCELL_X32 FILLER_195_897 ();
 FILLCELL_X32 FILLER_195_929 ();
 FILLCELL_X32 FILLER_195_961 ();
 FILLCELL_X32 FILLER_195_993 ();
 FILLCELL_X32 FILLER_195_1025 ();
 FILLCELL_X32 FILLER_195_1057 ();
 FILLCELL_X32 FILLER_195_1089 ();
 FILLCELL_X32 FILLER_195_1121 ();
 FILLCELL_X32 FILLER_195_1153 ();
 FILLCELL_X32 FILLER_195_1185 ();
 FILLCELL_X32 FILLER_195_1217 ();
 FILLCELL_X8 FILLER_195_1249 ();
 FILLCELL_X4 FILLER_195_1257 ();
 FILLCELL_X2 FILLER_195_1261 ();
 FILLCELL_X32 FILLER_195_1264 ();
 FILLCELL_X32 FILLER_195_1296 ();
 FILLCELL_X32 FILLER_195_1328 ();
 FILLCELL_X32 FILLER_195_1360 ();
 FILLCELL_X32 FILLER_195_1392 ();
 FILLCELL_X32 FILLER_195_1424 ();
 FILLCELL_X32 FILLER_195_1456 ();
 FILLCELL_X32 FILLER_195_1488 ();
 FILLCELL_X32 FILLER_195_1520 ();
 FILLCELL_X32 FILLER_195_1552 ();
 FILLCELL_X32 FILLER_195_1584 ();
 FILLCELL_X32 FILLER_195_1616 ();
 FILLCELL_X32 FILLER_195_1648 ();
 FILLCELL_X32 FILLER_195_1680 ();
 FILLCELL_X32 FILLER_195_1712 ();
 FILLCELL_X32 FILLER_195_1744 ();
 FILLCELL_X32 FILLER_195_1776 ();
 FILLCELL_X32 FILLER_195_1808 ();
 FILLCELL_X32 FILLER_195_1840 ();
 FILLCELL_X32 FILLER_195_1872 ();
 FILLCELL_X32 FILLER_195_1904 ();
 FILLCELL_X32 FILLER_195_1936 ();
 FILLCELL_X32 FILLER_195_1968 ();
 FILLCELL_X32 FILLER_195_2000 ();
 FILLCELL_X32 FILLER_195_2032 ();
 FILLCELL_X32 FILLER_195_2064 ();
 FILLCELL_X32 FILLER_195_2096 ();
 FILLCELL_X32 FILLER_195_2128 ();
 FILLCELL_X32 FILLER_195_2160 ();
 FILLCELL_X32 FILLER_195_2192 ();
 FILLCELL_X32 FILLER_195_2224 ();
 FILLCELL_X32 FILLER_195_2256 ();
 FILLCELL_X32 FILLER_195_2288 ();
 FILLCELL_X32 FILLER_195_2320 ();
 FILLCELL_X32 FILLER_195_2352 ();
 FILLCELL_X32 FILLER_195_2384 ();
 FILLCELL_X32 FILLER_195_2416 ();
 FILLCELL_X32 FILLER_195_2448 ();
 FILLCELL_X32 FILLER_195_2480 ();
 FILLCELL_X8 FILLER_195_2512 ();
 FILLCELL_X4 FILLER_195_2520 ();
 FILLCELL_X2 FILLER_195_2524 ();
 FILLCELL_X32 FILLER_195_2527 ();
 FILLCELL_X32 FILLER_195_2559 ();
 FILLCELL_X32 FILLER_195_2591 ();
 FILLCELL_X32 FILLER_195_2623 ();
 FILLCELL_X32 FILLER_195_2655 ();
 FILLCELL_X32 FILLER_195_2687 ();
 FILLCELL_X32 FILLER_195_2719 ();
 FILLCELL_X32 FILLER_195_2751 ();
 FILLCELL_X32 FILLER_195_2783 ();
 FILLCELL_X32 FILLER_195_2815 ();
 FILLCELL_X32 FILLER_195_2847 ();
 FILLCELL_X32 FILLER_195_2879 ();
 FILLCELL_X32 FILLER_195_2911 ();
 FILLCELL_X32 FILLER_195_2943 ();
 FILLCELL_X32 FILLER_195_2975 ();
 FILLCELL_X32 FILLER_195_3007 ();
 FILLCELL_X32 FILLER_195_3039 ();
 FILLCELL_X32 FILLER_195_3071 ();
 FILLCELL_X32 FILLER_195_3103 ();
 FILLCELL_X32 FILLER_195_3135 ();
 FILLCELL_X32 FILLER_195_3167 ();
 FILLCELL_X32 FILLER_195_3199 ();
 FILLCELL_X32 FILLER_195_3231 ();
 FILLCELL_X32 FILLER_195_3263 ();
 FILLCELL_X32 FILLER_195_3295 ();
 FILLCELL_X32 FILLER_195_3327 ();
 FILLCELL_X32 FILLER_195_3359 ();
 FILLCELL_X32 FILLER_195_3391 ();
 FILLCELL_X32 FILLER_195_3423 ();
 FILLCELL_X32 FILLER_195_3455 ();
 FILLCELL_X32 FILLER_195_3487 ();
 FILLCELL_X32 FILLER_195_3519 ();
 FILLCELL_X32 FILLER_195_3551 ();
 FILLCELL_X32 FILLER_195_3583 ();
 FILLCELL_X32 FILLER_195_3615 ();
 FILLCELL_X32 FILLER_195_3647 ();
 FILLCELL_X32 FILLER_195_3679 ();
 FILLCELL_X16 FILLER_195_3711 ();
 FILLCELL_X8 FILLER_195_3727 ();
 FILLCELL_X2 FILLER_195_3735 ();
 FILLCELL_X1 FILLER_195_3737 ();
 FILLCELL_X32 FILLER_196_1 ();
 FILLCELL_X32 FILLER_196_33 ();
 FILLCELL_X32 FILLER_196_65 ();
 FILLCELL_X32 FILLER_196_97 ();
 FILLCELL_X32 FILLER_196_129 ();
 FILLCELL_X32 FILLER_196_161 ();
 FILLCELL_X32 FILLER_196_193 ();
 FILLCELL_X32 FILLER_196_225 ();
 FILLCELL_X32 FILLER_196_257 ();
 FILLCELL_X32 FILLER_196_289 ();
 FILLCELL_X32 FILLER_196_321 ();
 FILLCELL_X32 FILLER_196_353 ();
 FILLCELL_X32 FILLER_196_385 ();
 FILLCELL_X32 FILLER_196_417 ();
 FILLCELL_X32 FILLER_196_449 ();
 FILLCELL_X32 FILLER_196_481 ();
 FILLCELL_X32 FILLER_196_513 ();
 FILLCELL_X32 FILLER_196_545 ();
 FILLCELL_X32 FILLER_196_577 ();
 FILLCELL_X16 FILLER_196_609 ();
 FILLCELL_X4 FILLER_196_625 ();
 FILLCELL_X2 FILLER_196_629 ();
 FILLCELL_X32 FILLER_196_632 ();
 FILLCELL_X32 FILLER_196_664 ();
 FILLCELL_X32 FILLER_196_696 ();
 FILLCELL_X32 FILLER_196_728 ();
 FILLCELL_X32 FILLER_196_760 ();
 FILLCELL_X32 FILLER_196_792 ();
 FILLCELL_X32 FILLER_196_824 ();
 FILLCELL_X32 FILLER_196_856 ();
 FILLCELL_X32 FILLER_196_888 ();
 FILLCELL_X32 FILLER_196_920 ();
 FILLCELL_X32 FILLER_196_952 ();
 FILLCELL_X32 FILLER_196_984 ();
 FILLCELL_X32 FILLER_196_1016 ();
 FILLCELL_X32 FILLER_196_1048 ();
 FILLCELL_X32 FILLER_196_1080 ();
 FILLCELL_X32 FILLER_196_1112 ();
 FILLCELL_X32 FILLER_196_1144 ();
 FILLCELL_X32 FILLER_196_1176 ();
 FILLCELL_X32 FILLER_196_1208 ();
 FILLCELL_X32 FILLER_196_1240 ();
 FILLCELL_X32 FILLER_196_1272 ();
 FILLCELL_X32 FILLER_196_1304 ();
 FILLCELL_X32 FILLER_196_1336 ();
 FILLCELL_X32 FILLER_196_1368 ();
 FILLCELL_X32 FILLER_196_1400 ();
 FILLCELL_X32 FILLER_196_1432 ();
 FILLCELL_X32 FILLER_196_1464 ();
 FILLCELL_X32 FILLER_196_1496 ();
 FILLCELL_X32 FILLER_196_1528 ();
 FILLCELL_X32 FILLER_196_1560 ();
 FILLCELL_X32 FILLER_196_1592 ();
 FILLCELL_X32 FILLER_196_1624 ();
 FILLCELL_X32 FILLER_196_1656 ();
 FILLCELL_X32 FILLER_196_1688 ();
 FILLCELL_X32 FILLER_196_1720 ();
 FILLCELL_X32 FILLER_196_1752 ();
 FILLCELL_X32 FILLER_196_1784 ();
 FILLCELL_X32 FILLER_196_1816 ();
 FILLCELL_X32 FILLER_196_1848 ();
 FILLCELL_X8 FILLER_196_1880 ();
 FILLCELL_X4 FILLER_196_1888 ();
 FILLCELL_X2 FILLER_196_1892 ();
 FILLCELL_X32 FILLER_196_1895 ();
 FILLCELL_X32 FILLER_196_1927 ();
 FILLCELL_X32 FILLER_196_1959 ();
 FILLCELL_X32 FILLER_196_1991 ();
 FILLCELL_X32 FILLER_196_2023 ();
 FILLCELL_X32 FILLER_196_2055 ();
 FILLCELL_X32 FILLER_196_2087 ();
 FILLCELL_X32 FILLER_196_2119 ();
 FILLCELL_X32 FILLER_196_2151 ();
 FILLCELL_X32 FILLER_196_2183 ();
 FILLCELL_X32 FILLER_196_2215 ();
 FILLCELL_X32 FILLER_196_2247 ();
 FILLCELL_X32 FILLER_196_2279 ();
 FILLCELL_X32 FILLER_196_2311 ();
 FILLCELL_X32 FILLER_196_2343 ();
 FILLCELL_X32 FILLER_196_2375 ();
 FILLCELL_X32 FILLER_196_2407 ();
 FILLCELL_X32 FILLER_196_2439 ();
 FILLCELL_X32 FILLER_196_2471 ();
 FILLCELL_X32 FILLER_196_2503 ();
 FILLCELL_X32 FILLER_196_2535 ();
 FILLCELL_X32 FILLER_196_2567 ();
 FILLCELL_X32 FILLER_196_2599 ();
 FILLCELL_X32 FILLER_196_2631 ();
 FILLCELL_X32 FILLER_196_2663 ();
 FILLCELL_X32 FILLER_196_2695 ();
 FILLCELL_X32 FILLER_196_2727 ();
 FILLCELL_X32 FILLER_196_2759 ();
 FILLCELL_X32 FILLER_196_2791 ();
 FILLCELL_X32 FILLER_196_2823 ();
 FILLCELL_X32 FILLER_196_2855 ();
 FILLCELL_X32 FILLER_196_2887 ();
 FILLCELL_X32 FILLER_196_2919 ();
 FILLCELL_X32 FILLER_196_2951 ();
 FILLCELL_X32 FILLER_196_2983 ();
 FILLCELL_X32 FILLER_196_3015 ();
 FILLCELL_X32 FILLER_196_3047 ();
 FILLCELL_X32 FILLER_196_3079 ();
 FILLCELL_X32 FILLER_196_3111 ();
 FILLCELL_X8 FILLER_196_3143 ();
 FILLCELL_X4 FILLER_196_3151 ();
 FILLCELL_X2 FILLER_196_3155 ();
 FILLCELL_X32 FILLER_196_3158 ();
 FILLCELL_X32 FILLER_196_3190 ();
 FILLCELL_X32 FILLER_196_3222 ();
 FILLCELL_X32 FILLER_196_3254 ();
 FILLCELL_X32 FILLER_196_3286 ();
 FILLCELL_X32 FILLER_196_3318 ();
 FILLCELL_X32 FILLER_196_3350 ();
 FILLCELL_X32 FILLER_196_3382 ();
 FILLCELL_X32 FILLER_196_3414 ();
 FILLCELL_X32 FILLER_196_3446 ();
 FILLCELL_X32 FILLER_196_3478 ();
 FILLCELL_X32 FILLER_196_3510 ();
 FILLCELL_X32 FILLER_196_3542 ();
 FILLCELL_X32 FILLER_196_3574 ();
 FILLCELL_X32 FILLER_196_3606 ();
 FILLCELL_X32 FILLER_196_3638 ();
 FILLCELL_X32 FILLER_196_3670 ();
 FILLCELL_X32 FILLER_196_3702 ();
 FILLCELL_X4 FILLER_196_3734 ();
 FILLCELL_X32 FILLER_197_1 ();
 FILLCELL_X32 FILLER_197_33 ();
 FILLCELL_X32 FILLER_197_65 ();
 FILLCELL_X32 FILLER_197_97 ();
 FILLCELL_X32 FILLER_197_129 ();
 FILLCELL_X32 FILLER_197_161 ();
 FILLCELL_X32 FILLER_197_193 ();
 FILLCELL_X32 FILLER_197_225 ();
 FILLCELL_X32 FILLER_197_257 ();
 FILLCELL_X32 FILLER_197_289 ();
 FILLCELL_X32 FILLER_197_321 ();
 FILLCELL_X32 FILLER_197_353 ();
 FILLCELL_X32 FILLER_197_385 ();
 FILLCELL_X32 FILLER_197_417 ();
 FILLCELL_X32 FILLER_197_449 ();
 FILLCELL_X32 FILLER_197_481 ();
 FILLCELL_X32 FILLER_197_513 ();
 FILLCELL_X32 FILLER_197_545 ();
 FILLCELL_X32 FILLER_197_577 ();
 FILLCELL_X32 FILLER_197_609 ();
 FILLCELL_X32 FILLER_197_641 ();
 FILLCELL_X32 FILLER_197_673 ();
 FILLCELL_X32 FILLER_197_705 ();
 FILLCELL_X32 FILLER_197_737 ();
 FILLCELL_X32 FILLER_197_769 ();
 FILLCELL_X32 FILLER_197_801 ();
 FILLCELL_X32 FILLER_197_833 ();
 FILLCELL_X32 FILLER_197_865 ();
 FILLCELL_X32 FILLER_197_897 ();
 FILLCELL_X32 FILLER_197_929 ();
 FILLCELL_X32 FILLER_197_961 ();
 FILLCELL_X32 FILLER_197_993 ();
 FILLCELL_X32 FILLER_197_1025 ();
 FILLCELL_X32 FILLER_197_1057 ();
 FILLCELL_X32 FILLER_197_1089 ();
 FILLCELL_X32 FILLER_197_1121 ();
 FILLCELL_X32 FILLER_197_1153 ();
 FILLCELL_X32 FILLER_197_1185 ();
 FILLCELL_X32 FILLER_197_1217 ();
 FILLCELL_X8 FILLER_197_1249 ();
 FILLCELL_X4 FILLER_197_1257 ();
 FILLCELL_X2 FILLER_197_1261 ();
 FILLCELL_X32 FILLER_197_1264 ();
 FILLCELL_X32 FILLER_197_1296 ();
 FILLCELL_X32 FILLER_197_1328 ();
 FILLCELL_X32 FILLER_197_1360 ();
 FILLCELL_X32 FILLER_197_1392 ();
 FILLCELL_X32 FILLER_197_1424 ();
 FILLCELL_X32 FILLER_197_1456 ();
 FILLCELL_X32 FILLER_197_1488 ();
 FILLCELL_X32 FILLER_197_1520 ();
 FILLCELL_X32 FILLER_197_1552 ();
 FILLCELL_X32 FILLER_197_1584 ();
 FILLCELL_X32 FILLER_197_1616 ();
 FILLCELL_X32 FILLER_197_1648 ();
 FILLCELL_X32 FILLER_197_1680 ();
 FILLCELL_X32 FILLER_197_1712 ();
 FILLCELL_X32 FILLER_197_1744 ();
 FILLCELL_X32 FILLER_197_1776 ();
 FILLCELL_X32 FILLER_197_1808 ();
 FILLCELL_X32 FILLER_197_1840 ();
 FILLCELL_X32 FILLER_197_1872 ();
 FILLCELL_X32 FILLER_197_1904 ();
 FILLCELL_X32 FILLER_197_1936 ();
 FILLCELL_X32 FILLER_197_1968 ();
 FILLCELL_X32 FILLER_197_2000 ();
 FILLCELL_X32 FILLER_197_2032 ();
 FILLCELL_X32 FILLER_197_2064 ();
 FILLCELL_X32 FILLER_197_2096 ();
 FILLCELL_X32 FILLER_197_2128 ();
 FILLCELL_X32 FILLER_197_2160 ();
 FILLCELL_X32 FILLER_197_2192 ();
 FILLCELL_X32 FILLER_197_2224 ();
 FILLCELL_X32 FILLER_197_2256 ();
 FILLCELL_X32 FILLER_197_2288 ();
 FILLCELL_X32 FILLER_197_2320 ();
 FILLCELL_X32 FILLER_197_2352 ();
 FILLCELL_X32 FILLER_197_2384 ();
 FILLCELL_X32 FILLER_197_2416 ();
 FILLCELL_X32 FILLER_197_2448 ();
 FILLCELL_X32 FILLER_197_2480 ();
 FILLCELL_X8 FILLER_197_2512 ();
 FILLCELL_X4 FILLER_197_2520 ();
 FILLCELL_X2 FILLER_197_2524 ();
 FILLCELL_X32 FILLER_197_2527 ();
 FILLCELL_X32 FILLER_197_2559 ();
 FILLCELL_X32 FILLER_197_2591 ();
 FILLCELL_X32 FILLER_197_2623 ();
 FILLCELL_X32 FILLER_197_2655 ();
 FILLCELL_X32 FILLER_197_2687 ();
 FILLCELL_X32 FILLER_197_2719 ();
 FILLCELL_X32 FILLER_197_2751 ();
 FILLCELL_X32 FILLER_197_2783 ();
 FILLCELL_X32 FILLER_197_2815 ();
 FILLCELL_X32 FILLER_197_2847 ();
 FILLCELL_X32 FILLER_197_2879 ();
 FILLCELL_X32 FILLER_197_2911 ();
 FILLCELL_X32 FILLER_197_2943 ();
 FILLCELL_X32 FILLER_197_2975 ();
 FILLCELL_X32 FILLER_197_3007 ();
 FILLCELL_X32 FILLER_197_3039 ();
 FILLCELL_X32 FILLER_197_3071 ();
 FILLCELL_X32 FILLER_197_3103 ();
 FILLCELL_X32 FILLER_197_3135 ();
 FILLCELL_X32 FILLER_197_3167 ();
 FILLCELL_X32 FILLER_197_3199 ();
 FILLCELL_X32 FILLER_197_3231 ();
 FILLCELL_X32 FILLER_197_3263 ();
 FILLCELL_X32 FILLER_197_3295 ();
 FILLCELL_X32 FILLER_197_3327 ();
 FILLCELL_X32 FILLER_197_3359 ();
 FILLCELL_X32 FILLER_197_3391 ();
 FILLCELL_X32 FILLER_197_3423 ();
 FILLCELL_X32 FILLER_197_3455 ();
 FILLCELL_X32 FILLER_197_3487 ();
 FILLCELL_X32 FILLER_197_3519 ();
 FILLCELL_X32 FILLER_197_3551 ();
 FILLCELL_X32 FILLER_197_3583 ();
 FILLCELL_X32 FILLER_197_3615 ();
 FILLCELL_X32 FILLER_197_3647 ();
 FILLCELL_X32 FILLER_197_3679 ();
 FILLCELL_X16 FILLER_197_3711 ();
 FILLCELL_X8 FILLER_197_3727 ();
 FILLCELL_X2 FILLER_197_3735 ();
 FILLCELL_X1 FILLER_197_3737 ();
 FILLCELL_X32 FILLER_198_1 ();
 FILLCELL_X32 FILLER_198_33 ();
 FILLCELL_X32 FILLER_198_65 ();
 FILLCELL_X32 FILLER_198_97 ();
 FILLCELL_X32 FILLER_198_129 ();
 FILLCELL_X32 FILLER_198_161 ();
 FILLCELL_X32 FILLER_198_193 ();
 FILLCELL_X32 FILLER_198_225 ();
 FILLCELL_X32 FILLER_198_257 ();
 FILLCELL_X32 FILLER_198_289 ();
 FILLCELL_X32 FILLER_198_321 ();
 FILLCELL_X32 FILLER_198_353 ();
 FILLCELL_X32 FILLER_198_385 ();
 FILLCELL_X32 FILLER_198_417 ();
 FILLCELL_X32 FILLER_198_449 ();
 FILLCELL_X32 FILLER_198_481 ();
 FILLCELL_X32 FILLER_198_513 ();
 FILLCELL_X32 FILLER_198_545 ();
 FILLCELL_X32 FILLER_198_577 ();
 FILLCELL_X16 FILLER_198_609 ();
 FILLCELL_X4 FILLER_198_625 ();
 FILLCELL_X2 FILLER_198_629 ();
 FILLCELL_X32 FILLER_198_632 ();
 FILLCELL_X32 FILLER_198_664 ();
 FILLCELL_X32 FILLER_198_696 ();
 FILLCELL_X32 FILLER_198_728 ();
 FILLCELL_X32 FILLER_198_760 ();
 FILLCELL_X32 FILLER_198_792 ();
 FILLCELL_X32 FILLER_198_824 ();
 FILLCELL_X32 FILLER_198_856 ();
 FILLCELL_X32 FILLER_198_888 ();
 FILLCELL_X32 FILLER_198_920 ();
 FILLCELL_X32 FILLER_198_952 ();
 FILLCELL_X32 FILLER_198_984 ();
 FILLCELL_X32 FILLER_198_1016 ();
 FILLCELL_X32 FILLER_198_1048 ();
 FILLCELL_X32 FILLER_198_1080 ();
 FILLCELL_X32 FILLER_198_1112 ();
 FILLCELL_X32 FILLER_198_1144 ();
 FILLCELL_X32 FILLER_198_1176 ();
 FILLCELL_X32 FILLER_198_1208 ();
 FILLCELL_X32 FILLER_198_1240 ();
 FILLCELL_X32 FILLER_198_1272 ();
 FILLCELL_X32 FILLER_198_1304 ();
 FILLCELL_X32 FILLER_198_1336 ();
 FILLCELL_X32 FILLER_198_1368 ();
 FILLCELL_X32 FILLER_198_1400 ();
 FILLCELL_X32 FILLER_198_1432 ();
 FILLCELL_X32 FILLER_198_1464 ();
 FILLCELL_X32 FILLER_198_1496 ();
 FILLCELL_X32 FILLER_198_1528 ();
 FILLCELL_X32 FILLER_198_1560 ();
 FILLCELL_X32 FILLER_198_1592 ();
 FILLCELL_X32 FILLER_198_1624 ();
 FILLCELL_X32 FILLER_198_1656 ();
 FILLCELL_X32 FILLER_198_1688 ();
 FILLCELL_X32 FILLER_198_1720 ();
 FILLCELL_X32 FILLER_198_1752 ();
 FILLCELL_X32 FILLER_198_1784 ();
 FILLCELL_X32 FILLER_198_1816 ();
 FILLCELL_X32 FILLER_198_1848 ();
 FILLCELL_X8 FILLER_198_1880 ();
 FILLCELL_X4 FILLER_198_1888 ();
 FILLCELL_X2 FILLER_198_1892 ();
 FILLCELL_X32 FILLER_198_1895 ();
 FILLCELL_X32 FILLER_198_1927 ();
 FILLCELL_X32 FILLER_198_1959 ();
 FILLCELL_X32 FILLER_198_1991 ();
 FILLCELL_X32 FILLER_198_2023 ();
 FILLCELL_X32 FILLER_198_2055 ();
 FILLCELL_X32 FILLER_198_2087 ();
 FILLCELL_X32 FILLER_198_2119 ();
 FILLCELL_X32 FILLER_198_2151 ();
 FILLCELL_X32 FILLER_198_2183 ();
 FILLCELL_X32 FILLER_198_2215 ();
 FILLCELL_X32 FILLER_198_2247 ();
 FILLCELL_X32 FILLER_198_2279 ();
 FILLCELL_X32 FILLER_198_2311 ();
 FILLCELL_X32 FILLER_198_2343 ();
 FILLCELL_X32 FILLER_198_2375 ();
 FILLCELL_X32 FILLER_198_2407 ();
 FILLCELL_X32 FILLER_198_2439 ();
 FILLCELL_X32 FILLER_198_2471 ();
 FILLCELL_X32 FILLER_198_2503 ();
 FILLCELL_X32 FILLER_198_2535 ();
 FILLCELL_X32 FILLER_198_2567 ();
 FILLCELL_X32 FILLER_198_2599 ();
 FILLCELL_X32 FILLER_198_2631 ();
 FILLCELL_X32 FILLER_198_2663 ();
 FILLCELL_X32 FILLER_198_2695 ();
 FILLCELL_X32 FILLER_198_2727 ();
 FILLCELL_X32 FILLER_198_2759 ();
 FILLCELL_X32 FILLER_198_2791 ();
 FILLCELL_X32 FILLER_198_2823 ();
 FILLCELL_X32 FILLER_198_2855 ();
 FILLCELL_X32 FILLER_198_2887 ();
 FILLCELL_X32 FILLER_198_2919 ();
 FILLCELL_X32 FILLER_198_2951 ();
 FILLCELL_X32 FILLER_198_2983 ();
 FILLCELL_X32 FILLER_198_3015 ();
 FILLCELL_X32 FILLER_198_3047 ();
 FILLCELL_X32 FILLER_198_3079 ();
 FILLCELL_X32 FILLER_198_3111 ();
 FILLCELL_X8 FILLER_198_3143 ();
 FILLCELL_X4 FILLER_198_3151 ();
 FILLCELL_X2 FILLER_198_3155 ();
 FILLCELL_X32 FILLER_198_3158 ();
 FILLCELL_X32 FILLER_198_3190 ();
 FILLCELL_X32 FILLER_198_3222 ();
 FILLCELL_X32 FILLER_198_3254 ();
 FILLCELL_X32 FILLER_198_3286 ();
 FILLCELL_X32 FILLER_198_3318 ();
 FILLCELL_X32 FILLER_198_3350 ();
 FILLCELL_X32 FILLER_198_3382 ();
 FILLCELL_X32 FILLER_198_3414 ();
 FILLCELL_X32 FILLER_198_3446 ();
 FILLCELL_X32 FILLER_198_3478 ();
 FILLCELL_X32 FILLER_198_3510 ();
 FILLCELL_X32 FILLER_198_3542 ();
 FILLCELL_X32 FILLER_198_3574 ();
 FILLCELL_X32 FILLER_198_3606 ();
 FILLCELL_X32 FILLER_198_3638 ();
 FILLCELL_X32 FILLER_198_3670 ();
 FILLCELL_X32 FILLER_198_3702 ();
 FILLCELL_X4 FILLER_198_3734 ();
 FILLCELL_X32 FILLER_199_1 ();
 FILLCELL_X32 FILLER_199_33 ();
 FILLCELL_X32 FILLER_199_65 ();
 FILLCELL_X32 FILLER_199_97 ();
 FILLCELL_X32 FILLER_199_129 ();
 FILLCELL_X32 FILLER_199_161 ();
 FILLCELL_X32 FILLER_199_193 ();
 FILLCELL_X32 FILLER_199_225 ();
 FILLCELL_X32 FILLER_199_257 ();
 FILLCELL_X32 FILLER_199_289 ();
 FILLCELL_X32 FILLER_199_321 ();
 FILLCELL_X32 FILLER_199_353 ();
 FILLCELL_X32 FILLER_199_385 ();
 FILLCELL_X32 FILLER_199_417 ();
 FILLCELL_X32 FILLER_199_449 ();
 FILLCELL_X32 FILLER_199_481 ();
 FILLCELL_X32 FILLER_199_513 ();
 FILLCELL_X32 FILLER_199_545 ();
 FILLCELL_X32 FILLER_199_577 ();
 FILLCELL_X32 FILLER_199_609 ();
 FILLCELL_X32 FILLER_199_641 ();
 FILLCELL_X32 FILLER_199_673 ();
 FILLCELL_X32 FILLER_199_705 ();
 FILLCELL_X32 FILLER_199_737 ();
 FILLCELL_X32 FILLER_199_769 ();
 FILLCELL_X32 FILLER_199_801 ();
 FILLCELL_X32 FILLER_199_833 ();
 FILLCELL_X32 FILLER_199_865 ();
 FILLCELL_X32 FILLER_199_897 ();
 FILLCELL_X32 FILLER_199_929 ();
 FILLCELL_X32 FILLER_199_961 ();
 FILLCELL_X32 FILLER_199_993 ();
 FILLCELL_X32 FILLER_199_1025 ();
 FILLCELL_X32 FILLER_199_1057 ();
 FILLCELL_X32 FILLER_199_1089 ();
 FILLCELL_X32 FILLER_199_1121 ();
 FILLCELL_X32 FILLER_199_1153 ();
 FILLCELL_X32 FILLER_199_1185 ();
 FILLCELL_X32 FILLER_199_1217 ();
 FILLCELL_X8 FILLER_199_1249 ();
 FILLCELL_X4 FILLER_199_1257 ();
 FILLCELL_X2 FILLER_199_1261 ();
 FILLCELL_X32 FILLER_199_1264 ();
 FILLCELL_X32 FILLER_199_1296 ();
 FILLCELL_X32 FILLER_199_1328 ();
 FILLCELL_X32 FILLER_199_1360 ();
 FILLCELL_X32 FILLER_199_1392 ();
 FILLCELL_X32 FILLER_199_1424 ();
 FILLCELL_X32 FILLER_199_1456 ();
 FILLCELL_X32 FILLER_199_1488 ();
 FILLCELL_X32 FILLER_199_1520 ();
 FILLCELL_X32 FILLER_199_1552 ();
 FILLCELL_X32 FILLER_199_1584 ();
 FILLCELL_X32 FILLER_199_1616 ();
 FILLCELL_X32 FILLER_199_1648 ();
 FILLCELL_X32 FILLER_199_1680 ();
 FILLCELL_X32 FILLER_199_1712 ();
 FILLCELL_X32 FILLER_199_1744 ();
 FILLCELL_X32 FILLER_199_1776 ();
 FILLCELL_X32 FILLER_199_1808 ();
 FILLCELL_X32 FILLER_199_1840 ();
 FILLCELL_X32 FILLER_199_1872 ();
 FILLCELL_X32 FILLER_199_1904 ();
 FILLCELL_X32 FILLER_199_1936 ();
 FILLCELL_X32 FILLER_199_1968 ();
 FILLCELL_X32 FILLER_199_2000 ();
 FILLCELL_X32 FILLER_199_2032 ();
 FILLCELL_X32 FILLER_199_2064 ();
 FILLCELL_X32 FILLER_199_2096 ();
 FILLCELL_X32 FILLER_199_2128 ();
 FILLCELL_X32 FILLER_199_2160 ();
 FILLCELL_X32 FILLER_199_2192 ();
 FILLCELL_X32 FILLER_199_2224 ();
 FILLCELL_X32 FILLER_199_2256 ();
 FILLCELL_X32 FILLER_199_2288 ();
 FILLCELL_X32 FILLER_199_2320 ();
 FILLCELL_X32 FILLER_199_2352 ();
 FILLCELL_X32 FILLER_199_2384 ();
 FILLCELL_X32 FILLER_199_2416 ();
 FILLCELL_X32 FILLER_199_2448 ();
 FILLCELL_X32 FILLER_199_2480 ();
 FILLCELL_X8 FILLER_199_2512 ();
 FILLCELL_X4 FILLER_199_2520 ();
 FILLCELL_X2 FILLER_199_2524 ();
 FILLCELL_X32 FILLER_199_2527 ();
 FILLCELL_X32 FILLER_199_2559 ();
 FILLCELL_X32 FILLER_199_2591 ();
 FILLCELL_X32 FILLER_199_2623 ();
 FILLCELL_X32 FILLER_199_2655 ();
 FILLCELL_X32 FILLER_199_2687 ();
 FILLCELL_X32 FILLER_199_2719 ();
 FILLCELL_X32 FILLER_199_2751 ();
 FILLCELL_X32 FILLER_199_2783 ();
 FILLCELL_X32 FILLER_199_2815 ();
 FILLCELL_X32 FILLER_199_2847 ();
 FILLCELL_X32 FILLER_199_2879 ();
 FILLCELL_X32 FILLER_199_2911 ();
 FILLCELL_X32 FILLER_199_2943 ();
 FILLCELL_X32 FILLER_199_2975 ();
 FILLCELL_X32 FILLER_199_3007 ();
 FILLCELL_X32 FILLER_199_3039 ();
 FILLCELL_X32 FILLER_199_3071 ();
 FILLCELL_X32 FILLER_199_3103 ();
 FILLCELL_X32 FILLER_199_3135 ();
 FILLCELL_X32 FILLER_199_3167 ();
 FILLCELL_X32 FILLER_199_3199 ();
 FILLCELL_X32 FILLER_199_3231 ();
 FILLCELL_X32 FILLER_199_3263 ();
 FILLCELL_X32 FILLER_199_3295 ();
 FILLCELL_X32 FILLER_199_3327 ();
 FILLCELL_X32 FILLER_199_3359 ();
 FILLCELL_X32 FILLER_199_3391 ();
 FILLCELL_X32 FILLER_199_3423 ();
 FILLCELL_X32 FILLER_199_3455 ();
 FILLCELL_X32 FILLER_199_3487 ();
 FILLCELL_X32 FILLER_199_3519 ();
 FILLCELL_X32 FILLER_199_3551 ();
 FILLCELL_X32 FILLER_199_3583 ();
 FILLCELL_X32 FILLER_199_3615 ();
 FILLCELL_X32 FILLER_199_3647 ();
 FILLCELL_X32 FILLER_199_3679 ();
 FILLCELL_X16 FILLER_199_3711 ();
 FILLCELL_X8 FILLER_199_3727 ();
 FILLCELL_X2 FILLER_199_3735 ();
 FILLCELL_X1 FILLER_199_3737 ();
 FILLCELL_X32 FILLER_200_1 ();
 FILLCELL_X32 FILLER_200_33 ();
 FILLCELL_X32 FILLER_200_65 ();
 FILLCELL_X32 FILLER_200_97 ();
 FILLCELL_X32 FILLER_200_129 ();
 FILLCELL_X32 FILLER_200_161 ();
 FILLCELL_X32 FILLER_200_193 ();
 FILLCELL_X32 FILLER_200_225 ();
 FILLCELL_X32 FILLER_200_257 ();
 FILLCELL_X32 FILLER_200_289 ();
 FILLCELL_X32 FILLER_200_321 ();
 FILLCELL_X32 FILLER_200_353 ();
 FILLCELL_X32 FILLER_200_385 ();
 FILLCELL_X32 FILLER_200_417 ();
 FILLCELL_X32 FILLER_200_449 ();
 FILLCELL_X32 FILLER_200_481 ();
 FILLCELL_X32 FILLER_200_513 ();
 FILLCELL_X32 FILLER_200_545 ();
 FILLCELL_X32 FILLER_200_577 ();
 FILLCELL_X16 FILLER_200_609 ();
 FILLCELL_X4 FILLER_200_625 ();
 FILLCELL_X2 FILLER_200_629 ();
 FILLCELL_X32 FILLER_200_632 ();
 FILLCELL_X32 FILLER_200_664 ();
 FILLCELL_X32 FILLER_200_696 ();
 FILLCELL_X32 FILLER_200_728 ();
 FILLCELL_X32 FILLER_200_760 ();
 FILLCELL_X32 FILLER_200_792 ();
 FILLCELL_X32 FILLER_200_824 ();
 FILLCELL_X32 FILLER_200_856 ();
 FILLCELL_X32 FILLER_200_888 ();
 FILLCELL_X32 FILLER_200_920 ();
 FILLCELL_X32 FILLER_200_952 ();
 FILLCELL_X32 FILLER_200_984 ();
 FILLCELL_X32 FILLER_200_1016 ();
 FILLCELL_X32 FILLER_200_1048 ();
 FILLCELL_X32 FILLER_200_1080 ();
 FILLCELL_X32 FILLER_200_1112 ();
 FILLCELL_X32 FILLER_200_1144 ();
 FILLCELL_X32 FILLER_200_1176 ();
 FILLCELL_X32 FILLER_200_1208 ();
 FILLCELL_X32 FILLER_200_1240 ();
 FILLCELL_X32 FILLER_200_1272 ();
 FILLCELL_X32 FILLER_200_1304 ();
 FILLCELL_X32 FILLER_200_1336 ();
 FILLCELL_X32 FILLER_200_1368 ();
 FILLCELL_X32 FILLER_200_1400 ();
 FILLCELL_X32 FILLER_200_1432 ();
 FILLCELL_X32 FILLER_200_1464 ();
 FILLCELL_X32 FILLER_200_1496 ();
 FILLCELL_X32 FILLER_200_1528 ();
 FILLCELL_X32 FILLER_200_1560 ();
 FILLCELL_X32 FILLER_200_1592 ();
 FILLCELL_X32 FILLER_200_1624 ();
 FILLCELL_X32 FILLER_200_1656 ();
 FILLCELL_X32 FILLER_200_1688 ();
 FILLCELL_X32 FILLER_200_1720 ();
 FILLCELL_X32 FILLER_200_1752 ();
 FILLCELL_X32 FILLER_200_1784 ();
 FILLCELL_X32 FILLER_200_1816 ();
 FILLCELL_X32 FILLER_200_1848 ();
 FILLCELL_X8 FILLER_200_1880 ();
 FILLCELL_X4 FILLER_200_1888 ();
 FILLCELL_X2 FILLER_200_1892 ();
 FILLCELL_X32 FILLER_200_1895 ();
 FILLCELL_X32 FILLER_200_1927 ();
 FILLCELL_X32 FILLER_200_1959 ();
 FILLCELL_X32 FILLER_200_1991 ();
 FILLCELL_X32 FILLER_200_2023 ();
 FILLCELL_X32 FILLER_200_2055 ();
 FILLCELL_X32 FILLER_200_2087 ();
 FILLCELL_X32 FILLER_200_2119 ();
 FILLCELL_X32 FILLER_200_2151 ();
 FILLCELL_X32 FILLER_200_2183 ();
 FILLCELL_X32 FILLER_200_2215 ();
 FILLCELL_X32 FILLER_200_2247 ();
 FILLCELL_X32 FILLER_200_2279 ();
 FILLCELL_X32 FILLER_200_2311 ();
 FILLCELL_X32 FILLER_200_2343 ();
 FILLCELL_X32 FILLER_200_2375 ();
 FILLCELL_X32 FILLER_200_2407 ();
 FILLCELL_X32 FILLER_200_2439 ();
 FILLCELL_X32 FILLER_200_2471 ();
 FILLCELL_X32 FILLER_200_2503 ();
 FILLCELL_X32 FILLER_200_2535 ();
 FILLCELL_X32 FILLER_200_2567 ();
 FILLCELL_X32 FILLER_200_2599 ();
 FILLCELL_X32 FILLER_200_2631 ();
 FILLCELL_X32 FILLER_200_2663 ();
 FILLCELL_X32 FILLER_200_2695 ();
 FILLCELL_X32 FILLER_200_2727 ();
 FILLCELL_X32 FILLER_200_2759 ();
 FILLCELL_X32 FILLER_200_2791 ();
 FILLCELL_X32 FILLER_200_2823 ();
 FILLCELL_X32 FILLER_200_2855 ();
 FILLCELL_X32 FILLER_200_2887 ();
 FILLCELL_X32 FILLER_200_2919 ();
 FILLCELL_X32 FILLER_200_2951 ();
 FILLCELL_X32 FILLER_200_2983 ();
 FILLCELL_X32 FILLER_200_3015 ();
 FILLCELL_X32 FILLER_200_3047 ();
 FILLCELL_X32 FILLER_200_3079 ();
 FILLCELL_X32 FILLER_200_3111 ();
 FILLCELL_X8 FILLER_200_3143 ();
 FILLCELL_X4 FILLER_200_3151 ();
 FILLCELL_X2 FILLER_200_3155 ();
 FILLCELL_X32 FILLER_200_3158 ();
 FILLCELL_X32 FILLER_200_3190 ();
 FILLCELL_X32 FILLER_200_3222 ();
 FILLCELL_X32 FILLER_200_3254 ();
 FILLCELL_X32 FILLER_200_3286 ();
 FILLCELL_X32 FILLER_200_3318 ();
 FILLCELL_X32 FILLER_200_3350 ();
 FILLCELL_X32 FILLER_200_3382 ();
 FILLCELL_X32 FILLER_200_3414 ();
 FILLCELL_X32 FILLER_200_3446 ();
 FILLCELL_X32 FILLER_200_3478 ();
 FILLCELL_X32 FILLER_200_3510 ();
 FILLCELL_X32 FILLER_200_3542 ();
 FILLCELL_X32 FILLER_200_3574 ();
 FILLCELL_X32 FILLER_200_3606 ();
 FILLCELL_X32 FILLER_200_3638 ();
 FILLCELL_X32 FILLER_200_3670 ();
 FILLCELL_X32 FILLER_200_3702 ();
 FILLCELL_X4 FILLER_200_3734 ();
 FILLCELL_X32 FILLER_201_1 ();
 FILLCELL_X32 FILLER_201_33 ();
 FILLCELL_X32 FILLER_201_65 ();
 FILLCELL_X32 FILLER_201_97 ();
 FILLCELL_X32 FILLER_201_129 ();
 FILLCELL_X32 FILLER_201_161 ();
 FILLCELL_X32 FILLER_201_193 ();
 FILLCELL_X32 FILLER_201_225 ();
 FILLCELL_X32 FILLER_201_257 ();
 FILLCELL_X32 FILLER_201_289 ();
 FILLCELL_X32 FILLER_201_321 ();
 FILLCELL_X32 FILLER_201_353 ();
 FILLCELL_X32 FILLER_201_385 ();
 FILLCELL_X32 FILLER_201_417 ();
 FILLCELL_X32 FILLER_201_449 ();
 FILLCELL_X32 FILLER_201_481 ();
 FILLCELL_X32 FILLER_201_513 ();
 FILLCELL_X32 FILLER_201_545 ();
 FILLCELL_X32 FILLER_201_577 ();
 FILLCELL_X32 FILLER_201_609 ();
 FILLCELL_X32 FILLER_201_641 ();
 FILLCELL_X32 FILLER_201_673 ();
 FILLCELL_X32 FILLER_201_705 ();
 FILLCELL_X32 FILLER_201_737 ();
 FILLCELL_X32 FILLER_201_769 ();
 FILLCELL_X32 FILLER_201_801 ();
 FILLCELL_X32 FILLER_201_833 ();
 FILLCELL_X32 FILLER_201_865 ();
 FILLCELL_X32 FILLER_201_897 ();
 FILLCELL_X32 FILLER_201_929 ();
 FILLCELL_X32 FILLER_201_961 ();
 FILLCELL_X32 FILLER_201_993 ();
 FILLCELL_X32 FILLER_201_1025 ();
 FILLCELL_X32 FILLER_201_1057 ();
 FILLCELL_X32 FILLER_201_1089 ();
 FILLCELL_X32 FILLER_201_1121 ();
 FILLCELL_X32 FILLER_201_1153 ();
 FILLCELL_X32 FILLER_201_1185 ();
 FILLCELL_X32 FILLER_201_1217 ();
 FILLCELL_X8 FILLER_201_1249 ();
 FILLCELL_X4 FILLER_201_1257 ();
 FILLCELL_X2 FILLER_201_1261 ();
 FILLCELL_X32 FILLER_201_1264 ();
 FILLCELL_X32 FILLER_201_1296 ();
 FILLCELL_X32 FILLER_201_1328 ();
 FILLCELL_X32 FILLER_201_1360 ();
 FILLCELL_X32 FILLER_201_1392 ();
 FILLCELL_X32 FILLER_201_1424 ();
 FILLCELL_X32 FILLER_201_1456 ();
 FILLCELL_X32 FILLER_201_1488 ();
 FILLCELL_X32 FILLER_201_1520 ();
 FILLCELL_X32 FILLER_201_1552 ();
 FILLCELL_X32 FILLER_201_1584 ();
 FILLCELL_X32 FILLER_201_1616 ();
 FILLCELL_X32 FILLER_201_1648 ();
 FILLCELL_X32 FILLER_201_1680 ();
 FILLCELL_X32 FILLER_201_1712 ();
 FILLCELL_X32 FILLER_201_1744 ();
 FILLCELL_X32 FILLER_201_1776 ();
 FILLCELL_X32 FILLER_201_1808 ();
 FILLCELL_X32 FILLER_201_1840 ();
 FILLCELL_X32 FILLER_201_1872 ();
 FILLCELL_X32 FILLER_201_1904 ();
 FILLCELL_X32 FILLER_201_1936 ();
 FILLCELL_X32 FILLER_201_1968 ();
 FILLCELL_X32 FILLER_201_2000 ();
 FILLCELL_X32 FILLER_201_2032 ();
 FILLCELL_X32 FILLER_201_2064 ();
 FILLCELL_X32 FILLER_201_2096 ();
 FILLCELL_X32 FILLER_201_2128 ();
 FILLCELL_X32 FILLER_201_2160 ();
 FILLCELL_X32 FILLER_201_2192 ();
 FILLCELL_X32 FILLER_201_2224 ();
 FILLCELL_X32 FILLER_201_2256 ();
 FILLCELL_X32 FILLER_201_2288 ();
 FILLCELL_X32 FILLER_201_2320 ();
 FILLCELL_X32 FILLER_201_2352 ();
 FILLCELL_X32 FILLER_201_2384 ();
 FILLCELL_X32 FILLER_201_2416 ();
 FILLCELL_X32 FILLER_201_2448 ();
 FILLCELL_X32 FILLER_201_2480 ();
 FILLCELL_X8 FILLER_201_2512 ();
 FILLCELL_X4 FILLER_201_2520 ();
 FILLCELL_X2 FILLER_201_2524 ();
 FILLCELL_X32 FILLER_201_2527 ();
 FILLCELL_X32 FILLER_201_2559 ();
 FILLCELL_X32 FILLER_201_2591 ();
 FILLCELL_X32 FILLER_201_2623 ();
 FILLCELL_X32 FILLER_201_2655 ();
 FILLCELL_X32 FILLER_201_2687 ();
 FILLCELL_X32 FILLER_201_2719 ();
 FILLCELL_X32 FILLER_201_2751 ();
 FILLCELL_X32 FILLER_201_2783 ();
 FILLCELL_X32 FILLER_201_2815 ();
 FILLCELL_X32 FILLER_201_2847 ();
 FILLCELL_X32 FILLER_201_2879 ();
 FILLCELL_X32 FILLER_201_2911 ();
 FILLCELL_X32 FILLER_201_2943 ();
 FILLCELL_X32 FILLER_201_2975 ();
 FILLCELL_X32 FILLER_201_3007 ();
 FILLCELL_X32 FILLER_201_3039 ();
 FILLCELL_X32 FILLER_201_3071 ();
 FILLCELL_X32 FILLER_201_3103 ();
 FILLCELL_X32 FILLER_201_3135 ();
 FILLCELL_X32 FILLER_201_3167 ();
 FILLCELL_X32 FILLER_201_3199 ();
 FILLCELL_X32 FILLER_201_3231 ();
 FILLCELL_X32 FILLER_201_3263 ();
 FILLCELL_X32 FILLER_201_3295 ();
 FILLCELL_X32 FILLER_201_3327 ();
 FILLCELL_X32 FILLER_201_3359 ();
 FILLCELL_X32 FILLER_201_3391 ();
 FILLCELL_X32 FILLER_201_3423 ();
 FILLCELL_X32 FILLER_201_3455 ();
 FILLCELL_X32 FILLER_201_3487 ();
 FILLCELL_X32 FILLER_201_3519 ();
 FILLCELL_X32 FILLER_201_3551 ();
 FILLCELL_X32 FILLER_201_3583 ();
 FILLCELL_X32 FILLER_201_3615 ();
 FILLCELL_X32 FILLER_201_3647 ();
 FILLCELL_X32 FILLER_201_3679 ();
 FILLCELL_X16 FILLER_201_3711 ();
 FILLCELL_X8 FILLER_201_3727 ();
 FILLCELL_X2 FILLER_201_3735 ();
 FILLCELL_X1 FILLER_201_3737 ();
 FILLCELL_X32 FILLER_202_1 ();
 FILLCELL_X32 FILLER_202_33 ();
 FILLCELL_X32 FILLER_202_65 ();
 FILLCELL_X32 FILLER_202_97 ();
 FILLCELL_X32 FILLER_202_129 ();
 FILLCELL_X32 FILLER_202_161 ();
 FILLCELL_X32 FILLER_202_193 ();
 FILLCELL_X32 FILLER_202_225 ();
 FILLCELL_X32 FILLER_202_257 ();
 FILLCELL_X32 FILLER_202_289 ();
 FILLCELL_X32 FILLER_202_321 ();
 FILLCELL_X32 FILLER_202_353 ();
 FILLCELL_X32 FILLER_202_385 ();
 FILLCELL_X32 FILLER_202_417 ();
 FILLCELL_X32 FILLER_202_449 ();
 FILLCELL_X32 FILLER_202_481 ();
 FILLCELL_X32 FILLER_202_513 ();
 FILLCELL_X32 FILLER_202_545 ();
 FILLCELL_X32 FILLER_202_577 ();
 FILLCELL_X16 FILLER_202_609 ();
 FILLCELL_X4 FILLER_202_625 ();
 FILLCELL_X2 FILLER_202_629 ();
 FILLCELL_X32 FILLER_202_632 ();
 FILLCELL_X32 FILLER_202_664 ();
 FILLCELL_X32 FILLER_202_696 ();
 FILLCELL_X32 FILLER_202_728 ();
 FILLCELL_X32 FILLER_202_760 ();
 FILLCELL_X32 FILLER_202_792 ();
 FILLCELL_X32 FILLER_202_824 ();
 FILLCELL_X32 FILLER_202_856 ();
 FILLCELL_X32 FILLER_202_888 ();
 FILLCELL_X32 FILLER_202_920 ();
 FILLCELL_X32 FILLER_202_952 ();
 FILLCELL_X32 FILLER_202_984 ();
 FILLCELL_X32 FILLER_202_1016 ();
 FILLCELL_X32 FILLER_202_1048 ();
 FILLCELL_X32 FILLER_202_1080 ();
 FILLCELL_X32 FILLER_202_1112 ();
 FILLCELL_X32 FILLER_202_1144 ();
 FILLCELL_X32 FILLER_202_1176 ();
 FILLCELL_X32 FILLER_202_1208 ();
 FILLCELL_X32 FILLER_202_1240 ();
 FILLCELL_X32 FILLER_202_1272 ();
 FILLCELL_X32 FILLER_202_1304 ();
 FILLCELL_X32 FILLER_202_1336 ();
 FILLCELL_X32 FILLER_202_1368 ();
 FILLCELL_X32 FILLER_202_1400 ();
 FILLCELL_X32 FILLER_202_1432 ();
 FILLCELL_X32 FILLER_202_1464 ();
 FILLCELL_X32 FILLER_202_1496 ();
 FILLCELL_X32 FILLER_202_1528 ();
 FILLCELL_X32 FILLER_202_1560 ();
 FILLCELL_X32 FILLER_202_1592 ();
 FILLCELL_X32 FILLER_202_1624 ();
 FILLCELL_X32 FILLER_202_1656 ();
 FILLCELL_X32 FILLER_202_1688 ();
 FILLCELL_X32 FILLER_202_1720 ();
 FILLCELL_X32 FILLER_202_1752 ();
 FILLCELL_X32 FILLER_202_1784 ();
 FILLCELL_X32 FILLER_202_1816 ();
 FILLCELL_X32 FILLER_202_1848 ();
 FILLCELL_X8 FILLER_202_1880 ();
 FILLCELL_X4 FILLER_202_1888 ();
 FILLCELL_X2 FILLER_202_1892 ();
 FILLCELL_X32 FILLER_202_1895 ();
 FILLCELL_X32 FILLER_202_1927 ();
 FILLCELL_X32 FILLER_202_1959 ();
 FILLCELL_X32 FILLER_202_1991 ();
 FILLCELL_X32 FILLER_202_2023 ();
 FILLCELL_X32 FILLER_202_2055 ();
 FILLCELL_X32 FILLER_202_2087 ();
 FILLCELL_X32 FILLER_202_2119 ();
 FILLCELL_X32 FILLER_202_2151 ();
 FILLCELL_X32 FILLER_202_2183 ();
 FILLCELL_X32 FILLER_202_2215 ();
 FILLCELL_X32 FILLER_202_2247 ();
 FILLCELL_X32 FILLER_202_2279 ();
 FILLCELL_X32 FILLER_202_2311 ();
 FILLCELL_X32 FILLER_202_2343 ();
 FILLCELL_X32 FILLER_202_2375 ();
 FILLCELL_X32 FILLER_202_2407 ();
 FILLCELL_X32 FILLER_202_2439 ();
 FILLCELL_X32 FILLER_202_2471 ();
 FILLCELL_X32 FILLER_202_2503 ();
 FILLCELL_X32 FILLER_202_2535 ();
 FILLCELL_X32 FILLER_202_2567 ();
 FILLCELL_X32 FILLER_202_2599 ();
 FILLCELL_X32 FILLER_202_2631 ();
 FILLCELL_X32 FILLER_202_2663 ();
 FILLCELL_X32 FILLER_202_2695 ();
 FILLCELL_X32 FILLER_202_2727 ();
 FILLCELL_X32 FILLER_202_2759 ();
 FILLCELL_X32 FILLER_202_2791 ();
 FILLCELL_X32 FILLER_202_2823 ();
 FILLCELL_X32 FILLER_202_2855 ();
 FILLCELL_X32 FILLER_202_2887 ();
 FILLCELL_X32 FILLER_202_2919 ();
 FILLCELL_X32 FILLER_202_2951 ();
 FILLCELL_X32 FILLER_202_2983 ();
 FILLCELL_X32 FILLER_202_3015 ();
 FILLCELL_X32 FILLER_202_3047 ();
 FILLCELL_X32 FILLER_202_3079 ();
 FILLCELL_X32 FILLER_202_3111 ();
 FILLCELL_X8 FILLER_202_3143 ();
 FILLCELL_X4 FILLER_202_3151 ();
 FILLCELL_X2 FILLER_202_3155 ();
 FILLCELL_X32 FILLER_202_3158 ();
 FILLCELL_X32 FILLER_202_3190 ();
 FILLCELL_X32 FILLER_202_3222 ();
 FILLCELL_X32 FILLER_202_3254 ();
 FILLCELL_X32 FILLER_202_3286 ();
 FILLCELL_X32 FILLER_202_3318 ();
 FILLCELL_X32 FILLER_202_3350 ();
 FILLCELL_X32 FILLER_202_3382 ();
 FILLCELL_X32 FILLER_202_3414 ();
 FILLCELL_X32 FILLER_202_3446 ();
 FILLCELL_X32 FILLER_202_3478 ();
 FILLCELL_X32 FILLER_202_3510 ();
 FILLCELL_X32 FILLER_202_3542 ();
 FILLCELL_X32 FILLER_202_3574 ();
 FILLCELL_X32 FILLER_202_3606 ();
 FILLCELL_X32 FILLER_202_3638 ();
 FILLCELL_X32 FILLER_202_3670 ();
 FILLCELL_X32 FILLER_202_3702 ();
 FILLCELL_X4 FILLER_202_3734 ();
 FILLCELL_X32 FILLER_203_1 ();
 FILLCELL_X32 FILLER_203_33 ();
 FILLCELL_X32 FILLER_203_65 ();
 FILLCELL_X32 FILLER_203_97 ();
 FILLCELL_X32 FILLER_203_129 ();
 FILLCELL_X32 FILLER_203_161 ();
 FILLCELL_X32 FILLER_203_193 ();
 FILLCELL_X32 FILLER_203_225 ();
 FILLCELL_X32 FILLER_203_257 ();
 FILLCELL_X32 FILLER_203_289 ();
 FILLCELL_X32 FILLER_203_321 ();
 FILLCELL_X32 FILLER_203_353 ();
 FILLCELL_X32 FILLER_203_385 ();
 FILLCELL_X32 FILLER_203_417 ();
 FILLCELL_X32 FILLER_203_449 ();
 FILLCELL_X32 FILLER_203_481 ();
 FILLCELL_X32 FILLER_203_513 ();
 FILLCELL_X32 FILLER_203_545 ();
 FILLCELL_X32 FILLER_203_577 ();
 FILLCELL_X32 FILLER_203_609 ();
 FILLCELL_X32 FILLER_203_641 ();
 FILLCELL_X32 FILLER_203_673 ();
 FILLCELL_X32 FILLER_203_705 ();
 FILLCELL_X32 FILLER_203_737 ();
 FILLCELL_X32 FILLER_203_769 ();
 FILLCELL_X32 FILLER_203_801 ();
 FILLCELL_X32 FILLER_203_833 ();
 FILLCELL_X32 FILLER_203_865 ();
 FILLCELL_X32 FILLER_203_897 ();
 FILLCELL_X32 FILLER_203_929 ();
 FILLCELL_X32 FILLER_203_961 ();
 FILLCELL_X32 FILLER_203_993 ();
 FILLCELL_X32 FILLER_203_1025 ();
 FILLCELL_X32 FILLER_203_1057 ();
 FILLCELL_X32 FILLER_203_1089 ();
 FILLCELL_X32 FILLER_203_1121 ();
 FILLCELL_X32 FILLER_203_1153 ();
 FILLCELL_X32 FILLER_203_1185 ();
 FILLCELL_X32 FILLER_203_1217 ();
 FILLCELL_X8 FILLER_203_1249 ();
 FILLCELL_X4 FILLER_203_1257 ();
 FILLCELL_X2 FILLER_203_1261 ();
 FILLCELL_X32 FILLER_203_1264 ();
 FILLCELL_X32 FILLER_203_1296 ();
 FILLCELL_X32 FILLER_203_1328 ();
 FILLCELL_X32 FILLER_203_1360 ();
 FILLCELL_X32 FILLER_203_1392 ();
 FILLCELL_X32 FILLER_203_1424 ();
 FILLCELL_X32 FILLER_203_1456 ();
 FILLCELL_X32 FILLER_203_1488 ();
 FILLCELL_X32 FILLER_203_1520 ();
 FILLCELL_X32 FILLER_203_1552 ();
 FILLCELL_X32 FILLER_203_1584 ();
 FILLCELL_X32 FILLER_203_1616 ();
 FILLCELL_X32 FILLER_203_1648 ();
 FILLCELL_X32 FILLER_203_1680 ();
 FILLCELL_X32 FILLER_203_1712 ();
 FILLCELL_X32 FILLER_203_1744 ();
 FILLCELL_X32 FILLER_203_1776 ();
 FILLCELL_X32 FILLER_203_1808 ();
 FILLCELL_X32 FILLER_203_1840 ();
 FILLCELL_X32 FILLER_203_1872 ();
 FILLCELL_X32 FILLER_203_1904 ();
 FILLCELL_X32 FILLER_203_1936 ();
 FILLCELL_X32 FILLER_203_1968 ();
 FILLCELL_X32 FILLER_203_2000 ();
 FILLCELL_X32 FILLER_203_2032 ();
 FILLCELL_X32 FILLER_203_2064 ();
 FILLCELL_X32 FILLER_203_2096 ();
 FILLCELL_X32 FILLER_203_2128 ();
 FILLCELL_X32 FILLER_203_2160 ();
 FILLCELL_X32 FILLER_203_2192 ();
 FILLCELL_X32 FILLER_203_2224 ();
 FILLCELL_X32 FILLER_203_2256 ();
 FILLCELL_X32 FILLER_203_2288 ();
 FILLCELL_X32 FILLER_203_2320 ();
 FILLCELL_X32 FILLER_203_2352 ();
 FILLCELL_X32 FILLER_203_2384 ();
 FILLCELL_X32 FILLER_203_2416 ();
 FILLCELL_X32 FILLER_203_2448 ();
 FILLCELL_X32 FILLER_203_2480 ();
 FILLCELL_X8 FILLER_203_2512 ();
 FILLCELL_X4 FILLER_203_2520 ();
 FILLCELL_X2 FILLER_203_2524 ();
 FILLCELL_X32 FILLER_203_2527 ();
 FILLCELL_X32 FILLER_203_2559 ();
 FILLCELL_X32 FILLER_203_2591 ();
 FILLCELL_X32 FILLER_203_2623 ();
 FILLCELL_X32 FILLER_203_2655 ();
 FILLCELL_X32 FILLER_203_2687 ();
 FILLCELL_X32 FILLER_203_2719 ();
 FILLCELL_X32 FILLER_203_2751 ();
 FILLCELL_X32 FILLER_203_2783 ();
 FILLCELL_X32 FILLER_203_2815 ();
 FILLCELL_X32 FILLER_203_2847 ();
 FILLCELL_X32 FILLER_203_2879 ();
 FILLCELL_X32 FILLER_203_2911 ();
 FILLCELL_X32 FILLER_203_2943 ();
 FILLCELL_X32 FILLER_203_2975 ();
 FILLCELL_X32 FILLER_203_3007 ();
 FILLCELL_X32 FILLER_203_3039 ();
 FILLCELL_X32 FILLER_203_3071 ();
 FILLCELL_X32 FILLER_203_3103 ();
 FILLCELL_X32 FILLER_203_3135 ();
 FILLCELL_X32 FILLER_203_3167 ();
 FILLCELL_X32 FILLER_203_3199 ();
 FILLCELL_X32 FILLER_203_3231 ();
 FILLCELL_X32 FILLER_203_3263 ();
 FILLCELL_X32 FILLER_203_3295 ();
 FILLCELL_X32 FILLER_203_3327 ();
 FILLCELL_X32 FILLER_203_3359 ();
 FILLCELL_X32 FILLER_203_3391 ();
 FILLCELL_X32 FILLER_203_3423 ();
 FILLCELL_X32 FILLER_203_3455 ();
 FILLCELL_X32 FILLER_203_3487 ();
 FILLCELL_X32 FILLER_203_3519 ();
 FILLCELL_X32 FILLER_203_3551 ();
 FILLCELL_X32 FILLER_203_3583 ();
 FILLCELL_X32 FILLER_203_3615 ();
 FILLCELL_X32 FILLER_203_3647 ();
 FILLCELL_X32 FILLER_203_3679 ();
 FILLCELL_X16 FILLER_203_3711 ();
 FILLCELL_X8 FILLER_203_3727 ();
 FILLCELL_X2 FILLER_203_3735 ();
 FILLCELL_X1 FILLER_203_3737 ();
 FILLCELL_X32 FILLER_204_1 ();
 FILLCELL_X32 FILLER_204_33 ();
 FILLCELL_X32 FILLER_204_65 ();
 FILLCELL_X32 FILLER_204_97 ();
 FILLCELL_X32 FILLER_204_129 ();
 FILLCELL_X32 FILLER_204_161 ();
 FILLCELL_X32 FILLER_204_193 ();
 FILLCELL_X32 FILLER_204_225 ();
 FILLCELL_X32 FILLER_204_257 ();
 FILLCELL_X32 FILLER_204_289 ();
 FILLCELL_X32 FILLER_204_321 ();
 FILLCELL_X32 FILLER_204_353 ();
 FILLCELL_X32 FILLER_204_385 ();
 FILLCELL_X32 FILLER_204_417 ();
 FILLCELL_X32 FILLER_204_449 ();
 FILLCELL_X32 FILLER_204_481 ();
 FILLCELL_X32 FILLER_204_513 ();
 FILLCELL_X32 FILLER_204_545 ();
 FILLCELL_X32 FILLER_204_577 ();
 FILLCELL_X16 FILLER_204_609 ();
 FILLCELL_X4 FILLER_204_625 ();
 FILLCELL_X2 FILLER_204_629 ();
 FILLCELL_X32 FILLER_204_632 ();
 FILLCELL_X32 FILLER_204_664 ();
 FILLCELL_X32 FILLER_204_696 ();
 FILLCELL_X32 FILLER_204_728 ();
 FILLCELL_X32 FILLER_204_760 ();
 FILLCELL_X32 FILLER_204_792 ();
 FILLCELL_X32 FILLER_204_824 ();
 FILLCELL_X32 FILLER_204_856 ();
 FILLCELL_X32 FILLER_204_888 ();
 FILLCELL_X32 FILLER_204_920 ();
 FILLCELL_X32 FILLER_204_952 ();
 FILLCELL_X32 FILLER_204_984 ();
 FILLCELL_X32 FILLER_204_1016 ();
 FILLCELL_X32 FILLER_204_1048 ();
 FILLCELL_X32 FILLER_204_1080 ();
 FILLCELL_X32 FILLER_204_1112 ();
 FILLCELL_X32 FILLER_204_1144 ();
 FILLCELL_X32 FILLER_204_1176 ();
 FILLCELL_X32 FILLER_204_1208 ();
 FILLCELL_X32 FILLER_204_1240 ();
 FILLCELL_X32 FILLER_204_1272 ();
 FILLCELL_X32 FILLER_204_1304 ();
 FILLCELL_X32 FILLER_204_1336 ();
 FILLCELL_X32 FILLER_204_1368 ();
 FILLCELL_X32 FILLER_204_1400 ();
 FILLCELL_X32 FILLER_204_1432 ();
 FILLCELL_X32 FILLER_204_1464 ();
 FILLCELL_X32 FILLER_204_1496 ();
 FILLCELL_X32 FILLER_204_1528 ();
 FILLCELL_X32 FILLER_204_1560 ();
 FILLCELL_X32 FILLER_204_1592 ();
 FILLCELL_X32 FILLER_204_1624 ();
 FILLCELL_X32 FILLER_204_1656 ();
 FILLCELL_X32 FILLER_204_1688 ();
 FILLCELL_X32 FILLER_204_1720 ();
 FILLCELL_X32 FILLER_204_1752 ();
 FILLCELL_X32 FILLER_204_1784 ();
 FILLCELL_X32 FILLER_204_1816 ();
 FILLCELL_X32 FILLER_204_1848 ();
 FILLCELL_X8 FILLER_204_1880 ();
 FILLCELL_X4 FILLER_204_1888 ();
 FILLCELL_X2 FILLER_204_1892 ();
 FILLCELL_X32 FILLER_204_1895 ();
 FILLCELL_X32 FILLER_204_1927 ();
 FILLCELL_X32 FILLER_204_1959 ();
 FILLCELL_X32 FILLER_204_1991 ();
 FILLCELL_X32 FILLER_204_2023 ();
 FILLCELL_X32 FILLER_204_2055 ();
 FILLCELL_X32 FILLER_204_2087 ();
 FILLCELL_X32 FILLER_204_2119 ();
 FILLCELL_X32 FILLER_204_2151 ();
 FILLCELL_X32 FILLER_204_2183 ();
 FILLCELL_X32 FILLER_204_2215 ();
 FILLCELL_X32 FILLER_204_2247 ();
 FILLCELL_X32 FILLER_204_2279 ();
 FILLCELL_X32 FILLER_204_2311 ();
 FILLCELL_X32 FILLER_204_2343 ();
 FILLCELL_X32 FILLER_204_2375 ();
 FILLCELL_X32 FILLER_204_2407 ();
 FILLCELL_X32 FILLER_204_2439 ();
 FILLCELL_X32 FILLER_204_2471 ();
 FILLCELL_X32 FILLER_204_2503 ();
 FILLCELL_X32 FILLER_204_2535 ();
 FILLCELL_X32 FILLER_204_2567 ();
 FILLCELL_X32 FILLER_204_2599 ();
 FILLCELL_X32 FILLER_204_2631 ();
 FILLCELL_X32 FILLER_204_2663 ();
 FILLCELL_X32 FILLER_204_2695 ();
 FILLCELL_X32 FILLER_204_2727 ();
 FILLCELL_X32 FILLER_204_2759 ();
 FILLCELL_X32 FILLER_204_2791 ();
 FILLCELL_X32 FILLER_204_2823 ();
 FILLCELL_X32 FILLER_204_2855 ();
 FILLCELL_X32 FILLER_204_2887 ();
 FILLCELL_X32 FILLER_204_2919 ();
 FILLCELL_X32 FILLER_204_2951 ();
 FILLCELL_X32 FILLER_204_2983 ();
 FILLCELL_X32 FILLER_204_3015 ();
 FILLCELL_X32 FILLER_204_3047 ();
 FILLCELL_X32 FILLER_204_3079 ();
 FILLCELL_X32 FILLER_204_3111 ();
 FILLCELL_X8 FILLER_204_3143 ();
 FILLCELL_X4 FILLER_204_3151 ();
 FILLCELL_X2 FILLER_204_3155 ();
 FILLCELL_X32 FILLER_204_3158 ();
 FILLCELL_X32 FILLER_204_3190 ();
 FILLCELL_X32 FILLER_204_3222 ();
 FILLCELL_X32 FILLER_204_3254 ();
 FILLCELL_X32 FILLER_204_3286 ();
 FILLCELL_X32 FILLER_204_3318 ();
 FILLCELL_X32 FILLER_204_3350 ();
 FILLCELL_X32 FILLER_204_3382 ();
 FILLCELL_X32 FILLER_204_3414 ();
 FILLCELL_X32 FILLER_204_3446 ();
 FILLCELL_X32 FILLER_204_3478 ();
 FILLCELL_X32 FILLER_204_3510 ();
 FILLCELL_X32 FILLER_204_3542 ();
 FILLCELL_X32 FILLER_204_3574 ();
 FILLCELL_X32 FILLER_204_3606 ();
 FILLCELL_X32 FILLER_204_3638 ();
 FILLCELL_X32 FILLER_204_3670 ();
 FILLCELL_X32 FILLER_204_3702 ();
 FILLCELL_X4 FILLER_204_3734 ();
 FILLCELL_X32 FILLER_205_1 ();
 FILLCELL_X32 FILLER_205_33 ();
 FILLCELL_X32 FILLER_205_65 ();
 FILLCELL_X32 FILLER_205_97 ();
 FILLCELL_X32 FILLER_205_129 ();
 FILLCELL_X32 FILLER_205_161 ();
 FILLCELL_X32 FILLER_205_193 ();
 FILLCELL_X32 FILLER_205_225 ();
 FILLCELL_X32 FILLER_205_257 ();
 FILLCELL_X32 FILLER_205_289 ();
 FILLCELL_X32 FILLER_205_321 ();
 FILLCELL_X32 FILLER_205_353 ();
 FILLCELL_X32 FILLER_205_385 ();
 FILLCELL_X32 FILLER_205_417 ();
 FILLCELL_X32 FILLER_205_449 ();
 FILLCELL_X32 FILLER_205_481 ();
 FILLCELL_X32 FILLER_205_513 ();
 FILLCELL_X32 FILLER_205_545 ();
 FILLCELL_X32 FILLER_205_577 ();
 FILLCELL_X32 FILLER_205_609 ();
 FILLCELL_X32 FILLER_205_641 ();
 FILLCELL_X32 FILLER_205_673 ();
 FILLCELL_X32 FILLER_205_705 ();
 FILLCELL_X32 FILLER_205_737 ();
 FILLCELL_X32 FILLER_205_769 ();
 FILLCELL_X32 FILLER_205_801 ();
 FILLCELL_X32 FILLER_205_833 ();
 FILLCELL_X32 FILLER_205_865 ();
 FILLCELL_X32 FILLER_205_897 ();
 FILLCELL_X32 FILLER_205_929 ();
 FILLCELL_X32 FILLER_205_961 ();
 FILLCELL_X32 FILLER_205_993 ();
 FILLCELL_X32 FILLER_205_1025 ();
 FILLCELL_X32 FILLER_205_1057 ();
 FILLCELL_X32 FILLER_205_1089 ();
 FILLCELL_X32 FILLER_205_1121 ();
 FILLCELL_X32 FILLER_205_1153 ();
 FILLCELL_X32 FILLER_205_1185 ();
 FILLCELL_X32 FILLER_205_1217 ();
 FILLCELL_X8 FILLER_205_1249 ();
 FILLCELL_X4 FILLER_205_1257 ();
 FILLCELL_X2 FILLER_205_1261 ();
 FILLCELL_X32 FILLER_205_1264 ();
 FILLCELL_X32 FILLER_205_1296 ();
 FILLCELL_X32 FILLER_205_1328 ();
 FILLCELL_X32 FILLER_205_1360 ();
 FILLCELL_X32 FILLER_205_1392 ();
 FILLCELL_X32 FILLER_205_1424 ();
 FILLCELL_X32 FILLER_205_1456 ();
 FILLCELL_X32 FILLER_205_1488 ();
 FILLCELL_X32 FILLER_205_1520 ();
 FILLCELL_X32 FILLER_205_1552 ();
 FILLCELL_X32 FILLER_205_1584 ();
 FILLCELL_X32 FILLER_205_1616 ();
 FILLCELL_X32 FILLER_205_1648 ();
 FILLCELL_X32 FILLER_205_1680 ();
 FILLCELL_X32 FILLER_205_1712 ();
 FILLCELL_X32 FILLER_205_1744 ();
 FILLCELL_X32 FILLER_205_1776 ();
 FILLCELL_X32 FILLER_205_1808 ();
 FILLCELL_X32 FILLER_205_1840 ();
 FILLCELL_X32 FILLER_205_1872 ();
 FILLCELL_X32 FILLER_205_1904 ();
 FILLCELL_X32 FILLER_205_1936 ();
 FILLCELL_X32 FILLER_205_1968 ();
 FILLCELL_X32 FILLER_205_2000 ();
 FILLCELL_X32 FILLER_205_2032 ();
 FILLCELL_X32 FILLER_205_2064 ();
 FILLCELL_X32 FILLER_205_2096 ();
 FILLCELL_X32 FILLER_205_2128 ();
 FILLCELL_X32 FILLER_205_2160 ();
 FILLCELL_X32 FILLER_205_2192 ();
 FILLCELL_X32 FILLER_205_2224 ();
 FILLCELL_X32 FILLER_205_2256 ();
 FILLCELL_X32 FILLER_205_2288 ();
 FILLCELL_X32 FILLER_205_2320 ();
 FILLCELL_X32 FILLER_205_2352 ();
 FILLCELL_X32 FILLER_205_2384 ();
 FILLCELL_X32 FILLER_205_2416 ();
 FILLCELL_X32 FILLER_205_2448 ();
 FILLCELL_X32 FILLER_205_2480 ();
 FILLCELL_X8 FILLER_205_2512 ();
 FILLCELL_X4 FILLER_205_2520 ();
 FILLCELL_X2 FILLER_205_2524 ();
 FILLCELL_X32 FILLER_205_2527 ();
 FILLCELL_X32 FILLER_205_2559 ();
 FILLCELL_X32 FILLER_205_2591 ();
 FILLCELL_X32 FILLER_205_2623 ();
 FILLCELL_X32 FILLER_205_2655 ();
 FILLCELL_X32 FILLER_205_2687 ();
 FILLCELL_X32 FILLER_205_2719 ();
 FILLCELL_X32 FILLER_205_2751 ();
 FILLCELL_X32 FILLER_205_2783 ();
 FILLCELL_X32 FILLER_205_2815 ();
 FILLCELL_X32 FILLER_205_2847 ();
 FILLCELL_X32 FILLER_205_2879 ();
 FILLCELL_X32 FILLER_205_2911 ();
 FILLCELL_X32 FILLER_205_2943 ();
 FILLCELL_X32 FILLER_205_2975 ();
 FILLCELL_X32 FILLER_205_3007 ();
 FILLCELL_X32 FILLER_205_3039 ();
 FILLCELL_X32 FILLER_205_3071 ();
 FILLCELL_X32 FILLER_205_3103 ();
 FILLCELL_X32 FILLER_205_3135 ();
 FILLCELL_X32 FILLER_205_3167 ();
 FILLCELL_X32 FILLER_205_3199 ();
 FILLCELL_X32 FILLER_205_3231 ();
 FILLCELL_X32 FILLER_205_3263 ();
 FILLCELL_X32 FILLER_205_3295 ();
 FILLCELL_X32 FILLER_205_3327 ();
 FILLCELL_X32 FILLER_205_3359 ();
 FILLCELL_X32 FILLER_205_3391 ();
 FILLCELL_X32 FILLER_205_3423 ();
 FILLCELL_X32 FILLER_205_3455 ();
 FILLCELL_X32 FILLER_205_3487 ();
 FILLCELL_X32 FILLER_205_3519 ();
 FILLCELL_X32 FILLER_205_3551 ();
 FILLCELL_X32 FILLER_205_3583 ();
 FILLCELL_X32 FILLER_205_3615 ();
 FILLCELL_X32 FILLER_205_3647 ();
 FILLCELL_X32 FILLER_205_3679 ();
 FILLCELL_X16 FILLER_205_3711 ();
 FILLCELL_X8 FILLER_205_3727 ();
 FILLCELL_X2 FILLER_205_3735 ();
 FILLCELL_X1 FILLER_205_3737 ();
 FILLCELL_X32 FILLER_206_1 ();
 FILLCELL_X32 FILLER_206_33 ();
 FILLCELL_X32 FILLER_206_65 ();
 FILLCELL_X32 FILLER_206_97 ();
 FILLCELL_X32 FILLER_206_129 ();
 FILLCELL_X32 FILLER_206_161 ();
 FILLCELL_X32 FILLER_206_193 ();
 FILLCELL_X32 FILLER_206_225 ();
 FILLCELL_X32 FILLER_206_257 ();
 FILLCELL_X32 FILLER_206_289 ();
 FILLCELL_X32 FILLER_206_321 ();
 FILLCELL_X32 FILLER_206_353 ();
 FILLCELL_X32 FILLER_206_385 ();
 FILLCELL_X32 FILLER_206_417 ();
 FILLCELL_X32 FILLER_206_449 ();
 FILLCELL_X32 FILLER_206_481 ();
 FILLCELL_X32 FILLER_206_513 ();
 FILLCELL_X32 FILLER_206_545 ();
 FILLCELL_X32 FILLER_206_577 ();
 FILLCELL_X16 FILLER_206_609 ();
 FILLCELL_X4 FILLER_206_625 ();
 FILLCELL_X2 FILLER_206_629 ();
 FILLCELL_X32 FILLER_206_632 ();
 FILLCELL_X32 FILLER_206_664 ();
 FILLCELL_X32 FILLER_206_696 ();
 FILLCELL_X32 FILLER_206_728 ();
 FILLCELL_X32 FILLER_206_760 ();
 FILLCELL_X32 FILLER_206_792 ();
 FILLCELL_X32 FILLER_206_824 ();
 FILLCELL_X32 FILLER_206_856 ();
 FILLCELL_X32 FILLER_206_888 ();
 FILLCELL_X32 FILLER_206_920 ();
 FILLCELL_X32 FILLER_206_952 ();
 FILLCELL_X32 FILLER_206_984 ();
 FILLCELL_X32 FILLER_206_1016 ();
 FILLCELL_X32 FILLER_206_1048 ();
 FILLCELL_X32 FILLER_206_1080 ();
 FILLCELL_X32 FILLER_206_1112 ();
 FILLCELL_X32 FILLER_206_1144 ();
 FILLCELL_X32 FILLER_206_1176 ();
 FILLCELL_X32 FILLER_206_1208 ();
 FILLCELL_X32 FILLER_206_1240 ();
 FILLCELL_X32 FILLER_206_1272 ();
 FILLCELL_X32 FILLER_206_1304 ();
 FILLCELL_X32 FILLER_206_1336 ();
 FILLCELL_X32 FILLER_206_1368 ();
 FILLCELL_X32 FILLER_206_1400 ();
 FILLCELL_X32 FILLER_206_1432 ();
 FILLCELL_X32 FILLER_206_1464 ();
 FILLCELL_X32 FILLER_206_1496 ();
 FILLCELL_X32 FILLER_206_1528 ();
 FILLCELL_X32 FILLER_206_1560 ();
 FILLCELL_X32 FILLER_206_1592 ();
 FILLCELL_X32 FILLER_206_1624 ();
 FILLCELL_X32 FILLER_206_1656 ();
 FILLCELL_X32 FILLER_206_1688 ();
 FILLCELL_X32 FILLER_206_1720 ();
 FILLCELL_X32 FILLER_206_1752 ();
 FILLCELL_X32 FILLER_206_1784 ();
 FILLCELL_X32 FILLER_206_1816 ();
 FILLCELL_X32 FILLER_206_1848 ();
 FILLCELL_X8 FILLER_206_1880 ();
 FILLCELL_X4 FILLER_206_1888 ();
 FILLCELL_X2 FILLER_206_1892 ();
 FILLCELL_X32 FILLER_206_1895 ();
 FILLCELL_X32 FILLER_206_1927 ();
 FILLCELL_X32 FILLER_206_1959 ();
 FILLCELL_X32 FILLER_206_1991 ();
 FILLCELL_X32 FILLER_206_2023 ();
 FILLCELL_X32 FILLER_206_2055 ();
 FILLCELL_X32 FILLER_206_2087 ();
 FILLCELL_X32 FILLER_206_2119 ();
 FILLCELL_X32 FILLER_206_2151 ();
 FILLCELL_X32 FILLER_206_2183 ();
 FILLCELL_X32 FILLER_206_2215 ();
 FILLCELL_X32 FILLER_206_2247 ();
 FILLCELL_X32 FILLER_206_2279 ();
 FILLCELL_X32 FILLER_206_2311 ();
 FILLCELL_X32 FILLER_206_2343 ();
 FILLCELL_X32 FILLER_206_2375 ();
 FILLCELL_X32 FILLER_206_2407 ();
 FILLCELL_X32 FILLER_206_2439 ();
 FILLCELL_X32 FILLER_206_2471 ();
 FILLCELL_X32 FILLER_206_2503 ();
 FILLCELL_X32 FILLER_206_2535 ();
 FILLCELL_X32 FILLER_206_2567 ();
 FILLCELL_X32 FILLER_206_2599 ();
 FILLCELL_X32 FILLER_206_2631 ();
 FILLCELL_X32 FILLER_206_2663 ();
 FILLCELL_X32 FILLER_206_2695 ();
 FILLCELL_X32 FILLER_206_2727 ();
 FILLCELL_X32 FILLER_206_2759 ();
 FILLCELL_X32 FILLER_206_2791 ();
 FILLCELL_X32 FILLER_206_2823 ();
 FILLCELL_X32 FILLER_206_2855 ();
 FILLCELL_X32 FILLER_206_2887 ();
 FILLCELL_X32 FILLER_206_2919 ();
 FILLCELL_X32 FILLER_206_2951 ();
 FILLCELL_X32 FILLER_206_2983 ();
 FILLCELL_X32 FILLER_206_3015 ();
 FILLCELL_X32 FILLER_206_3047 ();
 FILLCELL_X32 FILLER_206_3079 ();
 FILLCELL_X32 FILLER_206_3111 ();
 FILLCELL_X8 FILLER_206_3143 ();
 FILLCELL_X4 FILLER_206_3151 ();
 FILLCELL_X2 FILLER_206_3155 ();
 FILLCELL_X32 FILLER_206_3158 ();
 FILLCELL_X32 FILLER_206_3190 ();
 FILLCELL_X32 FILLER_206_3222 ();
 FILLCELL_X32 FILLER_206_3254 ();
 FILLCELL_X32 FILLER_206_3286 ();
 FILLCELL_X32 FILLER_206_3318 ();
 FILLCELL_X32 FILLER_206_3350 ();
 FILLCELL_X32 FILLER_206_3382 ();
 FILLCELL_X32 FILLER_206_3414 ();
 FILLCELL_X32 FILLER_206_3446 ();
 FILLCELL_X32 FILLER_206_3478 ();
 FILLCELL_X32 FILLER_206_3510 ();
 FILLCELL_X32 FILLER_206_3542 ();
 FILLCELL_X32 FILLER_206_3574 ();
 FILLCELL_X32 FILLER_206_3606 ();
 FILLCELL_X32 FILLER_206_3638 ();
 FILLCELL_X32 FILLER_206_3670 ();
 FILLCELL_X32 FILLER_206_3702 ();
 FILLCELL_X4 FILLER_206_3734 ();
 FILLCELL_X32 FILLER_207_1 ();
 FILLCELL_X32 FILLER_207_33 ();
 FILLCELL_X32 FILLER_207_65 ();
 FILLCELL_X32 FILLER_207_97 ();
 FILLCELL_X32 FILLER_207_129 ();
 FILLCELL_X32 FILLER_207_161 ();
 FILLCELL_X32 FILLER_207_193 ();
 FILLCELL_X32 FILLER_207_225 ();
 FILLCELL_X32 FILLER_207_257 ();
 FILLCELL_X32 FILLER_207_289 ();
 FILLCELL_X32 FILLER_207_321 ();
 FILLCELL_X32 FILLER_207_353 ();
 FILLCELL_X32 FILLER_207_385 ();
 FILLCELL_X32 FILLER_207_417 ();
 FILLCELL_X32 FILLER_207_449 ();
 FILLCELL_X32 FILLER_207_481 ();
 FILLCELL_X32 FILLER_207_513 ();
 FILLCELL_X32 FILLER_207_545 ();
 FILLCELL_X32 FILLER_207_577 ();
 FILLCELL_X32 FILLER_207_609 ();
 FILLCELL_X32 FILLER_207_641 ();
 FILLCELL_X32 FILLER_207_673 ();
 FILLCELL_X32 FILLER_207_705 ();
 FILLCELL_X32 FILLER_207_737 ();
 FILLCELL_X32 FILLER_207_769 ();
 FILLCELL_X32 FILLER_207_801 ();
 FILLCELL_X32 FILLER_207_833 ();
 FILLCELL_X32 FILLER_207_865 ();
 FILLCELL_X32 FILLER_207_897 ();
 FILLCELL_X32 FILLER_207_929 ();
 FILLCELL_X32 FILLER_207_961 ();
 FILLCELL_X32 FILLER_207_993 ();
 FILLCELL_X32 FILLER_207_1025 ();
 FILLCELL_X32 FILLER_207_1057 ();
 FILLCELL_X32 FILLER_207_1089 ();
 FILLCELL_X32 FILLER_207_1121 ();
 FILLCELL_X32 FILLER_207_1153 ();
 FILLCELL_X32 FILLER_207_1185 ();
 FILLCELL_X32 FILLER_207_1217 ();
 FILLCELL_X8 FILLER_207_1249 ();
 FILLCELL_X4 FILLER_207_1257 ();
 FILLCELL_X2 FILLER_207_1261 ();
 FILLCELL_X32 FILLER_207_1264 ();
 FILLCELL_X32 FILLER_207_1296 ();
 FILLCELL_X32 FILLER_207_1328 ();
 FILLCELL_X32 FILLER_207_1360 ();
 FILLCELL_X32 FILLER_207_1392 ();
 FILLCELL_X32 FILLER_207_1424 ();
 FILLCELL_X32 FILLER_207_1456 ();
 FILLCELL_X32 FILLER_207_1488 ();
 FILLCELL_X32 FILLER_207_1520 ();
 FILLCELL_X32 FILLER_207_1552 ();
 FILLCELL_X32 FILLER_207_1584 ();
 FILLCELL_X32 FILLER_207_1616 ();
 FILLCELL_X32 FILLER_207_1648 ();
 FILLCELL_X32 FILLER_207_1680 ();
 FILLCELL_X32 FILLER_207_1712 ();
 FILLCELL_X32 FILLER_207_1744 ();
 FILLCELL_X32 FILLER_207_1776 ();
 FILLCELL_X32 FILLER_207_1808 ();
 FILLCELL_X32 FILLER_207_1840 ();
 FILLCELL_X32 FILLER_207_1872 ();
 FILLCELL_X32 FILLER_207_1904 ();
 FILLCELL_X32 FILLER_207_1936 ();
 FILLCELL_X32 FILLER_207_1968 ();
 FILLCELL_X32 FILLER_207_2000 ();
 FILLCELL_X32 FILLER_207_2032 ();
 FILLCELL_X32 FILLER_207_2064 ();
 FILLCELL_X32 FILLER_207_2096 ();
 FILLCELL_X32 FILLER_207_2128 ();
 FILLCELL_X32 FILLER_207_2160 ();
 FILLCELL_X32 FILLER_207_2192 ();
 FILLCELL_X32 FILLER_207_2224 ();
 FILLCELL_X32 FILLER_207_2256 ();
 FILLCELL_X32 FILLER_207_2288 ();
 FILLCELL_X32 FILLER_207_2320 ();
 FILLCELL_X32 FILLER_207_2352 ();
 FILLCELL_X32 FILLER_207_2384 ();
 FILLCELL_X32 FILLER_207_2416 ();
 FILLCELL_X32 FILLER_207_2448 ();
 FILLCELL_X32 FILLER_207_2480 ();
 FILLCELL_X8 FILLER_207_2512 ();
 FILLCELL_X4 FILLER_207_2520 ();
 FILLCELL_X2 FILLER_207_2524 ();
 FILLCELL_X32 FILLER_207_2527 ();
 FILLCELL_X32 FILLER_207_2559 ();
 FILLCELL_X32 FILLER_207_2591 ();
 FILLCELL_X32 FILLER_207_2623 ();
 FILLCELL_X32 FILLER_207_2655 ();
 FILLCELL_X32 FILLER_207_2687 ();
 FILLCELL_X32 FILLER_207_2719 ();
 FILLCELL_X32 FILLER_207_2751 ();
 FILLCELL_X32 FILLER_207_2783 ();
 FILLCELL_X32 FILLER_207_2815 ();
 FILLCELL_X32 FILLER_207_2847 ();
 FILLCELL_X32 FILLER_207_2879 ();
 FILLCELL_X32 FILLER_207_2911 ();
 FILLCELL_X32 FILLER_207_2943 ();
 FILLCELL_X32 FILLER_207_2975 ();
 FILLCELL_X32 FILLER_207_3007 ();
 FILLCELL_X32 FILLER_207_3039 ();
 FILLCELL_X32 FILLER_207_3071 ();
 FILLCELL_X32 FILLER_207_3103 ();
 FILLCELL_X32 FILLER_207_3135 ();
 FILLCELL_X32 FILLER_207_3167 ();
 FILLCELL_X32 FILLER_207_3199 ();
 FILLCELL_X32 FILLER_207_3231 ();
 FILLCELL_X32 FILLER_207_3263 ();
 FILLCELL_X32 FILLER_207_3295 ();
 FILLCELL_X32 FILLER_207_3327 ();
 FILLCELL_X32 FILLER_207_3359 ();
 FILLCELL_X32 FILLER_207_3391 ();
 FILLCELL_X32 FILLER_207_3423 ();
 FILLCELL_X32 FILLER_207_3455 ();
 FILLCELL_X32 FILLER_207_3487 ();
 FILLCELL_X32 FILLER_207_3519 ();
 FILLCELL_X32 FILLER_207_3551 ();
 FILLCELL_X32 FILLER_207_3583 ();
 FILLCELL_X32 FILLER_207_3615 ();
 FILLCELL_X32 FILLER_207_3647 ();
 FILLCELL_X32 FILLER_207_3679 ();
 FILLCELL_X16 FILLER_207_3711 ();
 FILLCELL_X8 FILLER_207_3727 ();
 FILLCELL_X2 FILLER_207_3735 ();
 FILLCELL_X1 FILLER_207_3737 ();
 FILLCELL_X32 FILLER_208_1 ();
 FILLCELL_X32 FILLER_208_33 ();
 FILLCELL_X32 FILLER_208_65 ();
 FILLCELL_X32 FILLER_208_97 ();
 FILLCELL_X32 FILLER_208_129 ();
 FILLCELL_X32 FILLER_208_161 ();
 FILLCELL_X32 FILLER_208_193 ();
 FILLCELL_X32 FILLER_208_225 ();
 FILLCELL_X32 FILLER_208_257 ();
 FILLCELL_X32 FILLER_208_289 ();
 FILLCELL_X32 FILLER_208_321 ();
 FILLCELL_X32 FILLER_208_353 ();
 FILLCELL_X32 FILLER_208_385 ();
 FILLCELL_X32 FILLER_208_417 ();
 FILLCELL_X32 FILLER_208_449 ();
 FILLCELL_X32 FILLER_208_481 ();
 FILLCELL_X32 FILLER_208_513 ();
 FILLCELL_X32 FILLER_208_545 ();
 FILLCELL_X32 FILLER_208_577 ();
 FILLCELL_X16 FILLER_208_609 ();
 FILLCELL_X4 FILLER_208_625 ();
 FILLCELL_X2 FILLER_208_629 ();
 FILLCELL_X32 FILLER_208_632 ();
 FILLCELL_X32 FILLER_208_664 ();
 FILLCELL_X32 FILLER_208_696 ();
 FILLCELL_X32 FILLER_208_728 ();
 FILLCELL_X32 FILLER_208_760 ();
 FILLCELL_X32 FILLER_208_792 ();
 FILLCELL_X32 FILLER_208_824 ();
 FILLCELL_X32 FILLER_208_856 ();
 FILLCELL_X32 FILLER_208_888 ();
 FILLCELL_X32 FILLER_208_920 ();
 FILLCELL_X32 FILLER_208_952 ();
 FILLCELL_X32 FILLER_208_984 ();
 FILLCELL_X32 FILLER_208_1016 ();
 FILLCELL_X32 FILLER_208_1048 ();
 FILLCELL_X32 FILLER_208_1080 ();
 FILLCELL_X32 FILLER_208_1112 ();
 FILLCELL_X32 FILLER_208_1144 ();
 FILLCELL_X32 FILLER_208_1176 ();
 FILLCELL_X32 FILLER_208_1208 ();
 FILLCELL_X32 FILLER_208_1240 ();
 FILLCELL_X32 FILLER_208_1272 ();
 FILLCELL_X32 FILLER_208_1304 ();
 FILLCELL_X32 FILLER_208_1336 ();
 FILLCELL_X32 FILLER_208_1368 ();
 FILLCELL_X32 FILLER_208_1400 ();
 FILLCELL_X32 FILLER_208_1432 ();
 FILLCELL_X32 FILLER_208_1464 ();
 FILLCELL_X32 FILLER_208_1496 ();
 FILLCELL_X32 FILLER_208_1528 ();
 FILLCELL_X32 FILLER_208_1560 ();
 FILLCELL_X32 FILLER_208_1592 ();
 FILLCELL_X32 FILLER_208_1624 ();
 FILLCELL_X32 FILLER_208_1656 ();
 FILLCELL_X32 FILLER_208_1688 ();
 FILLCELL_X32 FILLER_208_1720 ();
 FILLCELL_X32 FILLER_208_1752 ();
 FILLCELL_X32 FILLER_208_1784 ();
 FILLCELL_X32 FILLER_208_1816 ();
 FILLCELL_X32 FILLER_208_1848 ();
 FILLCELL_X8 FILLER_208_1880 ();
 FILLCELL_X4 FILLER_208_1888 ();
 FILLCELL_X2 FILLER_208_1892 ();
 FILLCELL_X32 FILLER_208_1895 ();
 FILLCELL_X32 FILLER_208_1927 ();
 FILLCELL_X32 FILLER_208_1959 ();
 FILLCELL_X32 FILLER_208_1991 ();
 FILLCELL_X32 FILLER_208_2023 ();
 FILLCELL_X32 FILLER_208_2055 ();
 FILLCELL_X32 FILLER_208_2087 ();
 FILLCELL_X32 FILLER_208_2119 ();
 FILLCELL_X32 FILLER_208_2151 ();
 FILLCELL_X32 FILLER_208_2183 ();
 FILLCELL_X32 FILLER_208_2215 ();
 FILLCELL_X32 FILLER_208_2247 ();
 FILLCELL_X32 FILLER_208_2279 ();
 FILLCELL_X32 FILLER_208_2311 ();
 FILLCELL_X32 FILLER_208_2343 ();
 FILLCELL_X32 FILLER_208_2375 ();
 FILLCELL_X32 FILLER_208_2407 ();
 FILLCELL_X32 FILLER_208_2439 ();
 FILLCELL_X32 FILLER_208_2471 ();
 FILLCELL_X32 FILLER_208_2503 ();
 FILLCELL_X32 FILLER_208_2535 ();
 FILLCELL_X32 FILLER_208_2567 ();
 FILLCELL_X32 FILLER_208_2599 ();
 FILLCELL_X32 FILLER_208_2631 ();
 FILLCELL_X32 FILLER_208_2663 ();
 FILLCELL_X32 FILLER_208_2695 ();
 FILLCELL_X32 FILLER_208_2727 ();
 FILLCELL_X32 FILLER_208_2759 ();
 FILLCELL_X32 FILLER_208_2791 ();
 FILLCELL_X32 FILLER_208_2823 ();
 FILLCELL_X32 FILLER_208_2855 ();
 FILLCELL_X32 FILLER_208_2887 ();
 FILLCELL_X32 FILLER_208_2919 ();
 FILLCELL_X32 FILLER_208_2951 ();
 FILLCELL_X32 FILLER_208_2983 ();
 FILLCELL_X32 FILLER_208_3015 ();
 FILLCELL_X32 FILLER_208_3047 ();
 FILLCELL_X32 FILLER_208_3079 ();
 FILLCELL_X32 FILLER_208_3111 ();
 FILLCELL_X8 FILLER_208_3143 ();
 FILLCELL_X4 FILLER_208_3151 ();
 FILLCELL_X2 FILLER_208_3155 ();
 FILLCELL_X32 FILLER_208_3158 ();
 FILLCELL_X32 FILLER_208_3190 ();
 FILLCELL_X32 FILLER_208_3222 ();
 FILLCELL_X32 FILLER_208_3254 ();
 FILLCELL_X32 FILLER_208_3286 ();
 FILLCELL_X32 FILLER_208_3318 ();
 FILLCELL_X32 FILLER_208_3350 ();
 FILLCELL_X32 FILLER_208_3382 ();
 FILLCELL_X32 FILLER_208_3414 ();
 FILLCELL_X32 FILLER_208_3446 ();
 FILLCELL_X32 FILLER_208_3478 ();
 FILLCELL_X32 FILLER_208_3510 ();
 FILLCELL_X32 FILLER_208_3542 ();
 FILLCELL_X32 FILLER_208_3574 ();
 FILLCELL_X32 FILLER_208_3606 ();
 FILLCELL_X32 FILLER_208_3638 ();
 FILLCELL_X32 FILLER_208_3670 ();
 FILLCELL_X32 FILLER_208_3702 ();
 FILLCELL_X4 FILLER_208_3734 ();
 FILLCELL_X32 FILLER_209_1 ();
 FILLCELL_X32 FILLER_209_33 ();
 FILLCELL_X32 FILLER_209_65 ();
 FILLCELL_X32 FILLER_209_97 ();
 FILLCELL_X32 FILLER_209_129 ();
 FILLCELL_X32 FILLER_209_161 ();
 FILLCELL_X32 FILLER_209_193 ();
 FILLCELL_X32 FILLER_209_225 ();
 FILLCELL_X32 FILLER_209_257 ();
 FILLCELL_X32 FILLER_209_289 ();
 FILLCELL_X32 FILLER_209_321 ();
 FILLCELL_X32 FILLER_209_353 ();
 FILLCELL_X32 FILLER_209_385 ();
 FILLCELL_X32 FILLER_209_417 ();
 FILLCELL_X32 FILLER_209_449 ();
 FILLCELL_X32 FILLER_209_481 ();
 FILLCELL_X32 FILLER_209_513 ();
 FILLCELL_X32 FILLER_209_545 ();
 FILLCELL_X32 FILLER_209_577 ();
 FILLCELL_X32 FILLER_209_609 ();
 FILLCELL_X32 FILLER_209_641 ();
 FILLCELL_X32 FILLER_209_673 ();
 FILLCELL_X32 FILLER_209_705 ();
 FILLCELL_X32 FILLER_209_737 ();
 FILLCELL_X32 FILLER_209_769 ();
 FILLCELL_X32 FILLER_209_801 ();
 FILLCELL_X32 FILLER_209_833 ();
 FILLCELL_X32 FILLER_209_865 ();
 FILLCELL_X32 FILLER_209_897 ();
 FILLCELL_X32 FILLER_209_929 ();
 FILLCELL_X32 FILLER_209_961 ();
 FILLCELL_X32 FILLER_209_993 ();
 FILLCELL_X32 FILLER_209_1025 ();
 FILLCELL_X32 FILLER_209_1057 ();
 FILLCELL_X32 FILLER_209_1089 ();
 FILLCELL_X32 FILLER_209_1121 ();
 FILLCELL_X32 FILLER_209_1153 ();
 FILLCELL_X32 FILLER_209_1185 ();
 FILLCELL_X32 FILLER_209_1217 ();
 FILLCELL_X8 FILLER_209_1249 ();
 FILLCELL_X4 FILLER_209_1257 ();
 FILLCELL_X2 FILLER_209_1261 ();
 FILLCELL_X32 FILLER_209_1264 ();
 FILLCELL_X32 FILLER_209_1296 ();
 FILLCELL_X32 FILLER_209_1328 ();
 FILLCELL_X32 FILLER_209_1360 ();
 FILLCELL_X32 FILLER_209_1392 ();
 FILLCELL_X32 FILLER_209_1424 ();
 FILLCELL_X32 FILLER_209_1456 ();
 FILLCELL_X32 FILLER_209_1488 ();
 FILLCELL_X32 FILLER_209_1520 ();
 FILLCELL_X32 FILLER_209_1552 ();
 FILLCELL_X32 FILLER_209_1584 ();
 FILLCELL_X32 FILLER_209_1616 ();
 FILLCELL_X32 FILLER_209_1648 ();
 FILLCELL_X32 FILLER_209_1680 ();
 FILLCELL_X32 FILLER_209_1712 ();
 FILLCELL_X32 FILLER_209_1744 ();
 FILLCELL_X32 FILLER_209_1776 ();
 FILLCELL_X32 FILLER_209_1808 ();
 FILLCELL_X32 FILLER_209_1840 ();
 FILLCELL_X32 FILLER_209_1872 ();
 FILLCELL_X32 FILLER_209_1904 ();
 FILLCELL_X32 FILLER_209_1936 ();
 FILLCELL_X32 FILLER_209_1968 ();
 FILLCELL_X32 FILLER_209_2000 ();
 FILLCELL_X32 FILLER_209_2032 ();
 FILLCELL_X32 FILLER_209_2064 ();
 FILLCELL_X32 FILLER_209_2096 ();
 FILLCELL_X32 FILLER_209_2128 ();
 FILLCELL_X32 FILLER_209_2160 ();
 FILLCELL_X32 FILLER_209_2192 ();
 FILLCELL_X32 FILLER_209_2224 ();
 FILLCELL_X32 FILLER_209_2256 ();
 FILLCELL_X32 FILLER_209_2288 ();
 FILLCELL_X32 FILLER_209_2320 ();
 FILLCELL_X32 FILLER_209_2352 ();
 FILLCELL_X32 FILLER_209_2384 ();
 FILLCELL_X32 FILLER_209_2416 ();
 FILLCELL_X32 FILLER_209_2448 ();
 FILLCELL_X32 FILLER_209_2480 ();
 FILLCELL_X8 FILLER_209_2512 ();
 FILLCELL_X4 FILLER_209_2520 ();
 FILLCELL_X2 FILLER_209_2524 ();
 FILLCELL_X32 FILLER_209_2527 ();
 FILLCELL_X32 FILLER_209_2559 ();
 FILLCELL_X32 FILLER_209_2591 ();
 FILLCELL_X32 FILLER_209_2623 ();
 FILLCELL_X32 FILLER_209_2655 ();
 FILLCELL_X32 FILLER_209_2687 ();
 FILLCELL_X32 FILLER_209_2719 ();
 FILLCELL_X32 FILLER_209_2751 ();
 FILLCELL_X32 FILLER_209_2783 ();
 FILLCELL_X32 FILLER_209_2815 ();
 FILLCELL_X32 FILLER_209_2847 ();
 FILLCELL_X32 FILLER_209_2879 ();
 FILLCELL_X32 FILLER_209_2911 ();
 FILLCELL_X32 FILLER_209_2943 ();
 FILLCELL_X32 FILLER_209_2975 ();
 FILLCELL_X32 FILLER_209_3007 ();
 FILLCELL_X32 FILLER_209_3039 ();
 FILLCELL_X32 FILLER_209_3071 ();
 FILLCELL_X32 FILLER_209_3103 ();
 FILLCELL_X32 FILLER_209_3135 ();
 FILLCELL_X32 FILLER_209_3167 ();
 FILLCELL_X32 FILLER_209_3199 ();
 FILLCELL_X32 FILLER_209_3231 ();
 FILLCELL_X32 FILLER_209_3263 ();
 FILLCELL_X32 FILLER_209_3295 ();
 FILLCELL_X32 FILLER_209_3327 ();
 FILLCELL_X32 FILLER_209_3359 ();
 FILLCELL_X32 FILLER_209_3391 ();
 FILLCELL_X32 FILLER_209_3423 ();
 FILLCELL_X32 FILLER_209_3455 ();
 FILLCELL_X32 FILLER_209_3487 ();
 FILLCELL_X32 FILLER_209_3519 ();
 FILLCELL_X32 FILLER_209_3551 ();
 FILLCELL_X32 FILLER_209_3583 ();
 FILLCELL_X32 FILLER_209_3615 ();
 FILLCELL_X32 FILLER_209_3647 ();
 FILLCELL_X32 FILLER_209_3679 ();
 FILLCELL_X16 FILLER_209_3711 ();
 FILLCELL_X8 FILLER_209_3727 ();
 FILLCELL_X2 FILLER_209_3735 ();
 FILLCELL_X1 FILLER_209_3737 ();
 FILLCELL_X32 FILLER_210_1 ();
 FILLCELL_X32 FILLER_210_33 ();
 FILLCELL_X32 FILLER_210_65 ();
 FILLCELL_X32 FILLER_210_97 ();
 FILLCELL_X32 FILLER_210_129 ();
 FILLCELL_X32 FILLER_210_161 ();
 FILLCELL_X32 FILLER_210_193 ();
 FILLCELL_X32 FILLER_210_225 ();
 FILLCELL_X32 FILLER_210_257 ();
 FILLCELL_X32 FILLER_210_289 ();
 FILLCELL_X32 FILLER_210_321 ();
 FILLCELL_X32 FILLER_210_353 ();
 FILLCELL_X32 FILLER_210_385 ();
 FILLCELL_X32 FILLER_210_417 ();
 FILLCELL_X32 FILLER_210_449 ();
 FILLCELL_X32 FILLER_210_481 ();
 FILLCELL_X32 FILLER_210_513 ();
 FILLCELL_X32 FILLER_210_545 ();
 FILLCELL_X32 FILLER_210_577 ();
 FILLCELL_X16 FILLER_210_609 ();
 FILLCELL_X4 FILLER_210_625 ();
 FILLCELL_X2 FILLER_210_629 ();
 FILLCELL_X32 FILLER_210_632 ();
 FILLCELL_X32 FILLER_210_664 ();
 FILLCELL_X32 FILLER_210_696 ();
 FILLCELL_X32 FILLER_210_728 ();
 FILLCELL_X32 FILLER_210_760 ();
 FILLCELL_X32 FILLER_210_792 ();
 FILLCELL_X32 FILLER_210_824 ();
 FILLCELL_X32 FILLER_210_856 ();
 FILLCELL_X32 FILLER_210_888 ();
 FILLCELL_X32 FILLER_210_920 ();
 FILLCELL_X32 FILLER_210_952 ();
 FILLCELL_X32 FILLER_210_984 ();
 FILLCELL_X32 FILLER_210_1016 ();
 FILLCELL_X32 FILLER_210_1048 ();
 FILLCELL_X32 FILLER_210_1080 ();
 FILLCELL_X32 FILLER_210_1112 ();
 FILLCELL_X32 FILLER_210_1144 ();
 FILLCELL_X32 FILLER_210_1176 ();
 FILLCELL_X32 FILLER_210_1208 ();
 FILLCELL_X32 FILLER_210_1240 ();
 FILLCELL_X32 FILLER_210_1272 ();
 FILLCELL_X32 FILLER_210_1304 ();
 FILLCELL_X32 FILLER_210_1336 ();
 FILLCELL_X32 FILLER_210_1368 ();
 FILLCELL_X32 FILLER_210_1400 ();
 FILLCELL_X32 FILLER_210_1432 ();
 FILLCELL_X32 FILLER_210_1464 ();
 FILLCELL_X32 FILLER_210_1496 ();
 FILLCELL_X32 FILLER_210_1528 ();
 FILLCELL_X32 FILLER_210_1560 ();
 FILLCELL_X32 FILLER_210_1592 ();
 FILLCELL_X32 FILLER_210_1624 ();
 FILLCELL_X32 FILLER_210_1656 ();
 FILLCELL_X32 FILLER_210_1688 ();
 FILLCELL_X32 FILLER_210_1720 ();
 FILLCELL_X32 FILLER_210_1752 ();
 FILLCELL_X32 FILLER_210_1784 ();
 FILLCELL_X32 FILLER_210_1816 ();
 FILLCELL_X32 FILLER_210_1848 ();
 FILLCELL_X8 FILLER_210_1880 ();
 FILLCELL_X4 FILLER_210_1888 ();
 FILLCELL_X2 FILLER_210_1892 ();
 FILLCELL_X32 FILLER_210_1895 ();
 FILLCELL_X32 FILLER_210_1927 ();
 FILLCELL_X32 FILLER_210_1959 ();
 FILLCELL_X32 FILLER_210_1991 ();
 FILLCELL_X32 FILLER_210_2023 ();
 FILLCELL_X32 FILLER_210_2055 ();
 FILLCELL_X32 FILLER_210_2087 ();
 FILLCELL_X32 FILLER_210_2119 ();
 FILLCELL_X32 FILLER_210_2151 ();
 FILLCELL_X32 FILLER_210_2183 ();
 FILLCELL_X32 FILLER_210_2215 ();
 FILLCELL_X32 FILLER_210_2247 ();
 FILLCELL_X32 FILLER_210_2279 ();
 FILLCELL_X32 FILLER_210_2311 ();
 FILLCELL_X32 FILLER_210_2343 ();
 FILLCELL_X32 FILLER_210_2375 ();
 FILLCELL_X32 FILLER_210_2407 ();
 FILLCELL_X32 FILLER_210_2439 ();
 FILLCELL_X32 FILLER_210_2471 ();
 FILLCELL_X32 FILLER_210_2503 ();
 FILLCELL_X32 FILLER_210_2535 ();
 FILLCELL_X32 FILLER_210_2567 ();
 FILLCELL_X32 FILLER_210_2599 ();
 FILLCELL_X32 FILLER_210_2631 ();
 FILLCELL_X32 FILLER_210_2663 ();
 FILLCELL_X32 FILLER_210_2695 ();
 FILLCELL_X32 FILLER_210_2727 ();
 FILLCELL_X32 FILLER_210_2759 ();
 FILLCELL_X32 FILLER_210_2791 ();
 FILLCELL_X32 FILLER_210_2823 ();
 FILLCELL_X32 FILLER_210_2855 ();
 FILLCELL_X32 FILLER_210_2887 ();
 FILLCELL_X32 FILLER_210_2919 ();
 FILLCELL_X32 FILLER_210_2951 ();
 FILLCELL_X32 FILLER_210_2983 ();
 FILLCELL_X32 FILLER_210_3015 ();
 FILLCELL_X32 FILLER_210_3047 ();
 FILLCELL_X32 FILLER_210_3079 ();
 FILLCELL_X32 FILLER_210_3111 ();
 FILLCELL_X8 FILLER_210_3143 ();
 FILLCELL_X4 FILLER_210_3151 ();
 FILLCELL_X2 FILLER_210_3155 ();
 FILLCELL_X32 FILLER_210_3158 ();
 FILLCELL_X32 FILLER_210_3190 ();
 FILLCELL_X32 FILLER_210_3222 ();
 FILLCELL_X32 FILLER_210_3254 ();
 FILLCELL_X32 FILLER_210_3286 ();
 FILLCELL_X32 FILLER_210_3318 ();
 FILLCELL_X32 FILLER_210_3350 ();
 FILLCELL_X32 FILLER_210_3382 ();
 FILLCELL_X32 FILLER_210_3414 ();
 FILLCELL_X32 FILLER_210_3446 ();
 FILLCELL_X32 FILLER_210_3478 ();
 FILLCELL_X32 FILLER_210_3510 ();
 FILLCELL_X32 FILLER_210_3542 ();
 FILLCELL_X32 FILLER_210_3574 ();
 FILLCELL_X32 FILLER_210_3606 ();
 FILLCELL_X32 FILLER_210_3638 ();
 FILLCELL_X32 FILLER_210_3670 ();
 FILLCELL_X32 FILLER_210_3702 ();
 FILLCELL_X4 FILLER_210_3734 ();
 FILLCELL_X32 FILLER_211_1 ();
 FILLCELL_X32 FILLER_211_33 ();
 FILLCELL_X32 FILLER_211_65 ();
 FILLCELL_X32 FILLER_211_97 ();
 FILLCELL_X32 FILLER_211_129 ();
 FILLCELL_X32 FILLER_211_161 ();
 FILLCELL_X32 FILLER_211_193 ();
 FILLCELL_X32 FILLER_211_225 ();
 FILLCELL_X32 FILLER_211_257 ();
 FILLCELL_X32 FILLER_211_289 ();
 FILLCELL_X32 FILLER_211_321 ();
 FILLCELL_X32 FILLER_211_353 ();
 FILLCELL_X32 FILLER_211_385 ();
 FILLCELL_X32 FILLER_211_417 ();
 FILLCELL_X32 FILLER_211_449 ();
 FILLCELL_X32 FILLER_211_481 ();
 FILLCELL_X32 FILLER_211_513 ();
 FILLCELL_X32 FILLER_211_545 ();
 FILLCELL_X32 FILLER_211_577 ();
 FILLCELL_X32 FILLER_211_609 ();
 FILLCELL_X32 FILLER_211_641 ();
 FILLCELL_X32 FILLER_211_673 ();
 FILLCELL_X32 FILLER_211_705 ();
 FILLCELL_X32 FILLER_211_737 ();
 FILLCELL_X32 FILLER_211_769 ();
 FILLCELL_X32 FILLER_211_801 ();
 FILLCELL_X32 FILLER_211_833 ();
 FILLCELL_X32 FILLER_211_865 ();
 FILLCELL_X32 FILLER_211_897 ();
 FILLCELL_X32 FILLER_211_929 ();
 FILLCELL_X32 FILLER_211_961 ();
 FILLCELL_X32 FILLER_211_993 ();
 FILLCELL_X32 FILLER_211_1025 ();
 FILLCELL_X32 FILLER_211_1057 ();
 FILLCELL_X32 FILLER_211_1089 ();
 FILLCELL_X32 FILLER_211_1121 ();
 FILLCELL_X32 FILLER_211_1153 ();
 FILLCELL_X32 FILLER_211_1185 ();
 FILLCELL_X32 FILLER_211_1217 ();
 FILLCELL_X8 FILLER_211_1249 ();
 FILLCELL_X4 FILLER_211_1257 ();
 FILLCELL_X2 FILLER_211_1261 ();
 FILLCELL_X32 FILLER_211_1264 ();
 FILLCELL_X32 FILLER_211_1296 ();
 FILLCELL_X32 FILLER_211_1328 ();
 FILLCELL_X32 FILLER_211_1360 ();
 FILLCELL_X32 FILLER_211_1392 ();
 FILLCELL_X32 FILLER_211_1424 ();
 FILLCELL_X32 FILLER_211_1456 ();
 FILLCELL_X32 FILLER_211_1488 ();
 FILLCELL_X32 FILLER_211_1520 ();
 FILLCELL_X32 FILLER_211_1552 ();
 FILLCELL_X32 FILLER_211_1584 ();
 FILLCELL_X32 FILLER_211_1616 ();
 FILLCELL_X32 FILLER_211_1648 ();
 FILLCELL_X32 FILLER_211_1680 ();
 FILLCELL_X32 FILLER_211_1712 ();
 FILLCELL_X32 FILLER_211_1744 ();
 FILLCELL_X32 FILLER_211_1776 ();
 FILLCELL_X32 FILLER_211_1808 ();
 FILLCELL_X32 FILLER_211_1840 ();
 FILLCELL_X32 FILLER_211_1872 ();
 FILLCELL_X32 FILLER_211_1904 ();
 FILLCELL_X32 FILLER_211_1936 ();
 FILLCELL_X32 FILLER_211_1968 ();
 FILLCELL_X32 FILLER_211_2000 ();
 FILLCELL_X32 FILLER_211_2032 ();
 FILLCELL_X32 FILLER_211_2064 ();
 FILLCELL_X32 FILLER_211_2096 ();
 FILLCELL_X32 FILLER_211_2128 ();
 FILLCELL_X32 FILLER_211_2160 ();
 FILLCELL_X32 FILLER_211_2192 ();
 FILLCELL_X32 FILLER_211_2224 ();
 FILLCELL_X32 FILLER_211_2256 ();
 FILLCELL_X32 FILLER_211_2288 ();
 FILLCELL_X32 FILLER_211_2320 ();
 FILLCELL_X32 FILLER_211_2352 ();
 FILLCELL_X32 FILLER_211_2384 ();
 FILLCELL_X32 FILLER_211_2416 ();
 FILLCELL_X32 FILLER_211_2448 ();
 FILLCELL_X32 FILLER_211_2480 ();
 FILLCELL_X8 FILLER_211_2512 ();
 FILLCELL_X4 FILLER_211_2520 ();
 FILLCELL_X2 FILLER_211_2524 ();
 FILLCELL_X32 FILLER_211_2527 ();
 FILLCELL_X32 FILLER_211_2559 ();
 FILLCELL_X32 FILLER_211_2591 ();
 FILLCELL_X32 FILLER_211_2623 ();
 FILLCELL_X32 FILLER_211_2655 ();
 FILLCELL_X32 FILLER_211_2687 ();
 FILLCELL_X32 FILLER_211_2719 ();
 FILLCELL_X32 FILLER_211_2751 ();
 FILLCELL_X32 FILLER_211_2783 ();
 FILLCELL_X32 FILLER_211_2815 ();
 FILLCELL_X32 FILLER_211_2847 ();
 FILLCELL_X32 FILLER_211_2879 ();
 FILLCELL_X32 FILLER_211_2911 ();
 FILLCELL_X32 FILLER_211_2943 ();
 FILLCELL_X32 FILLER_211_2975 ();
 FILLCELL_X32 FILLER_211_3007 ();
 FILLCELL_X32 FILLER_211_3039 ();
 FILLCELL_X32 FILLER_211_3071 ();
 FILLCELL_X32 FILLER_211_3103 ();
 FILLCELL_X32 FILLER_211_3135 ();
 FILLCELL_X32 FILLER_211_3167 ();
 FILLCELL_X32 FILLER_211_3199 ();
 FILLCELL_X32 FILLER_211_3231 ();
 FILLCELL_X32 FILLER_211_3263 ();
 FILLCELL_X32 FILLER_211_3295 ();
 FILLCELL_X32 FILLER_211_3327 ();
 FILLCELL_X32 FILLER_211_3359 ();
 FILLCELL_X32 FILLER_211_3391 ();
 FILLCELL_X32 FILLER_211_3423 ();
 FILLCELL_X32 FILLER_211_3455 ();
 FILLCELL_X32 FILLER_211_3487 ();
 FILLCELL_X32 FILLER_211_3519 ();
 FILLCELL_X32 FILLER_211_3551 ();
 FILLCELL_X32 FILLER_211_3583 ();
 FILLCELL_X32 FILLER_211_3615 ();
 FILLCELL_X32 FILLER_211_3647 ();
 FILLCELL_X32 FILLER_211_3679 ();
 FILLCELL_X16 FILLER_211_3711 ();
 FILLCELL_X8 FILLER_211_3727 ();
 FILLCELL_X2 FILLER_211_3735 ();
 FILLCELL_X1 FILLER_211_3737 ();
 FILLCELL_X32 FILLER_212_1 ();
 FILLCELL_X32 FILLER_212_33 ();
 FILLCELL_X32 FILLER_212_65 ();
 FILLCELL_X32 FILLER_212_97 ();
 FILLCELL_X32 FILLER_212_129 ();
 FILLCELL_X32 FILLER_212_161 ();
 FILLCELL_X32 FILLER_212_193 ();
 FILLCELL_X32 FILLER_212_225 ();
 FILLCELL_X32 FILLER_212_257 ();
 FILLCELL_X32 FILLER_212_289 ();
 FILLCELL_X32 FILLER_212_321 ();
 FILLCELL_X32 FILLER_212_353 ();
 FILLCELL_X32 FILLER_212_385 ();
 FILLCELL_X32 FILLER_212_417 ();
 FILLCELL_X32 FILLER_212_449 ();
 FILLCELL_X32 FILLER_212_481 ();
 FILLCELL_X32 FILLER_212_513 ();
 FILLCELL_X32 FILLER_212_545 ();
 FILLCELL_X32 FILLER_212_577 ();
 FILLCELL_X16 FILLER_212_609 ();
 FILLCELL_X4 FILLER_212_625 ();
 FILLCELL_X2 FILLER_212_629 ();
 FILLCELL_X32 FILLER_212_632 ();
 FILLCELL_X32 FILLER_212_664 ();
 FILLCELL_X32 FILLER_212_696 ();
 FILLCELL_X32 FILLER_212_728 ();
 FILLCELL_X32 FILLER_212_760 ();
 FILLCELL_X32 FILLER_212_792 ();
 FILLCELL_X32 FILLER_212_824 ();
 FILLCELL_X32 FILLER_212_856 ();
 FILLCELL_X32 FILLER_212_888 ();
 FILLCELL_X32 FILLER_212_920 ();
 FILLCELL_X32 FILLER_212_952 ();
 FILLCELL_X32 FILLER_212_984 ();
 FILLCELL_X32 FILLER_212_1016 ();
 FILLCELL_X32 FILLER_212_1048 ();
 FILLCELL_X32 FILLER_212_1080 ();
 FILLCELL_X32 FILLER_212_1112 ();
 FILLCELL_X32 FILLER_212_1144 ();
 FILLCELL_X32 FILLER_212_1176 ();
 FILLCELL_X32 FILLER_212_1208 ();
 FILLCELL_X32 FILLER_212_1240 ();
 FILLCELL_X32 FILLER_212_1272 ();
 FILLCELL_X32 FILLER_212_1304 ();
 FILLCELL_X32 FILLER_212_1336 ();
 FILLCELL_X32 FILLER_212_1368 ();
 FILLCELL_X32 FILLER_212_1400 ();
 FILLCELL_X32 FILLER_212_1432 ();
 FILLCELL_X32 FILLER_212_1464 ();
 FILLCELL_X32 FILLER_212_1496 ();
 FILLCELL_X32 FILLER_212_1528 ();
 FILLCELL_X32 FILLER_212_1560 ();
 FILLCELL_X32 FILLER_212_1592 ();
 FILLCELL_X32 FILLER_212_1624 ();
 FILLCELL_X32 FILLER_212_1656 ();
 FILLCELL_X32 FILLER_212_1688 ();
 FILLCELL_X32 FILLER_212_1720 ();
 FILLCELL_X32 FILLER_212_1752 ();
 FILLCELL_X32 FILLER_212_1784 ();
 FILLCELL_X32 FILLER_212_1816 ();
 FILLCELL_X32 FILLER_212_1848 ();
 FILLCELL_X8 FILLER_212_1880 ();
 FILLCELL_X4 FILLER_212_1888 ();
 FILLCELL_X2 FILLER_212_1892 ();
 FILLCELL_X16 FILLER_212_1895 ();
 FILLCELL_X8 FILLER_212_1911 ();
 FILLCELL_X2 FILLER_212_1919 ();
 FILLCELL_X1 FILLER_212_1921 ();
 FILLCELL_X32 FILLER_212_1926 ();
 FILLCELL_X32 FILLER_212_1958 ();
 FILLCELL_X32 FILLER_212_1990 ();
 FILLCELL_X32 FILLER_212_2022 ();
 FILLCELL_X32 FILLER_212_2054 ();
 FILLCELL_X32 FILLER_212_2086 ();
 FILLCELL_X32 FILLER_212_2118 ();
 FILLCELL_X32 FILLER_212_2150 ();
 FILLCELL_X32 FILLER_212_2182 ();
 FILLCELL_X32 FILLER_212_2214 ();
 FILLCELL_X32 FILLER_212_2246 ();
 FILLCELL_X32 FILLER_212_2278 ();
 FILLCELL_X32 FILLER_212_2310 ();
 FILLCELL_X32 FILLER_212_2342 ();
 FILLCELL_X32 FILLER_212_2374 ();
 FILLCELL_X32 FILLER_212_2406 ();
 FILLCELL_X32 FILLER_212_2438 ();
 FILLCELL_X32 FILLER_212_2470 ();
 FILLCELL_X32 FILLER_212_2502 ();
 FILLCELL_X32 FILLER_212_2534 ();
 FILLCELL_X32 FILLER_212_2566 ();
 FILLCELL_X32 FILLER_212_2598 ();
 FILLCELL_X32 FILLER_212_2630 ();
 FILLCELL_X32 FILLER_212_2662 ();
 FILLCELL_X32 FILLER_212_2694 ();
 FILLCELL_X32 FILLER_212_2726 ();
 FILLCELL_X32 FILLER_212_2758 ();
 FILLCELL_X32 FILLER_212_2790 ();
 FILLCELL_X32 FILLER_212_2822 ();
 FILLCELL_X32 FILLER_212_2854 ();
 FILLCELL_X32 FILLER_212_2886 ();
 FILLCELL_X32 FILLER_212_2918 ();
 FILLCELL_X32 FILLER_212_2950 ();
 FILLCELL_X32 FILLER_212_2982 ();
 FILLCELL_X32 FILLER_212_3014 ();
 FILLCELL_X32 FILLER_212_3046 ();
 FILLCELL_X32 FILLER_212_3078 ();
 FILLCELL_X32 FILLER_212_3110 ();
 FILLCELL_X8 FILLER_212_3142 ();
 FILLCELL_X4 FILLER_212_3150 ();
 FILLCELL_X2 FILLER_212_3154 ();
 FILLCELL_X1 FILLER_212_3156 ();
 FILLCELL_X32 FILLER_212_3158 ();
 FILLCELL_X32 FILLER_212_3190 ();
 FILLCELL_X32 FILLER_212_3222 ();
 FILLCELL_X32 FILLER_212_3254 ();
 FILLCELL_X32 FILLER_212_3286 ();
 FILLCELL_X32 FILLER_212_3318 ();
 FILLCELL_X32 FILLER_212_3350 ();
 FILLCELL_X32 FILLER_212_3382 ();
 FILLCELL_X32 FILLER_212_3414 ();
 FILLCELL_X32 FILLER_212_3446 ();
 FILLCELL_X32 FILLER_212_3478 ();
 FILLCELL_X32 FILLER_212_3510 ();
 FILLCELL_X32 FILLER_212_3542 ();
 FILLCELL_X32 FILLER_212_3574 ();
 FILLCELL_X32 FILLER_212_3606 ();
 FILLCELL_X32 FILLER_212_3638 ();
 FILLCELL_X32 FILLER_212_3670 ();
 FILLCELL_X32 FILLER_212_3702 ();
 FILLCELL_X4 FILLER_212_3734 ();
 FILLCELL_X32 FILLER_213_1 ();
 FILLCELL_X32 FILLER_213_33 ();
 FILLCELL_X32 FILLER_213_65 ();
 FILLCELL_X32 FILLER_213_97 ();
 FILLCELL_X32 FILLER_213_129 ();
 FILLCELL_X32 FILLER_213_161 ();
 FILLCELL_X32 FILLER_213_193 ();
 FILLCELL_X32 FILLER_213_225 ();
 FILLCELL_X32 FILLER_213_257 ();
 FILLCELL_X32 FILLER_213_289 ();
 FILLCELL_X32 FILLER_213_321 ();
 FILLCELL_X32 FILLER_213_353 ();
 FILLCELL_X32 FILLER_213_385 ();
 FILLCELL_X32 FILLER_213_417 ();
 FILLCELL_X32 FILLER_213_449 ();
 FILLCELL_X32 FILLER_213_481 ();
 FILLCELL_X32 FILLER_213_513 ();
 FILLCELL_X32 FILLER_213_545 ();
 FILLCELL_X32 FILLER_213_577 ();
 FILLCELL_X32 FILLER_213_609 ();
 FILLCELL_X32 FILLER_213_641 ();
 FILLCELL_X32 FILLER_213_673 ();
 FILLCELL_X32 FILLER_213_705 ();
 FILLCELL_X32 FILLER_213_737 ();
 FILLCELL_X32 FILLER_213_769 ();
 FILLCELL_X32 FILLER_213_801 ();
 FILLCELL_X32 FILLER_213_833 ();
 FILLCELL_X32 FILLER_213_865 ();
 FILLCELL_X32 FILLER_213_897 ();
 FILLCELL_X32 FILLER_213_929 ();
 FILLCELL_X32 FILLER_213_961 ();
 FILLCELL_X32 FILLER_213_993 ();
 FILLCELL_X32 FILLER_213_1025 ();
 FILLCELL_X32 FILLER_213_1057 ();
 FILLCELL_X32 FILLER_213_1089 ();
 FILLCELL_X32 FILLER_213_1121 ();
 FILLCELL_X32 FILLER_213_1153 ();
 FILLCELL_X32 FILLER_213_1185 ();
 FILLCELL_X32 FILLER_213_1217 ();
 FILLCELL_X8 FILLER_213_1249 ();
 FILLCELL_X4 FILLER_213_1257 ();
 FILLCELL_X2 FILLER_213_1261 ();
 FILLCELL_X32 FILLER_213_1264 ();
 FILLCELL_X32 FILLER_213_1296 ();
 FILLCELL_X32 FILLER_213_1328 ();
 FILLCELL_X32 FILLER_213_1360 ();
 FILLCELL_X32 FILLER_213_1392 ();
 FILLCELL_X32 FILLER_213_1424 ();
 FILLCELL_X32 FILLER_213_1456 ();
 FILLCELL_X32 FILLER_213_1488 ();
 FILLCELL_X32 FILLER_213_1520 ();
 FILLCELL_X32 FILLER_213_1552 ();
 FILLCELL_X32 FILLER_213_1584 ();
 FILLCELL_X32 FILLER_213_1616 ();
 FILLCELL_X32 FILLER_213_1648 ();
 FILLCELL_X32 FILLER_213_1680 ();
 FILLCELL_X32 FILLER_213_1712 ();
 FILLCELL_X32 FILLER_213_1744 ();
 FILLCELL_X32 FILLER_213_1776 ();
 FILLCELL_X32 FILLER_213_1808 ();
 FILLCELL_X32 FILLER_213_1840 ();
 FILLCELL_X32 FILLER_213_1872 ();
 FILLCELL_X32 FILLER_213_1904 ();
 FILLCELL_X32 FILLER_213_1936 ();
 FILLCELL_X32 FILLER_213_1968 ();
 FILLCELL_X32 FILLER_213_2000 ();
 FILLCELL_X32 FILLER_213_2032 ();
 FILLCELL_X32 FILLER_213_2064 ();
 FILLCELL_X32 FILLER_213_2096 ();
 FILLCELL_X32 FILLER_213_2128 ();
 FILLCELL_X32 FILLER_213_2160 ();
 FILLCELL_X32 FILLER_213_2192 ();
 FILLCELL_X32 FILLER_213_2224 ();
 FILLCELL_X32 FILLER_213_2256 ();
 FILLCELL_X32 FILLER_213_2288 ();
 FILLCELL_X32 FILLER_213_2320 ();
 FILLCELL_X32 FILLER_213_2352 ();
 FILLCELL_X32 FILLER_213_2384 ();
 FILLCELL_X32 FILLER_213_2416 ();
 FILLCELL_X32 FILLER_213_2448 ();
 FILLCELL_X32 FILLER_213_2480 ();
 FILLCELL_X8 FILLER_213_2512 ();
 FILLCELL_X4 FILLER_213_2520 ();
 FILLCELL_X2 FILLER_213_2524 ();
 FILLCELL_X32 FILLER_213_2527 ();
 FILLCELL_X32 FILLER_213_2559 ();
 FILLCELL_X32 FILLER_213_2591 ();
 FILLCELL_X32 FILLER_213_2623 ();
 FILLCELL_X32 FILLER_213_2655 ();
 FILLCELL_X32 FILLER_213_2687 ();
 FILLCELL_X32 FILLER_213_2719 ();
 FILLCELL_X32 FILLER_213_2751 ();
 FILLCELL_X32 FILLER_213_2783 ();
 FILLCELL_X32 FILLER_213_2815 ();
 FILLCELL_X32 FILLER_213_2847 ();
 FILLCELL_X32 FILLER_213_2879 ();
 FILLCELL_X32 FILLER_213_2911 ();
 FILLCELL_X32 FILLER_213_2943 ();
 FILLCELL_X32 FILLER_213_2975 ();
 FILLCELL_X32 FILLER_213_3007 ();
 FILLCELL_X32 FILLER_213_3039 ();
 FILLCELL_X32 FILLER_213_3071 ();
 FILLCELL_X32 FILLER_213_3103 ();
 FILLCELL_X32 FILLER_213_3135 ();
 FILLCELL_X32 FILLER_213_3167 ();
 FILLCELL_X32 FILLER_213_3199 ();
 FILLCELL_X32 FILLER_213_3231 ();
 FILLCELL_X32 FILLER_213_3263 ();
 FILLCELL_X32 FILLER_213_3295 ();
 FILLCELL_X32 FILLER_213_3327 ();
 FILLCELL_X32 FILLER_213_3359 ();
 FILLCELL_X32 FILLER_213_3391 ();
 FILLCELL_X32 FILLER_213_3423 ();
 FILLCELL_X32 FILLER_213_3455 ();
 FILLCELL_X32 FILLER_213_3487 ();
 FILLCELL_X32 FILLER_213_3519 ();
 FILLCELL_X32 FILLER_213_3551 ();
 FILLCELL_X32 FILLER_213_3583 ();
 FILLCELL_X32 FILLER_213_3615 ();
 FILLCELL_X32 FILLER_213_3647 ();
 FILLCELL_X32 FILLER_213_3679 ();
 FILLCELL_X16 FILLER_213_3711 ();
 FILLCELL_X8 FILLER_213_3727 ();
 FILLCELL_X2 FILLER_213_3735 ();
 FILLCELL_X1 FILLER_213_3737 ();
 FILLCELL_X32 FILLER_214_1 ();
 FILLCELL_X32 FILLER_214_33 ();
 FILLCELL_X32 FILLER_214_65 ();
 FILLCELL_X32 FILLER_214_97 ();
 FILLCELL_X32 FILLER_214_129 ();
 FILLCELL_X32 FILLER_214_161 ();
 FILLCELL_X32 FILLER_214_193 ();
 FILLCELL_X32 FILLER_214_225 ();
 FILLCELL_X32 FILLER_214_257 ();
 FILLCELL_X32 FILLER_214_289 ();
 FILLCELL_X32 FILLER_214_321 ();
 FILLCELL_X32 FILLER_214_353 ();
 FILLCELL_X32 FILLER_214_385 ();
 FILLCELL_X32 FILLER_214_417 ();
 FILLCELL_X32 FILLER_214_449 ();
 FILLCELL_X32 FILLER_214_481 ();
 FILLCELL_X32 FILLER_214_513 ();
 FILLCELL_X32 FILLER_214_545 ();
 FILLCELL_X32 FILLER_214_577 ();
 FILLCELL_X16 FILLER_214_609 ();
 FILLCELL_X4 FILLER_214_625 ();
 FILLCELL_X2 FILLER_214_629 ();
 FILLCELL_X32 FILLER_214_632 ();
 FILLCELL_X32 FILLER_214_664 ();
 FILLCELL_X32 FILLER_214_696 ();
 FILLCELL_X32 FILLER_214_728 ();
 FILLCELL_X32 FILLER_214_760 ();
 FILLCELL_X32 FILLER_214_792 ();
 FILLCELL_X32 FILLER_214_824 ();
 FILLCELL_X32 FILLER_214_856 ();
 FILLCELL_X32 FILLER_214_888 ();
 FILLCELL_X32 FILLER_214_920 ();
 FILLCELL_X32 FILLER_214_952 ();
 FILLCELL_X32 FILLER_214_984 ();
 FILLCELL_X32 FILLER_214_1016 ();
 FILLCELL_X32 FILLER_214_1048 ();
 FILLCELL_X32 FILLER_214_1080 ();
 FILLCELL_X32 FILLER_214_1112 ();
 FILLCELL_X32 FILLER_214_1144 ();
 FILLCELL_X32 FILLER_214_1176 ();
 FILLCELL_X32 FILLER_214_1208 ();
 FILLCELL_X32 FILLER_214_1240 ();
 FILLCELL_X32 FILLER_214_1272 ();
 FILLCELL_X32 FILLER_214_1304 ();
 FILLCELL_X32 FILLER_214_1336 ();
 FILLCELL_X32 FILLER_214_1368 ();
 FILLCELL_X32 FILLER_214_1400 ();
 FILLCELL_X32 FILLER_214_1432 ();
 FILLCELL_X32 FILLER_214_1464 ();
 FILLCELL_X32 FILLER_214_1496 ();
 FILLCELL_X32 FILLER_214_1528 ();
 FILLCELL_X32 FILLER_214_1560 ();
 FILLCELL_X32 FILLER_214_1592 ();
 FILLCELL_X32 FILLER_214_1624 ();
 FILLCELL_X32 FILLER_214_1656 ();
 FILLCELL_X32 FILLER_214_1688 ();
 FILLCELL_X32 FILLER_214_1720 ();
 FILLCELL_X32 FILLER_214_1752 ();
 FILLCELL_X32 FILLER_214_1784 ();
 FILLCELL_X32 FILLER_214_1816 ();
 FILLCELL_X32 FILLER_214_1848 ();
 FILLCELL_X8 FILLER_214_1880 ();
 FILLCELL_X4 FILLER_214_1888 ();
 FILLCELL_X2 FILLER_214_1892 ();
 FILLCELL_X32 FILLER_214_1895 ();
 FILLCELL_X32 FILLER_214_1927 ();
 FILLCELL_X32 FILLER_214_1959 ();
 FILLCELL_X32 FILLER_214_1991 ();
 FILLCELL_X32 FILLER_214_2023 ();
 FILLCELL_X32 FILLER_214_2055 ();
 FILLCELL_X32 FILLER_214_2087 ();
 FILLCELL_X32 FILLER_214_2119 ();
 FILLCELL_X32 FILLER_214_2151 ();
 FILLCELL_X32 FILLER_214_2183 ();
 FILLCELL_X32 FILLER_214_2215 ();
 FILLCELL_X32 FILLER_214_2247 ();
 FILLCELL_X32 FILLER_214_2279 ();
 FILLCELL_X32 FILLER_214_2311 ();
 FILLCELL_X32 FILLER_214_2343 ();
 FILLCELL_X32 FILLER_214_2375 ();
 FILLCELL_X32 FILLER_214_2407 ();
 FILLCELL_X32 FILLER_214_2439 ();
 FILLCELL_X32 FILLER_214_2471 ();
 FILLCELL_X32 FILLER_214_2503 ();
 FILLCELL_X32 FILLER_214_2535 ();
 FILLCELL_X32 FILLER_214_2567 ();
 FILLCELL_X32 FILLER_214_2599 ();
 FILLCELL_X32 FILLER_214_2631 ();
 FILLCELL_X32 FILLER_214_2663 ();
 FILLCELL_X32 FILLER_214_2695 ();
 FILLCELL_X32 FILLER_214_2727 ();
 FILLCELL_X32 FILLER_214_2759 ();
 FILLCELL_X32 FILLER_214_2791 ();
 FILLCELL_X32 FILLER_214_2823 ();
 FILLCELL_X32 FILLER_214_2855 ();
 FILLCELL_X32 FILLER_214_2887 ();
 FILLCELL_X32 FILLER_214_2919 ();
 FILLCELL_X32 FILLER_214_2951 ();
 FILLCELL_X32 FILLER_214_2983 ();
 FILLCELL_X32 FILLER_214_3015 ();
 FILLCELL_X32 FILLER_214_3047 ();
 FILLCELL_X32 FILLER_214_3079 ();
 FILLCELL_X32 FILLER_214_3111 ();
 FILLCELL_X8 FILLER_214_3143 ();
 FILLCELL_X4 FILLER_214_3151 ();
 FILLCELL_X2 FILLER_214_3155 ();
 FILLCELL_X32 FILLER_214_3158 ();
 FILLCELL_X32 FILLER_214_3190 ();
 FILLCELL_X32 FILLER_214_3222 ();
 FILLCELL_X32 FILLER_214_3254 ();
 FILLCELL_X32 FILLER_214_3286 ();
 FILLCELL_X32 FILLER_214_3318 ();
 FILLCELL_X32 FILLER_214_3350 ();
 FILLCELL_X32 FILLER_214_3382 ();
 FILLCELL_X32 FILLER_214_3414 ();
 FILLCELL_X32 FILLER_214_3446 ();
 FILLCELL_X32 FILLER_214_3478 ();
 FILLCELL_X32 FILLER_214_3510 ();
 FILLCELL_X32 FILLER_214_3542 ();
 FILLCELL_X32 FILLER_214_3574 ();
 FILLCELL_X32 FILLER_214_3606 ();
 FILLCELL_X32 FILLER_214_3638 ();
 FILLCELL_X32 FILLER_214_3670 ();
 FILLCELL_X32 FILLER_214_3702 ();
 FILLCELL_X4 FILLER_214_3734 ();
 FILLCELL_X32 FILLER_215_1 ();
 FILLCELL_X32 FILLER_215_33 ();
 FILLCELL_X32 FILLER_215_65 ();
 FILLCELL_X32 FILLER_215_97 ();
 FILLCELL_X32 FILLER_215_129 ();
 FILLCELL_X32 FILLER_215_161 ();
 FILLCELL_X32 FILLER_215_193 ();
 FILLCELL_X32 FILLER_215_225 ();
 FILLCELL_X32 FILLER_215_257 ();
 FILLCELL_X32 FILLER_215_289 ();
 FILLCELL_X32 FILLER_215_321 ();
 FILLCELL_X32 FILLER_215_353 ();
 FILLCELL_X32 FILLER_215_385 ();
 FILLCELL_X32 FILLER_215_417 ();
 FILLCELL_X32 FILLER_215_449 ();
 FILLCELL_X32 FILLER_215_481 ();
 FILLCELL_X32 FILLER_215_513 ();
 FILLCELL_X32 FILLER_215_545 ();
 FILLCELL_X32 FILLER_215_577 ();
 FILLCELL_X32 FILLER_215_609 ();
 FILLCELL_X32 FILLER_215_641 ();
 FILLCELL_X32 FILLER_215_673 ();
 FILLCELL_X32 FILLER_215_705 ();
 FILLCELL_X32 FILLER_215_737 ();
 FILLCELL_X32 FILLER_215_769 ();
 FILLCELL_X32 FILLER_215_801 ();
 FILLCELL_X32 FILLER_215_833 ();
 FILLCELL_X32 FILLER_215_865 ();
 FILLCELL_X32 FILLER_215_897 ();
 FILLCELL_X32 FILLER_215_929 ();
 FILLCELL_X32 FILLER_215_961 ();
 FILLCELL_X32 FILLER_215_993 ();
 FILLCELL_X32 FILLER_215_1025 ();
 FILLCELL_X32 FILLER_215_1057 ();
 FILLCELL_X32 FILLER_215_1089 ();
 FILLCELL_X32 FILLER_215_1121 ();
 FILLCELL_X32 FILLER_215_1153 ();
 FILLCELL_X32 FILLER_215_1185 ();
 FILLCELL_X32 FILLER_215_1217 ();
 FILLCELL_X8 FILLER_215_1249 ();
 FILLCELL_X4 FILLER_215_1257 ();
 FILLCELL_X2 FILLER_215_1261 ();
 FILLCELL_X32 FILLER_215_1264 ();
 FILLCELL_X32 FILLER_215_1296 ();
 FILLCELL_X32 FILLER_215_1328 ();
 FILLCELL_X32 FILLER_215_1360 ();
 FILLCELL_X32 FILLER_215_1392 ();
 FILLCELL_X32 FILLER_215_1424 ();
 FILLCELL_X32 FILLER_215_1456 ();
 FILLCELL_X32 FILLER_215_1488 ();
 FILLCELL_X32 FILLER_215_1520 ();
 FILLCELL_X32 FILLER_215_1552 ();
 FILLCELL_X32 FILLER_215_1584 ();
 FILLCELL_X32 FILLER_215_1616 ();
 FILLCELL_X32 FILLER_215_1648 ();
 FILLCELL_X32 FILLER_215_1680 ();
 FILLCELL_X32 FILLER_215_1712 ();
 FILLCELL_X32 FILLER_215_1744 ();
 FILLCELL_X32 FILLER_215_1776 ();
 FILLCELL_X32 FILLER_215_1808 ();
 FILLCELL_X32 FILLER_215_1840 ();
 FILLCELL_X32 FILLER_215_1872 ();
 FILLCELL_X32 FILLER_215_1904 ();
 FILLCELL_X32 FILLER_215_1936 ();
 FILLCELL_X32 FILLER_215_1968 ();
 FILLCELL_X32 FILLER_215_2000 ();
 FILLCELL_X32 FILLER_215_2032 ();
 FILLCELL_X32 FILLER_215_2064 ();
 FILLCELL_X32 FILLER_215_2096 ();
 FILLCELL_X32 FILLER_215_2128 ();
 FILLCELL_X32 FILLER_215_2160 ();
 FILLCELL_X32 FILLER_215_2192 ();
 FILLCELL_X32 FILLER_215_2224 ();
 FILLCELL_X32 FILLER_215_2256 ();
 FILLCELL_X32 FILLER_215_2288 ();
 FILLCELL_X32 FILLER_215_2320 ();
 FILLCELL_X32 FILLER_215_2352 ();
 FILLCELL_X32 FILLER_215_2384 ();
 FILLCELL_X32 FILLER_215_2416 ();
 FILLCELL_X32 FILLER_215_2448 ();
 FILLCELL_X32 FILLER_215_2480 ();
 FILLCELL_X8 FILLER_215_2512 ();
 FILLCELL_X4 FILLER_215_2520 ();
 FILLCELL_X2 FILLER_215_2524 ();
 FILLCELL_X32 FILLER_215_2527 ();
 FILLCELL_X32 FILLER_215_2559 ();
 FILLCELL_X32 FILLER_215_2591 ();
 FILLCELL_X32 FILLER_215_2623 ();
 FILLCELL_X32 FILLER_215_2655 ();
 FILLCELL_X32 FILLER_215_2687 ();
 FILLCELL_X32 FILLER_215_2719 ();
 FILLCELL_X32 FILLER_215_2751 ();
 FILLCELL_X32 FILLER_215_2783 ();
 FILLCELL_X32 FILLER_215_2815 ();
 FILLCELL_X32 FILLER_215_2847 ();
 FILLCELL_X32 FILLER_215_2879 ();
 FILLCELL_X32 FILLER_215_2911 ();
 FILLCELL_X32 FILLER_215_2943 ();
 FILLCELL_X32 FILLER_215_2975 ();
 FILLCELL_X32 FILLER_215_3007 ();
 FILLCELL_X32 FILLER_215_3039 ();
 FILLCELL_X32 FILLER_215_3071 ();
 FILLCELL_X32 FILLER_215_3103 ();
 FILLCELL_X32 FILLER_215_3135 ();
 FILLCELL_X32 FILLER_215_3167 ();
 FILLCELL_X32 FILLER_215_3199 ();
 FILLCELL_X32 FILLER_215_3231 ();
 FILLCELL_X32 FILLER_215_3263 ();
 FILLCELL_X32 FILLER_215_3295 ();
 FILLCELL_X32 FILLER_215_3327 ();
 FILLCELL_X32 FILLER_215_3359 ();
 FILLCELL_X32 FILLER_215_3391 ();
 FILLCELL_X32 FILLER_215_3423 ();
 FILLCELL_X32 FILLER_215_3455 ();
 FILLCELL_X32 FILLER_215_3487 ();
 FILLCELL_X32 FILLER_215_3519 ();
 FILLCELL_X32 FILLER_215_3551 ();
 FILLCELL_X32 FILLER_215_3583 ();
 FILLCELL_X32 FILLER_215_3615 ();
 FILLCELL_X32 FILLER_215_3647 ();
 FILLCELL_X32 FILLER_215_3679 ();
 FILLCELL_X16 FILLER_215_3711 ();
 FILLCELL_X8 FILLER_215_3727 ();
 FILLCELL_X2 FILLER_215_3735 ();
 FILLCELL_X1 FILLER_215_3737 ();
 FILLCELL_X32 FILLER_216_1 ();
 FILLCELL_X32 FILLER_216_33 ();
 FILLCELL_X32 FILLER_216_65 ();
 FILLCELL_X32 FILLER_216_97 ();
 FILLCELL_X32 FILLER_216_129 ();
 FILLCELL_X32 FILLER_216_161 ();
 FILLCELL_X32 FILLER_216_193 ();
 FILLCELL_X32 FILLER_216_225 ();
 FILLCELL_X32 FILLER_216_257 ();
 FILLCELL_X32 FILLER_216_289 ();
 FILLCELL_X32 FILLER_216_321 ();
 FILLCELL_X32 FILLER_216_353 ();
 FILLCELL_X32 FILLER_216_385 ();
 FILLCELL_X32 FILLER_216_417 ();
 FILLCELL_X32 FILLER_216_449 ();
 FILLCELL_X32 FILLER_216_481 ();
 FILLCELL_X32 FILLER_216_513 ();
 FILLCELL_X32 FILLER_216_545 ();
 FILLCELL_X32 FILLER_216_577 ();
 FILLCELL_X16 FILLER_216_609 ();
 FILLCELL_X4 FILLER_216_625 ();
 FILLCELL_X2 FILLER_216_629 ();
 FILLCELL_X32 FILLER_216_632 ();
 FILLCELL_X32 FILLER_216_664 ();
 FILLCELL_X32 FILLER_216_696 ();
 FILLCELL_X32 FILLER_216_728 ();
 FILLCELL_X32 FILLER_216_760 ();
 FILLCELL_X32 FILLER_216_792 ();
 FILLCELL_X32 FILLER_216_824 ();
 FILLCELL_X32 FILLER_216_856 ();
 FILLCELL_X32 FILLER_216_888 ();
 FILLCELL_X32 FILLER_216_920 ();
 FILLCELL_X32 FILLER_216_952 ();
 FILLCELL_X32 FILLER_216_984 ();
 FILLCELL_X32 FILLER_216_1016 ();
 FILLCELL_X32 FILLER_216_1048 ();
 FILLCELL_X32 FILLER_216_1080 ();
 FILLCELL_X32 FILLER_216_1112 ();
 FILLCELL_X32 FILLER_216_1144 ();
 FILLCELL_X32 FILLER_216_1176 ();
 FILLCELL_X32 FILLER_216_1208 ();
 FILLCELL_X32 FILLER_216_1240 ();
 FILLCELL_X32 FILLER_216_1272 ();
 FILLCELL_X32 FILLER_216_1304 ();
 FILLCELL_X32 FILLER_216_1336 ();
 FILLCELL_X32 FILLER_216_1368 ();
 FILLCELL_X32 FILLER_216_1400 ();
 FILLCELL_X32 FILLER_216_1432 ();
 FILLCELL_X32 FILLER_216_1464 ();
 FILLCELL_X32 FILLER_216_1496 ();
 FILLCELL_X32 FILLER_216_1528 ();
 FILLCELL_X32 FILLER_216_1560 ();
 FILLCELL_X32 FILLER_216_1592 ();
 FILLCELL_X32 FILLER_216_1624 ();
 FILLCELL_X32 FILLER_216_1656 ();
 FILLCELL_X32 FILLER_216_1688 ();
 FILLCELL_X32 FILLER_216_1720 ();
 FILLCELL_X32 FILLER_216_1752 ();
 FILLCELL_X32 FILLER_216_1784 ();
 FILLCELL_X32 FILLER_216_1816 ();
 FILLCELL_X32 FILLER_216_1848 ();
 FILLCELL_X8 FILLER_216_1880 ();
 FILLCELL_X4 FILLER_216_1888 ();
 FILLCELL_X2 FILLER_216_1892 ();
 FILLCELL_X32 FILLER_216_1895 ();
 FILLCELL_X32 FILLER_216_1927 ();
 FILLCELL_X32 FILLER_216_1959 ();
 FILLCELL_X32 FILLER_216_1991 ();
 FILLCELL_X32 FILLER_216_2023 ();
 FILLCELL_X32 FILLER_216_2055 ();
 FILLCELL_X32 FILLER_216_2087 ();
 FILLCELL_X32 FILLER_216_2119 ();
 FILLCELL_X32 FILLER_216_2151 ();
 FILLCELL_X32 FILLER_216_2183 ();
 FILLCELL_X32 FILLER_216_2215 ();
 FILLCELL_X32 FILLER_216_2247 ();
 FILLCELL_X32 FILLER_216_2279 ();
 FILLCELL_X32 FILLER_216_2311 ();
 FILLCELL_X32 FILLER_216_2343 ();
 FILLCELL_X32 FILLER_216_2375 ();
 FILLCELL_X32 FILLER_216_2407 ();
 FILLCELL_X32 FILLER_216_2439 ();
 FILLCELL_X32 FILLER_216_2471 ();
 FILLCELL_X32 FILLER_216_2503 ();
 FILLCELL_X32 FILLER_216_2535 ();
 FILLCELL_X32 FILLER_216_2567 ();
 FILLCELL_X32 FILLER_216_2599 ();
 FILLCELL_X32 FILLER_216_2631 ();
 FILLCELL_X32 FILLER_216_2663 ();
 FILLCELL_X32 FILLER_216_2695 ();
 FILLCELL_X32 FILLER_216_2727 ();
 FILLCELL_X32 FILLER_216_2759 ();
 FILLCELL_X32 FILLER_216_2791 ();
 FILLCELL_X32 FILLER_216_2823 ();
 FILLCELL_X32 FILLER_216_2855 ();
 FILLCELL_X32 FILLER_216_2887 ();
 FILLCELL_X32 FILLER_216_2919 ();
 FILLCELL_X32 FILLER_216_2951 ();
 FILLCELL_X32 FILLER_216_2983 ();
 FILLCELL_X32 FILLER_216_3015 ();
 FILLCELL_X32 FILLER_216_3047 ();
 FILLCELL_X32 FILLER_216_3079 ();
 FILLCELL_X32 FILLER_216_3111 ();
 FILLCELL_X8 FILLER_216_3143 ();
 FILLCELL_X4 FILLER_216_3151 ();
 FILLCELL_X2 FILLER_216_3155 ();
 FILLCELL_X32 FILLER_216_3158 ();
 FILLCELL_X32 FILLER_216_3190 ();
 FILLCELL_X32 FILLER_216_3222 ();
 FILLCELL_X32 FILLER_216_3254 ();
 FILLCELL_X32 FILLER_216_3286 ();
 FILLCELL_X32 FILLER_216_3318 ();
 FILLCELL_X32 FILLER_216_3350 ();
 FILLCELL_X32 FILLER_216_3382 ();
 FILLCELL_X32 FILLER_216_3414 ();
 FILLCELL_X32 FILLER_216_3446 ();
 FILLCELL_X32 FILLER_216_3478 ();
 FILLCELL_X32 FILLER_216_3510 ();
 FILLCELL_X32 FILLER_216_3542 ();
 FILLCELL_X32 FILLER_216_3574 ();
 FILLCELL_X32 FILLER_216_3606 ();
 FILLCELL_X32 FILLER_216_3638 ();
 FILLCELL_X32 FILLER_216_3670 ();
 FILLCELL_X32 FILLER_216_3702 ();
 FILLCELL_X4 FILLER_216_3734 ();
 FILLCELL_X32 FILLER_217_1 ();
 FILLCELL_X32 FILLER_217_33 ();
 FILLCELL_X32 FILLER_217_65 ();
 FILLCELL_X32 FILLER_217_97 ();
 FILLCELL_X32 FILLER_217_129 ();
 FILLCELL_X32 FILLER_217_161 ();
 FILLCELL_X32 FILLER_217_193 ();
 FILLCELL_X32 FILLER_217_225 ();
 FILLCELL_X32 FILLER_217_257 ();
 FILLCELL_X32 FILLER_217_289 ();
 FILLCELL_X32 FILLER_217_321 ();
 FILLCELL_X32 FILLER_217_353 ();
 FILLCELL_X32 FILLER_217_385 ();
 FILLCELL_X32 FILLER_217_417 ();
 FILLCELL_X32 FILLER_217_449 ();
 FILLCELL_X32 FILLER_217_481 ();
 FILLCELL_X32 FILLER_217_513 ();
 FILLCELL_X32 FILLER_217_545 ();
 FILLCELL_X32 FILLER_217_577 ();
 FILLCELL_X32 FILLER_217_609 ();
 FILLCELL_X32 FILLER_217_641 ();
 FILLCELL_X32 FILLER_217_673 ();
 FILLCELL_X32 FILLER_217_705 ();
 FILLCELL_X32 FILLER_217_737 ();
 FILLCELL_X32 FILLER_217_769 ();
 FILLCELL_X32 FILLER_217_801 ();
 FILLCELL_X32 FILLER_217_833 ();
 FILLCELL_X32 FILLER_217_865 ();
 FILLCELL_X32 FILLER_217_897 ();
 FILLCELL_X32 FILLER_217_929 ();
 FILLCELL_X32 FILLER_217_961 ();
 FILLCELL_X32 FILLER_217_993 ();
 FILLCELL_X32 FILLER_217_1025 ();
 FILLCELL_X32 FILLER_217_1057 ();
 FILLCELL_X32 FILLER_217_1089 ();
 FILLCELL_X32 FILLER_217_1121 ();
 FILLCELL_X32 FILLER_217_1153 ();
 FILLCELL_X32 FILLER_217_1185 ();
 FILLCELL_X32 FILLER_217_1217 ();
 FILLCELL_X8 FILLER_217_1249 ();
 FILLCELL_X4 FILLER_217_1257 ();
 FILLCELL_X2 FILLER_217_1261 ();
 FILLCELL_X32 FILLER_217_1264 ();
 FILLCELL_X32 FILLER_217_1296 ();
 FILLCELL_X32 FILLER_217_1328 ();
 FILLCELL_X32 FILLER_217_1360 ();
 FILLCELL_X32 FILLER_217_1392 ();
 FILLCELL_X32 FILLER_217_1424 ();
 FILLCELL_X32 FILLER_217_1456 ();
 FILLCELL_X32 FILLER_217_1488 ();
 FILLCELL_X32 FILLER_217_1520 ();
 FILLCELL_X32 FILLER_217_1552 ();
 FILLCELL_X32 FILLER_217_1584 ();
 FILLCELL_X32 FILLER_217_1616 ();
 FILLCELL_X32 FILLER_217_1648 ();
 FILLCELL_X32 FILLER_217_1680 ();
 FILLCELL_X32 FILLER_217_1712 ();
 FILLCELL_X32 FILLER_217_1744 ();
 FILLCELL_X32 FILLER_217_1776 ();
 FILLCELL_X32 FILLER_217_1808 ();
 FILLCELL_X32 FILLER_217_1840 ();
 FILLCELL_X32 FILLER_217_1872 ();
 FILLCELL_X32 FILLER_217_1904 ();
 FILLCELL_X32 FILLER_217_1936 ();
 FILLCELL_X32 FILLER_217_1968 ();
 FILLCELL_X32 FILLER_217_2000 ();
 FILLCELL_X32 FILLER_217_2032 ();
 FILLCELL_X32 FILLER_217_2064 ();
 FILLCELL_X32 FILLER_217_2096 ();
 FILLCELL_X32 FILLER_217_2128 ();
 FILLCELL_X32 FILLER_217_2160 ();
 FILLCELL_X32 FILLER_217_2192 ();
 FILLCELL_X32 FILLER_217_2224 ();
 FILLCELL_X32 FILLER_217_2256 ();
 FILLCELL_X32 FILLER_217_2288 ();
 FILLCELL_X32 FILLER_217_2320 ();
 FILLCELL_X32 FILLER_217_2352 ();
 FILLCELL_X32 FILLER_217_2384 ();
 FILLCELL_X32 FILLER_217_2416 ();
 FILLCELL_X32 FILLER_217_2448 ();
 FILLCELL_X32 FILLER_217_2480 ();
 FILLCELL_X8 FILLER_217_2512 ();
 FILLCELL_X4 FILLER_217_2520 ();
 FILLCELL_X2 FILLER_217_2524 ();
 FILLCELL_X32 FILLER_217_2527 ();
 FILLCELL_X32 FILLER_217_2559 ();
 FILLCELL_X32 FILLER_217_2591 ();
 FILLCELL_X32 FILLER_217_2623 ();
 FILLCELL_X32 FILLER_217_2655 ();
 FILLCELL_X32 FILLER_217_2687 ();
 FILLCELL_X32 FILLER_217_2719 ();
 FILLCELL_X32 FILLER_217_2751 ();
 FILLCELL_X32 FILLER_217_2783 ();
 FILLCELL_X32 FILLER_217_2815 ();
 FILLCELL_X32 FILLER_217_2847 ();
 FILLCELL_X32 FILLER_217_2879 ();
 FILLCELL_X32 FILLER_217_2911 ();
 FILLCELL_X32 FILLER_217_2943 ();
 FILLCELL_X32 FILLER_217_2975 ();
 FILLCELL_X32 FILLER_217_3007 ();
 FILLCELL_X32 FILLER_217_3039 ();
 FILLCELL_X32 FILLER_217_3071 ();
 FILLCELL_X32 FILLER_217_3103 ();
 FILLCELL_X32 FILLER_217_3135 ();
 FILLCELL_X32 FILLER_217_3167 ();
 FILLCELL_X32 FILLER_217_3199 ();
 FILLCELL_X32 FILLER_217_3231 ();
 FILLCELL_X32 FILLER_217_3263 ();
 FILLCELL_X32 FILLER_217_3295 ();
 FILLCELL_X32 FILLER_217_3327 ();
 FILLCELL_X32 FILLER_217_3359 ();
 FILLCELL_X32 FILLER_217_3391 ();
 FILLCELL_X32 FILLER_217_3423 ();
 FILLCELL_X32 FILLER_217_3455 ();
 FILLCELL_X32 FILLER_217_3487 ();
 FILLCELL_X32 FILLER_217_3519 ();
 FILLCELL_X32 FILLER_217_3551 ();
 FILLCELL_X32 FILLER_217_3583 ();
 FILLCELL_X32 FILLER_217_3615 ();
 FILLCELL_X32 FILLER_217_3647 ();
 FILLCELL_X32 FILLER_217_3679 ();
 FILLCELL_X16 FILLER_217_3711 ();
 FILLCELL_X8 FILLER_217_3727 ();
 FILLCELL_X2 FILLER_217_3735 ();
 FILLCELL_X1 FILLER_217_3737 ();
 FILLCELL_X32 FILLER_218_1 ();
 FILLCELL_X32 FILLER_218_33 ();
 FILLCELL_X32 FILLER_218_65 ();
 FILLCELL_X32 FILLER_218_97 ();
 FILLCELL_X32 FILLER_218_129 ();
 FILLCELL_X32 FILLER_218_161 ();
 FILLCELL_X32 FILLER_218_193 ();
 FILLCELL_X32 FILLER_218_225 ();
 FILLCELL_X32 FILLER_218_257 ();
 FILLCELL_X32 FILLER_218_289 ();
 FILLCELL_X32 FILLER_218_321 ();
 FILLCELL_X32 FILLER_218_353 ();
 FILLCELL_X32 FILLER_218_385 ();
 FILLCELL_X32 FILLER_218_417 ();
 FILLCELL_X32 FILLER_218_449 ();
 FILLCELL_X32 FILLER_218_481 ();
 FILLCELL_X32 FILLER_218_513 ();
 FILLCELL_X32 FILLER_218_545 ();
 FILLCELL_X32 FILLER_218_577 ();
 FILLCELL_X16 FILLER_218_609 ();
 FILLCELL_X4 FILLER_218_625 ();
 FILLCELL_X2 FILLER_218_629 ();
 FILLCELL_X32 FILLER_218_632 ();
 FILLCELL_X32 FILLER_218_664 ();
 FILLCELL_X32 FILLER_218_696 ();
 FILLCELL_X32 FILLER_218_728 ();
 FILLCELL_X32 FILLER_218_760 ();
 FILLCELL_X32 FILLER_218_792 ();
 FILLCELL_X32 FILLER_218_824 ();
 FILLCELL_X32 FILLER_218_856 ();
 FILLCELL_X32 FILLER_218_888 ();
 FILLCELL_X32 FILLER_218_920 ();
 FILLCELL_X32 FILLER_218_952 ();
 FILLCELL_X32 FILLER_218_984 ();
 FILLCELL_X32 FILLER_218_1016 ();
 FILLCELL_X32 FILLER_218_1048 ();
 FILLCELL_X32 FILLER_218_1080 ();
 FILLCELL_X32 FILLER_218_1112 ();
 FILLCELL_X32 FILLER_218_1144 ();
 FILLCELL_X32 FILLER_218_1176 ();
 FILLCELL_X32 FILLER_218_1208 ();
 FILLCELL_X32 FILLER_218_1240 ();
 FILLCELL_X32 FILLER_218_1272 ();
 FILLCELL_X32 FILLER_218_1304 ();
 FILLCELL_X32 FILLER_218_1336 ();
 FILLCELL_X32 FILLER_218_1368 ();
 FILLCELL_X32 FILLER_218_1400 ();
 FILLCELL_X32 FILLER_218_1432 ();
 FILLCELL_X32 FILLER_218_1464 ();
 FILLCELL_X32 FILLER_218_1496 ();
 FILLCELL_X32 FILLER_218_1528 ();
 FILLCELL_X32 FILLER_218_1560 ();
 FILLCELL_X32 FILLER_218_1592 ();
 FILLCELL_X32 FILLER_218_1624 ();
 FILLCELL_X32 FILLER_218_1656 ();
 FILLCELL_X32 FILLER_218_1688 ();
 FILLCELL_X32 FILLER_218_1720 ();
 FILLCELL_X32 FILLER_218_1752 ();
 FILLCELL_X32 FILLER_218_1784 ();
 FILLCELL_X32 FILLER_218_1816 ();
 FILLCELL_X32 FILLER_218_1848 ();
 FILLCELL_X8 FILLER_218_1880 ();
 FILLCELL_X4 FILLER_218_1888 ();
 FILLCELL_X2 FILLER_218_1892 ();
 FILLCELL_X32 FILLER_218_1895 ();
 FILLCELL_X32 FILLER_218_1927 ();
 FILLCELL_X32 FILLER_218_1959 ();
 FILLCELL_X32 FILLER_218_1991 ();
 FILLCELL_X32 FILLER_218_2023 ();
 FILLCELL_X32 FILLER_218_2055 ();
 FILLCELL_X32 FILLER_218_2087 ();
 FILLCELL_X32 FILLER_218_2119 ();
 FILLCELL_X32 FILLER_218_2151 ();
 FILLCELL_X32 FILLER_218_2183 ();
 FILLCELL_X32 FILLER_218_2215 ();
 FILLCELL_X32 FILLER_218_2247 ();
 FILLCELL_X32 FILLER_218_2279 ();
 FILLCELL_X32 FILLER_218_2311 ();
 FILLCELL_X32 FILLER_218_2343 ();
 FILLCELL_X32 FILLER_218_2375 ();
 FILLCELL_X32 FILLER_218_2407 ();
 FILLCELL_X32 FILLER_218_2439 ();
 FILLCELL_X32 FILLER_218_2471 ();
 FILLCELL_X32 FILLER_218_2503 ();
 FILLCELL_X32 FILLER_218_2535 ();
 FILLCELL_X32 FILLER_218_2567 ();
 FILLCELL_X32 FILLER_218_2599 ();
 FILLCELL_X32 FILLER_218_2631 ();
 FILLCELL_X32 FILLER_218_2663 ();
 FILLCELL_X32 FILLER_218_2695 ();
 FILLCELL_X32 FILLER_218_2727 ();
 FILLCELL_X32 FILLER_218_2759 ();
 FILLCELL_X32 FILLER_218_2791 ();
 FILLCELL_X32 FILLER_218_2823 ();
 FILLCELL_X32 FILLER_218_2855 ();
 FILLCELL_X32 FILLER_218_2887 ();
 FILLCELL_X32 FILLER_218_2919 ();
 FILLCELL_X32 FILLER_218_2951 ();
 FILLCELL_X32 FILLER_218_2983 ();
 FILLCELL_X32 FILLER_218_3015 ();
 FILLCELL_X32 FILLER_218_3047 ();
 FILLCELL_X32 FILLER_218_3079 ();
 FILLCELL_X32 FILLER_218_3111 ();
 FILLCELL_X8 FILLER_218_3143 ();
 FILLCELL_X4 FILLER_218_3151 ();
 FILLCELL_X2 FILLER_218_3155 ();
 FILLCELL_X32 FILLER_218_3158 ();
 FILLCELL_X32 FILLER_218_3190 ();
 FILLCELL_X32 FILLER_218_3222 ();
 FILLCELL_X32 FILLER_218_3254 ();
 FILLCELL_X32 FILLER_218_3286 ();
 FILLCELL_X32 FILLER_218_3318 ();
 FILLCELL_X32 FILLER_218_3350 ();
 FILLCELL_X32 FILLER_218_3382 ();
 FILLCELL_X32 FILLER_218_3414 ();
 FILLCELL_X32 FILLER_218_3446 ();
 FILLCELL_X32 FILLER_218_3478 ();
 FILLCELL_X32 FILLER_218_3510 ();
 FILLCELL_X32 FILLER_218_3542 ();
 FILLCELL_X32 FILLER_218_3574 ();
 FILLCELL_X32 FILLER_218_3606 ();
 FILLCELL_X32 FILLER_218_3638 ();
 FILLCELL_X32 FILLER_218_3670 ();
 FILLCELL_X32 FILLER_218_3702 ();
 FILLCELL_X4 FILLER_218_3734 ();
 FILLCELL_X32 FILLER_219_1 ();
 FILLCELL_X32 FILLER_219_33 ();
 FILLCELL_X32 FILLER_219_65 ();
 FILLCELL_X32 FILLER_219_97 ();
 FILLCELL_X32 FILLER_219_129 ();
 FILLCELL_X32 FILLER_219_161 ();
 FILLCELL_X32 FILLER_219_193 ();
 FILLCELL_X32 FILLER_219_225 ();
 FILLCELL_X32 FILLER_219_257 ();
 FILLCELL_X32 FILLER_219_289 ();
 FILLCELL_X32 FILLER_219_321 ();
 FILLCELL_X32 FILLER_219_353 ();
 FILLCELL_X32 FILLER_219_385 ();
 FILLCELL_X32 FILLER_219_417 ();
 FILLCELL_X32 FILLER_219_449 ();
 FILLCELL_X32 FILLER_219_481 ();
 FILLCELL_X32 FILLER_219_513 ();
 FILLCELL_X32 FILLER_219_545 ();
 FILLCELL_X32 FILLER_219_577 ();
 FILLCELL_X32 FILLER_219_609 ();
 FILLCELL_X32 FILLER_219_641 ();
 FILLCELL_X32 FILLER_219_673 ();
 FILLCELL_X32 FILLER_219_705 ();
 FILLCELL_X32 FILLER_219_737 ();
 FILLCELL_X32 FILLER_219_769 ();
 FILLCELL_X32 FILLER_219_801 ();
 FILLCELL_X32 FILLER_219_833 ();
 FILLCELL_X32 FILLER_219_865 ();
 FILLCELL_X32 FILLER_219_897 ();
 FILLCELL_X32 FILLER_219_929 ();
 FILLCELL_X32 FILLER_219_961 ();
 FILLCELL_X32 FILLER_219_993 ();
 FILLCELL_X32 FILLER_219_1025 ();
 FILLCELL_X32 FILLER_219_1057 ();
 FILLCELL_X32 FILLER_219_1089 ();
 FILLCELL_X32 FILLER_219_1121 ();
 FILLCELL_X32 FILLER_219_1153 ();
 FILLCELL_X32 FILLER_219_1185 ();
 FILLCELL_X32 FILLER_219_1217 ();
 FILLCELL_X8 FILLER_219_1249 ();
 FILLCELL_X4 FILLER_219_1257 ();
 FILLCELL_X2 FILLER_219_1261 ();
 FILLCELL_X32 FILLER_219_1264 ();
 FILLCELL_X32 FILLER_219_1296 ();
 FILLCELL_X32 FILLER_219_1328 ();
 FILLCELL_X32 FILLER_219_1360 ();
 FILLCELL_X32 FILLER_219_1392 ();
 FILLCELL_X32 FILLER_219_1424 ();
 FILLCELL_X32 FILLER_219_1456 ();
 FILLCELL_X32 FILLER_219_1488 ();
 FILLCELL_X32 FILLER_219_1520 ();
 FILLCELL_X32 FILLER_219_1552 ();
 FILLCELL_X32 FILLER_219_1584 ();
 FILLCELL_X32 FILLER_219_1616 ();
 FILLCELL_X32 FILLER_219_1648 ();
 FILLCELL_X32 FILLER_219_1680 ();
 FILLCELL_X32 FILLER_219_1712 ();
 FILLCELL_X32 FILLER_219_1744 ();
 FILLCELL_X32 FILLER_219_1776 ();
 FILLCELL_X32 FILLER_219_1808 ();
 FILLCELL_X32 FILLER_219_1840 ();
 FILLCELL_X32 FILLER_219_1872 ();
 FILLCELL_X32 FILLER_219_1904 ();
 FILLCELL_X32 FILLER_219_1936 ();
 FILLCELL_X32 FILLER_219_1968 ();
 FILLCELL_X32 FILLER_219_2000 ();
 FILLCELL_X32 FILLER_219_2032 ();
 FILLCELL_X32 FILLER_219_2064 ();
 FILLCELL_X32 FILLER_219_2096 ();
 FILLCELL_X32 FILLER_219_2128 ();
 FILLCELL_X32 FILLER_219_2160 ();
 FILLCELL_X32 FILLER_219_2192 ();
 FILLCELL_X32 FILLER_219_2224 ();
 FILLCELL_X32 FILLER_219_2256 ();
 FILLCELL_X32 FILLER_219_2288 ();
 FILLCELL_X32 FILLER_219_2320 ();
 FILLCELL_X32 FILLER_219_2352 ();
 FILLCELL_X32 FILLER_219_2384 ();
 FILLCELL_X32 FILLER_219_2416 ();
 FILLCELL_X32 FILLER_219_2448 ();
 FILLCELL_X32 FILLER_219_2480 ();
 FILLCELL_X8 FILLER_219_2512 ();
 FILLCELL_X4 FILLER_219_2520 ();
 FILLCELL_X2 FILLER_219_2524 ();
 FILLCELL_X32 FILLER_219_2527 ();
 FILLCELL_X32 FILLER_219_2559 ();
 FILLCELL_X32 FILLER_219_2591 ();
 FILLCELL_X32 FILLER_219_2623 ();
 FILLCELL_X32 FILLER_219_2655 ();
 FILLCELL_X32 FILLER_219_2687 ();
 FILLCELL_X32 FILLER_219_2719 ();
 FILLCELL_X32 FILLER_219_2751 ();
 FILLCELL_X32 FILLER_219_2783 ();
 FILLCELL_X32 FILLER_219_2815 ();
 FILLCELL_X32 FILLER_219_2847 ();
 FILLCELL_X32 FILLER_219_2879 ();
 FILLCELL_X32 FILLER_219_2911 ();
 FILLCELL_X32 FILLER_219_2943 ();
 FILLCELL_X32 FILLER_219_2975 ();
 FILLCELL_X32 FILLER_219_3007 ();
 FILLCELL_X32 FILLER_219_3039 ();
 FILLCELL_X32 FILLER_219_3071 ();
 FILLCELL_X32 FILLER_219_3103 ();
 FILLCELL_X32 FILLER_219_3135 ();
 FILLCELL_X32 FILLER_219_3167 ();
 FILLCELL_X32 FILLER_219_3199 ();
 FILLCELL_X32 FILLER_219_3231 ();
 FILLCELL_X32 FILLER_219_3263 ();
 FILLCELL_X32 FILLER_219_3295 ();
 FILLCELL_X32 FILLER_219_3327 ();
 FILLCELL_X32 FILLER_219_3359 ();
 FILLCELL_X32 FILLER_219_3391 ();
 FILLCELL_X32 FILLER_219_3423 ();
 FILLCELL_X32 FILLER_219_3455 ();
 FILLCELL_X32 FILLER_219_3487 ();
 FILLCELL_X32 FILLER_219_3519 ();
 FILLCELL_X32 FILLER_219_3551 ();
 FILLCELL_X32 FILLER_219_3583 ();
 FILLCELL_X32 FILLER_219_3615 ();
 FILLCELL_X32 FILLER_219_3647 ();
 FILLCELL_X32 FILLER_219_3679 ();
 FILLCELL_X16 FILLER_219_3711 ();
 FILLCELL_X8 FILLER_219_3727 ();
 FILLCELL_X2 FILLER_219_3735 ();
 FILLCELL_X1 FILLER_219_3737 ();
 FILLCELL_X32 FILLER_220_1 ();
 FILLCELL_X32 FILLER_220_33 ();
 FILLCELL_X32 FILLER_220_65 ();
 FILLCELL_X32 FILLER_220_97 ();
 FILLCELL_X32 FILLER_220_129 ();
 FILLCELL_X32 FILLER_220_161 ();
 FILLCELL_X32 FILLER_220_193 ();
 FILLCELL_X32 FILLER_220_225 ();
 FILLCELL_X32 FILLER_220_257 ();
 FILLCELL_X32 FILLER_220_289 ();
 FILLCELL_X32 FILLER_220_321 ();
 FILLCELL_X32 FILLER_220_353 ();
 FILLCELL_X32 FILLER_220_385 ();
 FILLCELL_X32 FILLER_220_417 ();
 FILLCELL_X32 FILLER_220_449 ();
 FILLCELL_X32 FILLER_220_481 ();
 FILLCELL_X32 FILLER_220_513 ();
 FILLCELL_X32 FILLER_220_545 ();
 FILLCELL_X32 FILLER_220_577 ();
 FILLCELL_X16 FILLER_220_609 ();
 FILLCELL_X4 FILLER_220_625 ();
 FILLCELL_X2 FILLER_220_629 ();
 FILLCELL_X32 FILLER_220_632 ();
 FILLCELL_X32 FILLER_220_664 ();
 FILLCELL_X32 FILLER_220_696 ();
 FILLCELL_X32 FILLER_220_728 ();
 FILLCELL_X32 FILLER_220_760 ();
 FILLCELL_X32 FILLER_220_792 ();
 FILLCELL_X32 FILLER_220_824 ();
 FILLCELL_X32 FILLER_220_856 ();
 FILLCELL_X32 FILLER_220_888 ();
 FILLCELL_X32 FILLER_220_920 ();
 FILLCELL_X32 FILLER_220_952 ();
 FILLCELL_X32 FILLER_220_984 ();
 FILLCELL_X32 FILLER_220_1016 ();
 FILLCELL_X32 FILLER_220_1048 ();
 FILLCELL_X32 FILLER_220_1080 ();
 FILLCELL_X32 FILLER_220_1112 ();
 FILLCELL_X32 FILLER_220_1144 ();
 FILLCELL_X32 FILLER_220_1176 ();
 FILLCELL_X32 FILLER_220_1208 ();
 FILLCELL_X32 FILLER_220_1240 ();
 FILLCELL_X32 FILLER_220_1272 ();
 FILLCELL_X32 FILLER_220_1304 ();
 FILLCELL_X32 FILLER_220_1336 ();
 FILLCELL_X32 FILLER_220_1368 ();
 FILLCELL_X32 FILLER_220_1400 ();
 FILLCELL_X32 FILLER_220_1432 ();
 FILLCELL_X32 FILLER_220_1464 ();
 FILLCELL_X32 FILLER_220_1496 ();
 FILLCELL_X32 FILLER_220_1528 ();
 FILLCELL_X32 FILLER_220_1560 ();
 FILLCELL_X32 FILLER_220_1592 ();
 FILLCELL_X32 FILLER_220_1624 ();
 FILLCELL_X32 FILLER_220_1656 ();
 FILLCELL_X32 FILLER_220_1688 ();
 FILLCELL_X32 FILLER_220_1720 ();
 FILLCELL_X32 FILLER_220_1752 ();
 FILLCELL_X32 FILLER_220_1784 ();
 FILLCELL_X32 FILLER_220_1816 ();
 FILLCELL_X32 FILLER_220_1848 ();
 FILLCELL_X8 FILLER_220_1880 ();
 FILLCELL_X4 FILLER_220_1888 ();
 FILLCELL_X2 FILLER_220_1892 ();
 FILLCELL_X32 FILLER_220_1895 ();
 FILLCELL_X32 FILLER_220_1927 ();
 FILLCELL_X32 FILLER_220_1959 ();
 FILLCELL_X32 FILLER_220_1991 ();
 FILLCELL_X32 FILLER_220_2023 ();
 FILLCELL_X32 FILLER_220_2055 ();
 FILLCELL_X32 FILLER_220_2087 ();
 FILLCELL_X32 FILLER_220_2119 ();
 FILLCELL_X32 FILLER_220_2151 ();
 FILLCELL_X32 FILLER_220_2183 ();
 FILLCELL_X32 FILLER_220_2215 ();
 FILLCELL_X32 FILLER_220_2247 ();
 FILLCELL_X32 FILLER_220_2279 ();
 FILLCELL_X32 FILLER_220_2311 ();
 FILLCELL_X32 FILLER_220_2343 ();
 FILLCELL_X32 FILLER_220_2375 ();
 FILLCELL_X32 FILLER_220_2407 ();
 FILLCELL_X32 FILLER_220_2439 ();
 FILLCELL_X32 FILLER_220_2471 ();
 FILLCELL_X32 FILLER_220_2503 ();
 FILLCELL_X32 FILLER_220_2535 ();
 FILLCELL_X32 FILLER_220_2567 ();
 FILLCELL_X32 FILLER_220_2599 ();
 FILLCELL_X32 FILLER_220_2631 ();
 FILLCELL_X32 FILLER_220_2663 ();
 FILLCELL_X32 FILLER_220_2695 ();
 FILLCELL_X32 FILLER_220_2727 ();
 FILLCELL_X32 FILLER_220_2759 ();
 FILLCELL_X32 FILLER_220_2791 ();
 FILLCELL_X32 FILLER_220_2823 ();
 FILLCELL_X32 FILLER_220_2855 ();
 FILLCELL_X32 FILLER_220_2887 ();
 FILLCELL_X32 FILLER_220_2919 ();
 FILLCELL_X32 FILLER_220_2951 ();
 FILLCELL_X32 FILLER_220_2983 ();
 FILLCELL_X32 FILLER_220_3015 ();
 FILLCELL_X32 FILLER_220_3047 ();
 FILLCELL_X32 FILLER_220_3079 ();
 FILLCELL_X32 FILLER_220_3111 ();
 FILLCELL_X8 FILLER_220_3143 ();
 FILLCELL_X4 FILLER_220_3151 ();
 FILLCELL_X2 FILLER_220_3155 ();
 FILLCELL_X32 FILLER_220_3158 ();
 FILLCELL_X32 FILLER_220_3190 ();
 FILLCELL_X32 FILLER_220_3222 ();
 FILLCELL_X32 FILLER_220_3254 ();
 FILLCELL_X32 FILLER_220_3286 ();
 FILLCELL_X32 FILLER_220_3318 ();
 FILLCELL_X32 FILLER_220_3350 ();
 FILLCELL_X32 FILLER_220_3382 ();
 FILLCELL_X32 FILLER_220_3414 ();
 FILLCELL_X32 FILLER_220_3446 ();
 FILLCELL_X32 FILLER_220_3478 ();
 FILLCELL_X32 FILLER_220_3510 ();
 FILLCELL_X32 FILLER_220_3542 ();
 FILLCELL_X32 FILLER_220_3574 ();
 FILLCELL_X32 FILLER_220_3606 ();
 FILLCELL_X32 FILLER_220_3638 ();
 FILLCELL_X32 FILLER_220_3670 ();
 FILLCELL_X32 FILLER_220_3702 ();
 FILLCELL_X4 FILLER_220_3734 ();
 FILLCELL_X32 FILLER_221_1 ();
 FILLCELL_X32 FILLER_221_33 ();
 FILLCELL_X32 FILLER_221_65 ();
 FILLCELL_X32 FILLER_221_97 ();
 FILLCELL_X32 FILLER_221_129 ();
 FILLCELL_X32 FILLER_221_161 ();
 FILLCELL_X32 FILLER_221_193 ();
 FILLCELL_X32 FILLER_221_225 ();
 FILLCELL_X32 FILLER_221_257 ();
 FILLCELL_X32 FILLER_221_289 ();
 FILLCELL_X32 FILLER_221_321 ();
 FILLCELL_X32 FILLER_221_353 ();
 FILLCELL_X32 FILLER_221_385 ();
 FILLCELL_X32 FILLER_221_417 ();
 FILLCELL_X32 FILLER_221_449 ();
 FILLCELL_X32 FILLER_221_481 ();
 FILLCELL_X32 FILLER_221_513 ();
 FILLCELL_X32 FILLER_221_545 ();
 FILLCELL_X32 FILLER_221_577 ();
 FILLCELL_X32 FILLER_221_609 ();
 FILLCELL_X32 FILLER_221_641 ();
 FILLCELL_X32 FILLER_221_673 ();
 FILLCELL_X32 FILLER_221_705 ();
 FILLCELL_X32 FILLER_221_737 ();
 FILLCELL_X32 FILLER_221_769 ();
 FILLCELL_X32 FILLER_221_801 ();
 FILLCELL_X32 FILLER_221_833 ();
 FILLCELL_X32 FILLER_221_865 ();
 FILLCELL_X32 FILLER_221_897 ();
 FILLCELL_X32 FILLER_221_929 ();
 FILLCELL_X32 FILLER_221_961 ();
 FILLCELL_X32 FILLER_221_993 ();
 FILLCELL_X32 FILLER_221_1025 ();
 FILLCELL_X32 FILLER_221_1057 ();
 FILLCELL_X32 FILLER_221_1089 ();
 FILLCELL_X32 FILLER_221_1121 ();
 FILLCELL_X32 FILLER_221_1153 ();
 FILLCELL_X32 FILLER_221_1185 ();
 FILLCELL_X32 FILLER_221_1217 ();
 FILLCELL_X8 FILLER_221_1249 ();
 FILLCELL_X4 FILLER_221_1257 ();
 FILLCELL_X2 FILLER_221_1261 ();
 FILLCELL_X32 FILLER_221_1264 ();
 FILLCELL_X32 FILLER_221_1296 ();
 FILLCELL_X32 FILLER_221_1328 ();
 FILLCELL_X32 FILLER_221_1360 ();
 FILLCELL_X32 FILLER_221_1392 ();
 FILLCELL_X32 FILLER_221_1424 ();
 FILLCELL_X32 FILLER_221_1456 ();
 FILLCELL_X32 FILLER_221_1488 ();
 FILLCELL_X32 FILLER_221_1520 ();
 FILLCELL_X32 FILLER_221_1552 ();
 FILLCELL_X32 FILLER_221_1584 ();
 FILLCELL_X32 FILLER_221_1616 ();
 FILLCELL_X32 FILLER_221_1648 ();
 FILLCELL_X32 FILLER_221_1680 ();
 FILLCELL_X32 FILLER_221_1712 ();
 FILLCELL_X32 FILLER_221_1744 ();
 FILLCELL_X32 FILLER_221_1776 ();
 FILLCELL_X32 FILLER_221_1808 ();
 FILLCELL_X32 FILLER_221_1840 ();
 FILLCELL_X32 FILLER_221_1872 ();
 FILLCELL_X32 FILLER_221_1904 ();
 FILLCELL_X32 FILLER_221_1936 ();
 FILLCELL_X32 FILLER_221_1968 ();
 FILLCELL_X32 FILLER_221_2000 ();
 FILLCELL_X32 FILLER_221_2032 ();
 FILLCELL_X32 FILLER_221_2064 ();
 FILLCELL_X32 FILLER_221_2096 ();
 FILLCELL_X32 FILLER_221_2128 ();
 FILLCELL_X32 FILLER_221_2160 ();
 FILLCELL_X32 FILLER_221_2192 ();
 FILLCELL_X32 FILLER_221_2224 ();
 FILLCELL_X32 FILLER_221_2256 ();
 FILLCELL_X32 FILLER_221_2288 ();
 FILLCELL_X32 FILLER_221_2320 ();
 FILLCELL_X32 FILLER_221_2352 ();
 FILLCELL_X32 FILLER_221_2384 ();
 FILLCELL_X32 FILLER_221_2416 ();
 FILLCELL_X32 FILLER_221_2448 ();
 FILLCELL_X32 FILLER_221_2480 ();
 FILLCELL_X8 FILLER_221_2512 ();
 FILLCELL_X4 FILLER_221_2520 ();
 FILLCELL_X2 FILLER_221_2524 ();
 FILLCELL_X32 FILLER_221_2527 ();
 FILLCELL_X32 FILLER_221_2559 ();
 FILLCELL_X32 FILLER_221_2591 ();
 FILLCELL_X32 FILLER_221_2623 ();
 FILLCELL_X32 FILLER_221_2655 ();
 FILLCELL_X32 FILLER_221_2687 ();
 FILLCELL_X32 FILLER_221_2719 ();
 FILLCELL_X32 FILLER_221_2751 ();
 FILLCELL_X32 FILLER_221_2783 ();
 FILLCELL_X32 FILLER_221_2815 ();
 FILLCELL_X32 FILLER_221_2847 ();
 FILLCELL_X32 FILLER_221_2879 ();
 FILLCELL_X32 FILLER_221_2911 ();
 FILLCELL_X32 FILLER_221_2943 ();
 FILLCELL_X32 FILLER_221_2975 ();
 FILLCELL_X32 FILLER_221_3007 ();
 FILLCELL_X32 FILLER_221_3039 ();
 FILLCELL_X32 FILLER_221_3071 ();
 FILLCELL_X32 FILLER_221_3103 ();
 FILLCELL_X32 FILLER_221_3135 ();
 FILLCELL_X32 FILLER_221_3167 ();
 FILLCELL_X32 FILLER_221_3199 ();
 FILLCELL_X32 FILLER_221_3231 ();
 FILLCELL_X32 FILLER_221_3263 ();
 FILLCELL_X32 FILLER_221_3295 ();
 FILLCELL_X32 FILLER_221_3327 ();
 FILLCELL_X32 FILLER_221_3359 ();
 FILLCELL_X32 FILLER_221_3391 ();
 FILLCELL_X32 FILLER_221_3423 ();
 FILLCELL_X32 FILLER_221_3455 ();
 FILLCELL_X32 FILLER_221_3487 ();
 FILLCELL_X32 FILLER_221_3519 ();
 FILLCELL_X32 FILLER_221_3551 ();
 FILLCELL_X32 FILLER_221_3583 ();
 FILLCELL_X32 FILLER_221_3615 ();
 FILLCELL_X32 FILLER_221_3647 ();
 FILLCELL_X32 FILLER_221_3679 ();
 FILLCELL_X16 FILLER_221_3711 ();
 FILLCELL_X8 FILLER_221_3727 ();
 FILLCELL_X2 FILLER_221_3735 ();
 FILLCELL_X1 FILLER_221_3737 ();
 FILLCELL_X32 FILLER_222_1 ();
 FILLCELL_X32 FILLER_222_33 ();
 FILLCELL_X32 FILLER_222_65 ();
 FILLCELL_X32 FILLER_222_97 ();
 FILLCELL_X32 FILLER_222_129 ();
 FILLCELL_X32 FILLER_222_161 ();
 FILLCELL_X32 FILLER_222_193 ();
 FILLCELL_X32 FILLER_222_225 ();
 FILLCELL_X32 FILLER_222_257 ();
 FILLCELL_X32 FILLER_222_289 ();
 FILLCELL_X32 FILLER_222_321 ();
 FILLCELL_X32 FILLER_222_353 ();
 FILLCELL_X32 FILLER_222_385 ();
 FILLCELL_X32 FILLER_222_417 ();
 FILLCELL_X32 FILLER_222_449 ();
 FILLCELL_X32 FILLER_222_481 ();
 FILLCELL_X32 FILLER_222_513 ();
 FILLCELL_X32 FILLER_222_545 ();
 FILLCELL_X32 FILLER_222_577 ();
 FILLCELL_X16 FILLER_222_609 ();
 FILLCELL_X4 FILLER_222_625 ();
 FILLCELL_X2 FILLER_222_629 ();
 FILLCELL_X32 FILLER_222_632 ();
 FILLCELL_X32 FILLER_222_664 ();
 FILLCELL_X32 FILLER_222_696 ();
 FILLCELL_X32 FILLER_222_728 ();
 FILLCELL_X32 FILLER_222_760 ();
 FILLCELL_X32 FILLER_222_792 ();
 FILLCELL_X32 FILLER_222_824 ();
 FILLCELL_X32 FILLER_222_856 ();
 FILLCELL_X32 FILLER_222_888 ();
 FILLCELL_X32 FILLER_222_920 ();
 FILLCELL_X32 FILLER_222_952 ();
 FILLCELL_X32 FILLER_222_984 ();
 FILLCELL_X32 FILLER_222_1016 ();
 FILLCELL_X32 FILLER_222_1048 ();
 FILLCELL_X32 FILLER_222_1080 ();
 FILLCELL_X32 FILLER_222_1112 ();
 FILLCELL_X32 FILLER_222_1144 ();
 FILLCELL_X32 FILLER_222_1176 ();
 FILLCELL_X32 FILLER_222_1208 ();
 FILLCELL_X32 FILLER_222_1240 ();
 FILLCELL_X32 FILLER_222_1272 ();
 FILLCELL_X32 FILLER_222_1304 ();
 FILLCELL_X32 FILLER_222_1336 ();
 FILLCELL_X32 FILLER_222_1368 ();
 FILLCELL_X32 FILLER_222_1400 ();
 FILLCELL_X32 FILLER_222_1432 ();
 FILLCELL_X32 FILLER_222_1464 ();
 FILLCELL_X32 FILLER_222_1496 ();
 FILLCELL_X32 FILLER_222_1528 ();
 FILLCELL_X32 FILLER_222_1560 ();
 FILLCELL_X32 FILLER_222_1592 ();
 FILLCELL_X32 FILLER_222_1624 ();
 FILLCELL_X32 FILLER_222_1656 ();
 FILLCELL_X32 FILLER_222_1688 ();
 FILLCELL_X32 FILLER_222_1720 ();
 FILLCELL_X32 FILLER_222_1752 ();
 FILLCELL_X32 FILLER_222_1784 ();
 FILLCELL_X32 FILLER_222_1816 ();
 FILLCELL_X32 FILLER_222_1848 ();
 FILLCELL_X8 FILLER_222_1880 ();
 FILLCELL_X4 FILLER_222_1888 ();
 FILLCELL_X2 FILLER_222_1892 ();
 FILLCELL_X32 FILLER_222_1895 ();
 FILLCELL_X32 FILLER_222_1927 ();
 FILLCELL_X32 FILLER_222_1959 ();
 FILLCELL_X32 FILLER_222_1991 ();
 FILLCELL_X32 FILLER_222_2023 ();
 FILLCELL_X32 FILLER_222_2055 ();
 FILLCELL_X32 FILLER_222_2087 ();
 FILLCELL_X32 FILLER_222_2119 ();
 FILLCELL_X32 FILLER_222_2151 ();
 FILLCELL_X32 FILLER_222_2183 ();
 FILLCELL_X32 FILLER_222_2215 ();
 FILLCELL_X32 FILLER_222_2247 ();
 FILLCELL_X32 FILLER_222_2279 ();
 FILLCELL_X32 FILLER_222_2311 ();
 FILLCELL_X32 FILLER_222_2343 ();
 FILLCELL_X32 FILLER_222_2375 ();
 FILLCELL_X32 FILLER_222_2407 ();
 FILLCELL_X32 FILLER_222_2439 ();
 FILLCELL_X32 FILLER_222_2471 ();
 FILLCELL_X32 FILLER_222_2503 ();
 FILLCELL_X32 FILLER_222_2535 ();
 FILLCELL_X32 FILLER_222_2567 ();
 FILLCELL_X32 FILLER_222_2599 ();
 FILLCELL_X32 FILLER_222_2631 ();
 FILLCELL_X32 FILLER_222_2663 ();
 FILLCELL_X32 FILLER_222_2695 ();
 FILLCELL_X32 FILLER_222_2727 ();
 FILLCELL_X32 FILLER_222_2759 ();
 FILLCELL_X32 FILLER_222_2791 ();
 FILLCELL_X32 FILLER_222_2823 ();
 FILLCELL_X32 FILLER_222_2855 ();
 FILLCELL_X32 FILLER_222_2887 ();
 FILLCELL_X32 FILLER_222_2919 ();
 FILLCELL_X32 FILLER_222_2951 ();
 FILLCELL_X32 FILLER_222_2983 ();
 FILLCELL_X32 FILLER_222_3015 ();
 FILLCELL_X32 FILLER_222_3047 ();
 FILLCELL_X32 FILLER_222_3079 ();
 FILLCELL_X32 FILLER_222_3111 ();
 FILLCELL_X8 FILLER_222_3143 ();
 FILLCELL_X4 FILLER_222_3151 ();
 FILLCELL_X2 FILLER_222_3155 ();
 FILLCELL_X32 FILLER_222_3158 ();
 FILLCELL_X32 FILLER_222_3190 ();
 FILLCELL_X32 FILLER_222_3222 ();
 FILLCELL_X32 FILLER_222_3254 ();
 FILLCELL_X32 FILLER_222_3286 ();
 FILLCELL_X32 FILLER_222_3318 ();
 FILLCELL_X32 FILLER_222_3350 ();
 FILLCELL_X32 FILLER_222_3382 ();
 FILLCELL_X32 FILLER_222_3414 ();
 FILLCELL_X32 FILLER_222_3446 ();
 FILLCELL_X32 FILLER_222_3478 ();
 FILLCELL_X32 FILLER_222_3510 ();
 FILLCELL_X32 FILLER_222_3542 ();
 FILLCELL_X32 FILLER_222_3574 ();
 FILLCELL_X32 FILLER_222_3606 ();
 FILLCELL_X32 FILLER_222_3638 ();
 FILLCELL_X32 FILLER_222_3670 ();
 FILLCELL_X32 FILLER_222_3702 ();
 FILLCELL_X4 FILLER_222_3734 ();
 FILLCELL_X32 FILLER_223_1 ();
 FILLCELL_X32 FILLER_223_33 ();
 FILLCELL_X32 FILLER_223_65 ();
 FILLCELL_X32 FILLER_223_97 ();
 FILLCELL_X32 FILLER_223_129 ();
 FILLCELL_X32 FILLER_223_161 ();
 FILLCELL_X32 FILLER_223_193 ();
 FILLCELL_X32 FILLER_223_225 ();
 FILLCELL_X32 FILLER_223_257 ();
 FILLCELL_X32 FILLER_223_289 ();
 FILLCELL_X32 FILLER_223_321 ();
 FILLCELL_X32 FILLER_223_353 ();
 FILLCELL_X32 FILLER_223_385 ();
 FILLCELL_X32 FILLER_223_417 ();
 FILLCELL_X32 FILLER_223_449 ();
 FILLCELL_X32 FILLER_223_481 ();
 FILLCELL_X32 FILLER_223_513 ();
 FILLCELL_X32 FILLER_223_545 ();
 FILLCELL_X32 FILLER_223_577 ();
 FILLCELL_X32 FILLER_223_609 ();
 FILLCELL_X32 FILLER_223_641 ();
 FILLCELL_X32 FILLER_223_673 ();
 FILLCELL_X32 FILLER_223_705 ();
 FILLCELL_X32 FILLER_223_737 ();
 FILLCELL_X32 FILLER_223_769 ();
 FILLCELL_X32 FILLER_223_801 ();
 FILLCELL_X32 FILLER_223_833 ();
 FILLCELL_X32 FILLER_223_865 ();
 FILLCELL_X32 FILLER_223_897 ();
 FILLCELL_X32 FILLER_223_929 ();
 FILLCELL_X32 FILLER_223_961 ();
 FILLCELL_X32 FILLER_223_993 ();
 FILLCELL_X32 FILLER_223_1025 ();
 FILLCELL_X32 FILLER_223_1057 ();
 FILLCELL_X32 FILLER_223_1089 ();
 FILLCELL_X32 FILLER_223_1121 ();
 FILLCELL_X32 FILLER_223_1153 ();
 FILLCELL_X32 FILLER_223_1185 ();
 FILLCELL_X32 FILLER_223_1217 ();
 FILLCELL_X8 FILLER_223_1249 ();
 FILLCELL_X4 FILLER_223_1257 ();
 FILLCELL_X2 FILLER_223_1261 ();
 FILLCELL_X32 FILLER_223_1264 ();
 FILLCELL_X32 FILLER_223_1296 ();
 FILLCELL_X32 FILLER_223_1328 ();
 FILLCELL_X32 FILLER_223_1360 ();
 FILLCELL_X32 FILLER_223_1392 ();
 FILLCELL_X32 FILLER_223_1424 ();
 FILLCELL_X32 FILLER_223_1456 ();
 FILLCELL_X32 FILLER_223_1488 ();
 FILLCELL_X32 FILLER_223_1520 ();
 FILLCELL_X32 FILLER_223_1552 ();
 FILLCELL_X32 FILLER_223_1584 ();
 FILLCELL_X32 FILLER_223_1616 ();
 FILLCELL_X32 FILLER_223_1648 ();
 FILLCELL_X32 FILLER_223_1680 ();
 FILLCELL_X32 FILLER_223_1712 ();
 FILLCELL_X32 FILLER_223_1744 ();
 FILLCELL_X32 FILLER_223_1776 ();
 FILLCELL_X32 FILLER_223_1808 ();
 FILLCELL_X32 FILLER_223_1840 ();
 FILLCELL_X32 FILLER_223_1872 ();
 FILLCELL_X32 FILLER_223_1904 ();
 FILLCELL_X32 FILLER_223_1936 ();
 FILLCELL_X32 FILLER_223_1968 ();
 FILLCELL_X32 FILLER_223_2000 ();
 FILLCELL_X32 FILLER_223_2032 ();
 FILLCELL_X32 FILLER_223_2064 ();
 FILLCELL_X32 FILLER_223_2096 ();
 FILLCELL_X32 FILLER_223_2128 ();
 FILLCELL_X32 FILLER_223_2160 ();
 FILLCELL_X32 FILLER_223_2192 ();
 FILLCELL_X32 FILLER_223_2224 ();
 FILLCELL_X32 FILLER_223_2256 ();
 FILLCELL_X32 FILLER_223_2288 ();
 FILLCELL_X32 FILLER_223_2320 ();
 FILLCELL_X32 FILLER_223_2352 ();
 FILLCELL_X32 FILLER_223_2384 ();
 FILLCELL_X32 FILLER_223_2416 ();
 FILLCELL_X32 FILLER_223_2448 ();
 FILLCELL_X32 FILLER_223_2480 ();
 FILLCELL_X8 FILLER_223_2512 ();
 FILLCELL_X4 FILLER_223_2520 ();
 FILLCELL_X2 FILLER_223_2524 ();
 FILLCELL_X32 FILLER_223_2527 ();
 FILLCELL_X32 FILLER_223_2559 ();
 FILLCELL_X32 FILLER_223_2591 ();
 FILLCELL_X32 FILLER_223_2623 ();
 FILLCELL_X32 FILLER_223_2655 ();
 FILLCELL_X32 FILLER_223_2687 ();
 FILLCELL_X32 FILLER_223_2719 ();
 FILLCELL_X32 FILLER_223_2751 ();
 FILLCELL_X32 FILLER_223_2783 ();
 FILLCELL_X32 FILLER_223_2815 ();
 FILLCELL_X32 FILLER_223_2847 ();
 FILLCELL_X32 FILLER_223_2879 ();
 FILLCELL_X32 FILLER_223_2911 ();
 FILLCELL_X32 FILLER_223_2943 ();
 FILLCELL_X32 FILLER_223_2975 ();
 FILLCELL_X32 FILLER_223_3007 ();
 FILLCELL_X32 FILLER_223_3039 ();
 FILLCELL_X32 FILLER_223_3071 ();
 FILLCELL_X32 FILLER_223_3103 ();
 FILLCELL_X32 FILLER_223_3135 ();
 FILLCELL_X32 FILLER_223_3167 ();
 FILLCELL_X32 FILLER_223_3199 ();
 FILLCELL_X32 FILLER_223_3231 ();
 FILLCELL_X32 FILLER_223_3263 ();
 FILLCELL_X32 FILLER_223_3295 ();
 FILLCELL_X32 FILLER_223_3327 ();
 FILLCELL_X32 FILLER_223_3359 ();
 FILLCELL_X32 FILLER_223_3391 ();
 FILLCELL_X32 FILLER_223_3423 ();
 FILLCELL_X32 FILLER_223_3455 ();
 FILLCELL_X32 FILLER_223_3487 ();
 FILLCELL_X32 FILLER_223_3519 ();
 FILLCELL_X32 FILLER_223_3551 ();
 FILLCELL_X32 FILLER_223_3583 ();
 FILLCELL_X32 FILLER_223_3615 ();
 FILLCELL_X32 FILLER_223_3647 ();
 FILLCELL_X32 FILLER_223_3679 ();
 FILLCELL_X16 FILLER_223_3711 ();
 FILLCELL_X8 FILLER_223_3727 ();
 FILLCELL_X2 FILLER_223_3735 ();
 FILLCELL_X1 FILLER_223_3737 ();
 FILLCELL_X32 FILLER_224_1 ();
 FILLCELL_X32 FILLER_224_33 ();
 FILLCELL_X32 FILLER_224_65 ();
 FILLCELL_X32 FILLER_224_97 ();
 FILLCELL_X32 FILLER_224_129 ();
 FILLCELL_X32 FILLER_224_161 ();
 FILLCELL_X32 FILLER_224_193 ();
 FILLCELL_X32 FILLER_224_225 ();
 FILLCELL_X32 FILLER_224_257 ();
 FILLCELL_X32 FILLER_224_289 ();
 FILLCELL_X32 FILLER_224_321 ();
 FILLCELL_X32 FILLER_224_353 ();
 FILLCELL_X32 FILLER_224_385 ();
 FILLCELL_X32 FILLER_224_417 ();
 FILLCELL_X32 FILLER_224_449 ();
 FILLCELL_X32 FILLER_224_481 ();
 FILLCELL_X32 FILLER_224_513 ();
 FILLCELL_X32 FILLER_224_545 ();
 FILLCELL_X32 FILLER_224_577 ();
 FILLCELL_X16 FILLER_224_609 ();
 FILLCELL_X4 FILLER_224_625 ();
 FILLCELL_X2 FILLER_224_629 ();
 FILLCELL_X32 FILLER_224_632 ();
 FILLCELL_X32 FILLER_224_664 ();
 FILLCELL_X32 FILLER_224_696 ();
 FILLCELL_X32 FILLER_224_728 ();
 FILLCELL_X32 FILLER_224_760 ();
 FILLCELL_X32 FILLER_224_792 ();
 FILLCELL_X32 FILLER_224_824 ();
 FILLCELL_X32 FILLER_224_856 ();
 FILLCELL_X32 FILLER_224_888 ();
 FILLCELL_X32 FILLER_224_920 ();
 FILLCELL_X32 FILLER_224_952 ();
 FILLCELL_X32 FILLER_224_984 ();
 FILLCELL_X32 FILLER_224_1016 ();
 FILLCELL_X32 FILLER_224_1048 ();
 FILLCELL_X32 FILLER_224_1080 ();
 FILLCELL_X32 FILLER_224_1112 ();
 FILLCELL_X32 FILLER_224_1144 ();
 FILLCELL_X32 FILLER_224_1176 ();
 FILLCELL_X32 FILLER_224_1208 ();
 FILLCELL_X32 FILLER_224_1240 ();
 FILLCELL_X32 FILLER_224_1272 ();
 FILLCELL_X32 FILLER_224_1304 ();
 FILLCELL_X32 FILLER_224_1336 ();
 FILLCELL_X32 FILLER_224_1368 ();
 FILLCELL_X32 FILLER_224_1400 ();
 FILLCELL_X32 FILLER_224_1432 ();
 FILLCELL_X32 FILLER_224_1464 ();
 FILLCELL_X32 FILLER_224_1496 ();
 FILLCELL_X32 FILLER_224_1528 ();
 FILLCELL_X32 FILLER_224_1560 ();
 FILLCELL_X32 FILLER_224_1592 ();
 FILLCELL_X32 FILLER_224_1624 ();
 FILLCELL_X32 FILLER_224_1656 ();
 FILLCELL_X32 FILLER_224_1688 ();
 FILLCELL_X32 FILLER_224_1720 ();
 FILLCELL_X32 FILLER_224_1752 ();
 FILLCELL_X32 FILLER_224_1784 ();
 FILLCELL_X32 FILLER_224_1816 ();
 FILLCELL_X32 FILLER_224_1848 ();
 FILLCELL_X8 FILLER_224_1880 ();
 FILLCELL_X4 FILLER_224_1888 ();
 FILLCELL_X2 FILLER_224_1892 ();
 FILLCELL_X32 FILLER_224_1895 ();
 FILLCELL_X32 FILLER_224_1927 ();
 FILLCELL_X32 FILLER_224_1959 ();
 FILLCELL_X32 FILLER_224_1991 ();
 FILLCELL_X32 FILLER_224_2023 ();
 FILLCELL_X32 FILLER_224_2055 ();
 FILLCELL_X32 FILLER_224_2087 ();
 FILLCELL_X32 FILLER_224_2119 ();
 FILLCELL_X32 FILLER_224_2151 ();
 FILLCELL_X32 FILLER_224_2183 ();
 FILLCELL_X32 FILLER_224_2215 ();
 FILLCELL_X32 FILLER_224_2247 ();
 FILLCELL_X32 FILLER_224_2279 ();
 FILLCELL_X32 FILLER_224_2311 ();
 FILLCELL_X32 FILLER_224_2343 ();
 FILLCELL_X32 FILLER_224_2375 ();
 FILLCELL_X32 FILLER_224_2407 ();
 FILLCELL_X32 FILLER_224_2439 ();
 FILLCELL_X32 FILLER_224_2471 ();
 FILLCELL_X32 FILLER_224_2503 ();
 FILLCELL_X32 FILLER_224_2535 ();
 FILLCELL_X32 FILLER_224_2567 ();
 FILLCELL_X32 FILLER_224_2599 ();
 FILLCELL_X32 FILLER_224_2631 ();
 FILLCELL_X32 FILLER_224_2663 ();
 FILLCELL_X32 FILLER_224_2695 ();
 FILLCELL_X32 FILLER_224_2727 ();
 FILLCELL_X32 FILLER_224_2759 ();
 FILLCELL_X32 FILLER_224_2791 ();
 FILLCELL_X32 FILLER_224_2823 ();
 FILLCELL_X32 FILLER_224_2855 ();
 FILLCELL_X32 FILLER_224_2887 ();
 FILLCELL_X32 FILLER_224_2919 ();
 FILLCELL_X32 FILLER_224_2951 ();
 FILLCELL_X32 FILLER_224_2983 ();
 FILLCELL_X32 FILLER_224_3015 ();
 FILLCELL_X32 FILLER_224_3047 ();
 FILLCELL_X32 FILLER_224_3079 ();
 FILLCELL_X32 FILLER_224_3111 ();
 FILLCELL_X8 FILLER_224_3143 ();
 FILLCELL_X4 FILLER_224_3151 ();
 FILLCELL_X2 FILLER_224_3155 ();
 FILLCELL_X32 FILLER_224_3158 ();
 FILLCELL_X32 FILLER_224_3190 ();
 FILLCELL_X32 FILLER_224_3222 ();
 FILLCELL_X32 FILLER_224_3254 ();
 FILLCELL_X32 FILLER_224_3286 ();
 FILLCELL_X32 FILLER_224_3318 ();
 FILLCELL_X32 FILLER_224_3350 ();
 FILLCELL_X32 FILLER_224_3382 ();
 FILLCELL_X32 FILLER_224_3414 ();
 FILLCELL_X32 FILLER_224_3446 ();
 FILLCELL_X32 FILLER_224_3478 ();
 FILLCELL_X32 FILLER_224_3510 ();
 FILLCELL_X32 FILLER_224_3542 ();
 FILLCELL_X32 FILLER_224_3574 ();
 FILLCELL_X32 FILLER_224_3606 ();
 FILLCELL_X32 FILLER_224_3638 ();
 FILLCELL_X32 FILLER_224_3670 ();
 FILLCELL_X32 FILLER_224_3702 ();
 FILLCELL_X4 FILLER_224_3734 ();
 FILLCELL_X32 FILLER_225_1 ();
 FILLCELL_X32 FILLER_225_33 ();
 FILLCELL_X32 FILLER_225_65 ();
 FILLCELL_X32 FILLER_225_97 ();
 FILLCELL_X32 FILLER_225_129 ();
 FILLCELL_X32 FILLER_225_161 ();
 FILLCELL_X32 FILLER_225_193 ();
 FILLCELL_X32 FILLER_225_225 ();
 FILLCELL_X32 FILLER_225_257 ();
 FILLCELL_X32 FILLER_225_289 ();
 FILLCELL_X32 FILLER_225_321 ();
 FILLCELL_X32 FILLER_225_353 ();
 FILLCELL_X32 FILLER_225_385 ();
 FILLCELL_X32 FILLER_225_417 ();
 FILLCELL_X32 FILLER_225_449 ();
 FILLCELL_X32 FILLER_225_481 ();
 FILLCELL_X32 FILLER_225_513 ();
 FILLCELL_X32 FILLER_225_545 ();
 FILLCELL_X32 FILLER_225_577 ();
 FILLCELL_X32 FILLER_225_609 ();
 FILLCELL_X32 FILLER_225_641 ();
 FILLCELL_X32 FILLER_225_673 ();
 FILLCELL_X32 FILLER_225_705 ();
 FILLCELL_X32 FILLER_225_737 ();
 FILLCELL_X32 FILLER_225_769 ();
 FILLCELL_X32 FILLER_225_801 ();
 FILLCELL_X32 FILLER_225_833 ();
 FILLCELL_X32 FILLER_225_865 ();
 FILLCELL_X32 FILLER_225_897 ();
 FILLCELL_X32 FILLER_225_929 ();
 FILLCELL_X32 FILLER_225_961 ();
 FILLCELL_X32 FILLER_225_993 ();
 FILLCELL_X32 FILLER_225_1025 ();
 FILLCELL_X32 FILLER_225_1057 ();
 FILLCELL_X32 FILLER_225_1089 ();
 FILLCELL_X32 FILLER_225_1121 ();
 FILLCELL_X32 FILLER_225_1153 ();
 FILLCELL_X32 FILLER_225_1185 ();
 FILLCELL_X32 FILLER_225_1217 ();
 FILLCELL_X8 FILLER_225_1249 ();
 FILLCELL_X4 FILLER_225_1257 ();
 FILLCELL_X2 FILLER_225_1261 ();
 FILLCELL_X32 FILLER_225_1264 ();
 FILLCELL_X32 FILLER_225_1296 ();
 FILLCELL_X32 FILLER_225_1328 ();
 FILLCELL_X32 FILLER_225_1360 ();
 FILLCELL_X32 FILLER_225_1392 ();
 FILLCELL_X32 FILLER_225_1424 ();
 FILLCELL_X32 FILLER_225_1456 ();
 FILLCELL_X32 FILLER_225_1488 ();
 FILLCELL_X32 FILLER_225_1520 ();
 FILLCELL_X32 FILLER_225_1552 ();
 FILLCELL_X32 FILLER_225_1584 ();
 FILLCELL_X32 FILLER_225_1616 ();
 FILLCELL_X32 FILLER_225_1648 ();
 FILLCELL_X32 FILLER_225_1680 ();
 FILLCELL_X32 FILLER_225_1712 ();
 FILLCELL_X32 FILLER_225_1744 ();
 FILLCELL_X32 FILLER_225_1776 ();
 FILLCELL_X32 FILLER_225_1808 ();
 FILLCELL_X32 FILLER_225_1840 ();
 FILLCELL_X16 FILLER_225_1872 ();
 FILLCELL_X4 FILLER_225_1888 ();
 FILLCELL_X1 FILLER_225_1892 ();
 FILLCELL_X2 FILLER_225_1899 ();
 FILLCELL_X32 FILLER_225_1914 ();
 FILLCELL_X32 FILLER_225_1946 ();
 FILLCELL_X32 FILLER_225_1978 ();
 FILLCELL_X32 FILLER_225_2010 ();
 FILLCELL_X32 FILLER_225_2042 ();
 FILLCELL_X32 FILLER_225_2074 ();
 FILLCELL_X32 FILLER_225_2106 ();
 FILLCELL_X32 FILLER_225_2138 ();
 FILLCELL_X32 FILLER_225_2170 ();
 FILLCELL_X32 FILLER_225_2202 ();
 FILLCELL_X32 FILLER_225_2234 ();
 FILLCELL_X32 FILLER_225_2266 ();
 FILLCELL_X32 FILLER_225_2298 ();
 FILLCELL_X32 FILLER_225_2330 ();
 FILLCELL_X32 FILLER_225_2362 ();
 FILLCELL_X32 FILLER_225_2394 ();
 FILLCELL_X32 FILLER_225_2426 ();
 FILLCELL_X32 FILLER_225_2458 ();
 FILLCELL_X32 FILLER_225_2490 ();
 FILLCELL_X4 FILLER_225_2522 ();
 FILLCELL_X32 FILLER_225_2527 ();
 FILLCELL_X32 FILLER_225_2559 ();
 FILLCELL_X32 FILLER_225_2591 ();
 FILLCELL_X32 FILLER_225_2623 ();
 FILLCELL_X32 FILLER_225_2655 ();
 FILLCELL_X32 FILLER_225_2687 ();
 FILLCELL_X32 FILLER_225_2719 ();
 FILLCELL_X32 FILLER_225_2751 ();
 FILLCELL_X32 FILLER_225_2783 ();
 FILLCELL_X32 FILLER_225_2815 ();
 FILLCELL_X32 FILLER_225_2847 ();
 FILLCELL_X32 FILLER_225_2879 ();
 FILLCELL_X32 FILLER_225_2911 ();
 FILLCELL_X32 FILLER_225_2943 ();
 FILLCELL_X32 FILLER_225_2975 ();
 FILLCELL_X32 FILLER_225_3007 ();
 FILLCELL_X32 FILLER_225_3039 ();
 FILLCELL_X32 FILLER_225_3071 ();
 FILLCELL_X32 FILLER_225_3103 ();
 FILLCELL_X32 FILLER_225_3135 ();
 FILLCELL_X32 FILLER_225_3167 ();
 FILLCELL_X32 FILLER_225_3199 ();
 FILLCELL_X32 FILLER_225_3231 ();
 FILLCELL_X32 FILLER_225_3263 ();
 FILLCELL_X32 FILLER_225_3295 ();
 FILLCELL_X32 FILLER_225_3327 ();
 FILLCELL_X32 FILLER_225_3359 ();
 FILLCELL_X32 FILLER_225_3391 ();
 FILLCELL_X32 FILLER_225_3423 ();
 FILLCELL_X32 FILLER_225_3455 ();
 FILLCELL_X32 FILLER_225_3487 ();
 FILLCELL_X32 FILLER_225_3519 ();
 FILLCELL_X32 FILLER_225_3551 ();
 FILLCELL_X32 FILLER_225_3583 ();
 FILLCELL_X32 FILLER_225_3615 ();
 FILLCELL_X32 FILLER_225_3647 ();
 FILLCELL_X32 FILLER_225_3679 ();
 FILLCELL_X16 FILLER_225_3711 ();
 FILLCELL_X8 FILLER_225_3727 ();
 FILLCELL_X2 FILLER_225_3735 ();
 FILLCELL_X1 FILLER_225_3737 ();
 FILLCELL_X32 FILLER_226_1 ();
 FILLCELL_X32 FILLER_226_33 ();
 FILLCELL_X32 FILLER_226_65 ();
 FILLCELL_X32 FILLER_226_97 ();
 FILLCELL_X32 FILLER_226_129 ();
 FILLCELL_X32 FILLER_226_161 ();
 FILLCELL_X32 FILLER_226_193 ();
 FILLCELL_X32 FILLER_226_225 ();
 FILLCELL_X32 FILLER_226_257 ();
 FILLCELL_X32 FILLER_226_289 ();
 FILLCELL_X32 FILLER_226_321 ();
 FILLCELL_X32 FILLER_226_353 ();
 FILLCELL_X32 FILLER_226_385 ();
 FILLCELL_X32 FILLER_226_417 ();
 FILLCELL_X32 FILLER_226_449 ();
 FILLCELL_X32 FILLER_226_481 ();
 FILLCELL_X32 FILLER_226_513 ();
 FILLCELL_X32 FILLER_226_545 ();
 FILLCELL_X32 FILLER_226_577 ();
 FILLCELL_X16 FILLER_226_609 ();
 FILLCELL_X4 FILLER_226_625 ();
 FILLCELL_X2 FILLER_226_629 ();
 FILLCELL_X32 FILLER_226_632 ();
 FILLCELL_X32 FILLER_226_664 ();
 FILLCELL_X32 FILLER_226_696 ();
 FILLCELL_X32 FILLER_226_728 ();
 FILLCELL_X32 FILLER_226_760 ();
 FILLCELL_X32 FILLER_226_792 ();
 FILLCELL_X32 FILLER_226_824 ();
 FILLCELL_X32 FILLER_226_856 ();
 FILLCELL_X32 FILLER_226_888 ();
 FILLCELL_X32 FILLER_226_920 ();
 FILLCELL_X32 FILLER_226_952 ();
 FILLCELL_X32 FILLER_226_984 ();
 FILLCELL_X32 FILLER_226_1016 ();
 FILLCELL_X32 FILLER_226_1048 ();
 FILLCELL_X32 FILLER_226_1080 ();
 FILLCELL_X32 FILLER_226_1112 ();
 FILLCELL_X32 FILLER_226_1144 ();
 FILLCELL_X32 FILLER_226_1176 ();
 FILLCELL_X32 FILLER_226_1208 ();
 FILLCELL_X32 FILLER_226_1240 ();
 FILLCELL_X32 FILLER_226_1272 ();
 FILLCELL_X32 FILLER_226_1304 ();
 FILLCELL_X32 FILLER_226_1336 ();
 FILLCELL_X32 FILLER_226_1368 ();
 FILLCELL_X32 FILLER_226_1400 ();
 FILLCELL_X32 FILLER_226_1432 ();
 FILLCELL_X32 FILLER_226_1464 ();
 FILLCELL_X32 FILLER_226_1496 ();
 FILLCELL_X32 FILLER_226_1528 ();
 FILLCELL_X32 FILLER_226_1560 ();
 FILLCELL_X32 FILLER_226_1592 ();
 FILLCELL_X32 FILLER_226_1624 ();
 FILLCELL_X32 FILLER_226_1656 ();
 FILLCELL_X32 FILLER_226_1688 ();
 FILLCELL_X32 FILLER_226_1720 ();
 FILLCELL_X32 FILLER_226_1752 ();
 FILLCELL_X32 FILLER_226_1784 ();
 FILLCELL_X32 FILLER_226_1816 ();
 FILLCELL_X32 FILLER_226_1848 ();
 FILLCELL_X4 FILLER_226_1880 ();
 FILLCELL_X1 FILLER_226_1884 ();
 FILLCELL_X2 FILLER_226_1892 ();
 FILLCELL_X32 FILLER_226_1913 ();
 FILLCELL_X16 FILLER_226_1945 ();
 FILLCELL_X8 FILLER_226_1961 ();
 FILLCELL_X4 FILLER_226_1969 ();
 FILLCELL_X16 FILLER_226_1982 ();
 FILLCELL_X8 FILLER_226_1998 ();
 FILLCELL_X4 FILLER_226_2006 ();
 FILLCELL_X1 FILLER_226_2010 ();
 FILLCELL_X32 FILLER_226_2020 ();
 FILLCELL_X32 FILLER_226_2052 ();
 FILLCELL_X32 FILLER_226_2084 ();
 FILLCELL_X32 FILLER_226_2116 ();
 FILLCELL_X32 FILLER_226_2148 ();
 FILLCELL_X32 FILLER_226_2180 ();
 FILLCELL_X32 FILLER_226_2212 ();
 FILLCELL_X32 FILLER_226_2244 ();
 FILLCELL_X32 FILLER_226_2276 ();
 FILLCELL_X32 FILLER_226_2308 ();
 FILLCELL_X32 FILLER_226_2340 ();
 FILLCELL_X32 FILLER_226_2372 ();
 FILLCELL_X32 FILLER_226_2404 ();
 FILLCELL_X32 FILLER_226_2436 ();
 FILLCELL_X32 FILLER_226_2468 ();
 FILLCELL_X32 FILLER_226_2500 ();
 FILLCELL_X32 FILLER_226_2532 ();
 FILLCELL_X32 FILLER_226_2564 ();
 FILLCELL_X32 FILLER_226_2596 ();
 FILLCELL_X32 FILLER_226_2628 ();
 FILLCELL_X32 FILLER_226_2660 ();
 FILLCELL_X32 FILLER_226_2692 ();
 FILLCELL_X32 FILLER_226_2724 ();
 FILLCELL_X32 FILLER_226_2756 ();
 FILLCELL_X32 FILLER_226_2788 ();
 FILLCELL_X32 FILLER_226_2820 ();
 FILLCELL_X32 FILLER_226_2852 ();
 FILLCELL_X32 FILLER_226_2884 ();
 FILLCELL_X32 FILLER_226_2916 ();
 FILLCELL_X32 FILLER_226_2948 ();
 FILLCELL_X32 FILLER_226_2980 ();
 FILLCELL_X32 FILLER_226_3012 ();
 FILLCELL_X32 FILLER_226_3044 ();
 FILLCELL_X32 FILLER_226_3076 ();
 FILLCELL_X32 FILLER_226_3108 ();
 FILLCELL_X16 FILLER_226_3140 ();
 FILLCELL_X1 FILLER_226_3156 ();
 FILLCELL_X32 FILLER_226_3158 ();
 FILLCELL_X32 FILLER_226_3190 ();
 FILLCELL_X32 FILLER_226_3222 ();
 FILLCELL_X32 FILLER_226_3254 ();
 FILLCELL_X32 FILLER_226_3286 ();
 FILLCELL_X32 FILLER_226_3318 ();
 FILLCELL_X32 FILLER_226_3350 ();
 FILLCELL_X32 FILLER_226_3382 ();
 FILLCELL_X32 FILLER_226_3414 ();
 FILLCELL_X32 FILLER_226_3446 ();
 FILLCELL_X32 FILLER_226_3478 ();
 FILLCELL_X32 FILLER_226_3510 ();
 FILLCELL_X32 FILLER_226_3542 ();
 FILLCELL_X32 FILLER_226_3574 ();
 FILLCELL_X32 FILLER_226_3606 ();
 FILLCELL_X32 FILLER_226_3638 ();
 FILLCELL_X32 FILLER_226_3670 ();
 FILLCELL_X32 FILLER_226_3702 ();
 FILLCELL_X4 FILLER_226_3734 ();
 FILLCELL_X32 FILLER_227_1 ();
 FILLCELL_X32 FILLER_227_33 ();
 FILLCELL_X32 FILLER_227_65 ();
 FILLCELL_X32 FILLER_227_97 ();
 FILLCELL_X32 FILLER_227_129 ();
 FILLCELL_X32 FILLER_227_161 ();
 FILLCELL_X32 FILLER_227_193 ();
 FILLCELL_X32 FILLER_227_225 ();
 FILLCELL_X32 FILLER_227_257 ();
 FILLCELL_X32 FILLER_227_289 ();
 FILLCELL_X32 FILLER_227_321 ();
 FILLCELL_X32 FILLER_227_353 ();
 FILLCELL_X32 FILLER_227_385 ();
 FILLCELL_X32 FILLER_227_417 ();
 FILLCELL_X32 FILLER_227_449 ();
 FILLCELL_X32 FILLER_227_481 ();
 FILLCELL_X32 FILLER_227_513 ();
 FILLCELL_X32 FILLER_227_545 ();
 FILLCELL_X32 FILLER_227_577 ();
 FILLCELL_X32 FILLER_227_609 ();
 FILLCELL_X32 FILLER_227_641 ();
 FILLCELL_X32 FILLER_227_673 ();
 FILLCELL_X32 FILLER_227_705 ();
 FILLCELL_X32 FILLER_227_737 ();
 FILLCELL_X32 FILLER_227_769 ();
 FILLCELL_X32 FILLER_227_801 ();
 FILLCELL_X32 FILLER_227_833 ();
 FILLCELL_X32 FILLER_227_865 ();
 FILLCELL_X32 FILLER_227_897 ();
 FILLCELL_X32 FILLER_227_929 ();
 FILLCELL_X32 FILLER_227_961 ();
 FILLCELL_X32 FILLER_227_993 ();
 FILLCELL_X32 FILLER_227_1025 ();
 FILLCELL_X32 FILLER_227_1057 ();
 FILLCELL_X32 FILLER_227_1089 ();
 FILLCELL_X32 FILLER_227_1121 ();
 FILLCELL_X32 FILLER_227_1153 ();
 FILLCELL_X32 FILLER_227_1185 ();
 FILLCELL_X32 FILLER_227_1217 ();
 FILLCELL_X8 FILLER_227_1249 ();
 FILLCELL_X4 FILLER_227_1257 ();
 FILLCELL_X2 FILLER_227_1261 ();
 FILLCELL_X32 FILLER_227_1264 ();
 FILLCELL_X32 FILLER_227_1296 ();
 FILLCELL_X32 FILLER_227_1328 ();
 FILLCELL_X32 FILLER_227_1360 ();
 FILLCELL_X32 FILLER_227_1392 ();
 FILLCELL_X32 FILLER_227_1424 ();
 FILLCELL_X32 FILLER_227_1456 ();
 FILLCELL_X32 FILLER_227_1488 ();
 FILLCELL_X32 FILLER_227_1520 ();
 FILLCELL_X32 FILLER_227_1552 ();
 FILLCELL_X32 FILLER_227_1584 ();
 FILLCELL_X32 FILLER_227_1616 ();
 FILLCELL_X32 FILLER_227_1648 ();
 FILLCELL_X32 FILLER_227_1680 ();
 FILLCELL_X32 FILLER_227_1712 ();
 FILLCELL_X32 FILLER_227_1744 ();
 FILLCELL_X32 FILLER_227_1776 ();
 FILLCELL_X32 FILLER_227_1808 ();
 FILLCELL_X32 FILLER_227_1840 ();
 FILLCELL_X16 FILLER_227_1872 ();
 FILLCELL_X1 FILLER_227_1888 ();
 FILLCELL_X1 FILLER_227_1898 ();
 FILLCELL_X32 FILLER_227_1904 ();
 FILLCELL_X32 FILLER_227_1936 ();
 FILLCELL_X32 FILLER_227_1968 ();
 FILLCELL_X8 FILLER_227_2000 ();
 FILLCELL_X4 FILLER_227_2008 ();
 FILLCELL_X32 FILLER_227_2025 ();
 FILLCELL_X32 FILLER_227_2057 ();
 FILLCELL_X32 FILLER_227_2089 ();
 FILLCELL_X32 FILLER_227_2121 ();
 FILLCELL_X32 FILLER_227_2153 ();
 FILLCELL_X32 FILLER_227_2185 ();
 FILLCELL_X32 FILLER_227_2217 ();
 FILLCELL_X32 FILLER_227_2249 ();
 FILLCELL_X32 FILLER_227_2281 ();
 FILLCELL_X32 FILLER_227_2313 ();
 FILLCELL_X32 FILLER_227_2345 ();
 FILLCELL_X32 FILLER_227_2377 ();
 FILLCELL_X32 FILLER_227_2409 ();
 FILLCELL_X32 FILLER_227_2441 ();
 FILLCELL_X32 FILLER_227_2473 ();
 FILLCELL_X16 FILLER_227_2505 ();
 FILLCELL_X4 FILLER_227_2521 ();
 FILLCELL_X1 FILLER_227_2525 ();
 FILLCELL_X32 FILLER_227_2527 ();
 FILLCELL_X32 FILLER_227_2559 ();
 FILLCELL_X32 FILLER_227_2591 ();
 FILLCELL_X32 FILLER_227_2623 ();
 FILLCELL_X32 FILLER_227_2655 ();
 FILLCELL_X32 FILLER_227_2687 ();
 FILLCELL_X32 FILLER_227_2719 ();
 FILLCELL_X32 FILLER_227_2751 ();
 FILLCELL_X32 FILLER_227_2783 ();
 FILLCELL_X32 FILLER_227_2815 ();
 FILLCELL_X32 FILLER_227_2847 ();
 FILLCELL_X32 FILLER_227_2879 ();
 FILLCELL_X32 FILLER_227_2911 ();
 FILLCELL_X32 FILLER_227_2943 ();
 FILLCELL_X32 FILLER_227_2975 ();
 FILLCELL_X32 FILLER_227_3007 ();
 FILLCELL_X32 FILLER_227_3039 ();
 FILLCELL_X32 FILLER_227_3071 ();
 FILLCELL_X32 FILLER_227_3103 ();
 FILLCELL_X32 FILLER_227_3135 ();
 FILLCELL_X32 FILLER_227_3167 ();
 FILLCELL_X32 FILLER_227_3199 ();
 FILLCELL_X32 FILLER_227_3231 ();
 FILLCELL_X32 FILLER_227_3263 ();
 FILLCELL_X32 FILLER_227_3295 ();
 FILLCELL_X32 FILLER_227_3327 ();
 FILLCELL_X32 FILLER_227_3359 ();
 FILLCELL_X32 FILLER_227_3391 ();
 FILLCELL_X32 FILLER_227_3423 ();
 FILLCELL_X32 FILLER_227_3455 ();
 FILLCELL_X32 FILLER_227_3487 ();
 FILLCELL_X32 FILLER_227_3519 ();
 FILLCELL_X32 FILLER_227_3551 ();
 FILLCELL_X32 FILLER_227_3583 ();
 FILLCELL_X32 FILLER_227_3615 ();
 FILLCELL_X32 FILLER_227_3647 ();
 FILLCELL_X32 FILLER_227_3679 ();
 FILLCELL_X16 FILLER_227_3711 ();
 FILLCELL_X8 FILLER_227_3727 ();
 FILLCELL_X2 FILLER_227_3735 ();
 FILLCELL_X1 FILLER_227_3737 ();
 FILLCELL_X32 FILLER_228_1 ();
 FILLCELL_X32 FILLER_228_33 ();
 FILLCELL_X32 FILLER_228_65 ();
 FILLCELL_X32 FILLER_228_97 ();
 FILLCELL_X32 FILLER_228_129 ();
 FILLCELL_X32 FILLER_228_161 ();
 FILLCELL_X32 FILLER_228_193 ();
 FILLCELL_X32 FILLER_228_225 ();
 FILLCELL_X32 FILLER_228_257 ();
 FILLCELL_X32 FILLER_228_289 ();
 FILLCELL_X32 FILLER_228_321 ();
 FILLCELL_X32 FILLER_228_353 ();
 FILLCELL_X32 FILLER_228_385 ();
 FILLCELL_X32 FILLER_228_417 ();
 FILLCELL_X32 FILLER_228_449 ();
 FILLCELL_X32 FILLER_228_481 ();
 FILLCELL_X32 FILLER_228_513 ();
 FILLCELL_X32 FILLER_228_545 ();
 FILLCELL_X32 FILLER_228_577 ();
 FILLCELL_X16 FILLER_228_609 ();
 FILLCELL_X4 FILLER_228_625 ();
 FILLCELL_X2 FILLER_228_629 ();
 FILLCELL_X32 FILLER_228_632 ();
 FILLCELL_X32 FILLER_228_664 ();
 FILLCELL_X32 FILLER_228_696 ();
 FILLCELL_X32 FILLER_228_728 ();
 FILLCELL_X32 FILLER_228_760 ();
 FILLCELL_X32 FILLER_228_792 ();
 FILLCELL_X32 FILLER_228_824 ();
 FILLCELL_X32 FILLER_228_856 ();
 FILLCELL_X32 FILLER_228_888 ();
 FILLCELL_X32 FILLER_228_920 ();
 FILLCELL_X32 FILLER_228_952 ();
 FILLCELL_X32 FILLER_228_984 ();
 FILLCELL_X32 FILLER_228_1016 ();
 FILLCELL_X32 FILLER_228_1048 ();
 FILLCELL_X32 FILLER_228_1080 ();
 FILLCELL_X32 FILLER_228_1112 ();
 FILLCELL_X32 FILLER_228_1144 ();
 FILLCELL_X32 FILLER_228_1176 ();
 FILLCELL_X32 FILLER_228_1208 ();
 FILLCELL_X32 FILLER_228_1240 ();
 FILLCELL_X32 FILLER_228_1272 ();
 FILLCELL_X32 FILLER_228_1304 ();
 FILLCELL_X32 FILLER_228_1336 ();
 FILLCELL_X32 FILLER_228_1368 ();
 FILLCELL_X32 FILLER_228_1400 ();
 FILLCELL_X32 FILLER_228_1432 ();
 FILLCELL_X32 FILLER_228_1464 ();
 FILLCELL_X32 FILLER_228_1496 ();
 FILLCELL_X32 FILLER_228_1528 ();
 FILLCELL_X32 FILLER_228_1560 ();
 FILLCELL_X32 FILLER_228_1592 ();
 FILLCELL_X32 FILLER_228_1624 ();
 FILLCELL_X32 FILLER_228_1656 ();
 FILLCELL_X32 FILLER_228_1688 ();
 FILLCELL_X32 FILLER_228_1720 ();
 FILLCELL_X32 FILLER_228_1752 ();
 FILLCELL_X32 FILLER_228_1784 ();
 FILLCELL_X32 FILLER_228_1816 ();
 FILLCELL_X32 FILLER_228_1848 ();
 FILLCELL_X2 FILLER_228_1880 ();
 FILLCELL_X1 FILLER_228_1882 ();
 FILLCELL_X4 FILLER_228_1888 ();
 FILLCELL_X2 FILLER_228_1892 ();
 FILLCELL_X32 FILLER_228_1895 ();
 FILLCELL_X32 FILLER_228_1927 ();
 FILLCELL_X32 FILLER_228_1959 ();
 FILLCELL_X32 FILLER_228_1991 ();
 FILLCELL_X32 FILLER_228_2023 ();
 FILLCELL_X32 FILLER_228_2055 ();
 FILLCELL_X32 FILLER_228_2087 ();
 FILLCELL_X32 FILLER_228_2119 ();
 FILLCELL_X32 FILLER_228_2151 ();
 FILLCELL_X32 FILLER_228_2183 ();
 FILLCELL_X32 FILLER_228_2215 ();
 FILLCELL_X32 FILLER_228_2247 ();
 FILLCELL_X32 FILLER_228_2279 ();
 FILLCELL_X32 FILLER_228_2311 ();
 FILLCELL_X32 FILLER_228_2343 ();
 FILLCELL_X32 FILLER_228_2375 ();
 FILLCELL_X32 FILLER_228_2407 ();
 FILLCELL_X32 FILLER_228_2439 ();
 FILLCELL_X32 FILLER_228_2471 ();
 FILLCELL_X32 FILLER_228_2503 ();
 FILLCELL_X32 FILLER_228_2535 ();
 FILLCELL_X32 FILLER_228_2567 ();
 FILLCELL_X32 FILLER_228_2599 ();
 FILLCELL_X32 FILLER_228_2631 ();
 FILLCELL_X32 FILLER_228_2663 ();
 FILLCELL_X32 FILLER_228_2695 ();
 FILLCELL_X32 FILLER_228_2727 ();
 FILLCELL_X32 FILLER_228_2759 ();
 FILLCELL_X32 FILLER_228_2791 ();
 FILLCELL_X32 FILLER_228_2823 ();
 FILLCELL_X32 FILLER_228_2855 ();
 FILLCELL_X32 FILLER_228_2887 ();
 FILLCELL_X32 FILLER_228_2919 ();
 FILLCELL_X32 FILLER_228_2951 ();
 FILLCELL_X32 FILLER_228_2983 ();
 FILLCELL_X32 FILLER_228_3015 ();
 FILLCELL_X32 FILLER_228_3047 ();
 FILLCELL_X32 FILLER_228_3079 ();
 FILLCELL_X32 FILLER_228_3111 ();
 FILLCELL_X8 FILLER_228_3143 ();
 FILLCELL_X4 FILLER_228_3151 ();
 FILLCELL_X2 FILLER_228_3155 ();
 FILLCELL_X32 FILLER_228_3158 ();
 FILLCELL_X32 FILLER_228_3190 ();
 FILLCELL_X32 FILLER_228_3222 ();
 FILLCELL_X32 FILLER_228_3254 ();
 FILLCELL_X32 FILLER_228_3286 ();
 FILLCELL_X32 FILLER_228_3318 ();
 FILLCELL_X32 FILLER_228_3350 ();
 FILLCELL_X32 FILLER_228_3382 ();
 FILLCELL_X32 FILLER_228_3414 ();
 FILLCELL_X32 FILLER_228_3446 ();
 FILLCELL_X32 FILLER_228_3478 ();
 FILLCELL_X32 FILLER_228_3510 ();
 FILLCELL_X32 FILLER_228_3542 ();
 FILLCELL_X32 FILLER_228_3574 ();
 FILLCELL_X32 FILLER_228_3606 ();
 FILLCELL_X32 FILLER_228_3638 ();
 FILLCELL_X32 FILLER_228_3670 ();
 FILLCELL_X32 FILLER_228_3702 ();
 FILLCELL_X4 FILLER_228_3734 ();
 FILLCELL_X32 FILLER_229_1 ();
 FILLCELL_X32 FILLER_229_33 ();
 FILLCELL_X32 FILLER_229_65 ();
 FILLCELL_X32 FILLER_229_97 ();
 FILLCELL_X32 FILLER_229_129 ();
 FILLCELL_X32 FILLER_229_161 ();
 FILLCELL_X32 FILLER_229_193 ();
 FILLCELL_X32 FILLER_229_225 ();
 FILLCELL_X32 FILLER_229_257 ();
 FILLCELL_X32 FILLER_229_289 ();
 FILLCELL_X32 FILLER_229_321 ();
 FILLCELL_X32 FILLER_229_353 ();
 FILLCELL_X32 FILLER_229_385 ();
 FILLCELL_X32 FILLER_229_417 ();
 FILLCELL_X32 FILLER_229_449 ();
 FILLCELL_X32 FILLER_229_481 ();
 FILLCELL_X32 FILLER_229_513 ();
 FILLCELL_X32 FILLER_229_545 ();
 FILLCELL_X32 FILLER_229_577 ();
 FILLCELL_X32 FILLER_229_609 ();
 FILLCELL_X32 FILLER_229_641 ();
 FILLCELL_X32 FILLER_229_673 ();
 FILLCELL_X32 FILLER_229_705 ();
 FILLCELL_X32 FILLER_229_737 ();
 FILLCELL_X32 FILLER_229_769 ();
 FILLCELL_X32 FILLER_229_801 ();
 FILLCELL_X32 FILLER_229_833 ();
 FILLCELL_X32 FILLER_229_865 ();
 FILLCELL_X32 FILLER_229_897 ();
 FILLCELL_X32 FILLER_229_929 ();
 FILLCELL_X32 FILLER_229_961 ();
 FILLCELL_X32 FILLER_229_993 ();
 FILLCELL_X32 FILLER_229_1025 ();
 FILLCELL_X32 FILLER_229_1057 ();
 FILLCELL_X32 FILLER_229_1089 ();
 FILLCELL_X32 FILLER_229_1121 ();
 FILLCELL_X32 FILLER_229_1153 ();
 FILLCELL_X32 FILLER_229_1185 ();
 FILLCELL_X32 FILLER_229_1217 ();
 FILLCELL_X8 FILLER_229_1249 ();
 FILLCELL_X4 FILLER_229_1257 ();
 FILLCELL_X2 FILLER_229_1261 ();
 FILLCELL_X32 FILLER_229_1264 ();
 FILLCELL_X32 FILLER_229_1296 ();
 FILLCELL_X32 FILLER_229_1328 ();
 FILLCELL_X32 FILLER_229_1360 ();
 FILLCELL_X32 FILLER_229_1392 ();
 FILLCELL_X32 FILLER_229_1424 ();
 FILLCELL_X32 FILLER_229_1456 ();
 FILLCELL_X32 FILLER_229_1488 ();
 FILLCELL_X32 FILLER_229_1520 ();
 FILLCELL_X32 FILLER_229_1552 ();
 FILLCELL_X32 FILLER_229_1584 ();
 FILLCELL_X32 FILLER_229_1616 ();
 FILLCELL_X32 FILLER_229_1648 ();
 FILLCELL_X32 FILLER_229_1680 ();
 FILLCELL_X32 FILLER_229_1712 ();
 FILLCELL_X32 FILLER_229_1744 ();
 FILLCELL_X32 FILLER_229_1776 ();
 FILLCELL_X32 FILLER_229_1808 ();
 FILLCELL_X32 FILLER_229_1840 ();
 FILLCELL_X8 FILLER_229_1872 ();
 FILLCELL_X2 FILLER_229_1880 ();
 FILLCELL_X1 FILLER_229_1882 ();
 FILLCELL_X32 FILLER_229_1905 ();
 FILLCELL_X32 FILLER_229_1937 ();
 FILLCELL_X32 FILLER_229_1969 ();
 FILLCELL_X32 FILLER_229_2001 ();
 FILLCELL_X32 FILLER_229_2033 ();
 FILLCELL_X32 FILLER_229_2065 ();
 FILLCELL_X32 FILLER_229_2097 ();
 FILLCELL_X32 FILLER_229_2129 ();
 FILLCELL_X32 FILLER_229_2161 ();
 FILLCELL_X32 FILLER_229_2193 ();
 FILLCELL_X32 FILLER_229_2225 ();
 FILLCELL_X32 FILLER_229_2257 ();
 FILLCELL_X32 FILLER_229_2289 ();
 FILLCELL_X32 FILLER_229_2321 ();
 FILLCELL_X32 FILLER_229_2353 ();
 FILLCELL_X32 FILLER_229_2385 ();
 FILLCELL_X32 FILLER_229_2417 ();
 FILLCELL_X32 FILLER_229_2449 ();
 FILLCELL_X32 FILLER_229_2481 ();
 FILLCELL_X8 FILLER_229_2513 ();
 FILLCELL_X4 FILLER_229_2521 ();
 FILLCELL_X1 FILLER_229_2525 ();
 FILLCELL_X32 FILLER_229_2527 ();
 FILLCELL_X32 FILLER_229_2559 ();
 FILLCELL_X32 FILLER_229_2591 ();
 FILLCELL_X32 FILLER_229_2623 ();
 FILLCELL_X32 FILLER_229_2655 ();
 FILLCELL_X32 FILLER_229_2687 ();
 FILLCELL_X32 FILLER_229_2719 ();
 FILLCELL_X32 FILLER_229_2751 ();
 FILLCELL_X32 FILLER_229_2783 ();
 FILLCELL_X32 FILLER_229_2815 ();
 FILLCELL_X32 FILLER_229_2847 ();
 FILLCELL_X32 FILLER_229_2879 ();
 FILLCELL_X32 FILLER_229_2911 ();
 FILLCELL_X32 FILLER_229_2943 ();
 FILLCELL_X32 FILLER_229_2975 ();
 FILLCELL_X32 FILLER_229_3007 ();
 FILLCELL_X32 FILLER_229_3039 ();
 FILLCELL_X32 FILLER_229_3071 ();
 FILLCELL_X32 FILLER_229_3103 ();
 FILLCELL_X32 FILLER_229_3135 ();
 FILLCELL_X32 FILLER_229_3167 ();
 FILLCELL_X32 FILLER_229_3199 ();
 FILLCELL_X32 FILLER_229_3231 ();
 FILLCELL_X32 FILLER_229_3263 ();
 FILLCELL_X32 FILLER_229_3295 ();
 FILLCELL_X32 FILLER_229_3327 ();
 FILLCELL_X32 FILLER_229_3359 ();
 FILLCELL_X32 FILLER_229_3391 ();
 FILLCELL_X32 FILLER_229_3423 ();
 FILLCELL_X32 FILLER_229_3455 ();
 FILLCELL_X32 FILLER_229_3487 ();
 FILLCELL_X32 FILLER_229_3519 ();
 FILLCELL_X32 FILLER_229_3551 ();
 FILLCELL_X32 FILLER_229_3583 ();
 FILLCELL_X32 FILLER_229_3615 ();
 FILLCELL_X32 FILLER_229_3647 ();
 FILLCELL_X32 FILLER_229_3679 ();
 FILLCELL_X16 FILLER_229_3711 ();
 FILLCELL_X8 FILLER_229_3727 ();
 FILLCELL_X2 FILLER_229_3735 ();
 FILLCELL_X1 FILLER_229_3737 ();
 FILLCELL_X32 FILLER_230_1 ();
 FILLCELL_X32 FILLER_230_33 ();
 FILLCELL_X32 FILLER_230_65 ();
 FILLCELL_X32 FILLER_230_97 ();
 FILLCELL_X32 FILLER_230_129 ();
 FILLCELL_X32 FILLER_230_161 ();
 FILLCELL_X32 FILLER_230_193 ();
 FILLCELL_X32 FILLER_230_225 ();
 FILLCELL_X32 FILLER_230_257 ();
 FILLCELL_X32 FILLER_230_289 ();
 FILLCELL_X32 FILLER_230_321 ();
 FILLCELL_X32 FILLER_230_353 ();
 FILLCELL_X32 FILLER_230_385 ();
 FILLCELL_X32 FILLER_230_417 ();
 FILLCELL_X32 FILLER_230_449 ();
 FILLCELL_X32 FILLER_230_481 ();
 FILLCELL_X32 FILLER_230_513 ();
 FILLCELL_X32 FILLER_230_545 ();
 FILLCELL_X32 FILLER_230_577 ();
 FILLCELL_X16 FILLER_230_609 ();
 FILLCELL_X4 FILLER_230_625 ();
 FILLCELL_X2 FILLER_230_629 ();
 FILLCELL_X32 FILLER_230_632 ();
 FILLCELL_X32 FILLER_230_664 ();
 FILLCELL_X32 FILLER_230_696 ();
 FILLCELL_X32 FILLER_230_728 ();
 FILLCELL_X32 FILLER_230_760 ();
 FILLCELL_X32 FILLER_230_792 ();
 FILLCELL_X32 FILLER_230_824 ();
 FILLCELL_X32 FILLER_230_856 ();
 FILLCELL_X32 FILLER_230_888 ();
 FILLCELL_X32 FILLER_230_920 ();
 FILLCELL_X32 FILLER_230_952 ();
 FILLCELL_X32 FILLER_230_984 ();
 FILLCELL_X32 FILLER_230_1016 ();
 FILLCELL_X32 FILLER_230_1048 ();
 FILLCELL_X32 FILLER_230_1080 ();
 FILLCELL_X32 FILLER_230_1112 ();
 FILLCELL_X32 FILLER_230_1144 ();
 FILLCELL_X32 FILLER_230_1176 ();
 FILLCELL_X32 FILLER_230_1208 ();
 FILLCELL_X32 FILLER_230_1240 ();
 FILLCELL_X32 FILLER_230_1272 ();
 FILLCELL_X32 FILLER_230_1304 ();
 FILLCELL_X32 FILLER_230_1336 ();
 FILLCELL_X32 FILLER_230_1368 ();
 FILLCELL_X32 FILLER_230_1400 ();
 FILLCELL_X32 FILLER_230_1432 ();
 FILLCELL_X32 FILLER_230_1464 ();
 FILLCELL_X32 FILLER_230_1496 ();
 FILLCELL_X32 FILLER_230_1528 ();
 FILLCELL_X32 FILLER_230_1560 ();
 FILLCELL_X32 FILLER_230_1592 ();
 FILLCELL_X32 FILLER_230_1624 ();
 FILLCELL_X32 FILLER_230_1656 ();
 FILLCELL_X32 FILLER_230_1688 ();
 FILLCELL_X32 FILLER_230_1720 ();
 FILLCELL_X32 FILLER_230_1752 ();
 FILLCELL_X32 FILLER_230_1784 ();
 FILLCELL_X32 FILLER_230_1816 ();
 FILLCELL_X16 FILLER_230_1848 ();
 FILLCELL_X8 FILLER_230_1864 ();
 FILLCELL_X4 FILLER_230_1872 ();
 FILLCELL_X2 FILLER_230_1876 ();
 FILLCELL_X1 FILLER_230_1878 ();
 FILLCELL_X4 FILLER_230_1890 ();
 FILLCELL_X1 FILLER_230_1895 ();
 FILLCELL_X4 FILLER_230_1912 ();
 FILLCELL_X32 FILLER_230_1929 ();
 FILLCELL_X32 FILLER_230_1961 ();
 FILLCELL_X32 FILLER_230_1993 ();
 FILLCELL_X32 FILLER_230_2025 ();
 FILLCELL_X32 FILLER_230_2057 ();
 FILLCELL_X32 FILLER_230_2089 ();
 FILLCELL_X32 FILLER_230_2121 ();
 FILLCELL_X32 FILLER_230_2153 ();
 FILLCELL_X32 FILLER_230_2185 ();
 FILLCELL_X32 FILLER_230_2217 ();
 FILLCELL_X32 FILLER_230_2249 ();
 FILLCELL_X32 FILLER_230_2281 ();
 FILLCELL_X32 FILLER_230_2313 ();
 FILLCELL_X32 FILLER_230_2345 ();
 FILLCELL_X32 FILLER_230_2377 ();
 FILLCELL_X32 FILLER_230_2409 ();
 FILLCELL_X32 FILLER_230_2441 ();
 FILLCELL_X32 FILLER_230_2473 ();
 FILLCELL_X32 FILLER_230_2505 ();
 FILLCELL_X32 FILLER_230_2537 ();
 FILLCELL_X32 FILLER_230_2569 ();
 FILLCELL_X32 FILLER_230_2601 ();
 FILLCELL_X32 FILLER_230_2633 ();
 FILLCELL_X32 FILLER_230_2665 ();
 FILLCELL_X32 FILLER_230_2697 ();
 FILLCELL_X32 FILLER_230_2729 ();
 FILLCELL_X32 FILLER_230_2761 ();
 FILLCELL_X32 FILLER_230_2793 ();
 FILLCELL_X32 FILLER_230_2825 ();
 FILLCELL_X32 FILLER_230_2857 ();
 FILLCELL_X32 FILLER_230_2889 ();
 FILLCELL_X32 FILLER_230_2921 ();
 FILLCELL_X32 FILLER_230_2953 ();
 FILLCELL_X32 FILLER_230_2985 ();
 FILLCELL_X32 FILLER_230_3017 ();
 FILLCELL_X32 FILLER_230_3049 ();
 FILLCELL_X32 FILLER_230_3081 ();
 FILLCELL_X32 FILLER_230_3113 ();
 FILLCELL_X8 FILLER_230_3145 ();
 FILLCELL_X4 FILLER_230_3153 ();
 FILLCELL_X32 FILLER_230_3158 ();
 FILLCELL_X32 FILLER_230_3190 ();
 FILLCELL_X32 FILLER_230_3222 ();
 FILLCELL_X32 FILLER_230_3254 ();
 FILLCELL_X32 FILLER_230_3286 ();
 FILLCELL_X32 FILLER_230_3318 ();
 FILLCELL_X32 FILLER_230_3350 ();
 FILLCELL_X32 FILLER_230_3382 ();
 FILLCELL_X32 FILLER_230_3414 ();
 FILLCELL_X32 FILLER_230_3446 ();
 FILLCELL_X32 FILLER_230_3478 ();
 FILLCELL_X32 FILLER_230_3510 ();
 FILLCELL_X32 FILLER_230_3542 ();
 FILLCELL_X32 FILLER_230_3574 ();
 FILLCELL_X32 FILLER_230_3606 ();
 FILLCELL_X32 FILLER_230_3638 ();
 FILLCELL_X32 FILLER_230_3670 ();
 FILLCELL_X32 FILLER_230_3702 ();
 FILLCELL_X4 FILLER_230_3734 ();
 FILLCELL_X32 FILLER_231_1 ();
 FILLCELL_X32 FILLER_231_33 ();
 FILLCELL_X32 FILLER_231_65 ();
 FILLCELL_X32 FILLER_231_97 ();
 FILLCELL_X32 FILLER_231_129 ();
 FILLCELL_X32 FILLER_231_161 ();
 FILLCELL_X32 FILLER_231_193 ();
 FILLCELL_X32 FILLER_231_225 ();
 FILLCELL_X32 FILLER_231_257 ();
 FILLCELL_X32 FILLER_231_289 ();
 FILLCELL_X32 FILLER_231_321 ();
 FILLCELL_X32 FILLER_231_353 ();
 FILLCELL_X32 FILLER_231_385 ();
 FILLCELL_X32 FILLER_231_417 ();
 FILLCELL_X32 FILLER_231_449 ();
 FILLCELL_X32 FILLER_231_481 ();
 FILLCELL_X32 FILLER_231_513 ();
 FILLCELL_X32 FILLER_231_545 ();
 FILLCELL_X32 FILLER_231_577 ();
 FILLCELL_X32 FILLER_231_609 ();
 FILLCELL_X32 FILLER_231_641 ();
 FILLCELL_X32 FILLER_231_673 ();
 FILLCELL_X32 FILLER_231_705 ();
 FILLCELL_X32 FILLER_231_737 ();
 FILLCELL_X32 FILLER_231_769 ();
 FILLCELL_X32 FILLER_231_801 ();
 FILLCELL_X32 FILLER_231_833 ();
 FILLCELL_X32 FILLER_231_865 ();
 FILLCELL_X32 FILLER_231_897 ();
 FILLCELL_X32 FILLER_231_929 ();
 FILLCELL_X32 FILLER_231_961 ();
 FILLCELL_X32 FILLER_231_993 ();
 FILLCELL_X32 FILLER_231_1025 ();
 FILLCELL_X32 FILLER_231_1057 ();
 FILLCELL_X32 FILLER_231_1089 ();
 FILLCELL_X32 FILLER_231_1121 ();
 FILLCELL_X32 FILLER_231_1153 ();
 FILLCELL_X32 FILLER_231_1185 ();
 FILLCELL_X32 FILLER_231_1217 ();
 FILLCELL_X8 FILLER_231_1249 ();
 FILLCELL_X4 FILLER_231_1257 ();
 FILLCELL_X2 FILLER_231_1261 ();
 FILLCELL_X32 FILLER_231_1264 ();
 FILLCELL_X32 FILLER_231_1296 ();
 FILLCELL_X32 FILLER_231_1328 ();
 FILLCELL_X32 FILLER_231_1360 ();
 FILLCELL_X32 FILLER_231_1392 ();
 FILLCELL_X32 FILLER_231_1424 ();
 FILLCELL_X32 FILLER_231_1456 ();
 FILLCELL_X32 FILLER_231_1488 ();
 FILLCELL_X32 FILLER_231_1520 ();
 FILLCELL_X32 FILLER_231_1552 ();
 FILLCELL_X32 FILLER_231_1584 ();
 FILLCELL_X32 FILLER_231_1616 ();
 FILLCELL_X32 FILLER_231_1648 ();
 FILLCELL_X32 FILLER_231_1680 ();
 FILLCELL_X32 FILLER_231_1712 ();
 FILLCELL_X32 FILLER_231_1744 ();
 FILLCELL_X32 FILLER_231_1776 ();
 FILLCELL_X32 FILLER_231_1808 ();
 FILLCELL_X32 FILLER_231_1840 ();
 FILLCELL_X8 FILLER_231_1872 ();
 FILLCELL_X4 FILLER_231_1880 ();
 FILLCELL_X2 FILLER_231_1884 ();
 FILLCELL_X32 FILLER_231_1891 ();
 FILLCELL_X32 FILLER_231_1923 ();
 FILLCELL_X32 FILLER_231_1955 ();
 FILLCELL_X32 FILLER_231_1987 ();
 FILLCELL_X32 FILLER_231_2019 ();
 FILLCELL_X32 FILLER_231_2051 ();
 FILLCELL_X32 FILLER_231_2083 ();
 FILLCELL_X32 FILLER_231_2115 ();
 FILLCELL_X32 FILLER_231_2147 ();
 FILLCELL_X32 FILLER_231_2179 ();
 FILLCELL_X32 FILLER_231_2211 ();
 FILLCELL_X32 FILLER_231_2243 ();
 FILLCELL_X32 FILLER_231_2275 ();
 FILLCELL_X32 FILLER_231_2307 ();
 FILLCELL_X32 FILLER_231_2339 ();
 FILLCELL_X32 FILLER_231_2371 ();
 FILLCELL_X32 FILLER_231_2403 ();
 FILLCELL_X32 FILLER_231_2435 ();
 FILLCELL_X32 FILLER_231_2467 ();
 FILLCELL_X16 FILLER_231_2499 ();
 FILLCELL_X8 FILLER_231_2515 ();
 FILLCELL_X2 FILLER_231_2523 ();
 FILLCELL_X1 FILLER_231_2525 ();
 FILLCELL_X32 FILLER_231_2527 ();
 FILLCELL_X32 FILLER_231_2559 ();
 FILLCELL_X32 FILLER_231_2591 ();
 FILLCELL_X32 FILLER_231_2623 ();
 FILLCELL_X32 FILLER_231_2655 ();
 FILLCELL_X32 FILLER_231_2687 ();
 FILLCELL_X32 FILLER_231_2719 ();
 FILLCELL_X32 FILLER_231_2751 ();
 FILLCELL_X32 FILLER_231_2783 ();
 FILLCELL_X32 FILLER_231_2815 ();
 FILLCELL_X32 FILLER_231_2847 ();
 FILLCELL_X32 FILLER_231_2879 ();
 FILLCELL_X32 FILLER_231_2911 ();
 FILLCELL_X32 FILLER_231_2943 ();
 FILLCELL_X32 FILLER_231_2975 ();
 FILLCELL_X32 FILLER_231_3007 ();
 FILLCELL_X32 FILLER_231_3039 ();
 FILLCELL_X32 FILLER_231_3071 ();
 FILLCELL_X32 FILLER_231_3103 ();
 FILLCELL_X32 FILLER_231_3135 ();
 FILLCELL_X32 FILLER_231_3167 ();
 FILLCELL_X32 FILLER_231_3199 ();
 FILLCELL_X32 FILLER_231_3231 ();
 FILLCELL_X32 FILLER_231_3263 ();
 FILLCELL_X32 FILLER_231_3295 ();
 FILLCELL_X32 FILLER_231_3327 ();
 FILLCELL_X32 FILLER_231_3359 ();
 FILLCELL_X32 FILLER_231_3391 ();
 FILLCELL_X32 FILLER_231_3423 ();
 FILLCELL_X32 FILLER_231_3455 ();
 FILLCELL_X32 FILLER_231_3487 ();
 FILLCELL_X32 FILLER_231_3519 ();
 FILLCELL_X32 FILLER_231_3551 ();
 FILLCELL_X32 FILLER_231_3583 ();
 FILLCELL_X32 FILLER_231_3615 ();
 FILLCELL_X32 FILLER_231_3647 ();
 FILLCELL_X32 FILLER_231_3679 ();
 FILLCELL_X16 FILLER_231_3711 ();
 FILLCELL_X8 FILLER_231_3727 ();
 FILLCELL_X2 FILLER_231_3735 ();
 FILLCELL_X1 FILLER_231_3737 ();
 FILLCELL_X32 FILLER_232_1 ();
 FILLCELL_X32 FILLER_232_33 ();
 FILLCELL_X32 FILLER_232_65 ();
 FILLCELL_X32 FILLER_232_97 ();
 FILLCELL_X32 FILLER_232_129 ();
 FILLCELL_X32 FILLER_232_161 ();
 FILLCELL_X32 FILLER_232_193 ();
 FILLCELL_X32 FILLER_232_225 ();
 FILLCELL_X32 FILLER_232_257 ();
 FILLCELL_X32 FILLER_232_289 ();
 FILLCELL_X32 FILLER_232_321 ();
 FILLCELL_X32 FILLER_232_353 ();
 FILLCELL_X32 FILLER_232_385 ();
 FILLCELL_X32 FILLER_232_417 ();
 FILLCELL_X32 FILLER_232_449 ();
 FILLCELL_X32 FILLER_232_481 ();
 FILLCELL_X32 FILLER_232_513 ();
 FILLCELL_X32 FILLER_232_545 ();
 FILLCELL_X32 FILLER_232_577 ();
 FILLCELL_X16 FILLER_232_609 ();
 FILLCELL_X4 FILLER_232_625 ();
 FILLCELL_X2 FILLER_232_629 ();
 FILLCELL_X32 FILLER_232_632 ();
 FILLCELL_X32 FILLER_232_664 ();
 FILLCELL_X32 FILLER_232_696 ();
 FILLCELL_X32 FILLER_232_728 ();
 FILLCELL_X32 FILLER_232_760 ();
 FILLCELL_X32 FILLER_232_792 ();
 FILLCELL_X32 FILLER_232_824 ();
 FILLCELL_X32 FILLER_232_856 ();
 FILLCELL_X32 FILLER_232_888 ();
 FILLCELL_X32 FILLER_232_920 ();
 FILLCELL_X32 FILLER_232_952 ();
 FILLCELL_X32 FILLER_232_984 ();
 FILLCELL_X32 FILLER_232_1016 ();
 FILLCELL_X32 FILLER_232_1048 ();
 FILLCELL_X32 FILLER_232_1080 ();
 FILLCELL_X32 FILLER_232_1112 ();
 FILLCELL_X32 FILLER_232_1144 ();
 FILLCELL_X32 FILLER_232_1176 ();
 FILLCELL_X32 FILLER_232_1208 ();
 FILLCELL_X32 FILLER_232_1240 ();
 FILLCELL_X32 FILLER_232_1272 ();
 FILLCELL_X32 FILLER_232_1304 ();
 FILLCELL_X32 FILLER_232_1336 ();
 FILLCELL_X32 FILLER_232_1368 ();
 FILLCELL_X32 FILLER_232_1400 ();
 FILLCELL_X32 FILLER_232_1432 ();
 FILLCELL_X32 FILLER_232_1464 ();
 FILLCELL_X32 FILLER_232_1496 ();
 FILLCELL_X32 FILLER_232_1528 ();
 FILLCELL_X32 FILLER_232_1560 ();
 FILLCELL_X32 FILLER_232_1592 ();
 FILLCELL_X32 FILLER_232_1624 ();
 FILLCELL_X32 FILLER_232_1656 ();
 FILLCELL_X32 FILLER_232_1688 ();
 FILLCELL_X32 FILLER_232_1720 ();
 FILLCELL_X32 FILLER_232_1752 ();
 FILLCELL_X32 FILLER_232_1784 ();
 FILLCELL_X32 FILLER_232_1816 ();
 FILLCELL_X16 FILLER_232_1848 ();
 FILLCELL_X8 FILLER_232_1864 ();
 FILLCELL_X4 FILLER_232_1872 ();
 FILLCELL_X1 FILLER_232_1876 ();
 FILLCELL_X4 FILLER_232_1887 ();
 FILLCELL_X2 FILLER_232_1891 ();
 FILLCELL_X1 FILLER_232_1893 ();
 FILLCELL_X32 FILLER_232_1895 ();
 FILLCELL_X32 FILLER_232_1927 ();
 FILLCELL_X32 FILLER_232_1959 ();
 FILLCELL_X32 FILLER_232_1991 ();
 FILLCELL_X32 FILLER_232_2023 ();
 FILLCELL_X32 FILLER_232_2055 ();
 FILLCELL_X8 FILLER_232_2087 ();
 FILLCELL_X4 FILLER_232_2095 ();
 FILLCELL_X2 FILLER_232_2099 ();
 FILLCELL_X1 FILLER_232_2101 ();
 FILLCELL_X32 FILLER_232_2119 ();
 FILLCELL_X32 FILLER_232_2151 ();
 FILLCELL_X32 FILLER_232_2183 ();
 FILLCELL_X32 FILLER_232_2215 ();
 FILLCELL_X32 FILLER_232_2247 ();
 FILLCELL_X32 FILLER_232_2279 ();
 FILLCELL_X32 FILLER_232_2311 ();
 FILLCELL_X32 FILLER_232_2343 ();
 FILLCELL_X32 FILLER_232_2375 ();
 FILLCELL_X32 FILLER_232_2407 ();
 FILLCELL_X32 FILLER_232_2439 ();
 FILLCELL_X32 FILLER_232_2471 ();
 FILLCELL_X32 FILLER_232_2503 ();
 FILLCELL_X32 FILLER_232_2535 ();
 FILLCELL_X32 FILLER_232_2567 ();
 FILLCELL_X32 FILLER_232_2599 ();
 FILLCELL_X32 FILLER_232_2631 ();
 FILLCELL_X32 FILLER_232_2663 ();
 FILLCELL_X32 FILLER_232_2695 ();
 FILLCELL_X32 FILLER_232_2727 ();
 FILLCELL_X32 FILLER_232_2759 ();
 FILLCELL_X32 FILLER_232_2791 ();
 FILLCELL_X32 FILLER_232_2823 ();
 FILLCELL_X32 FILLER_232_2855 ();
 FILLCELL_X32 FILLER_232_2887 ();
 FILLCELL_X32 FILLER_232_2919 ();
 FILLCELL_X32 FILLER_232_2951 ();
 FILLCELL_X32 FILLER_232_2983 ();
 FILLCELL_X32 FILLER_232_3015 ();
 FILLCELL_X32 FILLER_232_3047 ();
 FILLCELL_X32 FILLER_232_3079 ();
 FILLCELL_X32 FILLER_232_3111 ();
 FILLCELL_X8 FILLER_232_3143 ();
 FILLCELL_X4 FILLER_232_3151 ();
 FILLCELL_X2 FILLER_232_3155 ();
 FILLCELL_X32 FILLER_232_3158 ();
 FILLCELL_X32 FILLER_232_3190 ();
 FILLCELL_X32 FILLER_232_3222 ();
 FILLCELL_X32 FILLER_232_3254 ();
 FILLCELL_X32 FILLER_232_3286 ();
 FILLCELL_X32 FILLER_232_3318 ();
 FILLCELL_X32 FILLER_232_3350 ();
 FILLCELL_X32 FILLER_232_3382 ();
 FILLCELL_X32 FILLER_232_3414 ();
 FILLCELL_X32 FILLER_232_3446 ();
 FILLCELL_X32 FILLER_232_3478 ();
 FILLCELL_X32 FILLER_232_3510 ();
 FILLCELL_X32 FILLER_232_3542 ();
 FILLCELL_X32 FILLER_232_3574 ();
 FILLCELL_X32 FILLER_232_3606 ();
 FILLCELL_X32 FILLER_232_3638 ();
 FILLCELL_X32 FILLER_232_3670 ();
 FILLCELL_X32 FILLER_232_3702 ();
 FILLCELL_X4 FILLER_232_3734 ();
 FILLCELL_X32 FILLER_233_1 ();
 FILLCELL_X32 FILLER_233_33 ();
 FILLCELL_X32 FILLER_233_65 ();
 FILLCELL_X32 FILLER_233_97 ();
 FILLCELL_X32 FILLER_233_129 ();
 FILLCELL_X32 FILLER_233_161 ();
 FILLCELL_X32 FILLER_233_193 ();
 FILLCELL_X32 FILLER_233_225 ();
 FILLCELL_X32 FILLER_233_257 ();
 FILLCELL_X32 FILLER_233_289 ();
 FILLCELL_X32 FILLER_233_321 ();
 FILLCELL_X32 FILLER_233_353 ();
 FILLCELL_X32 FILLER_233_385 ();
 FILLCELL_X32 FILLER_233_417 ();
 FILLCELL_X32 FILLER_233_449 ();
 FILLCELL_X32 FILLER_233_481 ();
 FILLCELL_X32 FILLER_233_513 ();
 FILLCELL_X32 FILLER_233_545 ();
 FILLCELL_X32 FILLER_233_577 ();
 FILLCELL_X32 FILLER_233_609 ();
 FILLCELL_X32 FILLER_233_641 ();
 FILLCELL_X32 FILLER_233_673 ();
 FILLCELL_X32 FILLER_233_705 ();
 FILLCELL_X32 FILLER_233_737 ();
 FILLCELL_X32 FILLER_233_769 ();
 FILLCELL_X32 FILLER_233_801 ();
 FILLCELL_X32 FILLER_233_833 ();
 FILLCELL_X32 FILLER_233_865 ();
 FILLCELL_X32 FILLER_233_897 ();
 FILLCELL_X32 FILLER_233_929 ();
 FILLCELL_X32 FILLER_233_961 ();
 FILLCELL_X32 FILLER_233_993 ();
 FILLCELL_X32 FILLER_233_1025 ();
 FILLCELL_X32 FILLER_233_1057 ();
 FILLCELL_X32 FILLER_233_1089 ();
 FILLCELL_X32 FILLER_233_1121 ();
 FILLCELL_X32 FILLER_233_1153 ();
 FILLCELL_X32 FILLER_233_1185 ();
 FILLCELL_X32 FILLER_233_1217 ();
 FILLCELL_X8 FILLER_233_1249 ();
 FILLCELL_X4 FILLER_233_1257 ();
 FILLCELL_X2 FILLER_233_1261 ();
 FILLCELL_X32 FILLER_233_1264 ();
 FILLCELL_X32 FILLER_233_1296 ();
 FILLCELL_X32 FILLER_233_1328 ();
 FILLCELL_X32 FILLER_233_1360 ();
 FILLCELL_X32 FILLER_233_1392 ();
 FILLCELL_X32 FILLER_233_1424 ();
 FILLCELL_X32 FILLER_233_1456 ();
 FILLCELL_X32 FILLER_233_1488 ();
 FILLCELL_X32 FILLER_233_1520 ();
 FILLCELL_X32 FILLER_233_1552 ();
 FILLCELL_X32 FILLER_233_1584 ();
 FILLCELL_X32 FILLER_233_1616 ();
 FILLCELL_X32 FILLER_233_1648 ();
 FILLCELL_X32 FILLER_233_1680 ();
 FILLCELL_X32 FILLER_233_1712 ();
 FILLCELL_X32 FILLER_233_1744 ();
 FILLCELL_X32 FILLER_233_1776 ();
 FILLCELL_X32 FILLER_233_1808 ();
 FILLCELL_X32 FILLER_233_1840 ();
 FILLCELL_X4 FILLER_233_1872 ();
 FILLCELL_X2 FILLER_233_1876 ();
 FILLCELL_X16 FILLER_233_1912 ();
 FILLCELL_X1 FILLER_233_1928 ();
 FILLCELL_X32 FILLER_233_1948 ();
 FILLCELL_X32 FILLER_233_1980 ();
 FILLCELL_X32 FILLER_233_2012 ();
 FILLCELL_X32 FILLER_233_2044 ();
 FILLCELL_X32 FILLER_233_2076 ();
 FILLCELL_X8 FILLER_233_2115 ();
 FILLCELL_X2 FILLER_233_2123 ();
 FILLCELL_X16 FILLER_233_2142 ();
 FILLCELL_X4 FILLER_233_2158 ();
 FILLCELL_X32 FILLER_233_2186 ();
 FILLCELL_X32 FILLER_233_2218 ();
 FILLCELL_X32 FILLER_233_2250 ();
 FILLCELL_X32 FILLER_233_2282 ();
 FILLCELL_X32 FILLER_233_2314 ();
 FILLCELL_X32 FILLER_233_2346 ();
 FILLCELL_X32 FILLER_233_2378 ();
 FILLCELL_X32 FILLER_233_2410 ();
 FILLCELL_X32 FILLER_233_2442 ();
 FILLCELL_X32 FILLER_233_2474 ();
 FILLCELL_X16 FILLER_233_2506 ();
 FILLCELL_X4 FILLER_233_2522 ();
 FILLCELL_X32 FILLER_233_2527 ();
 FILLCELL_X32 FILLER_233_2559 ();
 FILLCELL_X32 FILLER_233_2591 ();
 FILLCELL_X32 FILLER_233_2623 ();
 FILLCELL_X32 FILLER_233_2655 ();
 FILLCELL_X32 FILLER_233_2687 ();
 FILLCELL_X32 FILLER_233_2719 ();
 FILLCELL_X32 FILLER_233_2751 ();
 FILLCELL_X32 FILLER_233_2783 ();
 FILLCELL_X32 FILLER_233_2815 ();
 FILLCELL_X32 FILLER_233_2847 ();
 FILLCELL_X32 FILLER_233_2879 ();
 FILLCELL_X32 FILLER_233_2911 ();
 FILLCELL_X32 FILLER_233_2943 ();
 FILLCELL_X32 FILLER_233_2975 ();
 FILLCELL_X32 FILLER_233_3007 ();
 FILLCELL_X32 FILLER_233_3039 ();
 FILLCELL_X32 FILLER_233_3071 ();
 FILLCELL_X32 FILLER_233_3103 ();
 FILLCELL_X32 FILLER_233_3135 ();
 FILLCELL_X32 FILLER_233_3167 ();
 FILLCELL_X32 FILLER_233_3199 ();
 FILLCELL_X32 FILLER_233_3231 ();
 FILLCELL_X32 FILLER_233_3263 ();
 FILLCELL_X32 FILLER_233_3295 ();
 FILLCELL_X32 FILLER_233_3327 ();
 FILLCELL_X32 FILLER_233_3359 ();
 FILLCELL_X32 FILLER_233_3391 ();
 FILLCELL_X32 FILLER_233_3423 ();
 FILLCELL_X32 FILLER_233_3455 ();
 FILLCELL_X32 FILLER_233_3487 ();
 FILLCELL_X32 FILLER_233_3519 ();
 FILLCELL_X32 FILLER_233_3551 ();
 FILLCELL_X32 FILLER_233_3583 ();
 FILLCELL_X32 FILLER_233_3615 ();
 FILLCELL_X32 FILLER_233_3647 ();
 FILLCELL_X32 FILLER_233_3679 ();
 FILLCELL_X16 FILLER_233_3711 ();
 FILLCELL_X8 FILLER_233_3727 ();
 FILLCELL_X2 FILLER_233_3735 ();
 FILLCELL_X1 FILLER_233_3737 ();
 FILLCELL_X32 FILLER_234_1 ();
 FILLCELL_X32 FILLER_234_33 ();
 FILLCELL_X32 FILLER_234_65 ();
 FILLCELL_X32 FILLER_234_97 ();
 FILLCELL_X32 FILLER_234_129 ();
 FILLCELL_X32 FILLER_234_161 ();
 FILLCELL_X32 FILLER_234_193 ();
 FILLCELL_X32 FILLER_234_225 ();
 FILLCELL_X32 FILLER_234_257 ();
 FILLCELL_X32 FILLER_234_289 ();
 FILLCELL_X32 FILLER_234_321 ();
 FILLCELL_X32 FILLER_234_353 ();
 FILLCELL_X32 FILLER_234_385 ();
 FILLCELL_X32 FILLER_234_417 ();
 FILLCELL_X32 FILLER_234_449 ();
 FILLCELL_X32 FILLER_234_481 ();
 FILLCELL_X32 FILLER_234_513 ();
 FILLCELL_X32 FILLER_234_545 ();
 FILLCELL_X32 FILLER_234_577 ();
 FILLCELL_X16 FILLER_234_609 ();
 FILLCELL_X4 FILLER_234_625 ();
 FILLCELL_X2 FILLER_234_629 ();
 FILLCELL_X32 FILLER_234_632 ();
 FILLCELL_X32 FILLER_234_664 ();
 FILLCELL_X32 FILLER_234_696 ();
 FILLCELL_X32 FILLER_234_728 ();
 FILLCELL_X32 FILLER_234_760 ();
 FILLCELL_X32 FILLER_234_792 ();
 FILLCELL_X32 FILLER_234_824 ();
 FILLCELL_X32 FILLER_234_856 ();
 FILLCELL_X32 FILLER_234_888 ();
 FILLCELL_X32 FILLER_234_920 ();
 FILLCELL_X32 FILLER_234_952 ();
 FILLCELL_X32 FILLER_234_984 ();
 FILLCELL_X32 FILLER_234_1016 ();
 FILLCELL_X32 FILLER_234_1048 ();
 FILLCELL_X32 FILLER_234_1080 ();
 FILLCELL_X32 FILLER_234_1112 ();
 FILLCELL_X32 FILLER_234_1144 ();
 FILLCELL_X32 FILLER_234_1176 ();
 FILLCELL_X32 FILLER_234_1208 ();
 FILLCELL_X32 FILLER_234_1240 ();
 FILLCELL_X32 FILLER_234_1272 ();
 FILLCELL_X32 FILLER_234_1304 ();
 FILLCELL_X32 FILLER_234_1336 ();
 FILLCELL_X32 FILLER_234_1368 ();
 FILLCELL_X32 FILLER_234_1400 ();
 FILLCELL_X32 FILLER_234_1432 ();
 FILLCELL_X32 FILLER_234_1464 ();
 FILLCELL_X32 FILLER_234_1496 ();
 FILLCELL_X32 FILLER_234_1528 ();
 FILLCELL_X32 FILLER_234_1560 ();
 FILLCELL_X32 FILLER_234_1592 ();
 FILLCELL_X32 FILLER_234_1624 ();
 FILLCELL_X32 FILLER_234_1656 ();
 FILLCELL_X32 FILLER_234_1688 ();
 FILLCELL_X32 FILLER_234_1720 ();
 FILLCELL_X32 FILLER_234_1752 ();
 FILLCELL_X32 FILLER_234_1784 ();
 FILLCELL_X32 FILLER_234_1816 ();
 FILLCELL_X16 FILLER_234_1848 ();
 FILLCELL_X8 FILLER_234_1864 ();
 FILLCELL_X2 FILLER_234_1872 ();
 FILLCELL_X16 FILLER_234_1878 ();
 FILLCELL_X2 FILLER_234_1895 ();
 FILLCELL_X1 FILLER_234_1897 ();
 FILLCELL_X8 FILLER_234_1909 ();
 FILLCELL_X32 FILLER_234_1927 ();
 FILLCELL_X32 FILLER_234_1959 ();
 FILLCELL_X32 FILLER_234_1991 ();
 FILLCELL_X32 FILLER_234_2023 ();
 FILLCELL_X2 FILLER_234_2055 ();
 FILLCELL_X1 FILLER_234_2057 ();
 FILLCELL_X32 FILLER_234_2075 ();
 FILLCELL_X8 FILLER_234_2107 ();
 FILLCELL_X4 FILLER_234_2115 ();
 FILLCELL_X2 FILLER_234_2119 ();
 FILLCELL_X1 FILLER_234_2121 ();
 FILLCELL_X8 FILLER_234_2136 ();
 FILLCELL_X4 FILLER_234_2144 ();
 FILLCELL_X1 FILLER_234_2148 ();
 FILLCELL_X32 FILLER_234_2204 ();
 FILLCELL_X32 FILLER_234_2236 ();
 FILLCELL_X32 FILLER_234_2268 ();
 FILLCELL_X32 FILLER_234_2300 ();
 FILLCELL_X32 FILLER_234_2332 ();
 FILLCELL_X32 FILLER_234_2364 ();
 FILLCELL_X32 FILLER_234_2396 ();
 FILLCELL_X32 FILLER_234_2428 ();
 FILLCELL_X32 FILLER_234_2460 ();
 FILLCELL_X32 FILLER_234_2492 ();
 FILLCELL_X32 FILLER_234_2524 ();
 FILLCELL_X32 FILLER_234_2556 ();
 FILLCELL_X32 FILLER_234_2588 ();
 FILLCELL_X32 FILLER_234_2620 ();
 FILLCELL_X32 FILLER_234_2652 ();
 FILLCELL_X32 FILLER_234_2684 ();
 FILLCELL_X32 FILLER_234_2716 ();
 FILLCELL_X32 FILLER_234_2748 ();
 FILLCELL_X32 FILLER_234_2780 ();
 FILLCELL_X32 FILLER_234_2812 ();
 FILLCELL_X32 FILLER_234_2844 ();
 FILLCELL_X32 FILLER_234_2876 ();
 FILLCELL_X32 FILLER_234_2908 ();
 FILLCELL_X32 FILLER_234_2940 ();
 FILLCELL_X32 FILLER_234_2972 ();
 FILLCELL_X32 FILLER_234_3004 ();
 FILLCELL_X32 FILLER_234_3036 ();
 FILLCELL_X32 FILLER_234_3068 ();
 FILLCELL_X32 FILLER_234_3100 ();
 FILLCELL_X16 FILLER_234_3132 ();
 FILLCELL_X8 FILLER_234_3148 ();
 FILLCELL_X1 FILLER_234_3156 ();
 FILLCELL_X32 FILLER_234_3158 ();
 FILLCELL_X32 FILLER_234_3190 ();
 FILLCELL_X32 FILLER_234_3222 ();
 FILLCELL_X32 FILLER_234_3254 ();
 FILLCELL_X32 FILLER_234_3286 ();
 FILLCELL_X32 FILLER_234_3318 ();
 FILLCELL_X32 FILLER_234_3350 ();
 FILLCELL_X32 FILLER_234_3382 ();
 FILLCELL_X32 FILLER_234_3414 ();
 FILLCELL_X32 FILLER_234_3446 ();
 FILLCELL_X32 FILLER_234_3478 ();
 FILLCELL_X32 FILLER_234_3510 ();
 FILLCELL_X32 FILLER_234_3542 ();
 FILLCELL_X32 FILLER_234_3574 ();
 FILLCELL_X32 FILLER_234_3606 ();
 FILLCELL_X32 FILLER_234_3638 ();
 FILLCELL_X32 FILLER_234_3670 ();
 FILLCELL_X32 FILLER_234_3702 ();
 FILLCELL_X4 FILLER_234_3734 ();
 FILLCELL_X32 FILLER_235_1 ();
 FILLCELL_X32 FILLER_235_33 ();
 FILLCELL_X32 FILLER_235_65 ();
 FILLCELL_X32 FILLER_235_97 ();
 FILLCELL_X32 FILLER_235_129 ();
 FILLCELL_X32 FILLER_235_161 ();
 FILLCELL_X32 FILLER_235_193 ();
 FILLCELL_X32 FILLER_235_225 ();
 FILLCELL_X32 FILLER_235_257 ();
 FILLCELL_X32 FILLER_235_289 ();
 FILLCELL_X32 FILLER_235_321 ();
 FILLCELL_X32 FILLER_235_353 ();
 FILLCELL_X32 FILLER_235_385 ();
 FILLCELL_X32 FILLER_235_417 ();
 FILLCELL_X32 FILLER_235_449 ();
 FILLCELL_X32 FILLER_235_481 ();
 FILLCELL_X32 FILLER_235_513 ();
 FILLCELL_X32 FILLER_235_545 ();
 FILLCELL_X32 FILLER_235_577 ();
 FILLCELL_X32 FILLER_235_609 ();
 FILLCELL_X32 FILLER_235_641 ();
 FILLCELL_X32 FILLER_235_673 ();
 FILLCELL_X32 FILLER_235_705 ();
 FILLCELL_X32 FILLER_235_737 ();
 FILLCELL_X32 FILLER_235_769 ();
 FILLCELL_X32 FILLER_235_801 ();
 FILLCELL_X32 FILLER_235_833 ();
 FILLCELL_X32 FILLER_235_865 ();
 FILLCELL_X32 FILLER_235_897 ();
 FILLCELL_X32 FILLER_235_929 ();
 FILLCELL_X32 FILLER_235_961 ();
 FILLCELL_X32 FILLER_235_993 ();
 FILLCELL_X32 FILLER_235_1025 ();
 FILLCELL_X32 FILLER_235_1057 ();
 FILLCELL_X32 FILLER_235_1089 ();
 FILLCELL_X32 FILLER_235_1121 ();
 FILLCELL_X32 FILLER_235_1153 ();
 FILLCELL_X32 FILLER_235_1185 ();
 FILLCELL_X32 FILLER_235_1217 ();
 FILLCELL_X8 FILLER_235_1249 ();
 FILLCELL_X4 FILLER_235_1257 ();
 FILLCELL_X2 FILLER_235_1261 ();
 FILLCELL_X32 FILLER_235_1264 ();
 FILLCELL_X32 FILLER_235_1296 ();
 FILLCELL_X32 FILLER_235_1328 ();
 FILLCELL_X32 FILLER_235_1360 ();
 FILLCELL_X32 FILLER_235_1392 ();
 FILLCELL_X32 FILLER_235_1424 ();
 FILLCELL_X32 FILLER_235_1456 ();
 FILLCELL_X32 FILLER_235_1488 ();
 FILLCELL_X32 FILLER_235_1520 ();
 FILLCELL_X32 FILLER_235_1552 ();
 FILLCELL_X32 FILLER_235_1584 ();
 FILLCELL_X32 FILLER_235_1616 ();
 FILLCELL_X32 FILLER_235_1648 ();
 FILLCELL_X32 FILLER_235_1680 ();
 FILLCELL_X32 FILLER_235_1712 ();
 FILLCELL_X32 FILLER_235_1744 ();
 FILLCELL_X32 FILLER_235_1776 ();
 FILLCELL_X32 FILLER_235_1808 ();
 FILLCELL_X16 FILLER_235_1840 ();
 FILLCELL_X8 FILLER_235_1856 ();
 FILLCELL_X1 FILLER_235_1864 ();
 FILLCELL_X8 FILLER_235_1880 ();
 FILLCELL_X4 FILLER_235_1888 ();
 FILLCELL_X2 FILLER_235_1892 ();
 FILLCELL_X16 FILLER_235_1896 ();
 FILLCELL_X8 FILLER_235_1912 ();
 FILLCELL_X4 FILLER_235_1920 ();
 FILLCELL_X2 FILLER_235_1924 ();
 FILLCELL_X32 FILLER_235_1951 ();
 FILLCELL_X32 FILLER_235_1983 ();
 FILLCELL_X16 FILLER_235_2015 ();
 FILLCELL_X8 FILLER_235_2031 ();
 FILLCELL_X4 FILLER_235_2039 ();
 FILLCELL_X8 FILLER_235_2050 ();
 FILLCELL_X4 FILLER_235_2058 ();
 FILLCELL_X32 FILLER_235_2076 ();
 FILLCELL_X32 FILLER_235_2108 ();
 FILLCELL_X32 FILLER_235_2140 ();
 FILLCELL_X32 FILLER_235_2172 ();
 FILLCELL_X16 FILLER_235_2204 ();
 FILLCELL_X1 FILLER_235_2220 ();
 FILLCELL_X32 FILLER_235_2245 ();
 FILLCELL_X32 FILLER_235_2277 ();
 FILLCELL_X32 FILLER_235_2309 ();
 FILLCELL_X32 FILLER_235_2341 ();
 FILLCELL_X32 FILLER_235_2373 ();
 FILLCELL_X32 FILLER_235_2405 ();
 FILLCELL_X32 FILLER_235_2437 ();
 FILLCELL_X32 FILLER_235_2469 ();
 FILLCELL_X16 FILLER_235_2501 ();
 FILLCELL_X8 FILLER_235_2517 ();
 FILLCELL_X1 FILLER_235_2525 ();
 FILLCELL_X32 FILLER_235_2527 ();
 FILLCELL_X32 FILLER_235_2559 ();
 FILLCELL_X32 FILLER_235_2591 ();
 FILLCELL_X32 FILLER_235_2623 ();
 FILLCELL_X32 FILLER_235_2655 ();
 FILLCELL_X32 FILLER_235_2687 ();
 FILLCELL_X32 FILLER_235_2719 ();
 FILLCELL_X32 FILLER_235_2751 ();
 FILLCELL_X32 FILLER_235_2783 ();
 FILLCELL_X32 FILLER_235_2815 ();
 FILLCELL_X32 FILLER_235_2847 ();
 FILLCELL_X32 FILLER_235_2879 ();
 FILLCELL_X32 FILLER_235_2911 ();
 FILLCELL_X32 FILLER_235_2943 ();
 FILLCELL_X32 FILLER_235_2975 ();
 FILLCELL_X32 FILLER_235_3007 ();
 FILLCELL_X32 FILLER_235_3039 ();
 FILLCELL_X32 FILLER_235_3071 ();
 FILLCELL_X32 FILLER_235_3103 ();
 FILLCELL_X32 FILLER_235_3135 ();
 FILLCELL_X32 FILLER_235_3167 ();
 FILLCELL_X32 FILLER_235_3199 ();
 FILLCELL_X32 FILLER_235_3231 ();
 FILLCELL_X32 FILLER_235_3263 ();
 FILLCELL_X32 FILLER_235_3295 ();
 FILLCELL_X32 FILLER_235_3327 ();
 FILLCELL_X32 FILLER_235_3359 ();
 FILLCELL_X32 FILLER_235_3391 ();
 FILLCELL_X32 FILLER_235_3423 ();
 FILLCELL_X32 FILLER_235_3455 ();
 FILLCELL_X32 FILLER_235_3487 ();
 FILLCELL_X32 FILLER_235_3519 ();
 FILLCELL_X32 FILLER_235_3551 ();
 FILLCELL_X32 FILLER_235_3583 ();
 FILLCELL_X32 FILLER_235_3615 ();
 FILLCELL_X32 FILLER_235_3647 ();
 FILLCELL_X32 FILLER_235_3679 ();
 FILLCELL_X16 FILLER_235_3711 ();
 FILLCELL_X8 FILLER_235_3727 ();
 FILLCELL_X2 FILLER_235_3735 ();
 FILLCELL_X1 FILLER_235_3737 ();
 FILLCELL_X32 FILLER_236_1 ();
 FILLCELL_X32 FILLER_236_33 ();
 FILLCELL_X32 FILLER_236_65 ();
 FILLCELL_X32 FILLER_236_97 ();
 FILLCELL_X32 FILLER_236_129 ();
 FILLCELL_X32 FILLER_236_161 ();
 FILLCELL_X32 FILLER_236_193 ();
 FILLCELL_X32 FILLER_236_225 ();
 FILLCELL_X32 FILLER_236_257 ();
 FILLCELL_X32 FILLER_236_289 ();
 FILLCELL_X32 FILLER_236_321 ();
 FILLCELL_X32 FILLER_236_353 ();
 FILLCELL_X32 FILLER_236_385 ();
 FILLCELL_X32 FILLER_236_417 ();
 FILLCELL_X32 FILLER_236_449 ();
 FILLCELL_X32 FILLER_236_481 ();
 FILLCELL_X32 FILLER_236_513 ();
 FILLCELL_X32 FILLER_236_545 ();
 FILLCELL_X32 FILLER_236_577 ();
 FILLCELL_X16 FILLER_236_609 ();
 FILLCELL_X4 FILLER_236_625 ();
 FILLCELL_X2 FILLER_236_629 ();
 FILLCELL_X32 FILLER_236_632 ();
 FILLCELL_X32 FILLER_236_664 ();
 FILLCELL_X32 FILLER_236_696 ();
 FILLCELL_X32 FILLER_236_728 ();
 FILLCELL_X32 FILLER_236_760 ();
 FILLCELL_X32 FILLER_236_792 ();
 FILLCELL_X32 FILLER_236_824 ();
 FILLCELL_X32 FILLER_236_856 ();
 FILLCELL_X32 FILLER_236_888 ();
 FILLCELL_X32 FILLER_236_920 ();
 FILLCELL_X32 FILLER_236_952 ();
 FILLCELL_X32 FILLER_236_984 ();
 FILLCELL_X32 FILLER_236_1016 ();
 FILLCELL_X32 FILLER_236_1048 ();
 FILLCELL_X32 FILLER_236_1080 ();
 FILLCELL_X32 FILLER_236_1112 ();
 FILLCELL_X32 FILLER_236_1144 ();
 FILLCELL_X32 FILLER_236_1176 ();
 FILLCELL_X32 FILLER_236_1208 ();
 FILLCELL_X32 FILLER_236_1240 ();
 FILLCELL_X32 FILLER_236_1272 ();
 FILLCELL_X32 FILLER_236_1304 ();
 FILLCELL_X32 FILLER_236_1336 ();
 FILLCELL_X32 FILLER_236_1368 ();
 FILLCELL_X32 FILLER_236_1400 ();
 FILLCELL_X32 FILLER_236_1432 ();
 FILLCELL_X32 FILLER_236_1464 ();
 FILLCELL_X32 FILLER_236_1496 ();
 FILLCELL_X32 FILLER_236_1528 ();
 FILLCELL_X32 FILLER_236_1560 ();
 FILLCELL_X32 FILLER_236_1592 ();
 FILLCELL_X32 FILLER_236_1624 ();
 FILLCELL_X32 FILLER_236_1656 ();
 FILLCELL_X32 FILLER_236_1688 ();
 FILLCELL_X32 FILLER_236_1720 ();
 FILLCELL_X32 FILLER_236_1752 ();
 FILLCELL_X32 FILLER_236_1784 ();
 FILLCELL_X32 FILLER_236_1816 ();
 FILLCELL_X16 FILLER_236_1848 ();
 FILLCELL_X1 FILLER_236_1864 ();
 FILLCELL_X16 FILLER_236_1875 ();
 FILLCELL_X2 FILLER_236_1891 ();
 FILLCELL_X1 FILLER_236_1893 ();
 FILLCELL_X32 FILLER_236_1895 ();
 FILLCELL_X4 FILLER_236_1927 ();
 FILLCELL_X32 FILLER_236_1944 ();
 FILLCELL_X8 FILLER_236_1976 ();
 FILLCELL_X4 FILLER_236_1984 ();
 FILLCELL_X32 FILLER_236_2001 ();
 FILLCELL_X8 FILLER_236_2033 ();
 FILLCELL_X1 FILLER_236_2041 ();
 FILLCELL_X1 FILLER_236_2076 ();
 FILLCELL_X4 FILLER_236_2084 ();
 FILLCELL_X1 FILLER_236_2088 ();
 FILLCELL_X32 FILLER_236_2113 ();
 FILLCELL_X1 FILLER_236_2145 ();
 FILLCELL_X8 FILLER_236_2161 ();
 FILLCELL_X1 FILLER_236_2169 ();
 FILLCELL_X16 FILLER_236_2177 ();
 FILLCELL_X4 FILLER_236_2193 ();
 FILLCELL_X2 FILLER_236_2197 ();
 FILLCELL_X8 FILLER_236_2206 ();
 FILLCELL_X1 FILLER_236_2214 ();
 FILLCELL_X32 FILLER_236_2232 ();
 FILLCELL_X32 FILLER_236_2264 ();
 FILLCELL_X32 FILLER_236_2296 ();
 FILLCELL_X32 FILLER_236_2328 ();
 FILLCELL_X32 FILLER_236_2360 ();
 FILLCELL_X32 FILLER_236_2392 ();
 FILLCELL_X32 FILLER_236_2424 ();
 FILLCELL_X32 FILLER_236_2456 ();
 FILLCELL_X32 FILLER_236_2488 ();
 FILLCELL_X32 FILLER_236_2520 ();
 FILLCELL_X32 FILLER_236_2552 ();
 FILLCELL_X32 FILLER_236_2584 ();
 FILLCELL_X32 FILLER_236_2616 ();
 FILLCELL_X32 FILLER_236_2648 ();
 FILLCELL_X32 FILLER_236_2680 ();
 FILLCELL_X32 FILLER_236_2712 ();
 FILLCELL_X32 FILLER_236_2744 ();
 FILLCELL_X32 FILLER_236_2776 ();
 FILLCELL_X32 FILLER_236_2808 ();
 FILLCELL_X32 FILLER_236_2840 ();
 FILLCELL_X32 FILLER_236_2872 ();
 FILLCELL_X32 FILLER_236_2904 ();
 FILLCELL_X32 FILLER_236_2936 ();
 FILLCELL_X32 FILLER_236_2968 ();
 FILLCELL_X32 FILLER_236_3000 ();
 FILLCELL_X32 FILLER_236_3032 ();
 FILLCELL_X32 FILLER_236_3064 ();
 FILLCELL_X32 FILLER_236_3096 ();
 FILLCELL_X16 FILLER_236_3128 ();
 FILLCELL_X8 FILLER_236_3144 ();
 FILLCELL_X4 FILLER_236_3152 ();
 FILLCELL_X1 FILLER_236_3156 ();
 FILLCELL_X32 FILLER_236_3158 ();
 FILLCELL_X32 FILLER_236_3190 ();
 FILLCELL_X32 FILLER_236_3222 ();
 FILLCELL_X32 FILLER_236_3254 ();
 FILLCELL_X32 FILLER_236_3286 ();
 FILLCELL_X32 FILLER_236_3318 ();
 FILLCELL_X32 FILLER_236_3350 ();
 FILLCELL_X32 FILLER_236_3382 ();
 FILLCELL_X32 FILLER_236_3414 ();
 FILLCELL_X32 FILLER_236_3446 ();
 FILLCELL_X32 FILLER_236_3478 ();
 FILLCELL_X32 FILLER_236_3510 ();
 FILLCELL_X32 FILLER_236_3542 ();
 FILLCELL_X32 FILLER_236_3574 ();
 FILLCELL_X32 FILLER_236_3606 ();
 FILLCELL_X32 FILLER_236_3638 ();
 FILLCELL_X32 FILLER_236_3670 ();
 FILLCELL_X32 FILLER_236_3702 ();
 FILLCELL_X4 FILLER_236_3734 ();
 FILLCELL_X32 FILLER_237_1 ();
 FILLCELL_X32 FILLER_237_33 ();
 FILLCELL_X32 FILLER_237_65 ();
 FILLCELL_X32 FILLER_237_97 ();
 FILLCELL_X32 FILLER_237_129 ();
 FILLCELL_X32 FILLER_237_161 ();
 FILLCELL_X32 FILLER_237_193 ();
 FILLCELL_X32 FILLER_237_225 ();
 FILLCELL_X32 FILLER_237_257 ();
 FILLCELL_X32 FILLER_237_289 ();
 FILLCELL_X32 FILLER_237_321 ();
 FILLCELL_X32 FILLER_237_353 ();
 FILLCELL_X32 FILLER_237_385 ();
 FILLCELL_X32 FILLER_237_417 ();
 FILLCELL_X32 FILLER_237_449 ();
 FILLCELL_X32 FILLER_237_481 ();
 FILLCELL_X32 FILLER_237_513 ();
 FILLCELL_X32 FILLER_237_545 ();
 FILLCELL_X32 FILLER_237_577 ();
 FILLCELL_X32 FILLER_237_609 ();
 FILLCELL_X32 FILLER_237_641 ();
 FILLCELL_X32 FILLER_237_673 ();
 FILLCELL_X32 FILLER_237_705 ();
 FILLCELL_X32 FILLER_237_737 ();
 FILLCELL_X32 FILLER_237_769 ();
 FILLCELL_X32 FILLER_237_801 ();
 FILLCELL_X32 FILLER_237_833 ();
 FILLCELL_X32 FILLER_237_865 ();
 FILLCELL_X32 FILLER_237_897 ();
 FILLCELL_X32 FILLER_237_929 ();
 FILLCELL_X32 FILLER_237_961 ();
 FILLCELL_X32 FILLER_237_993 ();
 FILLCELL_X32 FILLER_237_1025 ();
 FILLCELL_X32 FILLER_237_1057 ();
 FILLCELL_X32 FILLER_237_1089 ();
 FILLCELL_X32 FILLER_237_1121 ();
 FILLCELL_X32 FILLER_237_1153 ();
 FILLCELL_X32 FILLER_237_1185 ();
 FILLCELL_X32 FILLER_237_1217 ();
 FILLCELL_X8 FILLER_237_1249 ();
 FILLCELL_X4 FILLER_237_1257 ();
 FILLCELL_X2 FILLER_237_1261 ();
 FILLCELL_X32 FILLER_237_1264 ();
 FILLCELL_X32 FILLER_237_1296 ();
 FILLCELL_X32 FILLER_237_1328 ();
 FILLCELL_X32 FILLER_237_1360 ();
 FILLCELL_X32 FILLER_237_1392 ();
 FILLCELL_X32 FILLER_237_1424 ();
 FILLCELL_X32 FILLER_237_1456 ();
 FILLCELL_X32 FILLER_237_1488 ();
 FILLCELL_X32 FILLER_237_1520 ();
 FILLCELL_X32 FILLER_237_1552 ();
 FILLCELL_X32 FILLER_237_1584 ();
 FILLCELL_X32 FILLER_237_1616 ();
 FILLCELL_X32 FILLER_237_1648 ();
 FILLCELL_X32 FILLER_237_1680 ();
 FILLCELL_X32 FILLER_237_1712 ();
 FILLCELL_X32 FILLER_237_1744 ();
 FILLCELL_X32 FILLER_237_1776 ();
 FILLCELL_X32 FILLER_237_1808 ();
 FILLCELL_X4 FILLER_237_1840 ();
 FILLCELL_X2 FILLER_237_1844 ();
 FILLCELL_X1 FILLER_237_1846 ();
 FILLCELL_X2 FILLER_237_1864 ();
 FILLCELL_X8 FILLER_237_1873 ();
 FILLCELL_X4 FILLER_237_1881 ();
 FILLCELL_X1 FILLER_237_1885 ();
 FILLCELL_X32 FILLER_237_1896 ();
 FILLCELL_X2 FILLER_237_1928 ();
 FILLCELL_X16 FILLER_237_1937 ();
 FILLCELL_X8 FILLER_237_1953 ();
 FILLCELL_X1 FILLER_237_1961 ();
 FILLCELL_X4 FILLER_237_1979 ();
 FILLCELL_X1 FILLER_237_1983 ();
 FILLCELL_X2 FILLER_237_1991 ();
 FILLCELL_X16 FILLER_237_2006 ();
 FILLCELL_X8 FILLER_237_2022 ();
 FILLCELL_X4 FILLER_237_2030 ();
 FILLCELL_X2 FILLER_237_2034 ();
 FILLCELL_X32 FILLER_237_2043 ();
 FILLCELL_X16 FILLER_237_2075 ();
 FILLCELL_X8 FILLER_237_2091 ();
 FILLCELL_X1 FILLER_237_2099 ();
 FILLCELL_X16 FILLER_237_2124 ();
 FILLCELL_X4 FILLER_237_2157 ();
 FILLCELL_X1 FILLER_237_2161 ();
 FILLCELL_X8 FILLER_237_2186 ();
 FILLCELL_X1 FILLER_237_2194 ();
 FILLCELL_X8 FILLER_237_2202 ();
 FILLCELL_X4 FILLER_237_2210 ();
 FILLCELL_X2 FILLER_237_2214 ();
 FILLCELL_X32 FILLER_237_2235 ();
 FILLCELL_X32 FILLER_237_2267 ();
 FILLCELL_X32 FILLER_237_2299 ();
 FILLCELL_X32 FILLER_237_2331 ();
 FILLCELL_X32 FILLER_237_2363 ();
 FILLCELL_X32 FILLER_237_2395 ();
 FILLCELL_X32 FILLER_237_2427 ();
 FILLCELL_X32 FILLER_237_2459 ();
 FILLCELL_X32 FILLER_237_2491 ();
 FILLCELL_X2 FILLER_237_2523 ();
 FILLCELL_X1 FILLER_237_2525 ();
 FILLCELL_X32 FILLER_237_2527 ();
 FILLCELL_X32 FILLER_237_2559 ();
 FILLCELL_X32 FILLER_237_2591 ();
 FILLCELL_X32 FILLER_237_2623 ();
 FILLCELL_X32 FILLER_237_2655 ();
 FILLCELL_X32 FILLER_237_2687 ();
 FILLCELL_X32 FILLER_237_2719 ();
 FILLCELL_X32 FILLER_237_2751 ();
 FILLCELL_X32 FILLER_237_2783 ();
 FILLCELL_X32 FILLER_237_2815 ();
 FILLCELL_X32 FILLER_237_2847 ();
 FILLCELL_X32 FILLER_237_2879 ();
 FILLCELL_X32 FILLER_237_2911 ();
 FILLCELL_X32 FILLER_237_2943 ();
 FILLCELL_X32 FILLER_237_2975 ();
 FILLCELL_X32 FILLER_237_3007 ();
 FILLCELL_X32 FILLER_237_3039 ();
 FILLCELL_X32 FILLER_237_3071 ();
 FILLCELL_X32 FILLER_237_3103 ();
 FILLCELL_X32 FILLER_237_3135 ();
 FILLCELL_X32 FILLER_237_3167 ();
 FILLCELL_X32 FILLER_237_3199 ();
 FILLCELL_X32 FILLER_237_3231 ();
 FILLCELL_X32 FILLER_237_3263 ();
 FILLCELL_X32 FILLER_237_3295 ();
 FILLCELL_X32 FILLER_237_3327 ();
 FILLCELL_X32 FILLER_237_3359 ();
 FILLCELL_X32 FILLER_237_3391 ();
 FILLCELL_X32 FILLER_237_3423 ();
 FILLCELL_X32 FILLER_237_3455 ();
 FILLCELL_X32 FILLER_237_3487 ();
 FILLCELL_X32 FILLER_237_3519 ();
 FILLCELL_X32 FILLER_237_3551 ();
 FILLCELL_X32 FILLER_237_3583 ();
 FILLCELL_X32 FILLER_237_3615 ();
 FILLCELL_X32 FILLER_237_3647 ();
 FILLCELL_X32 FILLER_237_3679 ();
 FILLCELL_X16 FILLER_237_3711 ();
 FILLCELL_X8 FILLER_237_3727 ();
 FILLCELL_X2 FILLER_237_3735 ();
 FILLCELL_X1 FILLER_237_3737 ();
 FILLCELL_X32 FILLER_238_1 ();
 FILLCELL_X32 FILLER_238_33 ();
 FILLCELL_X32 FILLER_238_65 ();
 FILLCELL_X32 FILLER_238_97 ();
 FILLCELL_X32 FILLER_238_129 ();
 FILLCELL_X32 FILLER_238_161 ();
 FILLCELL_X32 FILLER_238_193 ();
 FILLCELL_X32 FILLER_238_225 ();
 FILLCELL_X32 FILLER_238_257 ();
 FILLCELL_X32 FILLER_238_289 ();
 FILLCELL_X32 FILLER_238_321 ();
 FILLCELL_X32 FILLER_238_353 ();
 FILLCELL_X32 FILLER_238_385 ();
 FILLCELL_X32 FILLER_238_417 ();
 FILLCELL_X32 FILLER_238_449 ();
 FILLCELL_X32 FILLER_238_481 ();
 FILLCELL_X32 FILLER_238_513 ();
 FILLCELL_X32 FILLER_238_545 ();
 FILLCELL_X32 FILLER_238_577 ();
 FILLCELL_X16 FILLER_238_609 ();
 FILLCELL_X4 FILLER_238_625 ();
 FILLCELL_X2 FILLER_238_629 ();
 FILLCELL_X32 FILLER_238_632 ();
 FILLCELL_X32 FILLER_238_664 ();
 FILLCELL_X32 FILLER_238_696 ();
 FILLCELL_X32 FILLER_238_728 ();
 FILLCELL_X32 FILLER_238_760 ();
 FILLCELL_X32 FILLER_238_792 ();
 FILLCELL_X32 FILLER_238_824 ();
 FILLCELL_X32 FILLER_238_856 ();
 FILLCELL_X32 FILLER_238_888 ();
 FILLCELL_X32 FILLER_238_920 ();
 FILLCELL_X32 FILLER_238_952 ();
 FILLCELL_X32 FILLER_238_984 ();
 FILLCELL_X32 FILLER_238_1016 ();
 FILLCELL_X32 FILLER_238_1048 ();
 FILLCELL_X32 FILLER_238_1080 ();
 FILLCELL_X32 FILLER_238_1112 ();
 FILLCELL_X32 FILLER_238_1144 ();
 FILLCELL_X32 FILLER_238_1176 ();
 FILLCELL_X32 FILLER_238_1208 ();
 FILLCELL_X32 FILLER_238_1240 ();
 FILLCELL_X32 FILLER_238_1272 ();
 FILLCELL_X32 FILLER_238_1304 ();
 FILLCELL_X32 FILLER_238_1336 ();
 FILLCELL_X32 FILLER_238_1368 ();
 FILLCELL_X32 FILLER_238_1400 ();
 FILLCELL_X32 FILLER_238_1432 ();
 FILLCELL_X32 FILLER_238_1464 ();
 FILLCELL_X32 FILLER_238_1496 ();
 FILLCELL_X32 FILLER_238_1528 ();
 FILLCELL_X32 FILLER_238_1560 ();
 FILLCELL_X32 FILLER_238_1592 ();
 FILLCELL_X32 FILLER_238_1624 ();
 FILLCELL_X32 FILLER_238_1656 ();
 FILLCELL_X32 FILLER_238_1688 ();
 FILLCELL_X32 FILLER_238_1720 ();
 FILLCELL_X32 FILLER_238_1752 ();
 FILLCELL_X32 FILLER_238_1784 ();
 FILLCELL_X16 FILLER_238_1816 ();
 FILLCELL_X8 FILLER_238_1832 ();
 FILLCELL_X2 FILLER_238_1840 ();
 FILLCELL_X16 FILLER_238_1852 ();
 FILLCELL_X4 FILLER_238_1868 ();
 FILLCELL_X2 FILLER_238_1872 ();
 FILLCELL_X1 FILLER_238_1874 ();
 FILLCELL_X8 FILLER_238_1895 ();
 FILLCELL_X1 FILLER_238_1903 ();
 FILLCELL_X8 FILLER_238_1933 ();
 FILLCELL_X4 FILLER_238_1941 ();
 FILLCELL_X16 FILLER_238_1950 ();
 FILLCELL_X8 FILLER_238_1966 ();
 FILLCELL_X4 FILLER_238_1974 ();
 FILLCELL_X1 FILLER_238_1978 ();
 FILLCELL_X2 FILLER_238_2003 ();
 FILLCELL_X1 FILLER_238_2005 ();
 FILLCELL_X8 FILLER_238_2019 ();
 FILLCELL_X2 FILLER_238_2027 ();
 FILLCELL_X1 FILLER_238_2029 ();
 FILLCELL_X1 FILLER_238_2047 ();
 FILLCELL_X4 FILLER_238_2055 ();
 FILLCELL_X32 FILLER_238_2067 ();
 FILLCELL_X8 FILLER_238_2099 ();
 FILLCELL_X32 FILLER_238_2114 ();
 FILLCELL_X32 FILLER_238_2146 ();
 FILLCELL_X16 FILLER_238_2178 ();
 FILLCELL_X1 FILLER_238_2194 ();
 FILLCELL_X8 FILLER_238_2212 ();
 FILLCELL_X4 FILLER_238_2220 ();
 FILLCELL_X8 FILLER_238_2227 ();
 FILLCELL_X4 FILLER_238_2235 ();
 FILLCELL_X2 FILLER_238_2239 ();
 FILLCELL_X1 FILLER_238_2241 ();
 FILLCELL_X32 FILLER_238_2259 ();
 FILLCELL_X32 FILLER_238_2291 ();
 FILLCELL_X32 FILLER_238_2323 ();
 FILLCELL_X32 FILLER_238_2355 ();
 FILLCELL_X32 FILLER_238_2387 ();
 FILLCELL_X32 FILLER_238_2419 ();
 FILLCELL_X32 FILLER_238_2451 ();
 FILLCELL_X32 FILLER_238_2483 ();
 FILLCELL_X32 FILLER_238_2515 ();
 FILLCELL_X32 FILLER_238_2547 ();
 FILLCELL_X32 FILLER_238_2579 ();
 FILLCELL_X32 FILLER_238_2611 ();
 FILLCELL_X32 FILLER_238_2643 ();
 FILLCELL_X32 FILLER_238_2675 ();
 FILLCELL_X32 FILLER_238_2707 ();
 FILLCELL_X32 FILLER_238_2739 ();
 FILLCELL_X32 FILLER_238_2771 ();
 FILLCELL_X32 FILLER_238_2803 ();
 FILLCELL_X32 FILLER_238_2835 ();
 FILLCELL_X32 FILLER_238_2867 ();
 FILLCELL_X32 FILLER_238_2899 ();
 FILLCELL_X32 FILLER_238_2931 ();
 FILLCELL_X32 FILLER_238_2963 ();
 FILLCELL_X32 FILLER_238_2995 ();
 FILLCELL_X32 FILLER_238_3027 ();
 FILLCELL_X32 FILLER_238_3059 ();
 FILLCELL_X32 FILLER_238_3091 ();
 FILLCELL_X32 FILLER_238_3123 ();
 FILLCELL_X2 FILLER_238_3155 ();
 FILLCELL_X32 FILLER_238_3158 ();
 FILLCELL_X32 FILLER_238_3190 ();
 FILLCELL_X32 FILLER_238_3222 ();
 FILLCELL_X32 FILLER_238_3254 ();
 FILLCELL_X32 FILLER_238_3286 ();
 FILLCELL_X32 FILLER_238_3318 ();
 FILLCELL_X32 FILLER_238_3350 ();
 FILLCELL_X32 FILLER_238_3382 ();
 FILLCELL_X32 FILLER_238_3414 ();
 FILLCELL_X32 FILLER_238_3446 ();
 FILLCELL_X32 FILLER_238_3478 ();
 FILLCELL_X32 FILLER_238_3510 ();
 FILLCELL_X32 FILLER_238_3542 ();
 FILLCELL_X32 FILLER_238_3574 ();
 FILLCELL_X32 FILLER_238_3606 ();
 FILLCELL_X32 FILLER_238_3638 ();
 FILLCELL_X32 FILLER_238_3670 ();
 FILLCELL_X32 FILLER_238_3702 ();
 FILLCELL_X4 FILLER_238_3734 ();
 FILLCELL_X32 FILLER_239_1 ();
 FILLCELL_X32 FILLER_239_33 ();
 FILLCELL_X32 FILLER_239_65 ();
 FILLCELL_X32 FILLER_239_97 ();
 FILLCELL_X32 FILLER_239_129 ();
 FILLCELL_X32 FILLER_239_161 ();
 FILLCELL_X32 FILLER_239_193 ();
 FILLCELL_X32 FILLER_239_225 ();
 FILLCELL_X32 FILLER_239_257 ();
 FILLCELL_X32 FILLER_239_289 ();
 FILLCELL_X32 FILLER_239_321 ();
 FILLCELL_X32 FILLER_239_353 ();
 FILLCELL_X32 FILLER_239_385 ();
 FILLCELL_X32 FILLER_239_417 ();
 FILLCELL_X32 FILLER_239_449 ();
 FILLCELL_X32 FILLER_239_481 ();
 FILLCELL_X32 FILLER_239_513 ();
 FILLCELL_X32 FILLER_239_545 ();
 FILLCELL_X32 FILLER_239_577 ();
 FILLCELL_X32 FILLER_239_609 ();
 FILLCELL_X32 FILLER_239_641 ();
 FILLCELL_X32 FILLER_239_673 ();
 FILLCELL_X32 FILLER_239_705 ();
 FILLCELL_X32 FILLER_239_737 ();
 FILLCELL_X32 FILLER_239_769 ();
 FILLCELL_X32 FILLER_239_801 ();
 FILLCELL_X32 FILLER_239_833 ();
 FILLCELL_X32 FILLER_239_865 ();
 FILLCELL_X32 FILLER_239_897 ();
 FILLCELL_X32 FILLER_239_929 ();
 FILLCELL_X32 FILLER_239_961 ();
 FILLCELL_X32 FILLER_239_993 ();
 FILLCELL_X32 FILLER_239_1025 ();
 FILLCELL_X32 FILLER_239_1057 ();
 FILLCELL_X32 FILLER_239_1089 ();
 FILLCELL_X32 FILLER_239_1121 ();
 FILLCELL_X32 FILLER_239_1153 ();
 FILLCELL_X32 FILLER_239_1185 ();
 FILLCELL_X32 FILLER_239_1217 ();
 FILLCELL_X8 FILLER_239_1249 ();
 FILLCELL_X4 FILLER_239_1257 ();
 FILLCELL_X2 FILLER_239_1261 ();
 FILLCELL_X32 FILLER_239_1264 ();
 FILLCELL_X32 FILLER_239_1296 ();
 FILLCELL_X32 FILLER_239_1328 ();
 FILLCELL_X32 FILLER_239_1360 ();
 FILLCELL_X32 FILLER_239_1392 ();
 FILLCELL_X32 FILLER_239_1424 ();
 FILLCELL_X32 FILLER_239_1456 ();
 FILLCELL_X32 FILLER_239_1488 ();
 FILLCELL_X32 FILLER_239_1520 ();
 FILLCELL_X32 FILLER_239_1552 ();
 FILLCELL_X32 FILLER_239_1584 ();
 FILLCELL_X32 FILLER_239_1616 ();
 FILLCELL_X32 FILLER_239_1648 ();
 FILLCELL_X32 FILLER_239_1680 ();
 FILLCELL_X32 FILLER_239_1712 ();
 FILLCELL_X32 FILLER_239_1744 ();
 FILLCELL_X32 FILLER_239_1776 ();
 FILLCELL_X32 FILLER_239_1808 ();
 FILLCELL_X2 FILLER_239_1840 ();
 FILLCELL_X1 FILLER_239_1842 ();
 FILLCELL_X32 FILLER_239_1847 ();
 FILLCELL_X1 FILLER_239_1879 ();
 FILLCELL_X8 FILLER_239_1884 ();
 FILLCELL_X4 FILLER_239_1892 ();
 FILLCELL_X2 FILLER_239_1896 ();
 FILLCELL_X4 FILLER_239_1902 ();
 FILLCELL_X2 FILLER_239_1906 ();
 FILLCELL_X2 FILLER_239_1918 ();
 FILLCELL_X4 FILLER_239_1930 ();
 FILLCELL_X4 FILLER_239_1939 ();
 FILLCELL_X2 FILLER_239_1943 ();
 FILLCELL_X1 FILLER_239_1945 ();
 FILLCELL_X8 FILLER_239_1968 ();
 FILLCELL_X8 FILLER_239_1990 ();
 FILLCELL_X4 FILLER_239_1998 ();
 FILLCELL_X32 FILLER_239_2015 ();
 FILLCELL_X16 FILLER_239_2047 ();
 FILLCELL_X4 FILLER_239_2063 ();
 FILLCELL_X2 FILLER_239_2067 ();
 FILLCELL_X32 FILLER_239_2076 ();
 FILLCELL_X32 FILLER_239_2108 ();
 FILLCELL_X32 FILLER_239_2140 ();
 FILLCELL_X32 FILLER_239_2172 ();
 FILLCELL_X32 FILLER_239_2204 ();
 FILLCELL_X8 FILLER_239_2236 ();
 FILLCELL_X4 FILLER_239_2244 ();
 FILLCELL_X1 FILLER_239_2248 ();
 FILLCELL_X2 FILLER_239_2263 ();
 FILLCELL_X1 FILLER_239_2265 ();
 FILLCELL_X4 FILLER_239_2273 ();
 FILLCELL_X2 FILLER_239_2277 ();
 FILLCELL_X1 FILLER_239_2279 ();
 FILLCELL_X32 FILLER_239_2297 ();
 FILLCELL_X32 FILLER_239_2329 ();
 FILLCELL_X32 FILLER_239_2361 ();
 FILLCELL_X32 FILLER_239_2393 ();
 FILLCELL_X32 FILLER_239_2425 ();
 FILLCELL_X32 FILLER_239_2457 ();
 FILLCELL_X32 FILLER_239_2489 ();
 FILLCELL_X4 FILLER_239_2521 ();
 FILLCELL_X1 FILLER_239_2525 ();
 FILLCELL_X32 FILLER_239_2527 ();
 FILLCELL_X32 FILLER_239_2559 ();
 FILLCELL_X32 FILLER_239_2591 ();
 FILLCELL_X32 FILLER_239_2623 ();
 FILLCELL_X32 FILLER_239_2655 ();
 FILLCELL_X32 FILLER_239_2687 ();
 FILLCELL_X32 FILLER_239_2719 ();
 FILLCELL_X32 FILLER_239_2751 ();
 FILLCELL_X32 FILLER_239_2783 ();
 FILLCELL_X32 FILLER_239_2815 ();
 FILLCELL_X32 FILLER_239_2847 ();
 FILLCELL_X32 FILLER_239_2879 ();
 FILLCELL_X32 FILLER_239_2911 ();
 FILLCELL_X32 FILLER_239_2943 ();
 FILLCELL_X32 FILLER_239_2975 ();
 FILLCELL_X32 FILLER_239_3007 ();
 FILLCELL_X32 FILLER_239_3039 ();
 FILLCELL_X32 FILLER_239_3071 ();
 FILLCELL_X32 FILLER_239_3103 ();
 FILLCELL_X32 FILLER_239_3135 ();
 FILLCELL_X32 FILLER_239_3167 ();
 FILLCELL_X32 FILLER_239_3199 ();
 FILLCELL_X32 FILLER_239_3231 ();
 FILLCELL_X32 FILLER_239_3263 ();
 FILLCELL_X32 FILLER_239_3295 ();
 FILLCELL_X32 FILLER_239_3327 ();
 FILLCELL_X32 FILLER_239_3359 ();
 FILLCELL_X32 FILLER_239_3391 ();
 FILLCELL_X32 FILLER_239_3423 ();
 FILLCELL_X32 FILLER_239_3455 ();
 FILLCELL_X32 FILLER_239_3487 ();
 FILLCELL_X32 FILLER_239_3519 ();
 FILLCELL_X32 FILLER_239_3551 ();
 FILLCELL_X32 FILLER_239_3583 ();
 FILLCELL_X32 FILLER_239_3615 ();
 FILLCELL_X32 FILLER_239_3647 ();
 FILLCELL_X32 FILLER_239_3679 ();
 FILLCELL_X16 FILLER_239_3711 ();
 FILLCELL_X8 FILLER_239_3727 ();
 FILLCELL_X2 FILLER_239_3735 ();
 FILLCELL_X1 FILLER_239_3737 ();
 FILLCELL_X32 FILLER_240_1 ();
 FILLCELL_X32 FILLER_240_33 ();
 FILLCELL_X32 FILLER_240_65 ();
 FILLCELL_X32 FILLER_240_97 ();
 FILLCELL_X32 FILLER_240_129 ();
 FILLCELL_X32 FILLER_240_161 ();
 FILLCELL_X32 FILLER_240_193 ();
 FILLCELL_X32 FILLER_240_225 ();
 FILLCELL_X32 FILLER_240_257 ();
 FILLCELL_X32 FILLER_240_289 ();
 FILLCELL_X32 FILLER_240_321 ();
 FILLCELL_X32 FILLER_240_353 ();
 FILLCELL_X32 FILLER_240_385 ();
 FILLCELL_X32 FILLER_240_417 ();
 FILLCELL_X32 FILLER_240_449 ();
 FILLCELL_X32 FILLER_240_481 ();
 FILLCELL_X32 FILLER_240_513 ();
 FILLCELL_X32 FILLER_240_545 ();
 FILLCELL_X32 FILLER_240_577 ();
 FILLCELL_X16 FILLER_240_609 ();
 FILLCELL_X4 FILLER_240_625 ();
 FILLCELL_X2 FILLER_240_629 ();
 FILLCELL_X32 FILLER_240_632 ();
 FILLCELL_X32 FILLER_240_664 ();
 FILLCELL_X32 FILLER_240_696 ();
 FILLCELL_X32 FILLER_240_728 ();
 FILLCELL_X32 FILLER_240_760 ();
 FILLCELL_X32 FILLER_240_792 ();
 FILLCELL_X32 FILLER_240_824 ();
 FILLCELL_X32 FILLER_240_856 ();
 FILLCELL_X32 FILLER_240_888 ();
 FILLCELL_X32 FILLER_240_920 ();
 FILLCELL_X32 FILLER_240_952 ();
 FILLCELL_X32 FILLER_240_984 ();
 FILLCELL_X32 FILLER_240_1016 ();
 FILLCELL_X32 FILLER_240_1048 ();
 FILLCELL_X32 FILLER_240_1080 ();
 FILLCELL_X32 FILLER_240_1112 ();
 FILLCELL_X32 FILLER_240_1144 ();
 FILLCELL_X32 FILLER_240_1176 ();
 FILLCELL_X32 FILLER_240_1208 ();
 FILLCELL_X32 FILLER_240_1240 ();
 FILLCELL_X32 FILLER_240_1272 ();
 FILLCELL_X32 FILLER_240_1304 ();
 FILLCELL_X32 FILLER_240_1336 ();
 FILLCELL_X32 FILLER_240_1368 ();
 FILLCELL_X32 FILLER_240_1400 ();
 FILLCELL_X32 FILLER_240_1432 ();
 FILLCELL_X32 FILLER_240_1464 ();
 FILLCELL_X32 FILLER_240_1496 ();
 FILLCELL_X32 FILLER_240_1528 ();
 FILLCELL_X32 FILLER_240_1560 ();
 FILLCELL_X32 FILLER_240_1592 ();
 FILLCELL_X32 FILLER_240_1624 ();
 FILLCELL_X32 FILLER_240_1656 ();
 FILLCELL_X32 FILLER_240_1688 ();
 FILLCELL_X32 FILLER_240_1720 ();
 FILLCELL_X32 FILLER_240_1752 ();
 FILLCELL_X32 FILLER_240_1784 ();
 FILLCELL_X32 FILLER_240_1816 ();
 FILLCELL_X16 FILLER_240_1848 ();
 FILLCELL_X4 FILLER_240_1864 ();
 FILLCELL_X1 FILLER_240_1868 ();
 FILLCELL_X2 FILLER_240_1874 ();
 FILLCELL_X1 FILLER_240_1876 ();
 FILLCELL_X2 FILLER_240_1888 ();
 FILLCELL_X8 FILLER_240_1902 ();
 FILLCELL_X4 FILLER_240_1910 ();
 FILLCELL_X2 FILLER_240_1914 ();
 FILLCELL_X1 FILLER_240_1916 ();
 FILLCELL_X8 FILLER_240_1924 ();
 FILLCELL_X4 FILLER_240_1932 ();
 FILLCELL_X2 FILLER_240_1936 ();
 FILLCELL_X1 FILLER_240_1938 ();
 FILLCELL_X4 FILLER_240_1942 ();
 FILLCELL_X8 FILLER_240_1988 ();
 FILLCELL_X8 FILLER_240_2009 ();
 FILLCELL_X4 FILLER_240_2017 ();
 FILLCELL_X16 FILLER_240_2028 ();
 FILLCELL_X8 FILLER_240_2044 ();
 FILLCELL_X4 FILLER_240_2052 ();
 FILLCELL_X2 FILLER_240_2056 ();
 FILLCELL_X1 FILLER_240_2075 ();
 FILLCELL_X32 FILLER_240_2107 ();
 FILLCELL_X8 FILLER_240_2139 ();
 FILLCELL_X4 FILLER_240_2147 ();
 FILLCELL_X2 FILLER_240_2151 ();
 FILLCELL_X1 FILLER_240_2153 ();
 FILLCELL_X8 FILLER_240_2161 ();
 FILLCELL_X4 FILLER_240_2169 ();
 FILLCELL_X8 FILLER_240_2204 ();
 FILLCELL_X4 FILLER_240_2212 ();
 FILLCELL_X2 FILLER_240_2216 ();
 FILLCELL_X1 FILLER_240_2218 ();
 FILLCELL_X2 FILLER_240_2236 ();
 FILLCELL_X1 FILLER_240_2238 ();
 FILLCELL_X32 FILLER_240_2246 ();
 FILLCELL_X32 FILLER_240_2278 ();
 FILLCELL_X32 FILLER_240_2310 ();
 FILLCELL_X32 FILLER_240_2342 ();
 FILLCELL_X32 FILLER_240_2374 ();
 FILLCELL_X32 FILLER_240_2406 ();
 FILLCELL_X32 FILLER_240_2438 ();
 FILLCELL_X32 FILLER_240_2470 ();
 FILLCELL_X32 FILLER_240_2502 ();
 FILLCELL_X32 FILLER_240_2534 ();
 FILLCELL_X32 FILLER_240_2566 ();
 FILLCELL_X32 FILLER_240_2598 ();
 FILLCELL_X32 FILLER_240_2630 ();
 FILLCELL_X32 FILLER_240_2662 ();
 FILLCELL_X32 FILLER_240_2694 ();
 FILLCELL_X32 FILLER_240_2726 ();
 FILLCELL_X32 FILLER_240_2758 ();
 FILLCELL_X32 FILLER_240_2790 ();
 FILLCELL_X32 FILLER_240_2822 ();
 FILLCELL_X32 FILLER_240_2854 ();
 FILLCELL_X32 FILLER_240_2886 ();
 FILLCELL_X32 FILLER_240_2918 ();
 FILLCELL_X32 FILLER_240_2950 ();
 FILLCELL_X32 FILLER_240_2982 ();
 FILLCELL_X32 FILLER_240_3014 ();
 FILLCELL_X32 FILLER_240_3046 ();
 FILLCELL_X32 FILLER_240_3078 ();
 FILLCELL_X32 FILLER_240_3110 ();
 FILLCELL_X8 FILLER_240_3142 ();
 FILLCELL_X4 FILLER_240_3150 ();
 FILLCELL_X2 FILLER_240_3154 ();
 FILLCELL_X1 FILLER_240_3156 ();
 FILLCELL_X32 FILLER_240_3158 ();
 FILLCELL_X32 FILLER_240_3190 ();
 FILLCELL_X32 FILLER_240_3222 ();
 FILLCELL_X32 FILLER_240_3254 ();
 FILLCELL_X32 FILLER_240_3286 ();
 FILLCELL_X32 FILLER_240_3318 ();
 FILLCELL_X32 FILLER_240_3350 ();
 FILLCELL_X32 FILLER_240_3382 ();
 FILLCELL_X32 FILLER_240_3414 ();
 FILLCELL_X32 FILLER_240_3446 ();
 FILLCELL_X32 FILLER_240_3478 ();
 FILLCELL_X32 FILLER_240_3510 ();
 FILLCELL_X32 FILLER_240_3542 ();
 FILLCELL_X32 FILLER_240_3574 ();
 FILLCELL_X32 FILLER_240_3606 ();
 FILLCELL_X32 FILLER_240_3638 ();
 FILLCELL_X32 FILLER_240_3670 ();
 FILLCELL_X32 FILLER_240_3702 ();
 FILLCELL_X4 FILLER_240_3734 ();
 FILLCELL_X32 FILLER_241_1 ();
 FILLCELL_X32 FILLER_241_33 ();
 FILLCELL_X32 FILLER_241_65 ();
 FILLCELL_X32 FILLER_241_97 ();
 FILLCELL_X32 FILLER_241_129 ();
 FILLCELL_X32 FILLER_241_161 ();
 FILLCELL_X32 FILLER_241_193 ();
 FILLCELL_X32 FILLER_241_225 ();
 FILLCELL_X32 FILLER_241_257 ();
 FILLCELL_X32 FILLER_241_289 ();
 FILLCELL_X32 FILLER_241_321 ();
 FILLCELL_X32 FILLER_241_353 ();
 FILLCELL_X32 FILLER_241_385 ();
 FILLCELL_X32 FILLER_241_417 ();
 FILLCELL_X32 FILLER_241_449 ();
 FILLCELL_X32 FILLER_241_481 ();
 FILLCELL_X32 FILLER_241_513 ();
 FILLCELL_X32 FILLER_241_545 ();
 FILLCELL_X32 FILLER_241_577 ();
 FILLCELL_X32 FILLER_241_609 ();
 FILLCELL_X32 FILLER_241_641 ();
 FILLCELL_X32 FILLER_241_673 ();
 FILLCELL_X32 FILLER_241_705 ();
 FILLCELL_X32 FILLER_241_737 ();
 FILLCELL_X32 FILLER_241_769 ();
 FILLCELL_X32 FILLER_241_801 ();
 FILLCELL_X32 FILLER_241_833 ();
 FILLCELL_X32 FILLER_241_865 ();
 FILLCELL_X32 FILLER_241_897 ();
 FILLCELL_X32 FILLER_241_929 ();
 FILLCELL_X32 FILLER_241_961 ();
 FILLCELL_X32 FILLER_241_993 ();
 FILLCELL_X32 FILLER_241_1025 ();
 FILLCELL_X32 FILLER_241_1057 ();
 FILLCELL_X32 FILLER_241_1089 ();
 FILLCELL_X32 FILLER_241_1121 ();
 FILLCELL_X32 FILLER_241_1153 ();
 FILLCELL_X32 FILLER_241_1185 ();
 FILLCELL_X32 FILLER_241_1217 ();
 FILLCELL_X8 FILLER_241_1249 ();
 FILLCELL_X4 FILLER_241_1257 ();
 FILLCELL_X2 FILLER_241_1261 ();
 FILLCELL_X32 FILLER_241_1264 ();
 FILLCELL_X32 FILLER_241_1296 ();
 FILLCELL_X32 FILLER_241_1328 ();
 FILLCELL_X32 FILLER_241_1360 ();
 FILLCELL_X32 FILLER_241_1392 ();
 FILLCELL_X32 FILLER_241_1424 ();
 FILLCELL_X32 FILLER_241_1456 ();
 FILLCELL_X32 FILLER_241_1488 ();
 FILLCELL_X32 FILLER_241_1520 ();
 FILLCELL_X32 FILLER_241_1552 ();
 FILLCELL_X32 FILLER_241_1584 ();
 FILLCELL_X32 FILLER_241_1616 ();
 FILLCELL_X32 FILLER_241_1648 ();
 FILLCELL_X32 FILLER_241_1680 ();
 FILLCELL_X32 FILLER_241_1712 ();
 FILLCELL_X32 FILLER_241_1744 ();
 FILLCELL_X32 FILLER_241_1776 ();
 FILLCELL_X32 FILLER_241_1808 ();
 FILLCELL_X32 FILLER_241_1840 ();
 FILLCELL_X16 FILLER_241_1872 ();
 FILLCELL_X4 FILLER_241_1888 ();
 FILLCELL_X2 FILLER_241_1892 ();
 FILLCELL_X8 FILLER_241_1913 ();
 FILLCELL_X2 FILLER_241_1921 ();
 FILLCELL_X2 FILLER_241_1927 ();
 FILLCELL_X4 FILLER_241_1936 ();
 FILLCELL_X1 FILLER_241_1956 ();
 FILLCELL_X1 FILLER_241_1964 ();
 FILLCELL_X1 FILLER_241_1978 ();
 FILLCELL_X16 FILLER_241_1989 ();
 FILLCELL_X8 FILLER_241_2005 ();
 FILLCELL_X4 FILLER_241_2013 ();
 FILLCELL_X2 FILLER_241_2017 ();
 FILLCELL_X32 FILLER_241_2036 ();
 FILLCELL_X32 FILLER_241_2068 ();
 FILLCELL_X16 FILLER_241_2100 ();
 FILLCELL_X4 FILLER_241_2116 ();
 FILLCELL_X2 FILLER_241_2120 ();
 FILLCELL_X1 FILLER_241_2122 ();
 FILLCELL_X16 FILLER_241_2130 ();
 FILLCELL_X4 FILLER_241_2146 ();
 FILLCELL_X2 FILLER_241_2150 ();
 FILLCELL_X32 FILLER_241_2186 ();
 FILLCELL_X2 FILLER_241_2218 ();
 FILLCELL_X4 FILLER_241_2227 ();
 FILLCELL_X1 FILLER_241_2231 ();
 FILLCELL_X2 FILLER_241_2239 ();
 FILLCELL_X1 FILLER_241_2241 ();
 FILLCELL_X32 FILLER_241_2259 ();
 FILLCELL_X32 FILLER_241_2291 ();
 FILLCELL_X32 FILLER_241_2323 ();
 FILLCELL_X32 FILLER_241_2355 ();
 FILLCELL_X32 FILLER_241_2387 ();
 FILLCELL_X32 FILLER_241_2419 ();
 FILLCELL_X32 FILLER_241_2451 ();
 FILLCELL_X32 FILLER_241_2483 ();
 FILLCELL_X8 FILLER_241_2515 ();
 FILLCELL_X2 FILLER_241_2523 ();
 FILLCELL_X1 FILLER_241_2525 ();
 FILLCELL_X32 FILLER_241_2527 ();
 FILLCELL_X32 FILLER_241_2559 ();
 FILLCELL_X32 FILLER_241_2591 ();
 FILLCELL_X32 FILLER_241_2623 ();
 FILLCELL_X32 FILLER_241_2655 ();
 FILLCELL_X32 FILLER_241_2687 ();
 FILLCELL_X32 FILLER_241_2719 ();
 FILLCELL_X32 FILLER_241_2751 ();
 FILLCELL_X32 FILLER_241_2783 ();
 FILLCELL_X32 FILLER_241_2815 ();
 FILLCELL_X32 FILLER_241_2847 ();
 FILLCELL_X32 FILLER_241_2879 ();
 FILLCELL_X32 FILLER_241_2911 ();
 FILLCELL_X32 FILLER_241_2943 ();
 FILLCELL_X32 FILLER_241_2975 ();
 FILLCELL_X32 FILLER_241_3007 ();
 FILLCELL_X32 FILLER_241_3039 ();
 FILLCELL_X32 FILLER_241_3071 ();
 FILLCELL_X32 FILLER_241_3103 ();
 FILLCELL_X32 FILLER_241_3135 ();
 FILLCELL_X32 FILLER_241_3167 ();
 FILLCELL_X32 FILLER_241_3199 ();
 FILLCELL_X32 FILLER_241_3231 ();
 FILLCELL_X32 FILLER_241_3263 ();
 FILLCELL_X32 FILLER_241_3295 ();
 FILLCELL_X32 FILLER_241_3327 ();
 FILLCELL_X32 FILLER_241_3359 ();
 FILLCELL_X32 FILLER_241_3391 ();
 FILLCELL_X32 FILLER_241_3423 ();
 FILLCELL_X32 FILLER_241_3455 ();
 FILLCELL_X32 FILLER_241_3487 ();
 FILLCELL_X32 FILLER_241_3519 ();
 FILLCELL_X32 FILLER_241_3551 ();
 FILLCELL_X32 FILLER_241_3583 ();
 FILLCELL_X32 FILLER_241_3615 ();
 FILLCELL_X32 FILLER_241_3647 ();
 FILLCELL_X32 FILLER_241_3679 ();
 FILLCELL_X16 FILLER_241_3711 ();
 FILLCELL_X8 FILLER_241_3727 ();
 FILLCELL_X2 FILLER_241_3735 ();
 FILLCELL_X1 FILLER_241_3737 ();
 FILLCELL_X32 FILLER_242_1 ();
 FILLCELL_X32 FILLER_242_33 ();
 FILLCELL_X32 FILLER_242_65 ();
 FILLCELL_X32 FILLER_242_97 ();
 FILLCELL_X32 FILLER_242_129 ();
 FILLCELL_X32 FILLER_242_161 ();
 FILLCELL_X32 FILLER_242_193 ();
 FILLCELL_X32 FILLER_242_225 ();
 FILLCELL_X32 FILLER_242_257 ();
 FILLCELL_X32 FILLER_242_289 ();
 FILLCELL_X32 FILLER_242_321 ();
 FILLCELL_X32 FILLER_242_353 ();
 FILLCELL_X32 FILLER_242_385 ();
 FILLCELL_X32 FILLER_242_417 ();
 FILLCELL_X32 FILLER_242_449 ();
 FILLCELL_X32 FILLER_242_481 ();
 FILLCELL_X32 FILLER_242_513 ();
 FILLCELL_X32 FILLER_242_545 ();
 FILLCELL_X32 FILLER_242_577 ();
 FILLCELL_X16 FILLER_242_609 ();
 FILLCELL_X4 FILLER_242_625 ();
 FILLCELL_X2 FILLER_242_629 ();
 FILLCELL_X32 FILLER_242_632 ();
 FILLCELL_X32 FILLER_242_664 ();
 FILLCELL_X32 FILLER_242_696 ();
 FILLCELL_X32 FILLER_242_728 ();
 FILLCELL_X32 FILLER_242_760 ();
 FILLCELL_X32 FILLER_242_792 ();
 FILLCELL_X32 FILLER_242_824 ();
 FILLCELL_X32 FILLER_242_856 ();
 FILLCELL_X32 FILLER_242_888 ();
 FILLCELL_X32 FILLER_242_920 ();
 FILLCELL_X32 FILLER_242_952 ();
 FILLCELL_X32 FILLER_242_984 ();
 FILLCELL_X32 FILLER_242_1016 ();
 FILLCELL_X32 FILLER_242_1048 ();
 FILLCELL_X32 FILLER_242_1080 ();
 FILLCELL_X32 FILLER_242_1112 ();
 FILLCELL_X32 FILLER_242_1144 ();
 FILLCELL_X32 FILLER_242_1176 ();
 FILLCELL_X32 FILLER_242_1208 ();
 FILLCELL_X32 FILLER_242_1240 ();
 FILLCELL_X32 FILLER_242_1272 ();
 FILLCELL_X32 FILLER_242_1304 ();
 FILLCELL_X32 FILLER_242_1336 ();
 FILLCELL_X32 FILLER_242_1368 ();
 FILLCELL_X32 FILLER_242_1400 ();
 FILLCELL_X32 FILLER_242_1432 ();
 FILLCELL_X32 FILLER_242_1464 ();
 FILLCELL_X32 FILLER_242_1496 ();
 FILLCELL_X32 FILLER_242_1528 ();
 FILLCELL_X32 FILLER_242_1560 ();
 FILLCELL_X32 FILLER_242_1592 ();
 FILLCELL_X32 FILLER_242_1624 ();
 FILLCELL_X32 FILLER_242_1656 ();
 FILLCELL_X32 FILLER_242_1688 ();
 FILLCELL_X32 FILLER_242_1720 ();
 FILLCELL_X32 FILLER_242_1752 ();
 FILLCELL_X32 FILLER_242_1784 ();
 FILLCELL_X32 FILLER_242_1816 ();
 FILLCELL_X16 FILLER_242_1848 ();
 FILLCELL_X4 FILLER_242_1864 ();
 FILLCELL_X16 FILLER_242_1877 ();
 FILLCELL_X1 FILLER_242_1893 ();
 FILLCELL_X32 FILLER_242_1895 ();
 FILLCELL_X32 FILLER_242_1932 ();
 FILLCELL_X2 FILLER_242_1964 ();
 FILLCELL_X1 FILLER_242_1966 ();
 FILLCELL_X8 FILLER_242_1972 ();
 FILLCELL_X16 FILLER_242_1993 ();
 FILLCELL_X4 FILLER_242_2009 ();
 FILLCELL_X2 FILLER_242_2013 ();
 FILLCELL_X1 FILLER_242_2015 ();
 FILLCELL_X32 FILLER_242_2023 ();
 FILLCELL_X16 FILLER_242_2055 ();
 FILLCELL_X8 FILLER_242_2071 ();
 FILLCELL_X4 FILLER_242_2079 ();
 FILLCELL_X1 FILLER_242_2083 ();
 FILLCELL_X32 FILLER_242_2091 ();
 FILLCELL_X2 FILLER_242_2123 ();
 FILLCELL_X8 FILLER_242_2142 ();
 FILLCELL_X4 FILLER_242_2150 ();
 FILLCELL_X8 FILLER_242_2161 ();
 FILLCELL_X4 FILLER_242_2169 ();
 FILLCELL_X1 FILLER_242_2173 ();
 FILLCELL_X32 FILLER_242_2181 ();
 FILLCELL_X32 FILLER_242_2213 ();
 FILLCELL_X8 FILLER_242_2245 ();
 FILLCELL_X4 FILLER_242_2253 ();
 FILLCELL_X2 FILLER_242_2257 ();
 FILLCELL_X32 FILLER_242_2283 ();
 FILLCELL_X32 FILLER_242_2315 ();
 FILLCELL_X32 FILLER_242_2347 ();
 FILLCELL_X32 FILLER_242_2379 ();
 FILLCELL_X32 FILLER_242_2411 ();
 FILLCELL_X32 FILLER_242_2443 ();
 FILLCELL_X32 FILLER_242_2475 ();
 FILLCELL_X32 FILLER_242_2507 ();
 FILLCELL_X32 FILLER_242_2539 ();
 FILLCELL_X32 FILLER_242_2571 ();
 FILLCELL_X32 FILLER_242_2603 ();
 FILLCELL_X32 FILLER_242_2635 ();
 FILLCELL_X32 FILLER_242_2667 ();
 FILLCELL_X32 FILLER_242_2699 ();
 FILLCELL_X32 FILLER_242_2731 ();
 FILLCELL_X32 FILLER_242_2763 ();
 FILLCELL_X32 FILLER_242_2795 ();
 FILLCELL_X32 FILLER_242_2827 ();
 FILLCELL_X32 FILLER_242_2859 ();
 FILLCELL_X32 FILLER_242_2891 ();
 FILLCELL_X32 FILLER_242_2923 ();
 FILLCELL_X32 FILLER_242_2955 ();
 FILLCELL_X32 FILLER_242_2987 ();
 FILLCELL_X32 FILLER_242_3019 ();
 FILLCELL_X32 FILLER_242_3051 ();
 FILLCELL_X32 FILLER_242_3083 ();
 FILLCELL_X32 FILLER_242_3115 ();
 FILLCELL_X8 FILLER_242_3147 ();
 FILLCELL_X2 FILLER_242_3155 ();
 FILLCELL_X32 FILLER_242_3158 ();
 FILLCELL_X32 FILLER_242_3190 ();
 FILLCELL_X32 FILLER_242_3222 ();
 FILLCELL_X32 FILLER_242_3254 ();
 FILLCELL_X32 FILLER_242_3286 ();
 FILLCELL_X32 FILLER_242_3318 ();
 FILLCELL_X32 FILLER_242_3350 ();
 FILLCELL_X32 FILLER_242_3382 ();
 FILLCELL_X32 FILLER_242_3414 ();
 FILLCELL_X32 FILLER_242_3446 ();
 FILLCELL_X32 FILLER_242_3478 ();
 FILLCELL_X32 FILLER_242_3510 ();
 FILLCELL_X32 FILLER_242_3542 ();
 FILLCELL_X32 FILLER_242_3574 ();
 FILLCELL_X32 FILLER_242_3606 ();
 FILLCELL_X32 FILLER_242_3638 ();
 FILLCELL_X32 FILLER_242_3670 ();
 FILLCELL_X32 FILLER_242_3702 ();
 FILLCELL_X4 FILLER_242_3734 ();
 FILLCELL_X32 FILLER_243_1 ();
 FILLCELL_X32 FILLER_243_33 ();
 FILLCELL_X32 FILLER_243_65 ();
 FILLCELL_X32 FILLER_243_97 ();
 FILLCELL_X32 FILLER_243_129 ();
 FILLCELL_X32 FILLER_243_161 ();
 FILLCELL_X32 FILLER_243_193 ();
 FILLCELL_X32 FILLER_243_225 ();
 FILLCELL_X32 FILLER_243_257 ();
 FILLCELL_X32 FILLER_243_289 ();
 FILLCELL_X32 FILLER_243_321 ();
 FILLCELL_X32 FILLER_243_353 ();
 FILLCELL_X32 FILLER_243_385 ();
 FILLCELL_X32 FILLER_243_417 ();
 FILLCELL_X32 FILLER_243_449 ();
 FILLCELL_X32 FILLER_243_481 ();
 FILLCELL_X32 FILLER_243_513 ();
 FILLCELL_X32 FILLER_243_545 ();
 FILLCELL_X32 FILLER_243_577 ();
 FILLCELL_X32 FILLER_243_609 ();
 FILLCELL_X32 FILLER_243_641 ();
 FILLCELL_X32 FILLER_243_673 ();
 FILLCELL_X32 FILLER_243_705 ();
 FILLCELL_X32 FILLER_243_737 ();
 FILLCELL_X32 FILLER_243_769 ();
 FILLCELL_X32 FILLER_243_801 ();
 FILLCELL_X32 FILLER_243_833 ();
 FILLCELL_X32 FILLER_243_865 ();
 FILLCELL_X32 FILLER_243_897 ();
 FILLCELL_X32 FILLER_243_929 ();
 FILLCELL_X32 FILLER_243_961 ();
 FILLCELL_X32 FILLER_243_993 ();
 FILLCELL_X32 FILLER_243_1025 ();
 FILLCELL_X32 FILLER_243_1057 ();
 FILLCELL_X32 FILLER_243_1089 ();
 FILLCELL_X32 FILLER_243_1121 ();
 FILLCELL_X32 FILLER_243_1153 ();
 FILLCELL_X32 FILLER_243_1185 ();
 FILLCELL_X32 FILLER_243_1217 ();
 FILLCELL_X8 FILLER_243_1249 ();
 FILLCELL_X4 FILLER_243_1257 ();
 FILLCELL_X2 FILLER_243_1261 ();
 FILLCELL_X32 FILLER_243_1264 ();
 FILLCELL_X32 FILLER_243_1296 ();
 FILLCELL_X32 FILLER_243_1328 ();
 FILLCELL_X32 FILLER_243_1360 ();
 FILLCELL_X32 FILLER_243_1392 ();
 FILLCELL_X32 FILLER_243_1424 ();
 FILLCELL_X32 FILLER_243_1456 ();
 FILLCELL_X32 FILLER_243_1488 ();
 FILLCELL_X32 FILLER_243_1520 ();
 FILLCELL_X32 FILLER_243_1552 ();
 FILLCELL_X32 FILLER_243_1584 ();
 FILLCELL_X32 FILLER_243_1616 ();
 FILLCELL_X32 FILLER_243_1648 ();
 FILLCELL_X32 FILLER_243_1680 ();
 FILLCELL_X32 FILLER_243_1712 ();
 FILLCELL_X32 FILLER_243_1744 ();
 FILLCELL_X32 FILLER_243_1776 ();
 FILLCELL_X32 FILLER_243_1808 ();
 FILLCELL_X16 FILLER_243_1840 ();
 FILLCELL_X2 FILLER_243_1856 ();
 FILLCELL_X1 FILLER_243_1858 ();
 FILLCELL_X32 FILLER_243_1872 ();
 FILLCELL_X8 FILLER_243_1904 ();
 FILLCELL_X4 FILLER_243_1912 ();
 FILLCELL_X1 FILLER_243_1916 ();
 FILLCELL_X32 FILLER_243_1930 ();
 FILLCELL_X4 FILLER_243_1962 ();
 FILLCELL_X2 FILLER_243_1966 ();
 FILLCELL_X2 FILLER_243_1981 ();
 FILLCELL_X1 FILLER_243_1983 ();
 FILLCELL_X8 FILLER_243_1997 ();
 FILLCELL_X2 FILLER_243_2005 ();
 FILLCELL_X1 FILLER_243_2007 ();
 FILLCELL_X32 FILLER_243_2025 ();
 FILLCELL_X8 FILLER_243_2057 ();
 FILLCELL_X4 FILLER_243_2065 ();
 FILLCELL_X2 FILLER_243_2069 ();
 FILLCELL_X1 FILLER_243_2071 ();
 FILLCELL_X2 FILLER_243_2079 ();
 FILLCELL_X16 FILLER_243_2098 ();
 FILLCELL_X8 FILLER_243_2114 ();
 FILLCELL_X2 FILLER_243_2122 ();
 FILLCELL_X4 FILLER_243_2136 ();
 FILLCELL_X1 FILLER_243_2140 ();
 FILLCELL_X32 FILLER_243_2165 ();
 FILLCELL_X32 FILLER_243_2197 ();
 FILLCELL_X8 FILLER_243_2229 ();
 FILLCELL_X32 FILLER_243_2242 ();
 FILLCELL_X32 FILLER_243_2274 ();
 FILLCELL_X32 FILLER_243_2306 ();
 FILLCELL_X32 FILLER_243_2338 ();
 FILLCELL_X32 FILLER_243_2370 ();
 FILLCELL_X32 FILLER_243_2402 ();
 FILLCELL_X32 FILLER_243_2434 ();
 FILLCELL_X32 FILLER_243_2466 ();
 FILLCELL_X16 FILLER_243_2498 ();
 FILLCELL_X8 FILLER_243_2514 ();
 FILLCELL_X4 FILLER_243_2522 ();
 FILLCELL_X32 FILLER_243_2527 ();
 FILLCELL_X32 FILLER_243_2559 ();
 FILLCELL_X32 FILLER_243_2591 ();
 FILLCELL_X32 FILLER_243_2623 ();
 FILLCELL_X32 FILLER_243_2655 ();
 FILLCELL_X32 FILLER_243_2687 ();
 FILLCELL_X32 FILLER_243_2719 ();
 FILLCELL_X32 FILLER_243_2751 ();
 FILLCELL_X32 FILLER_243_2783 ();
 FILLCELL_X32 FILLER_243_2815 ();
 FILLCELL_X32 FILLER_243_2847 ();
 FILLCELL_X32 FILLER_243_2879 ();
 FILLCELL_X32 FILLER_243_2911 ();
 FILLCELL_X32 FILLER_243_2943 ();
 FILLCELL_X32 FILLER_243_2975 ();
 FILLCELL_X32 FILLER_243_3007 ();
 FILLCELL_X32 FILLER_243_3039 ();
 FILLCELL_X32 FILLER_243_3071 ();
 FILLCELL_X32 FILLER_243_3103 ();
 FILLCELL_X32 FILLER_243_3135 ();
 FILLCELL_X32 FILLER_243_3167 ();
 FILLCELL_X32 FILLER_243_3199 ();
 FILLCELL_X32 FILLER_243_3231 ();
 FILLCELL_X32 FILLER_243_3263 ();
 FILLCELL_X32 FILLER_243_3295 ();
 FILLCELL_X32 FILLER_243_3327 ();
 FILLCELL_X32 FILLER_243_3359 ();
 FILLCELL_X32 FILLER_243_3391 ();
 FILLCELL_X32 FILLER_243_3423 ();
 FILLCELL_X32 FILLER_243_3455 ();
 FILLCELL_X32 FILLER_243_3487 ();
 FILLCELL_X32 FILLER_243_3519 ();
 FILLCELL_X32 FILLER_243_3551 ();
 FILLCELL_X32 FILLER_243_3583 ();
 FILLCELL_X32 FILLER_243_3615 ();
 FILLCELL_X32 FILLER_243_3647 ();
 FILLCELL_X32 FILLER_243_3679 ();
 FILLCELL_X16 FILLER_243_3711 ();
 FILLCELL_X8 FILLER_243_3727 ();
 FILLCELL_X2 FILLER_243_3735 ();
 FILLCELL_X1 FILLER_243_3737 ();
 FILLCELL_X32 FILLER_244_1 ();
 FILLCELL_X32 FILLER_244_33 ();
 FILLCELL_X32 FILLER_244_65 ();
 FILLCELL_X32 FILLER_244_97 ();
 FILLCELL_X32 FILLER_244_129 ();
 FILLCELL_X32 FILLER_244_161 ();
 FILLCELL_X32 FILLER_244_193 ();
 FILLCELL_X32 FILLER_244_225 ();
 FILLCELL_X32 FILLER_244_257 ();
 FILLCELL_X32 FILLER_244_289 ();
 FILLCELL_X32 FILLER_244_321 ();
 FILLCELL_X32 FILLER_244_353 ();
 FILLCELL_X32 FILLER_244_385 ();
 FILLCELL_X32 FILLER_244_417 ();
 FILLCELL_X32 FILLER_244_449 ();
 FILLCELL_X32 FILLER_244_481 ();
 FILLCELL_X32 FILLER_244_513 ();
 FILLCELL_X32 FILLER_244_545 ();
 FILLCELL_X32 FILLER_244_577 ();
 FILLCELL_X16 FILLER_244_609 ();
 FILLCELL_X4 FILLER_244_625 ();
 FILLCELL_X2 FILLER_244_629 ();
 FILLCELL_X32 FILLER_244_632 ();
 FILLCELL_X32 FILLER_244_664 ();
 FILLCELL_X32 FILLER_244_696 ();
 FILLCELL_X32 FILLER_244_728 ();
 FILLCELL_X32 FILLER_244_760 ();
 FILLCELL_X32 FILLER_244_792 ();
 FILLCELL_X32 FILLER_244_824 ();
 FILLCELL_X32 FILLER_244_856 ();
 FILLCELL_X32 FILLER_244_888 ();
 FILLCELL_X32 FILLER_244_920 ();
 FILLCELL_X32 FILLER_244_952 ();
 FILLCELL_X32 FILLER_244_984 ();
 FILLCELL_X32 FILLER_244_1016 ();
 FILLCELL_X32 FILLER_244_1048 ();
 FILLCELL_X32 FILLER_244_1080 ();
 FILLCELL_X32 FILLER_244_1112 ();
 FILLCELL_X32 FILLER_244_1144 ();
 FILLCELL_X32 FILLER_244_1176 ();
 FILLCELL_X32 FILLER_244_1208 ();
 FILLCELL_X32 FILLER_244_1240 ();
 FILLCELL_X32 FILLER_244_1272 ();
 FILLCELL_X32 FILLER_244_1304 ();
 FILLCELL_X32 FILLER_244_1336 ();
 FILLCELL_X32 FILLER_244_1368 ();
 FILLCELL_X32 FILLER_244_1400 ();
 FILLCELL_X32 FILLER_244_1432 ();
 FILLCELL_X32 FILLER_244_1464 ();
 FILLCELL_X32 FILLER_244_1496 ();
 FILLCELL_X32 FILLER_244_1528 ();
 FILLCELL_X32 FILLER_244_1560 ();
 FILLCELL_X32 FILLER_244_1592 ();
 FILLCELL_X32 FILLER_244_1624 ();
 FILLCELL_X32 FILLER_244_1656 ();
 FILLCELL_X32 FILLER_244_1688 ();
 FILLCELL_X32 FILLER_244_1720 ();
 FILLCELL_X32 FILLER_244_1752 ();
 FILLCELL_X8 FILLER_244_1784 ();
 FILLCELL_X4 FILLER_244_1792 ();
 FILLCELL_X1 FILLER_244_1796 ();
 FILLCELL_X32 FILLER_244_1805 ();
 FILLCELL_X8 FILLER_244_1837 ();
 FILLCELL_X1 FILLER_244_1845 ();
 FILLCELL_X16 FILLER_244_1870 ();
 FILLCELL_X8 FILLER_244_1886 ();
 FILLCELL_X32 FILLER_244_1895 ();
 FILLCELL_X8 FILLER_244_1927 ();
 FILLCELL_X2 FILLER_244_1935 ();
 FILLCELL_X16 FILLER_244_1944 ();
 FILLCELL_X1 FILLER_244_1960 ();
 FILLCELL_X32 FILLER_244_1977 ();
 FILLCELL_X8 FILLER_244_2009 ();
 FILLCELL_X32 FILLER_244_2024 ();
 FILLCELL_X4 FILLER_244_2056 ();
 FILLCELL_X2 FILLER_244_2060 ();
 FILLCELL_X4 FILLER_244_2086 ();
 FILLCELL_X2 FILLER_244_2090 ();
 FILLCELL_X1 FILLER_244_2092 ();
 FILLCELL_X8 FILLER_244_2100 ();
 FILLCELL_X2 FILLER_244_2108 ();
 FILLCELL_X16 FILLER_244_2134 ();
 FILLCELL_X8 FILLER_244_2150 ();
 FILLCELL_X4 FILLER_244_2158 ();
 FILLCELL_X4 FILLER_244_2186 ();
 FILLCELL_X8 FILLER_244_2214 ();
 FILLCELL_X4 FILLER_244_2222 ();
 FILLCELL_X2 FILLER_244_2226 ();
 FILLCELL_X2 FILLER_244_2235 ();
 FILLCELL_X4 FILLER_244_2261 ();
 FILLCELL_X2 FILLER_244_2265 ();
 FILLCELL_X1 FILLER_244_2267 ();
 FILLCELL_X32 FILLER_244_2275 ();
 FILLCELL_X32 FILLER_244_2307 ();
 FILLCELL_X32 FILLER_244_2339 ();
 FILLCELL_X32 FILLER_244_2371 ();
 FILLCELL_X32 FILLER_244_2403 ();
 FILLCELL_X32 FILLER_244_2435 ();
 FILLCELL_X32 FILLER_244_2467 ();
 FILLCELL_X32 FILLER_244_2499 ();
 FILLCELL_X32 FILLER_244_2531 ();
 FILLCELL_X32 FILLER_244_2563 ();
 FILLCELL_X32 FILLER_244_2595 ();
 FILLCELL_X32 FILLER_244_2627 ();
 FILLCELL_X32 FILLER_244_2659 ();
 FILLCELL_X32 FILLER_244_2691 ();
 FILLCELL_X32 FILLER_244_2723 ();
 FILLCELL_X32 FILLER_244_2755 ();
 FILLCELL_X32 FILLER_244_2787 ();
 FILLCELL_X32 FILLER_244_2819 ();
 FILLCELL_X32 FILLER_244_2851 ();
 FILLCELL_X32 FILLER_244_2883 ();
 FILLCELL_X32 FILLER_244_2915 ();
 FILLCELL_X32 FILLER_244_2947 ();
 FILLCELL_X32 FILLER_244_2979 ();
 FILLCELL_X32 FILLER_244_3011 ();
 FILLCELL_X32 FILLER_244_3043 ();
 FILLCELL_X32 FILLER_244_3075 ();
 FILLCELL_X32 FILLER_244_3107 ();
 FILLCELL_X16 FILLER_244_3139 ();
 FILLCELL_X2 FILLER_244_3155 ();
 FILLCELL_X32 FILLER_244_3158 ();
 FILLCELL_X32 FILLER_244_3190 ();
 FILLCELL_X32 FILLER_244_3222 ();
 FILLCELL_X32 FILLER_244_3254 ();
 FILLCELL_X32 FILLER_244_3286 ();
 FILLCELL_X32 FILLER_244_3318 ();
 FILLCELL_X32 FILLER_244_3350 ();
 FILLCELL_X32 FILLER_244_3382 ();
 FILLCELL_X32 FILLER_244_3414 ();
 FILLCELL_X32 FILLER_244_3446 ();
 FILLCELL_X32 FILLER_244_3478 ();
 FILLCELL_X32 FILLER_244_3510 ();
 FILLCELL_X32 FILLER_244_3542 ();
 FILLCELL_X32 FILLER_244_3574 ();
 FILLCELL_X32 FILLER_244_3606 ();
 FILLCELL_X32 FILLER_244_3638 ();
 FILLCELL_X32 FILLER_244_3670 ();
 FILLCELL_X32 FILLER_244_3702 ();
 FILLCELL_X4 FILLER_244_3734 ();
 FILLCELL_X32 FILLER_245_1 ();
 FILLCELL_X32 FILLER_245_33 ();
 FILLCELL_X32 FILLER_245_65 ();
 FILLCELL_X32 FILLER_245_97 ();
 FILLCELL_X32 FILLER_245_129 ();
 FILLCELL_X32 FILLER_245_161 ();
 FILLCELL_X32 FILLER_245_193 ();
 FILLCELL_X32 FILLER_245_225 ();
 FILLCELL_X32 FILLER_245_257 ();
 FILLCELL_X32 FILLER_245_289 ();
 FILLCELL_X32 FILLER_245_321 ();
 FILLCELL_X32 FILLER_245_353 ();
 FILLCELL_X32 FILLER_245_385 ();
 FILLCELL_X32 FILLER_245_417 ();
 FILLCELL_X32 FILLER_245_449 ();
 FILLCELL_X32 FILLER_245_481 ();
 FILLCELL_X32 FILLER_245_513 ();
 FILLCELL_X32 FILLER_245_545 ();
 FILLCELL_X32 FILLER_245_577 ();
 FILLCELL_X32 FILLER_245_609 ();
 FILLCELL_X32 FILLER_245_641 ();
 FILLCELL_X32 FILLER_245_673 ();
 FILLCELL_X32 FILLER_245_705 ();
 FILLCELL_X32 FILLER_245_737 ();
 FILLCELL_X32 FILLER_245_769 ();
 FILLCELL_X32 FILLER_245_801 ();
 FILLCELL_X32 FILLER_245_833 ();
 FILLCELL_X32 FILLER_245_865 ();
 FILLCELL_X32 FILLER_245_897 ();
 FILLCELL_X32 FILLER_245_929 ();
 FILLCELL_X32 FILLER_245_961 ();
 FILLCELL_X32 FILLER_245_993 ();
 FILLCELL_X32 FILLER_245_1025 ();
 FILLCELL_X32 FILLER_245_1057 ();
 FILLCELL_X32 FILLER_245_1089 ();
 FILLCELL_X32 FILLER_245_1121 ();
 FILLCELL_X32 FILLER_245_1153 ();
 FILLCELL_X32 FILLER_245_1185 ();
 FILLCELL_X32 FILLER_245_1217 ();
 FILLCELL_X8 FILLER_245_1249 ();
 FILLCELL_X4 FILLER_245_1257 ();
 FILLCELL_X2 FILLER_245_1261 ();
 FILLCELL_X32 FILLER_245_1264 ();
 FILLCELL_X32 FILLER_245_1296 ();
 FILLCELL_X32 FILLER_245_1328 ();
 FILLCELL_X32 FILLER_245_1360 ();
 FILLCELL_X32 FILLER_245_1392 ();
 FILLCELL_X32 FILLER_245_1424 ();
 FILLCELL_X32 FILLER_245_1456 ();
 FILLCELL_X32 FILLER_245_1488 ();
 FILLCELL_X32 FILLER_245_1520 ();
 FILLCELL_X32 FILLER_245_1552 ();
 FILLCELL_X32 FILLER_245_1584 ();
 FILLCELL_X32 FILLER_245_1616 ();
 FILLCELL_X32 FILLER_245_1648 ();
 FILLCELL_X32 FILLER_245_1680 ();
 FILLCELL_X32 FILLER_245_1712 ();
 FILLCELL_X32 FILLER_245_1744 ();
 FILLCELL_X32 FILLER_245_1776 ();
 FILLCELL_X32 FILLER_245_1808 ();
 FILLCELL_X16 FILLER_245_1840 ();
 FILLCELL_X2 FILLER_245_1856 ();
 FILLCELL_X1 FILLER_245_1858 ();
 FILLCELL_X8 FILLER_245_1876 ();
 FILLCELL_X2 FILLER_245_1884 ();
 FILLCELL_X1 FILLER_245_1886 ();
 FILLCELL_X32 FILLER_245_1932 ();
 FILLCELL_X16 FILLER_245_1964 ();
 FILLCELL_X4 FILLER_245_1980 ();
 FILLCELL_X4 FILLER_245_1997 ();
 FILLCELL_X1 FILLER_245_2001 ();
 FILLCELL_X32 FILLER_245_2026 ();
 FILLCELL_X16 FILLER_245_2058 ();
 FILLCELL_X8 FILLER_245_2074 ();
 FILLCELL_X2 FILLER_245_2082 ();
 FILLCELL_X1 FILLER_245_2084 ();
 FILLCELL_X32 FILLER_245_2092 ();
 FILLCELL_X32 FILLER_245_2124 ();
 FILLCELL_X32 FILLER_245_2156 ();
 FILLCELL_X2 FILLER_245_2188 ();
 FILLCELL_X16 FILLER_245_2197 ();
 FILLCELL_X8 FILLER_245_2213 ();
 FILLCELL_X2 FILLER_245_2221 ();
 FILLCELL_X8 FILLER_245_2240 ();
 FILLCELL_X4 FILLER_245_2248 ();
 FILLCELL_X2 FILLER_245_2252 ();
 FILLCELL_X1 FILLER_245_2254 ();
 FILLCELL_X4 FILLER_245_2262 ();
 FILLCELL_X1 FILLER_245_2266 ();
 FILLCELL_X32 FILLER_245_2284 ();
 FILLCELL_X32 FILLER_245_2316 ();
 FILLCELL_X32 FILLER_245_2348 ();
 FILLCELL_X32 FILLER_245_2380 ();
 FILLCELL_X32 FILLER_245_2412 ();
 FILLCELL_X32 FILLER_245_2444 ();
 FILLCELL_X32 FILLER_245_2476 ();
 FILLCELL_X16 FILLER_245_2508 ();
 FILLCELL_X2 FILLER_245_2524 ();
 FILLCELL_X32 FILLER_245_2527 ();
 FILLCELL_X32 FILLER_245_2559 ();
 FILLCELL_X32 FILLER_245_2591 ();
 FILLCELL_X32 FILLER_245_2623 ();
 FILLCELL_X32 FILLER_245_2655 ();
 FILLCELL_X32 FILLER_245_2687 ();
 FILLCELL_X32 FILLER_245_2719 ();
 FILLCELL_X32 FILLER_245_2751 ();
 FILLCELL_X32 FILLER_245_2783 ();
 FILLCELL_X32 FILLER_245_2815 ();
 FILLCELL_X32 FILLER_245_2847 ();
 FILLCELL_X32 FILLER_245_2879 ();
 FILLCELL_X32 FILLER_245_2911 ();
 FILLCELL_X32 FILLER_245_2943 ();
 FILLCELL_X32 FILLER_245_2975 ();
 FILLCELL_X32 FILLER_245_3007 ();
 FILLCELL_X32 FILLER_245_3039 ();
 FILLCELL_X32 FILLER_245_3071 ();
 FILLCELL_X32 FILLER_245_3103 ();
 FILLCELL_X32 FILLER_245_3135 ();
 FILLCELL_X32 FILLER_245_3167 ();
 FILLCELL_X32 FILLER_245_3199 ();
 FILLCELL_X32 FILLER_245_3231 ();
 FILLCELL_X32 FILLER_245_3263 ();
 FILLCELL_X32 FILLER_245_3295 ();
 FILLCELL_X32 FILLER_245_3327 ();
 FILLCELL_X32 FILLER_245_3359 ();
 FILLCELL_X32 FILLER_245_3391 ();
 FILLCELL_X32 FILLER_245_3423 ();
 FILLCELL_X32 FILLER_245_3455 ();
 FILLCELL_X32 FILLER_245_3487 ();
 FILLCELL_X32 FILLER_245_3519 ();
 FILLCELL_X32 FILLER_245_3551 ();
 FILLCELL_X32 FILLER_245_3583 ();
 FILLCELL_X32 FILLER_245_3615 ();
 FILLCELL_X32 FILLER_245_3647 ();
 FILLCELL_X32 FILLER_245_3679 ();
 FILLCELL_X16 FILLER_245_3711 ();
 FILLCELL_X8 FILLER_245_3727 ();
 FILLCELL_X2 FILLER_245_3735 ();
 FILLCELL_X1 FILLER_245_3737 ();
 FILLCELL_X8 FILLER_246_1 ();
 FILLCELL_X32 FILLER_246_12 ();
 FILLCELL_X32 FILLER_246_44 ();
 FILLCELL_X32 FILLER_246_76 ();
 FILLCELL_X32 FILLER_246_108 ();
 FILLCELL_X32 FILLER_246_140 ();
 FILLCELL_X32 FILLER_246_172 ();
 FILLCELL_X32 FILLER_246_204 ();
 FILLCELL_X32 FILLER_246_236 ();
 FILLCELL_X32 FILLER_246_268 ();
 FILLCELL_X32 FILLER_246_300 ();
 FILLCELL_X32 FILLER_246_332 ();
 FILLCELL_X32 FILLER_246_364 ();
 FILLCELL_X32 FILLER_246_396 ();
 FILLCELL_X32 FILLER_246_428 ();
 FILLCELL_X32 FILLER_246_460 ();
 FILLCELL_X32 FILLER_246_492 ();
 FILLCELL_X32 FILLER_246_524 ();
 FILLCELL_X32 FILLER_246_556 ();
 FILLCELL_X32 FILLER_246_588 ();
 FILLCELL_X8 FILLER_246_620 ();
 FILLCELL_X2 FILLER_246_628 ();
 FILLCELL_X1 FILLER_246_630 ();
 FILLCELL_X32 FILLER_246_632 ();
 FILLCELL_X32 FILLER_246_664 ();
 FILLCELL_X32 FILLER_246_696 ();
 FILLCELL_X32 FILLER_246_728 ();
 FILLCELL_X32 FILLER_246_760 ();
 FILLCELL_X32 FILLER_246_792 ();
 FILLCELL_X32 FILLER_246_824 ();
 FILLCELL_X32 FILLER_246_856 ();
 FILLCELL_X32 FILLER_246_888 ();
 FILLCELL_X32 FILLER_246_920 ();
 FILLCELL_X32 FILLER_246_952 ();
 FILLCELL_X32 FILLER_246_984 ();
 FILLCELL_X32 FILLER_246_1016 ();
 FILLCELL_X32 FILLER_246_1048 ();
 FILLCELL_X32 FILLER_246_1080 ();
 FILLCELL_X32 FILLER_246_1112 ();
 FILLCELL_X32 FILLER_246_1144 ();
 FILLCELL_X32 FILLER_246_1176 ();
 FILLCELL_X32 FILLER_246_1208 ();
 FILLCELL_X32 FILLER_246_1240 ();
 FILLCELL_X32 FILLER_246_1272 ();
 FILLCELL_X32 FILLER_246_1304 ();
 FILLCELL_X32 FILLER_246_1336 ();
 FILLCELL_X32 FILLER_246_1368 ();
 FILLCELL_X32 FILLER_246_1400 ();
 FILLCELL_X32 FILLER_246_1432 ();
 FILLCELL_X32 FILLER_246_1464 ();
 FILLCELL_X32 FILLER_246_1496 ();
 FILLCELL_X32 FILLER_246_1528 ();
 FILLCELL_X32 FILLER_246_1560 ();
 FILLCELL_X32 FILLER_246_1592 ();
 FILLCELL_X32 FILLER_246_1624 ();
 FILLCELL_X32 FILLER_246_1656 ();
 FILLCELL_X32 FILLER_246_1688 ();
 FILLCELL_X32 FILLER_246_1720 ();
 FILLCELL_X32 FILLER_246_1752 ();
 FILLCELL_X32 FILLER_246_1784 ();
 FILLCELL_X32 FILLER_246_1816 ();
 FILLCELL_X8 FILLER_246_1848 ();
 FILLCELL_X2 FILLER_246_1856 ();
 FILLCELL_X8 FILLER_246_1872 ();
 FILLCELL_X4 FILLER_246_1880 ();
 FILLCELL_X4 FILLER_246_1888 ();
 FILLCELL_X2 FILLER_246_1892 ();
 FILLCELL_X4 FILLER_246_1895 ();
 FILLCELL_X1 FILLER_246_1899 ();
 FILLCELL_X4 FILLER_246_1910 ();
 FILLCELL_X8 FILLER_246_1918 ();
 FILLCELL_X1 FILLER_246_1931 ();
 FILLCELL_X8 FILLER_246_1936 ();
 FILLCELL_X2 FILLER_246_1944 ();
 FILLCELL_X1 FILLER_246_1946 ();
 FILLCELL_X1 FILLER_246_1960 ();
 FILLCELL_X8 FILLER_246_2000 ();
 FILLCELL_X2 FILLER_246_2008 ();
 FILLCELL_X1 FILLER_246_2010 ();
 FILLCELL_X8 FILLER_246_2018 ();
 FILLCELL_X2 FILLER_246_2026 ();
 FILLCELL_X1 FILLER_246_2028 ();
 FILLCELL_X8 FILLER_246_2036 ();
 FILLCELL_X4 FILLER_246_2044 ();
 FILLCELL_X8 FILLER_246_2072 ();
 FILLCELL_X4 FILLER_246_2080 ();
 FILLCELL_X2 FILLER_246_2084 ();
 FILLCELL_X16 FILLER_246_2093 ();
 FILLCELL_X8 FILLER_246_2109 ();
 FILLCELL_X4 FILLER_246_2117 ();
 FILLCELL_X2 FILLER_246_2121 ();
 FILLCELL_X1 FILLER_246_2123 ();
 FILLCELL_X4 FILLER_246_2131 ();
 FILLCELL_X2 FILLER_246_2135 ();
 FILLCELL_X1 FILLER_246_2137 ();
 FILLCELL_X32 FILLER_246_2145 ();
 FILLCELL_X32 FILLER_246_2177 ();
 FILLCELL_X16 FILLER_246_2209 ();
 FILLCELL_X8 FILLER_246_2225 ();
 FILLCELL_X2 FILLER_246_2233 ();
 FILLCELL_X32 FILLER_246_2242 ();
 FILLCELL_X32 FILLER_246_2274 ();
 FILLCELL_X32 FILLER_246_2306 ();
 FILLCELL_X32 FILLER_246_2338 ();
 FILLCELL_X32 FILLER_246_2370 ();
 FILLCELL_X32 FILLER_246_2402 ();
 FILLCELL_X32 FILLER_246_2434 ();
 FILLCELL_X32 FILLER_246_2466 ();
 FILLCELL_X32 FILLER_246_2498 ();
 FILLCELL_X32 FILLER_246_2530 ();
 FILLCELL_X32 FILLER_246_2562 ();
 FILLCELL_X32 FILLER_246_2594 ();
 FILLCELL_X32 FILLER_246_2626 ();
 FILLCELL_X32 FILLER_246_2658 ();
 FILLCELL_X32 FILLER_246_2690 ();
 FILLCELL_X32 FILLER_246_2722 ();
 FILLCELL_X32 FILLER_246_2754 ();
 FILLCELL_X32 FILLER_246_2786 ();
 FILLCELL_X32 FILLER_246_2818 ();
 FILLCELL_X32 FILLER_246_2850 ();
 FILLCELL_X32 FILLER_246_2882 ();
 FILLCELL_X32 FILLER_246_2914 ();
 FILLCELL_X32 FILLER_246_2946 ();
 FILLCELL_X32 FILLER_246_2978 ();
 FILLCELL_X32 FILLER_246_3010 ();
 FILLCELL_X32 FILLER_246_3042 ();
 FILLCELL_X32 FILLER_246_3074 ();
 FILLCELL_X32 FILLER_246_3106 ();
 FILLCELL_X16 FILLER_246_3138 ();
 FILLCELL_X2 FILLER_246_3154 ();
 FILLCELL_X1 FILLER_246_3156 ();
 FILLCELL_X32 FILLER_246_3158 ();
 FILLCELL_X32 FILLER_246_3190 ();
 FILLCELL_X32 FILLER_246_3222 ();
 FILLCELL_X32 FILLER_246_3254 ();
 FILLCELL_X32 FILLER_246_3286 ();
 FILLCELL_X32 FILLER_246_3318 ();
 FILLCELL_X32 FILLER_246_3350 ();
 FILLCELL_X32 FILLER_246_3382 ();
 FILLCELL_X32 FILLER_246_3414 ();
 FILLCELL_X32 FILLER_246_3446 ();
 FILLCELL_X32 FILLER_246_3478 ();
 FILLCELL_X32 FILLER_246_3510 ();
 FILLCELL_X32 FILLER_246_3542 ();
 FILLCELL_X32 FILLER_246_3574 ();
 FILLCELL_X32 FILLER_246_3606 ();
 FILLCELL_X32 FILLER_246_3638 ();
 FILLCELL_X32 FILLER_246_3670 ();
 FILLCELL_X32 FILLER_246_3702 ();
 FILLCELL_X4 FILLER_246_3734 ();
 FILLCELL_X8 FILLER_247_1 ();
 FILLCELL_X32 FILLER_247_12 ();
 FILLCELL_X32 FILLER_247_44 ();
 FILLCELL_X32 FILLER_247_76 ();
 FILLCELL_X32 FILLER_247_108 ();
 FILLCELL_X32 FILLER_247_140 ();
 FILLCELL_X32 FILLER_247_172 ();
 FILLCELL_X32 FILLER_247_204 ();
 FILLCELL_X32 FILLER_247_236 ();
 FILLCELL_X32 FILLER_247_268 ();
 FILLCELL_X32 FILLER_247_300 ();
 FILLCELL_X32 FILLER_247_332 ();
 FILLCELL_X32 FILLER_247_364 ();
 FILLCELL_X32 FILLER_247_396 ();
 FILLCELL_X32 FILLER_247_428 ();
 FILLCELL_X32 FILLER_247_460 ();
 FILLCELL_X32 FILLER_247_492 ();
 FILLCELL_X32 FILLER_247_524 ();
 FILLCELL_X32 FILLER_247_556 ();
 FILLCELL_X32 FILLER_247_588 ();
 FILLCELL_X32 FILLER_247_620 ();
 FILLCELL_X32 FILLER_247_652 ();
 FILLCELL_X32 FILLER_247_684 ();
 FILLCELL_X32 FILLER_247_716 ();
 FILLCELL_X32 FILLER_247_748 ();
 FILLCELL_X32 FILLER_247_780 ();
 FILLCELL_X32 FILLER_247_812 ();
 FILLCELL_X32 FILLER_247_844 ();
 FILLCELL_X32 FILLER_247_876 ();
 FILLCELL_X32 FILLER_247_908 ();
 FILLCELL_X32 FILLER_247_940 ();
 FILLCELL_X32 FILLER_247_972 ();
 FILLCELL_X32 FILLER_247_1004 ();
 FILLCELL_X32 FILLER_247_1036 ();
 FILLCELL_X32 FILLER_247_1068 ();
 FILLCELL_X32 FILLER_247_1100 ();
 FILLCELL_X32 FILLER_247_1132 ();
 FILLCELL_X32 FILLER_247_1164 ();
 FILLCELL_X32 FILLER_247_1196 ();
 FILLCELL_X32 FILLER_247_1228 ();
 FILLCELL_X2 FILLER_247_1260 ();
 FILLCELL_X1 FILLER_247_1262 ();
 FILLCELL_X32 FILLER_247_1264 ();
 FILLCELL_X32 FILLER_247_1296 ();
 FILLCELL_X32 FILLER_247_1328 ();
 FILLCELL_X32 FILLER_247_1360 ();
 FILLCELL_X32 FILLER_247_1392 ();
 FILLCELL_X32 FILLER_247_1424 ();
 FILLCELL_X32 FILLER_247_1456 ();
 FILLCELL_X32 FILLER_247_1488 ();
 FILLCELL_X32 FILLER_247_1520 ();
 FILLCELL_X32 FILLER_247_1552 ();
 FILLCELL_X16 FILLER_247_1584 ();
 FILLCELL_X1 FILLER_247_1600 ();
 FILLCELL_X32 FILLER_247_1620 ();
 FILLCELL_X32 FILLER_247_1652 ();
 FILLCELL_X32 FILLER_247_1684 ();
 FILLCELL_X32 FILLER_247_1716 ();
 FILLCELL_X32 FILLER_247_1748 ();
 FILLCELL_X32 FILLER_247_1780 ();
 FILLCELL_X32 FILLER_247_1816 ();
 FILLCELL_X16 FILLER_247_1848 ();
 FILLCELL_X8 FILLER_247_1864 ();
 FILLCELL_X1 FILLER_247_1872 ();
 FILLCELL_X8 FILLER_247_1890 ();
 FILLCELL_X8 FILLER_247_1903 ();
 FILLCELL_X2 FILLER_247_1911 ();
 FILLCELL_X2 FILLER_247_1924 ();
 FILLCELL_X32 FILLER_247_1933 ();
 FILLCELL_X32 FILLER_247_1965 ();
 FILLCELL_X1 FILLER_247_1997 ();
 FILLCELL_X4 FILLER_247_2005 ();
 FILLCELL_X1 FILLER_247_2009 ();
 FILLCELL_X4 FILLER_247_2017 ();
 FILLCELL_X1 FILLER_247_2021 ();
 FILLCELL_X16 FILLER_247_2046 ();
 FILLCELL_X8 FILLER_247_2062 ();
 FILLCELL_X16 FILLER_247_2094 ();
 FILLCELL_X1 FILLER_247_2110 ();
 FILLCELL_X4 FILLER_247_2128 ();
 FILLCELL_X2 FILLER_247_2132 ();
 FILLCELL_X2 FILLER_247_2158 ();
 FILLCELL_X32 FILLER_247_2215 ();
 FILLCELL_X32 FILLER_247_2247 ();
 FILLCELL_X32 FILLER_247_2279 ();
 FILLCELL_X32 FILLER_247_2311 ();
 FILLCELL_X32 FILLER_247_2343 ();
 FILLCELL_X32 FILLER_247_2375 ();
 FILLCELL_X32 FILLER_247_2407 ();
 FILLCELL_X32 FILLER_247_2439 ();
 FILLCELL_X32 FILLER_247_2471 ();
 FILLCELL_X16 FILLER_247_2503 ();
 FILLCELL_X4 FILLER_247_2519 ();
 FILLCELL_X2 FILLER_247_2523 ();
 FILLCELL_X1 FILLER_247_2525 ();
 FILLCELL_X32 FILLER_247_2527 ();
 FILLCELL_X32 FILLER_247_2559 ();
 FILLCELL_X32 FILLER_247_2591 ();
 FILLCELL_X32 FILLER_247_2623 ();
 FILLCELL_X32 FILLER_247_2655 ();
 FILLCELL_X32 FILLER_247_2687 ();
 FILLCELL_X32 FILLER_247_2719 ();
 FILLCELL_X32 FILLER_247_2751 ();
 FILLCELL_X32 FILLER_247_2783 ();
 FILLCELL_X32 FILLER_247_2815 ();
 FILLCELL_X32 FILLER_247_2847 ();
 FILLCELL_X32 FILLER_247_2879 ();
 FILLCELL_X32 FILLER_247_2911 ();
 FILLCELL_X32 FILLER_247_2943 ();
 FILLCELL_X32 FILLER_247_2975 ();
 FILLCELL_X32 FILLER_247_3007 ();
 FILLCELL_X32 FILLER_247_3039 ();
 FILLCELL_X32 FILLER_247_3071 ();
 FILLCELL_X32 FILLER_247_3103 ();
 FILLCELL_X32 FILLER_247_3135 ();
 FILLCELL_X32 FILLER_247_3167 ();
 FILLCELL_X32 FILLER_247_3199 ();
 FILLCELL_X32 FILLER_247_3231 ();
 FILLCELL_X32 FILLER_247_3263 ();
 FILLCELL_X32 FILLER_247_3295 ();
 FILLCELL_X32 FILLER_247_3327 ();
 FILLCELL_X32 FILLER_247_3359 ();
 FILLCELL_X32 FILLER_247_3391 ();
 FILLCELL_X32 FILLER_247_3423 ();
 FILLCELL_X32 FILLER_247_3455 ();
 FILLCELL_X32 FILLER_247_3487 ();
 FILLCELL_X32 FILLER_247_3519 ();
 FILLCELL_X32 FILLER_247_3551 ();
 FILLCELL_X32 FILLER_247_3583 ();
 FILLCELL_X32 FILLER_247_3615 ();
 FILLCELL_X32 FILLER_247_3647 ();
 FILLCELL_X32 FILLER_247_3679 ();
 FILLCELL_X2 FILLER_247_3711 ();
 FILLCELL_X1 FILLER_247_3713 ();
 FILLCELL_X16 FILLER_247_3717 ();
 FILLCELL_X4 FILLER_247_3733 ();
 FILLCELL_X1 FILLER_247_3737 ();
 FILLCELL_X4 FILLER_248_1 ();
 FILLCELL_X32 FILLER_248_8 ();
 FILLCELL_X32 FILLER_248_40 ();
 FILLCELL_X32 FILLER_248_72 ();
 FILLCELL_X32 FILLER_248_104 ();
 FILLCELL_X32 FILLER_248_136 ();
 FILLCELL_X32 FILLER_248_168 ();
 FILLCELL_X32 FILLER_248_200 ();
 FILLCELL_X32 FILLER_248_232 ();
 FILLCELL_X32 FILLER_248_264 ();
 FILLCELL_X32 FILLER_248_296 ();
 FILLCELL_X32 FILLER_248_328 ();
 FILLCELL_X32 FILLER_248_360 ();
 FILLCELL_X32 FILLER_248_392 ();
 FILLCELL_X32 FILLER_248_424 ();
 FILLCELL_X32 FILLER_248_456 ();
 FILLCELL_X32 FILLER_248_488 ();
 FILLCELL_X32 FILLER_248_520 ();
 FILLCELL_X32 FILLER_248_552 ();
 FILLCELL_X32 FILLER_248_584 ();
 FILLCELL_X8 FILLER_248_616 ();
 FILLCELL_X4 FILLER_248_624 ();
 FILLCELL_X2 FILLER_248_628 ();
 FILLCELL_X1 FILLER_248_630 ();
 FILLCELL_X32 FILLER_248_632 ();
 FILLCELL_X32 FILLER_248_664 ();
 FILLCELL_X32 FILLER_248_696 ();
 FILLCELL_X32 FILLER_248_728 ();
 FILLCELL_X32 FILLER_248_760 ();
 FILLCELL_X32 FILLER_248_792 ();
 FILLCELL_X32 FILLER_248_824 ();
 FILLCELL_X32 FILLER_248_856 ();
 FILLCELL_X32 FILLER_248_888 ();
 FILLCELL_X32 FILLER_248_920 ();
 FILLCELL_X32 FILLER_248_952 ();
 FILLCELL_X32 FILLER_248_984 ();
 FILLCELL_X32 FILLER_248_1016 ();
 FILLCELL_X32 FILLER_248_1048 ();
 FILLCELL_X32 FILLER_248_1080 ();
 FILLCELL_X32 FILLER_248_1112 ();
 FILLCELL_X32 FILLER_248_1144 ();
 FILLCELL_X32 FILLER_248_1176 ();
 FILLCELL_X32 FILLER_248_1208 ();
 FILLCELL_X32 FILLER_248_1240 ();
 FILLCELL_X32 FILLER_248_1272 ();
 FILLCELL_X32 FILLER_248_1304 ();
 FILLCELL_X32 FILLER_248_1336 ();
 FILLCELL_X32 FILLER_248_1368 ();
 FILLCELL_X32 FILLER_248_1400 ();
 FILLCELL_X32 FILLER_248_1432 ();
 FILLCELL_X32 FILLER_248_1464 ();
 FILLCELL_X32 FILLER_248_1496 ();
 FILLCELL_X32 FILLER_248_1528 ();
 FILLCELL_X32 FILLER_248_1560 ();
 FILLCELL_X8 FILLER_248_1592 ();
 FILLCELL_X2 FILLER_248_1600 ();
 FILLCELL_X1 FILLER_248_1602 ();
 FILLCELL_X32 FILLER_248_1607 ();
 FILLCELL_X8 FILLER_248_1639 ();
 FILLCELL_X1 FILLER_248_1647 ();
 FILLCELL_X32 FILLER_248_1667 ();
 FILLCELL_X32 FILLER_248_1699 ();
 FILLCELL_X32 FILLER_248_1731 ();
 FILLCELL_X32 FILLER_248_1763 ();
 FILLCELL_X32 FILLER_248_1795 ();
 FILLCELL_X16 FILLER_248_1827 ();
 FILLCELL_X8 FILLER_248_1843 ();
 FILLCELL_X4 FILLER_248_1851 ();
 FILLCELL_X2 FILLER_248_1855 ();
 FILLCELL_X1 FILLER_248_1857 ();
 FILLCELL_X16 FILLER_248_1863 ();
 FILLCELL_X8 FILLER_248_1879 ();
 FILLCELL_X4 FILLER_248_1887 ();
 FILLCELL_X2 FILLER_248_1891 ();
 FILLCELL_X1 FILLER_248_1893 ();
 FILLCELL_X8 FILLER_248_1895 ();
 FILLCELL_X4 FILLER_248_1903 ();
 FILLCELL_X2 FILLER_248_1907 ();
 FILLCELL_X1 FILLER_248_1909 ();
 FILLCELL_X8 FILLER_248_1913 ();
 FILLCELL_X2 FILLER_248_1921 ();
 FILLCELL_X1 FILLER_248_1923 ();
 FILLCELL_X32 FILLER_248_1931 ();
 FILLCELL_X32 FILLER_248_1963 ();
 FILLCELL_X32 FILLER_248_1995 ();
 FILLCELL_X32 FILLER_248_2034 ();
 FILLCELL_X32 FILLER_248_2066 ();
 FILLCELL_X32 FILLER_248_2098 ();
 FILLCELL_X32 FILLER_248_2130 ();
 FILLCELL_X32 FILLER_248_2162 ();
 FILLCELL_X16 FILLER_248_2194 ();
 FILLCELL_X2 FILLER_248_2210 ();
 FILLCELL_X1 FILLER_248_2212 ();
 FILLCELL_X32 FILLER_248_2220 ();
 FILLCELL_X8 FILLER_248_2252 ();
 FILLCELL_X4 FILLER_248_2260 ();
 FILLCELL_X1 FILLER_248_2264 ();
 FILLCELL_X2 FILLER_248_2276 ();
 FILLCELL_X16 FILLER_248_2295 ();
 FILLCELL_X8 FILLER_248_2311 ();
 FILLCELL_X4 FILLER_248_2319 ();
 FILLCELL_X2 FILLER_248_2323 ();
 FILLCELL_X32 FILLER_248_2329 ();
 FILLCELL_X32 FILLER_248_2361 ();
 FILLCELL_X32 FILLER_248_2393 ();
 FILLCELL_X32 FILLER_248_2425 ();
 FILLCELL_X32 FILLER_248_2457 ();
 FILLCELL_X32 FILLER_248_2489 ();
 FILLCELL_X32 FILLER_248_2521 ();
 FILLCELL_X32 FILLER_248_2553 ();
 FILLCELL_X32 FILLER_248_2585 ();
 FILLCELL_X32 FILLER_248_2617 ();
 FILLCELL_X32 FILLER_248_2649 ();
 FILLCELL_X32 FILLER_248_2681 ();
 FILLCELL_X32 FILLER_248_2713 ();
 FILLCELL_X32 FILLER_248_2745 ();
 FILLCELL_X32 FILLER_248_2777 ();
 FILLCELL_X32 FILLER_248_2809 ();
 FILLCELL_X32 FILLER_248_2841 ();
 FILLCELL_X32 FILLER_248_2873 ();
 FILLCELL_X32 FILLER_248_2905 ();
 FILLCELL_X32 FILLER_248_2937 ();
 FILLCELL_X32 FILLER_248_2969 ();
 FILLCELL_X32 FILLER_248_3001 ();
 FILLCELL_X32 FILLER_248_3033 ();
 FILLCELL_X32 FILLER_248_3065 ();
 FILLCELL_X32 FILLER_248_3097 ();
 FILLCELL_X16 FILLER_248_3129 ();
 FILLCELL_X8 FILLER_248_3145 ();
 FILLCELL_X4 FILLER_248_3153 ();
 FILLCELL_X32 FILLER_248_3158 ();
 FILLCELL_X32 FILLER_248_3190 ();
 FILLCELL_X32 FILLER_248_3222 ();
 FILLCELL_X32 FILLER_248_3254 ();
 FILLCELL_X32 FILLER_248_3286 ();
 FILLCELL_X32 FILLER_248_3318 ();
 FILLCELL_X32 FILLER_248_3350 ();
 FILLCELL_X32 FILLER_248_3382 ();
 FILLCELL_X32 FILLER_248_3414 ();
 FILLCELL_X32 FILLER_248_3446 ();
 FILLCELL_X32 FILLER_248_3478 ();
 FILLCELL_X32 FILLER_248_3510 ();
 FILLCELL_X32 FILLER_248_3542 ();
 FILLCELL_X32 FILLER_248_3574 ();
 FILLCELL_X32 FILLER_248_3606 ();
 FILLCELL_X32 FILLER_248_3638 ();
 FILLCELL_X32 FILLER_248_3670 ();
 FILLCELL_X32 FILLER_248_3702 ();
 FILLCELL_X4 FILLER_248_3734 ();
 FILLCELL_X32 FILLER_249_4 ();
 FILLCELL_X32 FILLER_249_36 ();
 FILLCELL_X32 FILLER_249_68 ();
 FILLCELL_X32 FILLER_249_100 ();
 FILLCELL_X32 FILLER_249_132 ();
 FILLCELL_X32 FILLER_249_164 ();
 FILLCELL_X32 FILLER_249_196 ();
 FILLCELL_X32 FILLER_249_228 ();
 FILLCELL_X32 FILLER_249_260 ();
 FILLCELL_X32 FILLER_249_292 ();
 FILLCELL_X32 FILLER_249_324 ();
 FILLCELL_X32 FILLER_249_356 ();
 FILLCELL_X32 FILLER_249_388 ();
 FILLCELL_X32 FILLER_249_420 ();
 FILLCELL_X32 FILLER_249_452 ();
 FILLCELL_X32 FILLER_249_484 ();
 FILLCELL_X32 FILLER_249_516 ();
 FILLCELL_X32 FILLER_249_548 ();
 FILLCELL_X32 FILLER_249_580 ();
 FILLCELL_X32 FILLER_249_612 ();
 FILLCELL_X32 FILLER_249_644 ();
 FILLCELL_X32 FILLER_249_676 ();
 FILLCELL_X32 FILLER_249_708 ();
 FILLCELL_X32 FILLER_249_740 ();
 FILLCELL_X32 FILLER_249_772 ();
 FILLCELL_X32 FILLER_249_804 ();
 FILLCELL_X32 FILLER_249_836 ();
 FILLCELL_X32 FILLER_249_868 ();
 FILLCELL_X32 FILLER_249_900 ();
 FILLCELL_X32 FILLER_249_932 ();
 FILLCELL_X32 FILLER_249_964 ();
 FILLCELL_X32 FILLER_249_996 ();
 FILLCELL_X32 FILLER_249_1028 ();
 FILLCELL_X32 FILLER_249_1060 ();
 FILLCELL_X32 FILLER_249_1092 ();
 FILLCELL_X32 FILLER_249_1124 ();
 FILLCELL_X32 FILLER_249_1156 ();
 FILLCELL_X32 FILLER_249_1188 ();
 FILLCELL_X32 FILLER_249_1220 ();
 FILLCELL_X8 FILLER_249_1252 ();
 FILLCELL_X2 FILLER_249_1260 ();
 FILLCELL_X1 FILLER_249_1262 ();
 FILLCELL_X32 FILLER_249_1264 ();
 FILLCELL_X32 FILLER_249_1296 ();
 FILLCELL_X32 FILLER_249_1328 ();
 FILLCELL_X32 FILLER_249_1360 ();
 FILLCELL_X32 FILLER_249_1392 ();
 FILLCELL_X32 FILLER_249_1424 ();
 FILLCELL_X32 FILLER_249_1456 ();
 FILLCELL_X32 FILLER_249_1488 ();
 FILLCELL_X32 FILLER_249_1520 ();
 FILLCELL_X32 FILLER_249_1552 ();
 FILLCELL_X8 FILLER_249_1584 ();
 FILLCELL_X4 FILLER_249_1592 ();
 FILLCELL_X1 FILLER_249_1596 ();
 FILLCELL_X4 FILLER_249_1615 ();
 FILLCELL_X2 FILLER_249_1619 ();
 FILLCELL_X1 FILLER_249_1621 ();
 FILLCELL_X1 FILLER_249_1626 ();
 FILLCELL_X16 FILLER_249_1632 ();
 FILLCELL_X4 FILLER_249_1648 ();
 FILLCELL_X2 FILLER_249_1652 ();
 FILLCELL_X32 FILLER_249_1667 ();
 FILLCELL_X32 FILLER_249_1699 ();
 FILLCELL_X32 FILLER_249_1731 ();
 FILLCELL_X32 FILLER_249_1763 ();
 FILLCELL_X32 FILLER_249_1795 ();
 FILLCELL_X8 FILLER_249_1827 ();
 FILLCELL_X2 FILLER_249_1835 ();
 FILLCELL_X1 FILLER_249_1837 ();
 FILLCELL_X2 FILLER_249_1841 ();
 FILLCELL_X8 FILLER_249_1847 ();
 FILLCELL_X2 FILLER_249_1855 ();
 FILLCELL_X32 FILLER_249_1862 ();
 FILLCELL_X8 FILLER_249_1894 ();
 FILLCELL_X2 FILLER_249_1902 ();
 FILLCELL_X1 FILLER_249_1904 ();
 FILLCELL_X4 FILLER_249_1912 ();
 FILLCELL_X2 FILLER_249_1916 ();
 FILLCELL_X4 FILLER_249_1925 ();
 FILLCELL_X32 FILLER_249_1953 ();
 FILLCELL_X16 FILLER_249_1985 ();
 FILLCELL_X4 FILLER_249_2001 ();
 FILLCELL_X2 FILLER_249_2005 ();
 FILLCELL_X1 FILLER_249_2007 ();
 FILLCELL_X32 FILLER_249_2015 ();
 FILLCELL_X4 FILLER_249_2047 ();
 FILLCELL_X2 FILLER_249_2051 ();
 FILLCELL_X32 FILLER_249_2060 ();
 FILLCELL_X16 FILLER_249_2092 ();
 FILLCELL_X8 FILLER_249_2115 ();
 FILLCELL_X2 FILLER_249_2123 ();
 FILLCELL_X1 FILLER_249_2125 ();
 FILLCELL_X32 FILLER_249_2133 ();
 FILLCELL_X16 FILLER_249_2165 ();
 FILLCELL_X8 FILLER_249_2181 ();
 FILLCELL_X2 FILLER_249_2189 ();
 FILLCELL_X1 FILLER_249_2191 ();
 FILLCELL_X8 FILLER_249_2200 ();
 FILLCELL_X2 FILLER_249_2232 ();
 FILLCELL_X32 FILLER_249_2241 ();
 FILLCELL_X16 FILLER_249_2273 ();
 FILLCELL_X8 FILLER_249_2289 ();
 FILLCELL_X2 FILLER_249_2297 ();
 FILLCELL_X1 FILLER_249_2299 ();
 FILLCELL_X32 FILLER_249_2324 ();
 FILLCELL_X32 FILLER_249_2356 ();
 FILLCELL_X32 FILLER_249_2388 ();
 FILLCELL_X32 FILLER_249_2420 ();
 FILLCELL_X32 FILLER_249_2452 ();
 FILLCELL_X32 FILLER_249_2484 ();
 FILLCELL_X8 FILLER_249_2516 ();
 FILLCELL_X2 FILLER_249_2524 ();
 FILLCELL_X32 FILLER_249_2527 ();
 FILLCELL_X32 FILLER_249_2559 ();
 FILLCELL_X32 FILLER_249_2591 ();
 FILLCELL_X32 FILLER_249_2623 ();
 FILLCELL_X32 FILLER_249_2655 ();
 FILLCELL_X32 FILLER_249_2687 ();
 FILLCELL_X32 FILLER_249_2719 ();
 FILLCELL_X32 FILLER_249_2751 ();
 FILLCELL_X32 FILLER_249_2783 ();
 FILLCELL_X32 FILLER_249_2815 ();
 FILLCELL_X32 FILLER_249_2847 ();
 FILLCELL_X32 FILLER_249_2879 ();
 FILLCELL_X32 FILLER_249_2911 ();
 FILLCELL_X32 FILLER_249_2943 ();
 FILLCELL_X32 FILLER_249_2975 ();
 FILLCELL_X32 FILLER_249_3007 ();
 FILLCELL_X32 FILLER_249_3039 ();
 FILLCELL_X32 FILLER_249_3071 ();
 FILLCELL_X32 FILLER_249_3103 ();
 FILLCELL_X32 FILLER_249_3135 ();
 FILLCELL_X32 FILLER_249_3167 ();
 FILLCELL_X32 FILLER_249_3199 ();
 FILLCELL_X32 FILLER_249_3231 ();
 FILLCELL_X32 FILLER_249_3263 ();
 FILLCELL_X32 FILLER_249_3295 ();
 FILLCELL_X32 FILLER_249_3327 ();
 FILLCELL_X32 FILLER_249_3359 ();
 FILLCELL_X32 FILLER_249_3391 ();
 FILLCELL_X32 FILLER_249_3423 ();
 FILLCELL_X32 FILLER_249_3455 ();
 FILLCELL_X32 FILLER_249_3487 ();
 FILLCELL_X32 FILLER_249_3519 ();
 FILLCELL_X32 FILLER_249_3551 ();
 FILLCELL_X32 FILLER_249_3583 ();
 FILLCELL_X32 FILLER_249_3615 ();
 FILLCELL_X32 FILLER_249_3647 ();
 FILLCELL_X32 FILLER_249_3679 ();
 FILLCELL_X16 FILLER_249_3711 ();
 FILLCELL_X8 FILLER_249_3727 ();
 FILLCELL_X2 FILLER_249_3735 ();
 FILLCELL_X1 FILLER_249_3737 ();
 FILLCELL_X32 FILLER_250_1 ();
 FILLCELL_X32 FILLER_250_33 ();
 FILLCELL_X32 FILLER_250_65 ();
 FILLCELL_X32 FILLER_250_97 ();
 FILLCELL_X32 FILLER_250_129 ();
 FILLCELL_X32 FILLER_250_161 ();
 FILLCELL_X32 FILLER_250_193 ();
 FILLCELL_X32 FILLER_250_225 ();
 FILLCELL_X32 FILLER_250_257 ();
 FILLCELL_X32 FILLER_250_289 ();
 FILLCELL_X32 FILLER_250_321 ();
 FILLCELL_X32 FILLER_250_353 ();
 FILLCELL_X32 FILLER_250_385 ();
 FILLCELL_X32 FILLER_250_417 ();
 FILLCELL_X32 FILLER_250_449 ();
 FILLCELL_X32 FILLER_250_481 ();
 FILLCELL_X32 FILLER_250_513 ();
 FILLCELL_X32 FILLER_250_545 ();
 FILLCELL_X32 FILLER_250_577 ();
 FILLCELL_X16 FILLER_250_609 ();
 FILLCELL_X4 FILLER_250_625 ();
 FILLCELL_X2 FILLER_250_629 ();
 FILLCELL_X32 FILLER_250_632 ();
 FILLCELL_X32 FILLER_250_664 ();
 FILLCELL_X32 FILLER_250_696 ();
 FILLCELL_X32 FILLER_250_728 ();
 FILLCELL_X32 FILLER_250_760 ();
 FILLCELL_X32 FILLER_250_792 ();
 FILLCELL_X32 FILLER_250_824 ();
 FILLCELL_X32 FILLER_250_856 ();
 FILLCELL_X32 FILLER_250_888 ();
 FILLCELL_X32 FILLER_250_920 ();
 FILLCELL_X32 FILLER_250_952 ();
 FILLCELL_X32 FILLER_250_984 ();
 FILLCELL_X32 FILLER_250_1016 ();
 FILLCELL_X32 FILLER_250_1048 ();
 FILLCELL_X32 FILLER_250_1080 ();
 FILLCELL_X32 FILLER_250_1112 ();
 FILLCELL_X32 FILLER_250_1144 ();
 FILLCELL_X32 FILLER_250_1176 ();
 FILLCELL_X32 FILLER_250_1208 ();
 FILLCELL_X32 FILLER_250_1240 ();
 FILLCELL_X32 FILLER_250_1272 ();
 FILLCELL_X32 FILLER_250_1304 ();
 FILLCELL_X32 FILLER_250_1336 ();
 FILLCELL_X32 FILLER_250_1368 ();
 FILLCELL_X32 FILLER_250_1400 ();
 FILLCELL_X32 FILLER_250_1432 ();
 FILLCELL_X4 FILLER_250_1464 ();
 FILLCELL_X2 FILLER_250_1468 ();
 FILLCELL_X1 FILLER_250_1470 ();
 FILLCELL_X32 FILLER_250_1495 ();
 FILLCELL_X32 FILLER_250_1527 ();
 FILLCELL_X4 FILLER_250_1559 ();
 FILLCELL_X2 FILLER_250_1563 ();
 FILLCELL_X4 FILLER_250_1582 ();
 FILLCELL_X1 FILLER_250_1586 ();
 FILLCELL_X32 FILLER_250_1633 ();
 FILLCELL_X2 FILLER_250_1665 ();
 FILLCELL_X1 FILLER_250_1667 ();
 FILLCELL_X32 FILLER_250_1675 ();
 FILLCELL_X32 FILLER_250_1707 ();
 FILLCELL_X32 FILLER_250_1739 ();
 FILLCELL_X16 FILLER_250_1771 ();
 FILLCELL_X2 FILLER_250_1787 ();
 FILLCELL_X32 FILLER_250_1806 ();
 FILLCELL_X16 FILLER_250_1838 ();
 FILLCELL_X4 FILLER_250_1854 ();
 FILLCELL_X2 FILLER_250_1858 ();
 FILLCELL_X1 FILLER_250_1860 ();
 FILLCELL_X4 FILLER_250_1866 ();
 FILLCELL_X1 FILLER_250_1870 ();
 FILLCELL_X16 FILLER_250_1902 ();
 FILLCELL_X1 FILLER_250_1918 ();
 FILLCELL_X8 FILLER_250_1927 ();
 FILLCELL_X1 FILLER_250_1953 ();
 FILLCELL_X8 FILLER_250_1959 ();
 FILLCELL_X4 FILLER_250_1967 ();
 FILLCELL_X1 FILLER_250_1971 ();
 FILLCELL_X8 FILLER_250_1981 ();
 FILLCELL_X4 FILLER_250_1989 ();
 FILLCELL_X1 FILLER_250_1993 ();
 FILLCELL_X8 FILLER_250_2011 ();
 FILLCELL_X4 FILLER_250_2019 ();
 FILLCELL_X2 FILLER_250_2023 ();
 FILLCELL_X16 FILLER_250_2032 ();
 FILLCELL_X1 FILLER_250_2048 ();
 FILLCELL_X1 FILLER_250_2066 ();
 FILLCELL_X4 FILLER_250_2074 ();
 FILLCELL_X16 FILLER_250_2083 ();
 FILLCELL_X2 FILLER_250_2099 ();
 FILLCELL_X1 FILLER_250_2101 ();
 FILLCELL_X1 FILLER_250_2126 ();
 FILLCELL_X16 FILLER_250_2144 ();
 FILLCELL_X8 FILLER_250_2160 ();
 FILLCELL_X2 FILLER_250_2171 ();
 FILLCELL_X1 FILLER_250_2173 ();
 FILLCELL_X8 FILLER_250_2177 ();
 FILLCELL_X2 FILLER_250_2185 ();
 FILLCELL_X4 FILLER_250_2190 ();
 FILLCELL_X1 FILLER_250_2194 ();
 FILLCELL_X2 FILLER_250_2204 ();
 FILLCELL_X1 FILLER_250_2206 ();
 FILLCELL_X16 FILLER_250_2216 ();
 FILLCELL_X2 FILLER_250_2232 ();
 FILLCELL_X8 FILLER_250_2251 ();
 FILLCELL_X2 FILLER_250_2259 ();
 FILLCELL_X32 FILLER_250_2275 ();
 FILLCELL_X32 FILLER_250_2307 ();
 FILLCELL_X32 FILLER_250_2339 ();
 FILLCELL_X32 FILLER_250_2371 ();
 FILLCELL_X32 FILLER_250_2403 ();
 FILLCELL_X32 FILLER_250_2435 ();
 FILLCELL_X32 FILLER_250_2467 ();
 FILLCELL_X32 FILLER_250_2499 ();
 FILLCELL_X32 FILLER_250_2531 ();
 FILLCELL_X32 FILLER_250_2563 ();
 FILLCELL_X32 FILLER_250_2595 ();
 FILLCELL_X32 FILLER_250_2627 ();
 FILLCELL_X32 FILLER_250_2659 ();
 FILLCELL_X32 FILLER_250_2691 ();
 FILLCELL_X32 FILLER_250_2723 ();
 FILLCELL_X32 FILLER_250_2755 ();
 FILLCELL_X32 FILLER_250_2787 ();
 FILLCELL_X32 FILLER_250_2819 ();
 FILLCELL_X32 FILLER_250_2851 ();
 FILLCELL_X32 FILLER_250_2883 ();
 FILLCELL_X32 FILLER_250_2915 ();
 FILLCELL_X32 FILLER_250_2947 ();
 FILLCELL_X32 FILLER_250_2979 ();
 FILLCELL_X32 FILLER_250_3011 ();
 FILLCELL_X32 FILLER_250_3043 ();
 FILLCELL_X32 FILLER_250_3075 ();
 FILLCELL_X32 FILLER_250_3107 ();
 FILLCELL_X16 FILLER_250_3139 ();
 FILLCELL_X2 FILLER_250_3155 ();
 FILLCELL_X32 FILLER_250_3158 ();
 FILLCELL_X32 FILLER_250_3190 ();
 FILLCELL_X32 FILLER_250_3222 ();
 FILLCELL_X32 FILLER_250_3254 ();
 FILLCELL_X32 FILLER_250_3286 ();
 FILLCELL_X32 FILLER_250_3318 ();
 FILLCELL_X32 FILLER_250_3350 ();
 FILLCELL_X32 FILLER_250_3382 ();
 FILLCELL_X32 FILLER_250_3414 ();
 FILLCELL_X32 FILLER_250_3446 ();
 FILLCELL_X32 FILLER_250_3478 ();
 FILLCELL_X32 FILLER_250_3510 ();
 FILLCELL_X32 FILLER_250_3542 ();
 FILLCELL_X32 FILLER_250_3574 ();
 FILLCELL_X32 FILLER_250_3606 ();
 FILLCELL_X32 FILLER_250_3638 ();
 FILLCELL_X32 FILLER_250_3670 ();
 FILLCELL_X32 FILLER_250_3702 ();
 FILLCELL_X4 FILLER_250_3734 ();
 FILLCELL_X8 FILLER_251_1 ();
 FILLCELL_X4 FILLER_251_9 ();
 FILLCELL_X4 FILLER_251_16 ();
 FILLCELL_X2 FILLER_251_20 ();
 FILLCELL_X32 FILLER_251_25 ();
 FILLCELL_X32 FILLER_251_57 ();
 FILLCELL_X32 FILLER_251_89 ();
 FILLCELL_X32 FILLER_251_121 ();
 FILLCELL_X32 FILLER_251_153 ();
 FILLCELL_X32 FILLER_251_185 ();
 FILLCELL_X32 FILLER_251_217 ();
 FILLCELL_X32 FILLER_251_249 ();
 FILLCELL_X32 FILLER_251_281 ();
 FILLCELL_X32 FILLER_251_313 ();
 FILLCELL_X32 FILLER_251_345 ();
 FILLCELL_X32 FILLER_251_377 ();
 FILLCELL_X32 FILLER_251_409 ();
 FILLCELL_X32 FILLER_251_441 ();
 FILLCELL_X32 FILLER_251_473 ();
 FILLCELL_X32 FILLER_251_505 ();
 FILLCELL_X32 FILLER_251_537 ();
 FILLCELL_X32 FILLER_251_569 ();
 FILLCELL_X32 FILLER_251_601 ();
 FILLCELL_X32 FILLER_251_633 ();
 FILLCELL_X32 FILLER_251_665 ();
 FILLCELL_X32 FILLER_251_697 ();
 FILLCELL_X32 FILLER_251_729 ();
 FILLCELL_X32 FILLER_251_761 ();
 FILLCELL_X32 FILLER_251_793 ();
 FILLCELL_X32 FILLER_251_825 ();
 FILLCELL_X32 FILLER_251_857 ();
 FILLCELL_X32 FILLER_251_889 ();
 FILLCELL_X32 FILLER_251_921 ();
 FILLCELL_X32 FILLER_251_953 ();
 FILLCELL_X32 FILLER_251_985 ();
 FILLCELL_X32 FILLER_251_1017 ();
 FILLCELL_X32 FILLER_251_1049 ();
 FILLCELL_X32 FILLER_251_1081 ();
 FILLCELL_X32 FILLER_251_1113 ();
 FILLCELL_X32 FILLER_251_1145 ();
 FILLCELL_X32 FILLER_251_1177 ();
 FILLCELL_X32 FILLER_251_1209 ();
 FILLCELL_X16 FILLER_251_1241 ();
 FILLCELL_X4 FILLER_251_1257 ();
 FILLCELL_X2 FILLER_251_1261 ();
 FILLCELL_X32 FILLER_251_1264 ();
 FILLCELL_X32 FILLER_251_1296 ();
 FILLCELL_X32 FILLER_251_1328 ();
 FILLCELL_X32 FILLER_251_1360 ();
 FILLCELL_X32 FILLER_251_1392 ();
 FILLCELL_X32 FILLER_251_1424 ();
 FILLCELL_X8 FILLER_251_1456 ();
 FILLCELL_X4 FILLER_251_1464 ();
 FILLCELL_X2 FILLER_251_1468 ();
 FILLCELL_X16 FILLER_251_1487 ();
 FILLCELL_X4 FILLER_251_1503 ();
 FILLCELL_X2 FILLER_251_1507 ();
 FILLCELL_X1 FILLER_251_1509 ();
 FILLCELL_X8 FILLER_251_1534 ();
 FILLCELL_X2 FILLER_251_1542 ();
 FILLCELL_X1 FILLER_251_1551 ();
 FILLCELL_X1 FILLER_251_1569 ();
 FILLCELL_X32 FILLER_251_1577 ();
 FILLCELL_X32 FILLER_251_1609 ();
 FILLCELL_X8 FILLER_251_1641 ();
 FILLCELL_X4 FILLER_251_1649 ();
 FILLCELL_X2 FILLER_251_1653 ();
 FILLCELL_X1 FILLER_251_1655 ();
 FILLCELL_X16 FILLER_251_1680 ();
 FILLCELL_X1 FILLER_251_1696 ();
 FILLCELL_X32 FILLER_251_1725 ();
 FILLCELL_X32 FILLER_251_1757 ();
 FILLCELL_X1 FILLER_251_1789 ();
 FILLCELL_X1 FILLER_251_1800 ();
 FILLCELL_X32 FILLER_251_1805 ();
 FILLCELL_X32 FILLER_251_1837 ();
 FILLCELL_X8 FILLER_251_1869 ();
 FILLCELL_X16 FILLER_251_1882 ();
 FILLCELL_X2 FILLER_251_1898 ();
 FILLCELL_X1 FILLER_251_1900 ();
 FILLCELL_X8 FILLER_251_1904 ();
 FILLCELL_X2 FILLER_251_1912 ();
 FILLCELL_X16 FILLER_251_1918 ();
 FILLCELL_X1 FILLER_251_1934 ();
 FILLCELL_X1 FILLER_251_1962 ();
 FILLCELL_X16 FILLER_251_1986 ();
 FILLCELL_X8 FILLER_251_2002 ();
 FILLCELL_X4 FILLER_251_2010 ();
 FILLCELL_X2 FILLER_251_2014 ();
 FILLCELL_X16 FILLER_251_2040 ();
 FILLCELL_X4 FILLER_251_2056 ();
 FILLCELL_X1 FILLER_251_2060 ();
 FILLCELL_X32 FILLER_251_2090 ();
 FILLCELL_X16 FILLER_251_2122 ();
 FILLCELL_X1 FILLER_251_2138 ();
 FILLCELL_X4 FILLER_251_2161 ();
 FILLCELL_X1 FILLER_251_2165 ();
 FILLCELL_X16 FILLER_251_2180 ();
 FILLCELL_X2 FILLER_251_2196 ();
 FILLCELL_X1 FILLER_251_2205 ();
 FILLCELL_X1 FILLER_251_2216 ();
 FILLCELL_X16 FILLER_251_2244 ();
 FILLCELL_X2 FILLER_251_2260 ();
 FILLCELL_X1 FILLER_251_2262 ();
 FILLCELL_X16 FILLER_251_2280 ();
 FILLCELL_X4 FILLER_251_2296 ();
 FILLCELL_X1 FILLER_251_2300 ();
 FILLCELL_X32 FILLER_251_2308 ();
 FILLCELL_X32 FILLER_251_2340 ();
 FILLCELL_X32 FILLER_251_2372 ();
 FILLCELL_X32 FILLER_251_2404 ();
 FILLCELL_X32 FILLER_251_2436 ();
 FILLCELL_X32 FILLER_251_2468 ();
 FILLCELL_X16 FILLER_251_2500 ();
 FILLCELL_X8 FILLER_251_2516 ();
 FILLCELL_X2 FILLER_251_2524 ();
 FILLCELL_X32 FILLER_251_2527 ();
 FILLCELL_X32 FILLER_251_2559 ();
 FILLCELL_X32 FILLER_251_2591 ();
 FILLCELL_X32 FILLER_251_2623 ();
 FILLCELL_X32 FILLER_251_2655 ();
 FILLCELL_X32 FILLER_251_2687 ();
 FILLCELL_X32 FILLER_251_2719 ();
 FILLCELL_X32 FILLER_251_2751 ();
 FILLCELL_X32 FILLER_251_2783 ();
 FILLCELL_X32 FILLER_251_2815 ();
 FILLCELL_X32 FILLER_251_2847 ();
 FILLCELL_X32 FILLER_251_2879 ();
 FILLCELL_X32 FILLER_251_2911 ();
 FILLCELL_X32 FILLER_251_2943 ();
 FILLCELL_X32 FILLER_251_2975 ();
 FILLCELL_X32 FILLER_251_3007 ();
 FILLCELL_X32 FILLER_251_3039 ();
 FILLCELL_X32 FILLER_251_3071 ();
 FILLCELL_X32 FILLER_251_3103 ();
 FILLCELL_X32 FILLER_251_3135 ();
 FILLCELL_X32 FILLER_251_3167 ();
 FILLCELL_X32 FILLER_251_3199 ();
 FILLCELL_X32 FILLER_251_3231 ();
 FILLCELL_X32 FILLER_251_3263 ();
 FILLCELL_X32 FILLER_251_3295 ();
 FILLCELL_X32 FILLER_251_3327 ();
 FILLCELL_X32 FILLER_251_3359 ();
 FILLCELL_X32 FILLER_251_3391 ();
 FILLCELL_X32 FILLER_251_3423 ();
 FILLCELL_X32 FILLER_251_3455 ();
 FILLCELL_X32 FILLER_251_3487 ();
 FILLCELL_X32 FILLER_251_3519 ();
 FILLCELL_X32 FILLER_251_3551 ();
 FILLCELL_X32 FILLER_251_3583 ();
 FILLCELL_X32 FILLER_251_3615 ();
 FILLCELL_X32 FILLER_251_3647 ();
 FILLCELL_X32 FILLER_251_3679 ();
 FILLCELL_X16 FILLER_251_3711 ();
 FILLCELL_X8 FILLER_251_3727 ();
 FILLCELL_X2 FILLER_251_3735 ();
 FILLCELL_X1 FILLER_251_3737 ();
 FILLCELL_X8 FILLER_252_1 ();
 FILLCELL_X2 FILLER_252_9 ();
 FILLCELL_X32 FILLER_252_14 ();
 FILLCELL_X32 FILLER_252_46 ();
 FILLCELL_X32 FILLER_252_78 ();
 FILLCELL_X32 FILLER_252_110 ();
 FILLCELL_X32 FILLER_252_142 ();
 FILLCELL_X32 FILLER_252_174 ();
 FILLCELL_X32 FILLER_252_206 ();
 FILLCELL_X32 FILLER_252_238 ();
 FILLCELL_X32 FILLER_252_270 ();
 FILLCELL_X32 FILLER_252_302 ();
 FILLCELL_X32 FILLER_252_334 ();
 FILLCELL_X32 FILLER_252_366 ();
 FILLCELL_X32 FILLER_252_398 ();
 FILLCELL_X32 FILLER_252_430 ();
 FILLCELL_X32 FILLER_252_462 ();
 FILLCELL_X32 FILLER_252_494 ();
 FILLCELL_X32 FILLER_252_526 ();
 FILLCELL_X32 FILLER_252_558 ();
 FILLCELL_X32 FILLER_252_590 ();
 FILLCELL_X8 FILLER_252_622 ();
 FILLCELL_X1 FILLER_252_630 ();
 FILLCELL_X32 FILLER_252_632 ();
 FILLCELL_X32 FILLER_252_664 ();
 FILLCELL_X32 FILLER_252_696 ();
 FILLCELL_X32 FILLER_252_728 ();
 FILLCELL_X32 FILLER_252_760 ();
 FILLCELL_X32 FILLER_252_792 ();
 FILLCELL_X32 FILLER_252_824 ();
 FILLCELL_X32 FILLER_252_856 ();
 FILLCELL_X32 FILLER_252_888 ();
 FILLCELL_X32 FILLER_252_920 ();
 FILLCELL_X32 FILLER_252_952 ();
 FILLCELL_X32 FILLER_252_984 ();
 FILLCELL_X32 FILLER_252_1016 ();
 FILLCELL_X32 FILLER_252_1048 ();
 FILLCELL_X32 FILLER_252_1080 ();
 FILLCELL_X32 FILLER_252_1112 ();
 FILLCELL_X32 FILLER_252_1144 ();
 FILLCELL_X32 FILLER_252_1176 ();
 FILLCELL_X32 FILLER_252_1208 ();
 FILLCELL_X32 FILLER_252_1240 ();
 FILLCELL_X32 FILLER_252_1272 ();
 FILLCELL_X32 FILLER_252_1304 ();
 FILLCELL_X32 FILLER_252_1336 ();
 FILLCELL_X32 FILLER_252_1368 ();
 FILLCELL_X32 FILLER_252_1400 ();
 FILLCELL_X32 FILLER_252_1432 ();
 FILLCELL_X4 FILLER_252_1464 ();
 FILLCELL_X2 FILLER_252_1468 ();
 FILLCELL_X8 FILLER_252_1477 ();
 FILLCELL_X2 FILLER_252_1485 ();
 FILLCELL_X1 FILLER_252_1487 ();
 FILLCELL_X8 FILLER_252_1495 ();
 FILLCELL_X4 FILLER_252_1503 ();
 FILLCELL_X2 FILLER_252_1507 ();
 FILLCELL_X1 FILLER_252_1509 ();
 FILLCELL_X32 FILLER_252_1518 ();
 FILLCELL_X8 FILLER_252_1550 ();
 FILLCELL_X4 FILLER_252_1558 ();
 FILLCELL_X2 FILLER_252_1562 ();
 FILLCELL_X8 FILLER_252_1571 ();
 FILLCELL_X4 FILLER_252_1579 ();
 FILLCELL_X2 FILLER_252_1583 ();
 FILLCELL_X1 FILLER_252_1585 ();
 FILLCELL_X8 FILLER_252_1593 ();
 FILLCELL_X8 FILLER_252_1610 ();
 FILLCELL_X2 FILLER_252_1618 ();
 FILLCELL_X1 FILLER_252_1620 ();
 FILLCELL_X4 FILLER_252_1640 ();
 FILLCELL_X2 FILLER_252_1644 ();
 FILLCELL_X1 FILLER_252_1646 ();
 FILLCELL_X1 FILLER_252_1664 ();
 FILLCELL_X32 FILLER_252_1672 ();
 FILLCELL_X2 FILLER_252_1704 ();
 FILLCELL_X1 FILLER_252_1706 ();
 FILLCELL_X16 FILLER_252_1711 ();
 FILLCELL_X4 FILLER_252_1727 ();
 FILLCELL_X2 FILLER_252_1731 ();
 FILLCELL_X16 FILLER_252_1738 ();
 FILLCELL_X1 FILLER_252_1754 ();
 FILLCELL_X32 FILLER_252_1764 ();
 FILLCELL_X8 FILLER_252_1796 ();
 FILLCELL_X4 FILLER_252_1804 ();
 FILLCELL_X2 FILLER_252_1808 ();
 FILLCELL_X1 FILLER_252_1810 ();
 FILLCELL_X1 FILLER_252_1821 ();
 FILLCELL_X32 FILLER_252_1829 ();
 FILLCELL_X32 FILLER_252_1861 ();
 FILLCELL_X1 FILLER_252_1893 ();
 FILLCELL_X16 FILLER_252_1895 ();
 FILLCELL_X8 FILLER_252_1911 ();
 FILLCELL_X1 FILLER_252_1919 ();
 FILLCELL_X8 FILLER_252_1925 ();
 FILLCELL_X4 FILLER_252_1933 ();
 FILLCELL_X2 FILLER_252_1937 ();
 FILLCELL_X1 FILLER_252_1939 ();
 FILLCELL_X8 FILLER_252_1949 ();
 FILLCELL_X2 FILLER_252_1957 ();
 FILLCELL_X32 FILLER_252_1964 ();
 FILLCELL_X32 FILLER_252_1996 ();
 FILLCELL_X32 FILLER_252_2028 ();
 FILLCELL_X8 FILLER_252_2060 ();
 FILLCELL_X8 FILLER_252_2070 ();
 FILLCELL_X4 FILLER_252_2078 ();
 FILLCELL_X4 FILLER_252_2085 ();
 FILLCELL_X1 FILLER_252_2092 ();
 FILLCELL_X8 FILLER_252_2096 ();
 FILLCELL_X2 FILLER_252_2104 ();
 FILLCELL_X8 FILLER_252_2111 ();
 FILLCELL_X4 FILLER_252_2119 ();
 FILLCELL_X2 FILLER_252_2123 ();
 FILLCELL_X4 FILLER_252_2128 ();
 FILLCELL_X2 FILLER_252_2132 ();
 FILLCELL_X4 FILLER_252_2137 ();
 FILLCELL_X2 FILLER_252_2141 ();
 FILLCELL_X1 FILLER_252_2143 ();
 FILLCELL_X16 FILLER_252_2147 ();
 FILLCELL_X8 FILLER_252_2163 ();
 FILLCELL_X4 FILLER_252_2171 ();
 FILLCELL_X2 FILLER_252_2175 ();
 FILLCELL_X1 FILLER_252_2177 ();
 FILLCELL_X16 FILLER_252_2181 ();
 FILLCELL_X4 FILLER_252_2197 ();
 FILLCELL_X2 FILLER_252_2201 ();
 FILLCELL_X4 FILLER_252_2206 ();
 FILLCELL_X2 FILLER_252_2210 ();
 FILLCELL_X8 FILLER_252_2215 ();
 FILLCELL_X32 FILLER_252_2230 ();
 FILLCELL_X32 FILLER_252_2262 ();
 FILLCELL_X32 FILLER_252_2299 ();
 FILLCELL_X32 FILLER_252_2331 ();
 FILLCELL_X32 FILLER_252_2363 ();
 FILLCELL_X32 FILLER_252_2395 ();
 FILLCELL_X32 FILLER_252_2427 ();
 FILLCELL_X32 FILLER_252_2459 ();
 FILLCELL_X32 FILLER_252_2491 ();
 FILLCELL_X32 FILLER_252_2523 ();
 FILLCELL_X32 FILLER_252_2555 ();
 FILLCELL_X32 FILLER_252_2587 ();
 FILLCELL_X32 FILLER_252_2619 ();
 FILLCELL_X32 FILLER_252_2651 ();
 FILLCELL_X32 FILLER_252_2683 ();
 FILLCELL_X32 FILLER_252_2715 ();
 FILLCELL_X32 FILLER_252_2747 ();
 FILLCELL_X32 FILLER_252_2779 ();
 FILLCELL_X32 FILLER_252_2811 ();
 FILLCELL_X32 FILLER_252_2843 ();
 FILLCELL_X32 FILLER_252_2875 ();
 FILLCELL_X32 FILLER_252_2907 ();
 FILLCELL_X32 FILLER_252_2939 ();
 FILLCELL_X32 FILLER_252_2971 ();
 FILLCELL_X32 FILLER_252_3003 ();
 FILLCELL_X32 FILLER_252_3035 ();
 FILLCELL_X32 FILLER_252_3067 ();
 FILLCELL_X32 FILLER_252_3099 ();
 FILLCELL_X16 FILLER_252_3131 ();
 FILLCELL_X8 FILLER_252_3147 ();
 FILLCELL_X2 FILLER_252_3155 ();
 FILLCELL_X32 FILLER_252_3158 ();
 FILLCELL_X32 FILLER_252_3190 ();
 FILLCELL_X32 FILLER_252_3222 ();
 FILLCELL_X32 FILLER_252_3254 ();
 FILLCELL_X32 FILLER_252_3286 ();
 FILLCELL_X32 FILLER_252_3318 ();
 FILLCELL_X32 FILLER_252_3350 ();
 FILLCELL_X32 FILLER_252_3382 ();
 FILLCELL_X32 FILLER_252_3414 ();
 FILLCELL_X32 FILLER_252_3446 ();
 FILLCELL_X32 FILLER_252_3478 ();
 FILLCELL_X32 FILLER_252_3510 ();
 FILLCELL_X32 FILLER_252_3542 ();
 FILLCELL_X32 FILLER_252_3574 ();
 FILLCELL_X32 FILLER_252_3606 ();
 FILLCELL_X32 FILLER_252_3638 ();
 FILLCELL_X32 FILLER_252_3670 ();
 FILLCELL_X32 FILLER_252_3702 ();
 FILLCELL_X4 FILLER_252_3734 ();
 FILLCELL_X32 FILLER_253_1 ();
 FILLCELL_X32 FILLER_253_33 ();
 FILLCELL_X32 FILLER_253_65 ();
 FILLCELL_X32 FILLER_253_97 ();
 FILLCELL_X32 FILLER_253_129 ();
 FILLCELL_X32 FILLER_253_161 ();
 FILLCELL_X32 FILLER_253_193 ();
 FILLCELL_X32 FILLER_253_225 ();
 FILLCELL_X32 FILLER_253_257 ();
 FILLCELL_X32 FILLER_253_289 ();
 FILLCELL_X32 FILLER_253_321 ();
 FILLCELL_X32 FILLER_253_353 ();
 FILLCELL_X32 FILLER_253_385 ();
 FILLCELL_X32 FILLER_253_417 ();
 FILLCELL_X32 FILLER_253_449 ();
 FILLCELL_X32 FILLER_253_481 ();
 FILLCELL_X32 FILLER_253_513 ();
 FILLCELL_X32 FILLER_253_545 ();
 FILLCELL_X32 FILLER_253_577 ();
 FILLCELL_X32 FILLER_253_609 ();
 FILLCELL_X32 FILLER_253_641 ();
 FILLCELL_X32 FILLER_253_673 ();
 FILLCELL_X32 FILLER_253_705 ();
 FILLCELL_X32 FILLER_253_737 ();
 FILLCELL_X32 FILLER_253_769 ();
 FILLCELL_X32 FILLER_253_801 ();
 FILLCELL_X32 FILLER_253_833 ();
 FILLCELL_X32 FILLER_253_865 ();
 FILLCELL_X32 FILLER_253_897 ();
 FILLCELL_X32 FILLER_253_929 ();
 FILLCELL_X32 FILLER_253_961 ();
 FILLCELL_X32 FILLER_253_993 ();
 FILLCELL_X32 FILLER_253_1025 ();
 FILLCELL_X32 FILLER_253_1057 ();
 FILLCELL_X32 FILLER_253_1089 ();
 FILLCELL_X32 FILLER_253_1121 ();
 FILLCELL_X32 FILLER_253_1153 ();
 FILLCELL_X32 FILLER_253_1185 ();
 FILLCELL_X32 FILLER_253_1217 ();
 FILLCELL_X8 FILLER_253_1249 ();
 FILLCELL_X4 FILLER_253_1257 ();
 FILLCELL_X2 FILLER_253_1261 ();
 FILLCELL_X32 FILLER_253_1264 ();
 FILLCELL_X32 FILLER_253_1296 ();
 FILLCELL_X32 FILLER_253_1328 ();
 FILLCELL_X32 FILLER_253_1360 ();
 FILLCELL_X32 FILLER_253_1392 ();
 FILLCELL_X32 FILLER_253_1424 ();
 FILLCELL_X4 FILLER_253_1463 ();
 FILLCELL_X4 FILLER_253_1474 ();
 FILLCELL_X2 FILLER_253_1478 ();
 FILLCELL_X1 FILLER_253_1480 ();
 FILLCELL_X32 FILLER_253_1505 ();
 FILLCELL_X16 FILLER_253_1537 ();
 FILLCELL_X4 FILLER_253_1553 ();
 FILLCELL_X2 FILLER_253_1557 ();
 FILLCELL_X8 FILLER_253_1566 ();
 FILLCELL_X2 FILLER_253_1574 ();
 FILLCELL_X1 FILLER_253_1576 ();
 FILLCELL_X4 FILLER_253_1613 ();
 FILLCELL_X2 FILLER_253_1617 ();
 FILLCELL_X2 FILLER_253_1623 ();
 FILLCELL_X1 FILLER_253_1625 ();
 FILLCELL_X16 FILLER_253_1631 ();
 FILLCELL_X8 FILLER_253_1647 ();
 FILLCELL_X2 FILLER_253_1655 ();
 FILLCELL_X1 FILLER_253_1657 ();
 FILLCELL_X8 FILLER_253_1666 ();
 FILLCELL_X1 FILLER_253_1674 ();
 FILLCELL_X32 FILLER_253_1699 ();
 FILLCELL_X32 FILLER_253_1731 ();
 FILLCELL_X16 FILLER_253_1763 ();
 FILLCELL_X8 FILLER_253_1779 ();
 FILLCELL_X1 FILLER_253_1787 ();
 FILLCELL_X4 FILLER_253_1799 ();
 FILLCELL_X32 FILLER_253_1827 ();
 FILLCELL_X32 FILLER_253_1859 ();
 FILLCELL_X8 FILLER_253_1891 ();
 FILLCELL_X2 FILLER_253_1899 ();
 FILLCELL_X32 FILLER_253_1933 ();
 FILLCELL_X16 FILLER_253_1965 ();
 FILLCELL_X8 FILLER_253_1981 ();
 FILLCELL_X4 FILLER_253_1989 ();
 FILLCELL_X8 FILLER_253_2012 ();
 FILLCELL_X1 FILLER_253_2020 ();
 FILLCELL_X16 FILLER_253_2024 ();
 FILLCELL_X8 FILLER_253_2040 ();
 FILLCELL_X4 FILLER_253_2048 ();
 FILLCELL_X2 FILLER_253_2052 ();
 FILLCELL_X1 FILLER_253_2054 ();
 FILLCELL_X2 FILLER_253_2058 ();
 FILLCELL_X1 FILLER_253_2060 ();
 FILLCELL_X32 FILLER_253_2066 ();
 FILLCELL_X1 FILLER_253_2098 ();
 FILLCELL_X16 FILLER_253_2102 ();
 FILLCELL_X8 FILLER_253_2118 ();
 FILLCELL_X2 FILLER_253_2126 ();
 FILLCELL_X32 FILLER_253_2131 ();
 FILLCELL_X1 FILLER_253_2163 ();
 FILLCELL_X16 FILLER_253_2167 ();
 FILLCELL_X8 FILLER_253_2200 ();
 FILLCELL_X4 FILLER_253_2208 ();
 FILLCELL_X2 FILLER_253_2212 ();
 FILLCELL_X32 FILLER_253_2217 ();
 FILLCELL_X16 FILLER_253_2249 ();
 FILLCELL_X8 FILLER_253_2265 ();
 FILLCELL_X2 FILLER_253_2273 ();
 FILLCELL_X4 FILLER_253_2306 ();
 FILLCELL_X2 FILLER_253_2310 ();
 FILLCELL_X32 FILLER_253_2336 ();
 FILLCELL_X32 FILLER_253_2368 ();
 FILLCELL_X32 FILLER_253_2400 ();
 FILLCELL_X32 FILLER_253_2432 ();
 FILLCELL_X32 FILLER_253_2464 ();
 FILLCELL_X16 FILLER_253_2496 ();
 FILLCELL_X8 FILLER_253_2512 ();
 FILLCELL_X4 FILLER_253_2520 ();
 FILLCELL_X2 FILLER_253_2524 ();
 FILLCELL_X32 FILLER_253_2527 ();
 FILLCELL_X32 FILLER_253_2559 ();
 FILLCELL_X32 FILLER_253_2591 ();
 FILLCELL_X32 FILLER_253_2623 ();
 FILLCELL_X32 FILLER_253_2655 ();
 FILLCELL_X32 FILLER_253_2687 ();
 FILLCELL_X32 FILLER_253_2719 ();
 FILLCELL_X32 FILLER_253_2751 ();
 FILLCELL_X32 FILLER_253_2783 ();
 FILLCELL_X32 FILLER_253_2815 ();
 FILLCELL_X32 FILLER_253_2847 ();
 FILLCELL_X32 FILLER_253_2879 ();
 FILLCELL_X32 FILLER_253_2911 ();
 FILLCELL_X32 FILLER_253_2943 ();
 FILLCELL_X32 FILLER_253_2975 ();
 FILLCELL_X32 FILLER_253_3007 ();
 FILLCELL_X32 FILLER_253_3039 ();
 FILLCELL_X32 FILLER_253_3071 ();
 FILLCELL_X32 FILLER_253_3103 ();
 FILLCELL_X32 FILLER_253_3135 ();
 FILLCELL_X32 FILLER_253_3167 ();
 FILLCELL_X32 FILLER_253_3199 ();
 FILLCELL_X32 FILLER_253_3231 ();
 FILLCELL_X32 FILLER_253_3263 ();
 FILLCELL_X32 FILLER_253_3295 ();
 FILLCELL_X32 FILLER_253_3327 ();
 FILLCELL_X32 FILLER_253_3359 ();
 FILLCELL_X32 FILLER_253_3391 ();
 FILLCELL_X32 FILLER_253_3423 ();
 FILLCELL_X32 FILLER_253_3455 ();
 FILLCELL_X32 FILLER_253_3487 ();
 FILLCELL_X32 FILLER_253_3519 ();
 FILLCELL_X32 FILLER_253_3551 ();
 FILLCELL_X32 FILLER_253_3583 ();
 FILLCELL_X32 FILLER_253_3615 ();
 FILLCELL_X32 FILLER_253_3647 ();
 FILLCELL_X32 FILLER_253_3679 ();
 FILLCELL_X16 FILLER_253_3711 ();
 FILLCELL_X8 FILLER_253_3727 ();
 FILLCELL_X2 FILLER_253_3735 ();
 FILLCELL_X1 FILLER_253_3737 ();
 FILLCELL_X32 FILLER_254_1 ();
 FILLCELL_X32 FILLER_254_33 ();
 FILLCELL_X32 FILLER_254_65 ();
 FILLCELL_X32 FILLER_254_97 ();
 FILLCELL_X32 FILLER_254_129 ();
 FILLCELL_X32 FILLER_254_161 ();
 FILLCELL_X32 FILLER_254_193 ();
 FILLCELL_X32 FILLER_254_225 ();
 FILLCELL_X32 FILLER_254_257 ();
 FILLCELL_X32 FILLER_254_289 ();
 FILLCELL_X32 FILLER_254_321 ();
 FILLCELL_X32 FILLER_254_353 ();
 FILLCELL_X32 FILLER_254_385 ();
 FILLCELL_X32 FILLER_254_417 ();
 FILLCELL_X32 FILLER_254_449 ();
 FILLCELL_X32 FILLER_254_481 ();
 FILLCELL_X32 FILLER_254_513 ();
 FILLCELL_X32 FILLER_254_545 ();
 FILLCELL_X32 FILLER_254_577 ();
 FILLCELL_X16 FILLER_254_609 ();
 FILLCELL_X4 FILLER_254_625 ();
 FILLCELL_X2 FILLER_254_629 ();
 FILLCELL_X32 FILLER_254_632 ();
 FILLCELL_X32 FILLER_254_664 ();
 FILLCELL_X32 FILLER_254_696 ();
 FILLCELL_X32 FILLER_254_728 ();
 FILLCELL_X32 FILLER_254_760 ();
 FILLCELL_X32 FILLER_254_792 ();
 FILLCELL_X32 FILLER_254_824 ();
 FILLCELL_X32 FILLER_254_856 ();
 FILLCELL_X32 FILLER_254_888 ();
 FILLCELL_X32 FILLER_254_920 ();
 FILLCELL_X32 FILLER_254_952 ();
 FILLCELL_X32 FILLER_254_984 ();
 FILLCELL_X32 FILLER_254_1016 ();
 FILLCELL_X32 FILLER_254_1048 ();
 FILLCELL_X32 FILLER_254_1080 ();
 FILLCELL_X32 FILLER_254_1112 ();
 FILLCELL_X32 FILLER_254_1144 ();
 FILLCELL_X32 FILLER_254_1176 ();
 FILLCELL_X32 FILLER_254_1208 ();
 FILLCELL_X32 FILLER_254_1240 ();
 FILLCELL_X32 FILLER_254_1272 ();
 FILLCELL_X32 FILLER_254_1304 ();
 FILLCELL_X32 FILLER_254_1336 ();
 FILLCELL_X32 FILLER_254_1368 ();
 FILLCELL_X32 FILLER_254_1400 ();
 FILLCELL_X16 FILLER_254_1432 ();
 FILLCELL_X8 FILLER_254_1448 ();
 FILLCELL_X32 FILLER_254_1473 ();
 FILLCELL_X8 FILLER_254_1505 ();
 FILLCELL_X4 FILLER_254_1513 ();
 FILLCELL_X1 FILLER_254_1517 ();
 FILLCELL_X16 FILLER_254_1525 ();
 FILLCELL_X8 FILLER_254_1541 ();
 FILLCELL_X32 FILLER_254_1566 ();
 FILLCELL_X16 FILLER_254_1602 ();
 FILLCELL_X2 FILLER_254_1618 ();
 FILLCELL_X1 FILLER_254_1620 ();
 FILLCELL_X32 FILLER_254_1625 ();
 FILLCELL_X4 FILLER_254_1657 ();
 FILLCELL_X2 FILLER_254_1661 ();
 FILLCELL_X2 FILLER_254_1670 ();
 FILLCELL_X32 FILLER_254_1679 ();
 FILLCELL_X32 FILLER_254_1711 ();
 FILLCELL_X2 FILLER_254_1743 ();
 FILLCELL_X1 FILLER_254_1745 ();
 FILLCELL_X4 FILLER_254_1755 ();
 FILLCELL_X8 FILLER_254_1778 ();
 FILLCELL_X2 FILLER_254_1786 ();
 FILLCELL_X32 FILLER_254_1807 ();
 FILLCELL_X32 FILLER_254_1839 ();
 FILLCELL_X16 FILLER_254_1871 ();
 FILLCELL_X4 FILLER_254_1887 ();
 FILLCELL_X2 FILLER_254_1891 ();
 FILLCELL_X1 FILLER_254_1893 ();
 FILLCELL_X16 FILLER_254_1895 ();
 FILLCELL_X8 FILLER_254_1911 ();
 FILLCELL_X8 FILLER_254_1927 ();
 FILLCELL_X1 FILLER_254_1935 ();
 FILLCELL_X8 FILLER_254_1941 ();
 FILLCELL_X16 FILLER_254_1990 ();
 FILLCELL_X8 FILLER_254_2006 ();
 FILLCELL_X1 FILLER_254_2014 ();
 FILLCELL_X4 FILLER_254_2022 ();
 FILLCELL_X16 FILLER_254_2029 ();
 FILLCELL_X4 FILLER_254_2045 ();
 FILLCELL_X2 FILLER_254_2049 ();
 FILLCELL_X1 FILLER_254_2051 ();
 FILLCELL_X1 FILLER_254_2059 ();
 FILLCELL_X1 FILLER_254_2071 ();
 FILLCELL_X2 FILLER_254_2082 ();
 FILLCELL_X8 FILLER_254_2087 ();
 FILLCELL_X1 FILLER_254_2095 ();
 FILLCELL_X16 FILLER_254_2106 ();
 FILLCELL_X2 FILLER_254_2122 ();
 FILLCELL_X1 FILLER_254_2124 ();
 FILLCELL_X8 FILLER_254_2132 ();
 FILLCELL_X2 FILLER_254_2147 ();
 FILLCELL_X2 FILLER_254_2170 ();
 FILLCELL_X1 FILLER_254_2172 ();
 FILLCELL_X2 FILLER_254_2176 ();
 FILLCELL_X1 FILLER_254_2178 ();
 FILLCELL_X1 FILLER_254_2182 ();
 FILLCELL_X1 FILLER_254_2197 ();
 FILLCELL_X16 FILLER_254_2205 ();
 FILLCELL_X4 FILLER_254_2221 ();
 FILLCELL_X1 FILLER_254_2225 ();
 FILLCELL_X32 FILLER_254_2233 ();
 FILLCELL_X2 FILLER_254_2265 ();
 FILLCELL_X16 FILLER_254_2278 ();
 FILLCELL_X32 FILLER_254_2297 ();
 FILLCELL_X32 FILLER_254_2329 ();
 FILLCELL_X32 FILLER_254_2361 ();
 FILLCELL_X32 FILLER_254_2393 ();
 FILLCELL_X32 FILLER_254_2425 ();
 FILLCELL_X32 FILLER_254_2457 ();
 FILLCELL_X32 FILLER_254_2489 ();
 FILLCELL_X32 FILLER_254_2521 ();
 FILLCELL_X32 FILLER_254_2553 ();
 FILLCELL_X32 FILLER_254_2585 ();
 FILLCELL_X32 FILLER_254_2617 ();
 FILLCELL_X32 FILLER_254_2649 ();
 FILLCELL_X32 FILLER_254_2681 ();
 FILLCELL_X32 FILLER_254_2713 ();
 FILLCELL_X32 FILLER_254_2745 ();
 FILLCELL_X32 FILLER_254_2777 ();
 FILLCELL_X32 FILLER_254_2809 ();
 FILLCELL_X32 FILLER_254_2841 ();
 FILLCELL_X32 FILLER_254_2873 ();
 FILLCELL_X32 FILLER_254_2905 ();
 FILLCELL_X32 FILLER_254_2937 ();
 FILLCELL_X32 FILLER_254_2969 ();
 FILLCELL_X32 FILLER_254_3001 ();
 FILLCELL_X32 FILLER_254_3033 ();
 FILLCELL_X32 FILLER_254_3065 ();
 FILLCELL_X32 FILLER_254_3097 ();
 FILLCELL_X16 FILLER_254_3129 ();
 FILLCELL_X8 FILLER_254_3145 ();
 FILLCELL_X4 FILLER_254_3153 ();
 FILLCELL_X32 FILLER_254_3158 ();
 FILLCELL_X32 FILLER_254_3190 ();
 FILLCELL_X32 FILLER_254_3222 ();
 FILLCELL_X32 FILLER_254_3254 ();
 FILLCELL_X32 FILLER_254_3286 ();
 FILLCELL_X32 FILLER_254_3318 ();
 FILLCELL_X32 FILLER_254_3350 ();
 FILLCELL_X32 FILLER_254_3382 ();
 FILLCELL_X32 FILLER_254_3414 ();
 FILLCELL_X32 FILLER_254_3446 ();
 FILLCELL_X32 FILLER_254_3478 ();
 FILLCELL_X32 FILLER_254_3510 ();
 FILLCELL_X32 FILLER_254_3542 ();
 FILLCELL_X32 FILLER_254_3574 ();
 FILLCELL_X32 FILLER_254_3606 ();
 FILLCELL_X32 FILLER_254_3638 ();
 FILLCELL_X32 FILLER_254_3670 ();
 FILLCELL_X2 FILLER_254_3702 ();
 FILLCELL_X1 FILLER_254_3704 ();
 FILLCELL_X16 FILLER_254_3708 ();
 FILLCELL_X4 FILLER_254_3724 ();
 FILLCELL_X2 FILLER_254_3728 ();
 FILLCELL_X1 FILLER_254_3730 ();
 FILLCELL_X1 FILLER_254_3734 ();
 FILLCELL_X32 FILLER_255_1 ();
 FILLCELL_X32 FILLER_255_33 ();
 FILLCELL_X32 FILLER_255_65 ();
 FILLCELL_X32 FILLER_255_97 ();
 FILLCELL_X32 FILLER_255_129 ();
 FILLCELL_X32 FILLER_255_161 ();
 FILLCELL_X32 FILLER_255_193 ();
 FILLCELL_X32 FILLER_255_225 ();
 FILLCELL_X32 FILLER_255_257 ();
 FILLCELL_X32 FILLER_255_289 ();
 FILLCELL_X32 FILLER_255_321 ();
 FILLCELL_X32 FILLER_255_353 ();
 FILLCELL_X32 FILLER_255_385 ();
 FILLCELL_X32 FILLER_255_417 ();
 FILLCELL_X32 FILLER_255_449 ();
 FILLCELL_X32 FILLER_255_481 ();
 FILLCELL_X32 FILLER_255_513 ();
 FILLCELL_X32 FILLER_255_545 ();
 FILLCELL_X32 FILLER_255_577 ();
 FILLCELL_X32 FILLER_255_609 ();
 FILLCELL_X32 FILLER_255_641 ();
 FILLCELL_X32 FILLER_255_673 ();
 FILLCELL_X32 FILLER_255_705 ();
 FILLCELL_X32 FILLER_255_737 ();
 FILLCELL_X32 FILLER_255_769 ();
 FILLCELL_X32 FILLER_255_801 ();
 FILLCELL_X32 FILLER_255_833 ();
 FILLCELL_X32 FILLER_255_865 ();
 FILLCELL_X32 FILLER_255_897 ();
 FILLCELL_X32 FILLER_255_929 ();
 FILLCELL_X32 FILLER_255_961 ();
 FILLCELL_X32 FILLER_255_993 ();
 FILLCELL_X32 FILLER_255_1025 ();
 FILLCELL_X32 FILLER_255_1057 ();
 FILLCELL_X32 FILLER_255_1089 ();
 FILLCELL_X32 FILLER_255_1121 ();
 FILLCELL_X32 FILLER_255_1153 ();
 FILLCELL_X32 FILLER_255_1185 ();
 FILLCELL_X32 FILLER_255_1217 ();
 FILLCELL_X8 FILLER_255_1249 ();
 FILLCELL_X4 FILLER_255_1257 ();
 FILLCELL_X2 FILLER_255_1261 ();
 FILLCELL_X32 FILLER_255_1264 ();
 FILLCELL_X32 FILLER_255_1296 ();
 FILLCELL_X32 FILLER_255_1328 ();
 FILLCELL_X32 FILLER_255_1360 ();
 FILLCELL_X32 FILLER_255_1392 ();
 FILLCELL_X32 FILLER_255_1424 ();
 FILLCELL_X32 FILLER_255_1456 ();
 FILLCELL_X8 FILLER_255_1488 ();
 FILLCELL_X4 FILLER_255_1496 ();
 FILLCELL_X2 FILLER_255_1500 ();
 FILLCELL_X16 FILLER_255_1526 ();
 FILLCELL_X8 FILLER_255_1542 ();
 FILLCELL_X16 FILLER_255_1557 ();
 FILLCELL_X4 FILLER_255_1573 ();
 FILLCELL_X1 FILLER_255_1577 ();
 FILLCELL_X16 FILLER_255_1585 ();
 FILLCELL_X8 FILLER_255_1601 ();
 FILLCELL_X4 FILLER_255_1609 ();
 FILLCELL_X8 FILLER_255_1620 ();
 FILLCELL_X4 FILLER_255_1628 ();
 FILLCELL_X16 FILLER_255_1639 ();
 FILLCELL_X8 FILLER_255_1655 ();
 FILLCELL_X4 FILLER_255_1680 ();
 FILLCELL_X2 FILLER_255_1684 ();
 FILLCELL_X1 FILLER_255_1686 ();
 FILLCELL_X8 FILLER_255_1711 ();
 FILLCELL_X4 FILLER_255_1719 ();
 FILLCELL_X1 FILLER_255_1723 ();
 FILLCELL_X1 FILLER_255_1731 ();
 FILLCELL_X32 FILLER_255_1753 ();
 FILLCELL_X8 FILLER_255_1785 ();
 FILLCELL_X8 FILLER_255_1804 ();
 FILLCELL_X4 FILLER_255_1812 ();
 FILLCELL_X2 FILLER_255_1816 ();
 FILLCELL_X32 FILLER_255_1822 ();
 FILLCELL_X32 FILLER_255_1854 ();
 FILLCELL_X8 FILLER_255_1886 ();
 FILLCELL_X4 FILLER_255_1894 ();
 FILLCELL_X1 FILLER_255_1898 ();
 FILLCELL_X4 FILLER_255_1926 ();
 FILLCELL_X1 FILLER_255_1930 ();
 FILLCELL_X2 FILLER_255_1935 ();
 FILLCELL_X1 FILLER_255_1937 ();
 FILLCELL_X8 FILLER_255_1942 ();
 FILLCELL_X4 FILLER_255_1950 ();
 FILLCELL_X2 FILLER_255_1954 ();
 FILLCELL_X16 FILLER_255_1960 ();
 FILLCELL_X1 FILLER_255_1976 ();
 FILLCELL_X16 FILLER_255_1990 ();
 FILLCELL_X8 FILLER_255_2006 ();
 FILLCELL_X1 FILLER_255_2020 ();
 FILLCELL_X16 FILLER_255_2024 ();
 FILLCELL_X2 FILLER_255_2040 ();
 FILLCELL_X1 FILLER_255_2042 ();
 FILLCELL_X16 FILLER_255_2060 ();
 FILLCELL_X1 FILLER_255_2076 ();
 FILLCELL_X8 FILLER_255_2088 ();
 FILLCELL_X2 FILLER_255_2096 ();
 FILLCELL_X2 FILLER_255_2101 ();
 FILLCELL_X8 FILLER_255_2106 ();
 FILLCELL_X4 FILLER_255_2114 ();
 FILLCELL_X1 FILLER_255_2132 ();
 FILLCELL_X16 FILLER_255_2144 ();
 FILLCELL_X8 FILLER_255_2160 ();
 FILLCELL_X4 FILLER_255_2171 ();
 FILLCELL_X1 FILLER_255_2175 ();
 FILLCELL_X8 FILLER_255_2182 ();
 FILLCELL_X4 FILLER_255_2190 ();
 FILLCELL_X2 FILLER_255_2194 ();
 FILLCELL_X1 FILLER_255_2196 ();
 FILLCELL_X32 FILLER_255_2231 ();
 FILLCELL_X2 FILLER_255_2280 ();
 FILLCELL_X1 FILLER_255_2282 ();
 FILLCELL_X32 FILLER_255_2311 ();
 FILLCELL_X32 FILLER_255_2343 ();
 FILLCELL_X32 FILLER_255_2375 ();
 FILLCELL_X32 FILLER_255_2407 ();
 FILLCELL_X32 FILLER_255_2439 ();
 FILLCELL_X32 FILLER_255_2471 ();
 FILLCELL_X16 FILLER_255_2503 ();
 FILLCELL_X4 FILLER_255_2519 ();
 FILLCELL_X2 FILLER_255_2523 ();
 FILLCELL_X1 FILLER_255_2525 ();
 FILLCELL_X32 FILLER_255_2527 ();
 FILLCELL_X32 FILLER_255_2559 ();
 FILLCELL_X32 FILLER_255_2591 ();
 FILLCELL_X32 FILLER_255_2623 ();
 FILLCELL_X32 FILLER_255_2655 ();
 FILLCELL_X32 FILLER_255_2687 ();
 FILLCELL_X32 FILLER_255_2719 ();
 FILLCELL_X32 FILLER_255_2751 ();
 FILLCELL_X32 FILLER_255_2783 ();
 FILLCELL_X32 FILLER_255_2815 ();
 FILLCELL_X32 FILLER_255_2847 ();
 FILLCELL_X32 FILLER_255_2879 ();
 FILLCELL_X32 FILLER_255_2911 ();
 FILLCELL_X32 FILLER_255_2943 ();
 FILLCELL_X32 FILLER_255_2975 ();
 FILLCELL_X32 FILLER_255_3007 ();
 FILLCELL_X32 FILLER_255_3039 ();
 FILLCELL_X32 FILLER_255_3071 ();
 FILLCELL_X32 FILLER_255_3103 ();
 FILLCELL_X32 FILLER_255_3135 ();
 FILLCELL_X32 FILLER_255_3167 ();
 FILLCELL_X32 FILLER_255_3199 ();
 FILLCELL_X32 FILLER_255_3231 ();
 FILLCELL_X32 FILLER_255_3263 ();
 FILLCELL_X32 FILLER_255_3295 ();
 FILLCELL_X32 FILLER_255_3327 ();
 FILLCELL_X32 FILLER_255_3359 ();
 FILLCELL_X32 FILLER_255_3391 ();
 FILLCELL_X32 FILLER_255_3423 ();
 FILLCELL_X32 FILLER_255_3455 ();
 FILLCELL_X32 FILLER_255_3487 ();
 FILLCELL_X32 FILLER_255_3519 ();
 FILLCELL_X32 FILLER_255_3551 ();
 FILLCELL_X32 FILLER_255_3583 ();
 FILLCELL_X32 FILLER_255_3615 ();
 FILLCELL_X32 FILLER_255_3647 ();
 FILLCELL_X32 FILLER_255_3679 ();
 FILLCELL_X4 FILLER_255_3711 ();
 FILLCELL_X2 FILLER_255_3715 ();
 FILLCELL_X1 FILLER_255_3717 ();
 FILLCELL_X16 FILLER_255_3721 ();
 FILLCELL_X1 FILLER_255_3737 ();
 FILLCELL_X32 FILLER_256_1 ();
 FILLCELL_X32 FILLER_256_33 ();
 FILLCELL_X32 FILLER_256_65 ();
 FILLCELL_X32 FILLER_256_97 ();
 FILLCELL_X32 FILLER_256_129 ();
 FILLCELL_X32 FILLER_256_161 ();
 FILLCELL_X32 FILLER_256_193 ();
 FILLCELL_X32 FILLER_256_225 ();
 FILLCELL_X32 FILLER_256_257 ();
 FILLCELL_X32 FILLER_256_289 ();
 FILLCELL_X32 FILLER_256_321 ();
 FILLCELL_X32 FILLER_256_353 ();
 FILLCELL_X32 FILLER_256_385 ();
 FILLCELL_X32 FILLER_256_417 ();
 FILLCELL_X32 FILLER_256_449 ();
 FILLCELL_X32 FILLER_256_481 ();
 FILLCELL_X32 FILLER_256_513 ();
 FILLCELL_X32 FILLER_256_545 ();
 FILLCELL_X32 FILLER_256_577 ();
 FILLCELL_X16 FILLER_256_609 ();
 FILLCELL_X4 FILLER_256_625 ();
 FILLCELL_X2 FILLER_256_629 ();
 FILLCELL_X32 FILLER_256_632 ();
 FILLCELL_X32 FILLER_256_664 ();
 FILLCELL_X32 FILLER_256_696 ();
 FILLCELL_X32 FILLER_256_728 ();
 FILLCELL_X32 FILLER_256_760 ();
 FILLCELL_X32 FILLER_256_792 ();
 FILLCELL_X32 FILLER_256_824 ();
 FILLCELL_X32 FILLER_256_856 ();
 FILLCELL_X32 FILLER_256_888 ();
 FILLCELL_X32 FILLER_256_920 ();
 FILLCELL_X32 FILLER_256_952 ();
 FILLCELL_X32 FILLER_256_984 ();
 FILLCELL_X32 FILLER_256_1016 ();
 FILLCELL_X32 FILLER_256_1048 ();
 FILLCELL_X32 FILLER_256_1080 ();
 FILLCELL_X32 FILLER_256_1112 ();
 FILLCELL_X32 FILLER_256_1144 ();
 FILLCELL_X32 FILLER_256_1176 ();
 FILLCELL_X32 FILLER_256_1208 ();
 FILLCELL_X32 FILLER_256_1240 ();
 FILLCELL_X32 FILLER_256_1272 ();
 FILLCELL_X32 FILLER_256_1304 ();
 FILLCELL_X32 FILLER_256_1336 ();
 FILLCELL_X32 FILLER_256_1368 ();
 FILLCELL_X16 FILLER_256_1400 ();
 FILLCELL_X8 FILLER_256_1416 ();
 FILLCELL_X1 FILLER_256_1424 ();
 FILLCELL_X8 FILLER_256_1449 ();
 FILLCELL_X4 FILLER_256_1457 ();
 FILLCELL_X2 FILLER_256_1461 ();
 FILLCELL_X32 FILLER_256_1487 ();
 FILLCELL_X16 FILLER_256_1519 ();
 FILLCELL_X4 FILLER_256_1535 ();
 FILLCELL_X8 FILLER_256_1563 ();
 FILLCELL_X4 FILLER_256_1571 ();
 FILLCELL_X2 FILLER_256_1575 ();
 FILLCELL_X4 FILLER_256_1594 ();
 FILLCELL_X2 FILLER_256_1598 ();
 FILLCELL_X4 FILLER_256_1622 ();
 FILLCELL_X1 FILLER_256_1626 ();
 FILLCELL_X32 FILLER_256_1651 ();
 FILLCELL_X16 FILLER_256_1683 ();
 FILLCELL_X4 FILLER_256_1699 ();
 FILLCELL_X2 FILLER_256_1703 ();
 FILLCELL_X1 FILLER_256_1705 ();
 FILLCELL_X32 FILLER_256_1713 ();
 FILLCELL_X16 FILLER_256_1745 ();
 FILLCELL_X8 FILLER_256_1761 ();
 FILLCELL_X4 FILLER_256_1769 ();
 FILLCELL_X16 FILLER_256_1778 ();
 FILLCELL_X8 FILLER_256_1804 ();
 FILLCELL_X1 FILLER_256_1812 ();
 FILLCELL_X32 FILLER_256_1853 ();
 FILLCELL_X8 FILLER_256_1885 ();
 FILLCELL_X1 FILLER_256_1893 ();
 FILLCELL_X16 FILLER_256_1895 ();
 FILLCELL_X8 FILLER_256_1911 ();
 FILLCELL_X4 FILLER_256_1919 ();
 FILLCELL_X2 FILLER_256_1923 ();
 FILLCELL_X1 FILLER_256_1925 ();
 FILLCELL_X32 FILLER_256_1945 ();
 FILLCELL_X4 FILLER_256_1977 ();
 FILLCELL_X2 FILLER_256_1981 ();
 FILLCELL_X8 FILLER_256_2002 ();
 FILLCELL_X4 FILLER_256_2010 ();
 FILLCELL_X1 FILLER_256_2014 ();
 FILLCELL_X8 FILLER_256_2021 ();
 FILLCELL_X4 FILLER_256_2029 ();
 FILLCELL_X2 FILLER_256_2033 ();
 FILLCELL_X1 FILLER_256_2035 ();
 FILLCELL_X2 FILLER_256_2041 ();
 FILLCELL_X32 FILLER_256_2060 ();
 FILLCELL_X8 FILLER_256_2092 ();
 FILLCELL_X4 FILLER_256_2100 ();
 FILLCELL_X8 FILLER_256_2107 ();
 FILLCELL_X4 FILLER_256_2127 ();
 FILLCELL_X2 FILLER_256_2131 ();
 FILLCELL_X1 FILLER_256_2133 ();
 FILLCELL_X4 FILLER_256_2137 ();
 FILLCELL_X16 FILLER_256_2144 ();
 FILLCELL_X4 FILLER_256_2160 ();
 FILLCELL_X16 FILLER_256_2167 ();
 FILLCELL_X8 FILLER_256_2183 ();
 FILLCELL_X4 FILLER_256_2191 ();
 FILLCELL_X2 FILLER_256_2195 ();
 FILLCELL_X1 FILLER_256_2197 ();
 FILLCELL_X8 FILLER_256_2201 ();
 FILLCELL_X32 FILLER_256_2216 ();
 FILLCELL_X32 FILLER_256_2248 ();
 FILLCELL_X8 FILLER_256_2280 ();
 FILLCELL_X1 FILLER_256_2288 ();
 FILLCELL_X1 FILLER_256_2296 ();
 FILLCELL_X32 FILLER_256_2304 ();
 FILLCELL_X32 FILLER_256_2336 ();
 FILLCELL_X32 FILLER_256_2368 ();
 FILLCELL_X32 FILLER_256_2400 ();
 FILLCELL_X32 FILLER_256_2432 ();
 FILLCELL_X32 FILLER_256_2464 ();
 FILLCELL_X32 FILLER_256_2496 ();
 FILLCELL_X32 FILLER_256_2528 ();
 FILLCELL_X32 FILLER_256_2560 ();
 FILLCELL_X32 FILLER_256_2592 ();
 FILLCELL_X32 FILLER_256_2624 ();
 FILLCELL_X32 FILLER_256_2656 ();
 FILLCELL_X32 FILLER_256_2688 ();
 FILLCELL_X32 FILLER_256_2720 ();
 FILLCELL_X32 FILLER_256_2752 ();
 FILLCELL_X32 FILLER_256_2784 ();
 FILLCELL_X32 FILLER_256_2816 ();
 FILLCELL_X32 FILLER_256_2848 ();
 FILLCELL_X32 FILLER_256_2880 ();
 FILLCELL_X32 FILLER_256_2912 ();
 FILLCELL_X32 FILLER_256_2944 ();
 FILLCELL_X32 FILLER_256_2976 ();
 FILLCELL_X32 FILLER_256_3008 ();
 FILLCELL_X32 FILLER_256_3040 ();
 FILLCELL_X32 FILLER_256_3072 ();
 FILLCELL_X32 FILLER_256_3104 ();
 FILLCELL_X16 FILLER_256_3136 ();
 FILLCELL_X4 FILLER_256_3152 ();
 FILLCELL_X1 FILLER_256_3156 ();
 FILLCELL_X32 FILLER_256_3158 ();
 FILLCELL_X32 FILLER_256_3190 ();
 FILLCELL_X32 FILLER_256_3222 ();
 FILLCELL_X32 FILLER_256_3254 ();
 FILLCELL_X32 FILLER_256_3286 ();
 FILLCELL_X32 FILLER_256_3318 ();
 FILLCELL_X32 FILLER_256_3350 ();
 FILLCELL_X32 FILLER_256_3382 ();
 FILLCELL_X32 FILLER_256_3414 ();
 FILLCELL_X32 FILLER_256_3446 ();
 FILLCELL_X32 FILLER_256_3478 ();
 FILLCELL_X32 FILLER_256_3510 ();
 FILLCELL_X32 FILLER_256_3542 ();
 FILLCELL_X32 FILLER_256_3574 ();
 FILLCELL_X32 FILLER_256_3606 ();
 FILLCELL_X32 FILLER_256_3638 ();
 FILLCELL_X32 FILLER_256_3670 ();
 FILLCELL_X32 FILLER_256_3702 ();
 FILLCELL_X4 FILLER_256_3734 ();
 FILLCELL_X32 FILLER_257_1 ();
 FILLCELL_X32 FILLER_257_33 ();
 FILLCELL_X32 FILLER_257_65 ();
 FILLCELL_X32 FILLER_257_97 ();
 FILLCELL_X32 FILLER_257_129 ();
 FILLCELL_X32 FILLER_257_161 ();
 FILLCELL_X32 FILLER_257_193 ();
 FILLCELL_X32 FILLER_257_225 ();
 FILLCELL_X32 FILLER_257_257 ();
 FILLCELL_X32 FILLER_257_289 ();
 FILLCELL_X32 FILLER_257_321 ();
 FILLCELL_X32 FILLER_257_353 ();
 FILLCELL_X32 FILLER_257_385 ();
 FILLCELL_X32 FILLER_257_417 ();
 FILLCELL_X32 FILLER_257_449 ();
 FILLCELL_X32 FILLER_257_481 ();
 FILLCELL_X32 FILLER_257_513 ();
 FILLCELL_X32 FILLER_257_545 ();
 FILLCELL_X32 FILLER_257_577 ();
 FILLCELL_X32 FILLER_257_609 ();
 FILLCELL_X32 FILLER_257_641 ();
 FILLCELL_X32 FILLER_257_673 ();
 FILLCELL_X32 FILLER_257_705 ();
 FILLCELL_X32 FILLER_257_737 ();
 FILLCELL_X32 FILLER_257_769 ();
 FILLCELL_X32 FILLER_257_801 ();
 FILLCELL_X32 FILLER_257_833 ();
 FILLCELL_X32 FILLER_257_865 ();
 FILLCELL_X32 FILLER_257_897 ();
 FILLCELL_X32 FILLER_257_929 ();
 FILLCELL_X32 FILLER_257_961 ();
 FILLCELL_X32 FILLER_257_993 ();
 FILLCELL_X32 FILLER_257_1025 ();
 FILLCELL_X32 FILLER_257_1057 ();
 FILLCELL_X32 FILLER_257_1089 ();
 FILLCELL_X32 FILLER_257_1121 ();
 FILLCELL_X32 FILLER_257_1153 ();
 FILLCELL_X32 FILLER_257_1185 ();
 FILLCELL_X32 FILLER_257_1217 ();
 FILLCELL_X8 FILLER_257_1249 ();
 FILLCELL_X4 FILLER_257_1257 ();
 FILLCELL_X2 FILLER_257_1261 ();
 FILLCELL_X32 FILLER_257_1264 ();
 FILLCELL_X32 FILLER_257_1296 ();
 FILLCELL_X32 FILLER_257_1328 ();
 FILLCELL_X32 FILLER_257_1360 ();
 FILLCELL_X32 FILLER_257_1392 ();
 FILLCELL_X8 FILLER_257_1424 ();
 FILLCELL_X4 FILLER_257_1432 ();
 FILLCELL_X1 FILLER_257_1436 ();
 FILLCELL_X8 FILLER_257_1461 ();
 FILLCELL_X4 FILLER_257_1469 ();
 FILLCELL_X1 FILLER_257_1473 ();
 FILLCELL_X32 FILLER_257_1505 ();
 FILLCELL_X32 FILLER_257_1537 ();
 FILLCELL_X8 FILLER_257_1569 ();
 FILLCELL_X4 FILLER_257_1577 ();
 FILLCELL_X32 FILLER_257_1588 ();
 FILLCELL_X32 FILLER_257_1620 ();
 FILLCELL_X32 FILLER_257_1652 ();
 FILLCELL_X16 FILLER_257_1684 ();
 FILLCELL_X4 FILLER_257_1700 ();
 FILLCELL_X1 FILLER_257_1704 ();
 FILLCELL_X16 FILLER_257_1712 ();
 FILLCELL_X4 FILLER_257_1728 ();
 FILLCELL_X1 FILLER_257_1732 ();
 FILLCELL_X8 FILLER_257_1740 ();
 FILLCELL_X4 FILLER_257_1748 ();
 FILLCELL_X2 FILLER_257_1752 ();
 FILLCELL_X1 FILLER_257_1754 ();
 FILLCELL_X32 FILLER_257_1759 ();
 FILLCELL_X32 FILLER_257_1791 ();
 FILLCELL_X32 FILLER_257_1823 ();
 FILLCELL_X32 FILLER_257_1855 ();
 FILLCELL_X32 FILLER_257_1887 ();
 FILLCELL_X32 FILLER_257_1919 ();
 FILLCELL_X32 FILLER_257_1951 ();
 FILLCELL_X8 FILLER_257_1983 ();
 FILLCELL_X4 FILLER_257_1991 ();
 FILLCELL_X2 FILLER_257_1995 ();
 FILLCELL_X1 FILLER_257_1997 ();
 FILLCELL_X8 FILLER_257_2001 ();
 FILLCELL_X4 FILLER_257_2009 ();
 FILLCELL_X8 FILLER_257_2023 ();
 FILLCELL_X4 FILLER_257_2031 ();
 FILLCELL_X2 FILLER_257_2035 ();
 FILLCELL_X8 FILLER_257_2044 ();
 FILLCELL_X4 FILLER_257_2052 ();
 FILLCELL_X2 FILLER_257_2062 ();
 FILLCELL_X1 FILLER_257_2064 ();
 FILLCELL_X8 FILLER_257_2070 ();
 FILLCELL_X2 FILLER_257_2078 ();
 FILLCELL_X1 FILLER_257_2080 ();
 FILLCELL_X16 FILLER_257_2091 ();
 FILLCELL_X8 FILLER_257_2107 ();
 FILLCELL_X4 FILLER_257_2115 ();
 FILLCELL_X1 FILLER_257_2119 ();
 FILLCELL_X2 FILLER_257_2123 ();
 FILLCELL_X1 FILLER_257_2125 ();
 FILLCELL_X8 FILLER_257_2129 ();
 FILLCELL_X4 FILLER_257_2137 ();
 FILLCELL_X16 FILLER_257_2144 ();
 FILLCELL_X8 FILLER_257_2160 ();
 FILLCELL_X4 FILLER_257_2168 ();
 FILLCELL_X1 FILLER_257_2172 ();
 FILLCELL_X2 FILLER_257_2176 ();
 FILLCELL_X8 FILLER_257_2185 ();
 FILLCELL_X4 FILLER_257_2193 ();
 FILLCELL_X1 FILLER_257_2197 ();
 FILLCELL_X4 FILLER_257_2201 ();
 FILLCELL_X2 FILLER_257_2205 ();
 FILLCELL_X1 FILLER_257_2207 ();
 FILLCELL_X32 FILLER_257_2211 ();
 FILLCELL_X32 FILLER_257_2243 ();
 FILLCELL_X8 FILLER_257_2275 ();
 FILLCELL_X2 FILLER_257_2283 ();
 FILLCELL_X32 FILLER_257_2302 ();
 FILLCELL_X32 FILLER_257_2334 ();
 FILLCELL_X32 FILLER_257_2366 ();
 FILLCELL_X32 FILLER_257_2398 ();
 FILLCELL_X32 FILLER_257_2430 ();
 FILLCELL_X32 FILLER_257_2462 ();
 FILLCELL_X32 FILLER_257_2494 ();
 FILLCELL_X32 FILLER_257_2527 ();
 FILLCELL_X32 FILLER_257_2559 ();
 FILLCELL_X32 FILLER_257_2591 ();
 FILLCELL_X32 FILLER_257_2623 ();
 FILLCELL_X32 FILLER_257_2655 ();
 FILLCELL_X32 FILLER_257_2687 ();
 FILLCELL_X32 FILLER_257_2719 ();
 FILLCELL_X32 FILLER_257_2751 ();
 FILLCELL_X32 FILLER_257_2783 ();
 FILLCELL_X32 FILLER_257_2815 ();
 FILLCELL_X32 FILLER_257_2847 ();
 FILLCELL_X32 FILLER_257_2879 ();
 FILLCELL_X32 FILLER_257_2911 ();
 FILLCELL_X32 FILLER_257_2943 ();
 FILLCELL_X32 FILLER_257_2975 ();
 FILLCELL_X32 FILLER_257_3007 ();
 FILLCELL_X32 FILLER_257_3039 ();
 FILLCELL_X32 FILLER_257_3071 ();
 FILLCELL_X32 FILLER_257_3103 ();
 FILLCELL_X32 FILLER_257_3135 ();
 FILLCELL_X32 FILLER_257_3167 ();
 FILLCELL_X32 FILLER_257_3199 ();
 FILLCELL_X32 FILLER_257_3231 ();
 FILLCELL_X32 FILLER_257_3263 ();
 FILLCELL_X32 FILLER_257_3295 ();
 FILLCELL_X32 FILLER_257_3327 ();
 FILLCELL_X32 FILLER_257_3359 ();
 FILLCELL_X32 FILLER_257_3391 ();
 FILLCELL_X32 FILLER_257_3423 ();
 FILLCELL_X32 FILLER_257_3455 ();
 FILLCELL_X32 FILLER_257_3487 ();
 FILLCELL_X32 FILLER_257_3519 ();
 FILLCELL_X32 FILLER_257_3551 ();
 FILLCELL_X32 FILLER_257_3583 ();
 FILLCELL_X32 FILLER_257_3615 ();
 FILLCELL_X32 FILLER_257_3647 ();
 FILLCELL_X32 FILLER_257_3679 ();
 FILLCELL_X16 FILLER_257_3711 ();
 FILLCELL_X8 FILLER_257_3727 ();
 FILLCELL_X2 FILLER_257_3735 ();
 FILLCELL_X1 FILLER_257_3737 ();
 FILLCELL_X32 FILLER_258_1 ();
 FILLCELL_X32 FILLER_258_33 ();
 FILLCELL_X32 FILLER_258_65 ();
 FILLCELL_X32 FILLER_258_97 ();
 FILLCELL_X32 FILLER_258_129 ();
 FILLCELL_X32 FILLER_258_161 ();
 FILLCELL_X32 FILLER_258_193 ();
 FILLCELL_X32 FILLER_258_225 ();
 FILLCELL_X32 FILLER_258_257 ();
 FILLCELL_X32 FILLER_258_289 ();
 FILLCELL_X32 FILLER_258_321 ();
 FILLCELL_X32 FILLER_258_353 ();
 FILLCELL_X32 FILLER_258_385 ();
 FILLCELL_X32 FILLER_258_417 ();
 FILLCELL_X32 FILLER_258_449 ();
 FILLCELL_X32 FILLER_258_481 ();
 FILLCELL_X32 FILLER_258_513 ();
 FILLCELL_X32 FILLER_258_545 ();
 FILLCELL_X32 FILLER_258_577 ();
 FILLCELL_X16 FILLER_258_609 ();
 FILLCELL_X4 FILLER_258_625 ();
 FILLCELL_X2 FILLER_258_629 ();
 FILLCELL_X32 FILLER_258_632 ();
 FILLCELL_X32 FILLER_258_664 ();
 FILLCELL_X32 FILLER_258_696 ();
 FILLCELL_X32 FILLER_258_728 ();
 FILLCELL_X32 FILLER_258_760 ();
 FILLCELL_X32 FILLER_258_792 ();
 FILLCELL_X32 FILLER_258_824 ();
 FILLCELL_X32 FILLER_258_856 ();
 FILLCELL_X32 FILLER_258_888 ();
 FILLCELL_X32 FILLER_258_920 ();
 FILLCELL_X32 FILLER_258_952 ();
 FILLCELL_X32 FILLER_258_984 ();
 FILLCELL_X32 FILLER_258_1016 ();
 FILLCELL_X32 FILLER_258_1048 ();
 FILLCELL_X32 FILLER_258_1080 ();
 FILLCELL_X32 FILLER_258_1112 ();
 FILLCELL_X32 FILLER_258_1144 ();
 FILLCELL_X32 FILLER_258_1176 ();
 FILLCELL_X32 FILLER_258_1208 ();
 FILLCELL_X32 FILLER_258_1240 ();
 FILLCELL_X32 FILLER_258_1272 ();
 FILLCELL_X32 FILLER_258_1304 ();
 FILLCELL_X32 FILLER_258_1336 ();
 FILLCELL_X32 FILLER_258_1368 ();
 FILLCELL_X32 FILLER_258_1400 ();
 FILLCELL_X16 FILLER_258_1432 ();
 FILLCELL_X2 FILLER_258_1448 ();
 FILLCELL_X32 FILLER_258_1457 ();
 FILLCELL_X16 FILLER_258_1489 ();
 FILLCELL_X8 FILLER_258_1505 ();
 FILLCELL_X4 FILLER_258_1513 ();
 FILLCELL_X2 FILLER_258_1517 ();
 FILLCELL_X1 FILLER_258_1519 ();
 FILLCELL_X8 FILLER_258_1527 ();
 FILLCELL_X4 FILLER_258_1535 ();
 FILLCELL_X2 FILLER_258_1539 ();
 FILLCELL_X1 FILLER_258_1541 ();
 FILLCELL_X4 FILLER_258_1550 ();
 FILLCELL_X32 FILLER_258_1571 ();
 FILLCELL_X16 FILLER_258_1603 ();
 FILLCELL_X4 FILLER_258_1619 ();
 FILLCELL_X16 FILLER_258_1630 ();
 FILLCELL_X8 FILLER_258_1646 ();
 FILLCELL_X32 FILLER_258_1661 ();
 FILLCELL_X8 FILLER_258_1693 ();
 FILLCELL_X2 FILLER_258_1701 ();
 FILLCELL_X4 FILLER_258_1720 ();
 FILLCELL_X1 FILLER_258_1724 ();
 FILLCELL_X16 FILLER_258_1738 ();
 FILLCELL_X1 FILLER_258_1754 ();
 FILLCELL_X8 FILLER_258_1768 ();
 FILLCELL_X2 FILLER_258_1776 ();
 FILLCELL_X4 FILLER_258_1783 ();
 FILLCELL_X2 FILLER_258_1787 ();
 FILLCELL_X32 FILLER_258_1799 ();
 FILLCELL_X32 FILLER_258_1831 ();
 FILLCELL_X16 FILLER_258_1863 ();
 FILLCELL_X8 FILLER_258_1879 ();
 FILLCELL_X4 FILLER_258_1887 ();
 FILLCELL_X2 FILLER_258_1891 ();
 FILLCELL_X1 FILLER_258_1893 ();
 FILLCELL_X32 FILLER_258_1895 ();
 FILLCELL_X32 FILLER_258_1927 ();
 FILLCELL_X32 FILLER_258_1959 ();
 FILLCELL_X16 FILLER_258_1991 ();
 FILLCELL_X8 FILLER_258_2007 ();
 FILLCELL_X1 FILLER_258_2015 ();
 FILLCELL_X8 FILLER_258_2019 ();
 FILLCELL_X2 FILLER_258_2027 ();
 FILLCELL_X1 FILLER_258_2029 ();
 FILLCELL_X16 FILLER_258_2047 ();
 FILLCELL_X2 FILLER_258_2070 ();
 FILLCELL_X1 FILLER_258_2072 ();
 FILLCELL_X8 FILLER_258_2080 ();
 FILLCELL_X2 FILLER_258_2091 ();
 FILLCELL_X1 FILLER_258_2093 ();
 FILLCELL_X8 FILLER_258_2097 ();
 FILLCELL_X4 FILLER_258_2105 ();
 FILLCELL_X8 FILLER_258_2116 ();
 FILLCELL_X1 FILLER_258_2124 ();
 FILLCELL_X16 FILLER_258_2128 ();
 FILLCELL_X8 FILLER_258_2144 ();
 FILLCELL_X4 FILLER_258_2152 ();
 FILLCELL_X1 FILLER_258_2156 ();
 FILLCELL_X16 FILLER_258_2195 ();
 FILLCELL_X2 FILLER_258_2211 ();
 FILLCELL_X1 FILLER_258_2213 ();
 FILLCELL_X8 FILLER_258_2220 ();
 FILLCELL_X2 FILLER_258_2228 ();
 FILLCELL_X1 FILLER_258_2230 ();
 FILLCELL_X8 FILLER_258_2238 ();
 FILLCELL_X1 FILLER_258_2246 ();
 FILLCELL_X32 FILLER_258_2271 ();
 FILLCELL_X32 FILLER_258_2303 ();
 FILLCELL_X32 FILLER_258_2335 ();
 FILLCELL_X32 FILLER_258_2367 ();
 FILLCELL_X32 FILLER_258_2399 ();
 FILLCELL_X32 FILLER_258_2431 ();
 FILLCELL_X32 FILLER_258_2463 ();
 FILLCELL_X32 FILLER_258_2495 ();
 FILLCELL_X32 FILLER_258_2527 ();
 FILLCELL_X32 FILLER_258_2559 ();
 FILLCELL_X32 FILLER_258_2591 ();
 FILLCELL_X32 FILLER_258_2623 ();
 FILLCELL_X32 FILLER_258_2655 ();
 FILLCELL_X32 FILLER_258_2687 ();
 FILLCELL_X32 FILLER_258_2719 ();
 FILLCELL_X32 FILLER_258_2751 ();
 FILLCELL_X32 FILLER_258_2783 ();
 FILLCELL_X32 FILLER_258_2815 ();
 FILLCELL_X32 FILLER_258_2847 ();
 FILLCELL_X32 FILLER_258_2879 ();
 FILLCELL_X32 FILLER_258_2911 ();
 FILLCELL_X32 FILLER_258_2943 ();
 FILLCELL_X32 FILLER_258_2975 ();
 FILLCELL_X32 FILLER_258_3007 ();
 FILLCELL_X32 FILLER_258_3039 ();
 FILLCELL_X32 FILLER_258_3071 ();
 FILLCELL_X32 FILLER_258_3103 ();
 FILLCELL_X16 FILLER_258_3135 ();
 FILLCELL_X4 FILLER_258_3151 ();
 FILLCELL_X2 FILLER_258_3155 ();
 FILLCELL_X32 FILLER_258_3158 ();
 FILLCELL_X32 FILLER_258_3190 ();
 FILLCELL_X32 FILLER_258_3222 ();
 FILLCELL_X32 FILLER_258_3254 ();
 FILLCELL_X32 FILLER_258_3286 ();
 FILLCELL_X32 FILLER_258_3318 ();
 FILLCELL_X32 FILLER_258_3350 ();
 FILLCELL_X32 FILLER_258_3382 ();
 FILLCELL_X32 FILLER_258_3414 ();
 FILLCELL_X32 FILLER_258_3446 ();
 FILLCELL_X32 FILLER_258_3478 ();
 FILLCELL_X32 FILLER_258_3510 ();
 FILLCELL_X32 FILLER_258_3542 ();
 FILLCELL_X32 FILLER_258_3574 ();
 FILLCELL_X32 FILLER_258_3606 ();
 FILLCELL_X32 FILLER_258_3638 ();
 FILLCELL_X32 FILLER_258_3670 ();
 FILLCELL_X32 FILLER_258_3702 ();
 FILLCELL_X4 FILLER_258_3734 ();
 FILLCELL_X32 FILLER_259_1 ();
 FILLCELL_X32 FILLER_259_33 ();
 FILLCELL_X32 FILLER_259_65 ();
 FILLCELL_X32 FILLER_259_97 ();
 FILLCELL_X32 FILLER_259_129 ();
 FILLCELL_X32 FILLER_259_161 ();
 FILLCELL_X32 FILLER_259_193 ();
 FILLCELL_X32 FILLER_259_225 ();
 FILLCELL_X32 FILLER_259_257 ();
 FILLCELL_X32 FILLER_259_289 ();
 FILLCELL_X32 FILLER_259_321 ();
 FILLCELL_X32 FILLER_259_353 ();
 FILLCELL_X32 FILLER_259_385 ();
 FILLCELL_X32 FILLER_259_417 ();
 FILLCELL_X32 FILLER_259_449 ();
 FILLCELL_X32 FILLER_259_481 ();
 FILLCELL_X32 FILLER_259_513 ();
 FILLCELL_X32 FILLER_259_545 ();
 FILLCELL_X32 FILLER_259_577 ();
 FILLCELL_X32 FILLER_259_609 ();
 FILLCELL_X32 FILLER_259_641 ();
 FILLCELL_X32 FILLER_259_673 ();
 FILLCELL_X32 FILLER_259_705 ();
 FILLCELL_X32 FILLER_259_737 ();
 FILLCELL_X32 FILLER_259_769 ();
 FILLCELL_X32 FILLER_259_801 ();
 FILLCELL_X32 FILLER_259_833 ();
 FILLCELL_X32 FILLER_259_865 ();
 FILLCELL_X32 FILLER_259_897 ();
 FILLCELL_X32 FILLER_259_929 ();
 FILLCELL_X32 FILLER_259_961 ();
 FILLCELL_X32 FILLER_259_993 ();
 FILLCELL_X32 FILLER_259_1025 ();
 FILLCELL_X32 FILLER_259_1057 ();
 FILLCELL_X32 FILLER_259_1089 ();
 FILLCELL_X32 FILLER_259_1121 ();
 FILLCELL_X32 FILLER_259_1153 ();
 FILLCELL_X32 FILLER_259_1185 ();
 FILLCELL_X32 FILLER_259_1217 ();
 FILLCELL_X8 FILLER_259_1249 ();
 FILLCELL_X4 FILLER_259_1257 ();
 FILLCELL_X2 FILLER_259_1261 ();
 FILLCELL_X32 FILLER_259_1264 ();
 FILLCELL_X32 FILLER_259_1296 ();
 FILLCELL_X32 FILLER_259_1328 ();
 FILLCELL_X32 FILLER_259_1360 ();
 FILLCELL_X32 FILLER_259_1392 ();
 FILLCELL_X4 FILLER_259_1424 ();
 FILLCELL_X1 FILLER_259_1428 ();
 FILLCELL_X2 FILLER_259_1453 ();
 FILLCELL_X32 FILLER_259_1463 ();
 FILLCELL_X16 FILLER_259_1495 ();
 FILLCELL_X4 FILLER_259_1511 ();
 FILLCELL_X16 FILLER_259_1532 ();
 FILLCELL_X1 FILLER_259_1548 ();
 FILLCELL_X2 FILLER_259_1556 ();
 FILLCELL_X32 FILLER_259_1572 ();
 FILLCELL_X8 FILLER_259_1604 ();
 FILLCELL_X4 FILLER_259_1612 ();
 FILLCELL_X1 FILLER_259_1616 ();
 FILLCELL_X16 FILLER_259_1634 ();
 FILLCELL_X16 FILLER_259_1667 ();
 FILLCELL_X2 FILLER_259_1683 ();
 FILLCELL_X16 FILLER_259_1692 ();
 FILLCELL_X8 FILLER_259_1708 ();
 FILLCELL_X4 FILLER_259_1716 ();
 FILLCELL_X16 FILLER_259_1740 ();
 FILLCELL_X8 FILLER_259_1756 ();
 FILLCELL_X4 FILLER_259_1764 ();
 FILLCELL_X2 FILLER_259_1768 ();
 FILLCELL_X1 FILLER_259_1790 ();
 FILLCELL_X8 FILLER_259_1796 ();
 FILLCELL_X1 FILLER_259_1804 ();
 FILLCELL_X2 FILLER_259_1818 ();
 FILLCELL_X32 FILLER_259_1827 ();
 FILLCELL_X32 FILLER_259_1859 ();
 FILLCELL_X32 FILLER_259_1891 ();
 FILLCELL_X32 FILLER_259_1923 ();
 FILLCELL_X16 FILLER_259_1955 ();
 FILLCELL_X1 FILLER_259_1971 ();
 FILLCELL_X8 FILLER_259_1979 ();
 FILLCELL_X2 FILLER_259_1987 ();
 FILLCELL_X1 FILLER_259_1989 ();
 FILLCELL_X16 FILLER_259_2029 ();
 FILLCELL_X8 FILLER_259_2045 ();
 FILLCELL_X4 FILLER_259_2053 ();
 FILLCELL_X16 FILLER_259_2074 ();
 FILLCELL_X8 FILLER_259_2090 ();
 FILLCELL_X1 FILLER_259_2098 ();
 FILLCELL_X16 FILLER_259_2123 ();
 FILLCELL_X2 FILLER_259_2139 ();
 FILLCELL_X1 FILLER_259_2141 ();
 FILLCELL_X2 FILLER_259_2149 ();
 FILLCELL_X1 FILLER_259_2151 ();
 FILLCELL_X1 FILLER_259_2159 ();
 FILLCELL_X8 FILLER_259_2168 ();
 FILLCELL_X4 FILLER_259_2176 ();
 FILLCELL_X1 FILLER_259_2180 ();
 FILLCELL_X16 FILLER_259_2198 ();
 FILLCELL_X8 FILLER_259_2214 ();
 FILLCELL_X2 FILLER_259_2222 ();
 FILLCELL_X1 FILLER_259_2224 ();
 FILLCELL_X2 FILLER_259_2253 ();
 FILLCELL_X16 FILLER_259_2267 ();
 FILLCELL_X4 FILLER_259_2283 ();
 FILLCELL_X2 FILLER_259_2294 ();
 FILLCELL_X2 FILLER_259_2303 ();
 FILLCELL_X1 FILLER_259_2305 ();
 FILLCELL_X32 FILLER_259_2330 ();
 FILLCELL_X32 FILLER_259_2362 ();
 FILLCELL_X32 FILLER_259_2394 ();
 FILLCELL_X32 FILLER_259_2426 ();
 FILLCELL_X32 FILLER_259_2458 ();
 FILLCELL_X32 FILLER_259_2490 ();
 FILLCELL_X4 FILLER_259_2522 ();
 FILLCELL_X32 FILLER_259_2527 ();
 FILLCELL_X32 FILLER_259_2559 ();
 FILLCELL_X32 FILLER_259_2591 ();
 FILLCELL_X32 FILLER_259_2623 ();
 FILLCELL_X32 FILLER_259_2655 ();
 FILLCELL_X32 FILLER_259_2687 ();
 FILLCELL_X32 FILLER_259_2719 ();
 FILLCELL_X32 FILLER_259_2751 ();
 FILLCELL_X32 FILLER_259_2783 ();
 FILLCELL_X32 FILLER_259_2815 ();
 FILLCELL_X32 FILLER_259_2847 ();
 FILLCELL_X32 FILLER_259_2879 ();
 FILLCELL_X32 FILLER_259_2911 ();
 FILLCELL_X32 FILLER_259_2943 ();
 FILLCELL_X32 FILLER_259_2975 ();
 FILLCELL_X32 FILLER_259_3007 ();
 FILLCELL_X32 FILLER_259_3039 ();
 FILLCELL_X32 FILLER_259_3071 ();
 FILLCELL_X32 FILLER_259_3103 ();
 FILLCELL_X32 FILLER_259_3135 ();
 FILLCELL_X32 FILLER_259_3167 ();
 FILLCELL_X32 FILLER_259_3199 ();
 FILLCELL_X32 FILLER_259_3231 ();
 FILLCELL_X32 FILLER_259_3263 ();
 FILLCELL_X32 FILLER_259_3295 ();
 FILLCELL_X32 FILLER_259_3327 ();
 FILLCELL_X32 FILLER_259_3359 ();
 FILLCELL_X32 FILLER_259_3391 ();
 FILLCELL_X32 FILLER_259_3423 ();
 FILLCELL_X32 FILLER_259_3455 ();
 FILLCELL_X32 FILLER_259_3487 ();
 FILLCELL_X32 FILLER_259_3519 ();
 FILLCELL_X32 FILLER_259_3551 ();
 FILLCELL_X32 FILLER_259_3583 ();
 FILLCELL_X32 FILLER_259_3615 ();
 FILLCELL_X32 FILLER_259_3647 ();
 FILLCELL_X32 FILLER_259_3679 ();
 FILLCELL_X8 FILLER_259_3711 ();
 FILLCELL_X4 FILLER_259_3719 ();
 FILLCELL_X1 FILLER_259_3723 ();
 FILLCELL_X8 FILLER_259_3727 ();
 FILLCELL_X2 FILLER_259_3735 ();
 FILLCELL_X1 FILLER_259_3737 ();
 FILLCELL_X32 FILLER_260_1 ();
 FILLCELL_X32 FILLER_260_33 ();
 FILLCELL_X32 FILLER_260_65 ();
 FILLCELL_X32 FILLER_260_97 ();
 FILLCELL_X32 FILLER_260_129 ();
 FILLCELL_X32 FILLER_260_161 ();
 FILLCELL_X32 FILLER_260_193 ();
 FILLCELL_X32 FILLER_260_225 ();
 FILLCELL_X32 FILLER_260_257 ();
 FILLCELL_X32 FILLER_260_289 ();
 FILLCELL_X32 FILLER_260_321 ();
 FILLCELL_X32 FILLER_260_353 ();
 FILLCELL_X32 FILLER_260_385 ();
 FILLCELL_X32 FILLER_260_417 ();
 FILLCELL_X32 FILLER_260_449 ();
 FILLCELL_X32 FILLER_260_481 ();
 FILLCELL_X32 FILLER_260_513 ();
 FILLCELL_X32 FILLER_260_545 ();
 FILLCELL_X32 FILLER_260_577 ();
 FILLCELL_X16 FILLER_260_609 ();
 FILLCELL_X4 FILLER_260_625 ();
 FILLCELL_X2 FILLER_260_629 ();
 FILLCELL_X32 FILLER_260_632 ();
 FILLCELL_X32 FILLER_260_664 ();
 FILLCELL_X32 FILLER_260_696 ();
 FILLCELL_X32 FILLER_260_728 ();
 FILLCELL_X32 FILLER_260_760 ();
 FILLCELL_X32 FILLER_260_792 ();
 FILLCELL_X32 FILLER_260_824 ();
 FILLCELL_X32 FILLER_260_856 ();
 FILLCELL_X32 FILLER_260_888 ();
 FILLCELL_X32 FILLER_260_920 ();
 FILLCELL_X32 FILLER_260_952 ();
 FILLCELL_X32 FILLER_260_984 ();
 FILLCELL_X32 FILLER_260_1016 ();
 FILLCELL_X32 FILLER_260_1048 ();
 FILLCELL_X32 FILLER_260_1080 ();
 FILLCELL_X32 FILLER_260_1112 ();
 FILLCELL_X32 FILLER_260_1144 ();
 FILLCELL_X32 FILLER_260_1176 ();
 FILLCELL_X32 FILLER_260_1208 ();
 FILLCELL_X32 FILLER_260_1240 ();
 FILLCELL_X32 FILLER_260_1272 ();
 FILLCELL_X32 FILLER_260_1304 ();
 FILLCELL_X32 FILLER_260_1336 ();
 FILLCELL_X32 FILLER_260_1368 ();
 FILLCELL_X16 FILLER_260_1400 ();
 FILLCELL_X8 FILLER_260_1416 ();
 FILLCELL_X4 FILLER_260_1424 ();
 FILLCELL_X2 FILLER_260_1428 ();
 FILLCELL_X1 FILLER_260_1430 ();
 FILLCELL_X32 FILLER_260_1438 ();
 FILLCELL_X2 FILLER_260_1470 ();
 FILLCELL_X1 FILLER_260_1479 ();
 FILLCELL_X32 FILLER_260_1487 ();
 FILLCELL_X16 FILLER_260_1519 ();
 FILLCELL_X8 FILLER_260_1535 ();
 FILLCELL_X2 FILLER_260_1543 ();
 FILLCELL_X16 FILLER_260_1562 ();
 FILLCELL_X4 FILLER_260_1578 ();
 FILLCELL_X4 FILLER_260_1606 ();
 FILLCELL_X1 FILLER_260_1610 ();
 FILLCELL_X8 FILLER_260_1635 ();
 FILLCELL_X4 FILLER_260_1643 ();
 FILLCELL_X32 FILLER_260_1664 ();
 FILLCELL_X16 FILLER_260_1696 ();
 FILLCELL_X8 FILLER_260_1712 ();
 FILLCELL_X1 FILLER_260_1720 ();
 FILLCELL_X1 FILLER_260_1734 ();
 FILLCELL_X32 FILLER_260_1742 ();
 FILLCELL_X4 FILLER_260_1774 ();
 FILLCELL_X1 FILLER_260_1778 ();
 FILLCELL_X1 FILLER_260_1786 ();
 FILLCELL_X1 FILLER_260_1791 ();
 FILLCELL_X8 FILLER_260_1802 ();
 FILLCELL_X4 FILLER_260_1810 ();
 FILLCELL_X2 FILLER_260_1814 ();
 FILLCELL_X1 FILLER_260_1816 ();
 FILLCELL_X16 FILLER_260_1836 ();
 FILLCELL_X2 FILLER_260_1852 ();
 FILLCELL_X16 FILLER_260_1868 ();
 FILLCELL_X8 FILLER_260_1884 ();
 FILLCELL_X2 FILLER_260_1892 ();
 FILLCELL_X8 FILLER_260_1895 ();
 FILLCELL_X2 FILLER_260_1903 ();
 FILLCELL_X1 FILLER_260_1905 ();
 FILLCELL_X32 FILLER_260_1924 ();
 FILLCELL_X8 FILLER_260_1956 ();
 FILLCELL_X2 FILLER_260_1964 ();
 FILLCELL_X1 FILLER_260_1966 ();
 FILLCELL_X8 FILLER_260_1984 ();
 FILLCELL_X2 FILLER_260_1992 ();
 FILLCELL_X1 FILLER_260_1994 ();
 FILLCELL_X32 FILLER_260_2019 ();
 FILLCELL_X32 FILLER_260_2051 ();
 FILLCELL_X16 FILLER_260_2083 ();
 FILLCELL_X8 FILLER_260_2099 ();
 FILLCELL_X2 FILLER_260_2107 ();
 FILLCELL_X16 FILLER_260_2116 ();
 FILLCELL_X4 FILLER_260_2132 ();
 FILLCELL_X1 FILLER_260_2136 ();
 FILLCELL_X32 FILLER_260_2154 ();
 FILLCELL_X32 FILLER_260_2186 ();
 FILLCELL_X4 FILLER_260_2218 ();
 FILLCELL_X32 FILLER_260_2229 ();
 FILLCELL_X16 FILLER_260_2261 ();
 FILLCELL_X4 FILLER_260_2277 ();
 FILLCELL_X1 FILLER_260_2281 ();
 FILLCELL_X32 FILLER_260_2299 ();
 FILLCELL_X32 FILLER_260_2331 ();
 FILLCELL_X32 FILLER_260_2363 ();
 FILLCELL_X32 FILLER_260_2395 ();
 FILLCELL_X32 FILLER_260_2427 ();
 FILLCELL_X32 FILLER_260_2459 ();
 FILLCELL_X32 FILLER_260_2491 ();
 FILLCELL_X32 FILLER_260_2523 ();
 FILLCELL_X32 FILLER_260_2555 ();
 FILLCELL_X32 FILLER_260_2587 ();
 FILLCELL_X32 FILLER_260_2619 ();
 FILLCELL_X32 FILLER_260_2651 ();
 FILLCELL_X32 FILLER_260_2683 ();
 FILLCELL_X32 FILLER_260_2715 ();
 FILLCELL_X32 FILLER_260_2747 ();
 FILLCELL_X32 FILLER_260_2779 ();
 FILLCELL_X32 FILLER_260_2811 ();
 FILLCELL_X32 FILLER_260_2843 ();
 FILLCELL_X32 FILLER_260_2875 ();
 FILLCELL_X32 FILLER_260_2907 ();
 FILLCELL_X32 FILLER_260_2939 ();
 FILLCELL_X32 FILLER_260_2971 ();
 FILLCELL_X32 FILLER_260_3003 ();
 FILLCELL_X32 FILLER_260_3035 ();
 FILLCELL_X32 FILLER_260_3067 ();
 FILLCELL_X32 FILLER_260_3099 ();
 FILLCELL_X16 FILLER_260_3131 ();
 FILLCELL_X8 FILLER_260_3147 ();
 FILLCELL_X2 FILLER_260_3155 ();
 FILLCELL_X32 FILLER_260_3158 ();
 FILLCELL_X32 FILLER_260_3190 ();
 FILLCELL_X32 FILLER_260_3222 ();
 FILLCELL_X32 FILLER_260_3254 ();
 FILLCELL_X32 FILLER_260_3286 ();
 FILLCELL_X32 FILLER_260_3318 ();
 FILLCELL_X32 FILLER_260_3350 ();
 FILLCELL_X32 FILLER_260_3382 ();
 FILLCELL_X32 FILLER_260_3414 ();
 FILLCELL_X32 FILLER_260_3446 ();
 FILLCELL_X32 FILLER_260_3478 ();
 FILLCELL_X32 FILLER_260_3510 ();
 FILLCELL_X32 FILLER_260_3542 ();
 FILLCELL_X32 FILLER_260_3574 ();
 FILLCELL_X32 FILLER_260_3606 ();
 FILLCELL_X32 FILLER_260_3638 ();
 FILLCELL_X32 FILLER_260_3670 ();
 FILLCELL_X16 FILLER_260_3702 ();
 FILLCELL_X8 FILLER_260_3718 ();
 FILLCELL_X8 FILLER_260_3729 ();
 FILLCELL_X1 FILLER_260_3737 ();
 FILLCELL_X32 FILLER_261_1 ();
 FILLCELL_X32 FILLER_261_33 ();
 FILLCELL_X32 FILLER_261_65 ();
 FILLCELL_X32 FILLER_261_97 ();
 FILLCELL_X32 FILLER_261_129 ();
 FILLCELL_X32 FILLER_261_161 ();
 FILLCELL_X32 FILLER_261_193 ();
 FILLCELL_X32 FILLER_261_225 ();
 FILLCELL_X32 FILLER_261_257 ();
 FILLCELL_X32 FILLER_261_289 ();
 FILLCELL_X32 FILLER_261_321 ();
 FILLCELL_X32 FILLER_261_353 ();
 FILLCELL_X32 FILLER_261_385 ();
 FILLCELL_X32 FILLER_261_417 ();
 FILLCELL_X32 FILLER_261_449 ();
 FILLCELL_X32 FILLER_261_481 ();
 FILLCELL_X32 FILLER_261_513 ();
 FILLCELL_X32 FILLER_261_545 ();
 FILLCELL_X32 FILLER_261_577 ();
 FILLCELL_X32 FILLER_261_609 ();
 FILLCELL_X32 FILLER_261_641 ();
 FILLCELL_X32 FILLER_261_673 ();
 FILLCELL_X32 FILLER_261_705 ();
 FILLCELL_X32 FILLER_261_737 ();
 FILLCELL_X32 FILLER_261_769 ();
 FILLCELL_X32 FILLER_261_801 ();
 FILLCELL_X32 FILLER_261_833 ();
 FILLCELL_X32 FILLER_261_865 ();
 FILLCELL_X32 FILLER_261_897 ();
 FILLCELL_X32 FILLER_261_929 ();
 FILLCELL_X32 FILLER_261_961 ();
 FILLCELL_X32 FILLER_261_993 ();
 FILLCELL_X32 FILLER_261_1025 ();
 FILLCELL_X32 FILLER_261_1057 ();
 FILLCELL_X32 FILLER_261_1089 ();
 FILLCELL_X32 FILLER_261_1121 ();
 FILLCELL_X32 FILLER_261_1153 ();
 FILLCELL_X32 FILLER_261_1185 ();
 FILLCELL_X32 FILLER_261_1217 ();
 FILLCELL_X8 FILLER_261_1249 ();
 FILLCELL_X4 FILLER_261_1257 ();
 FILLCELL_X2 FILLER_261_1261 ();
 FILLCELL_X32 FILLER_261_1264 ();
 FILLCELL_X32 FILLER_261_1296 ();
 FILLCELL_X32 FILLER_261_1328 ();
 FILLCELL_X32 FILLER_261_1360 ();
 FILLCELL_X16 FILLER_261_1392 ();
 FILLCELL_X8 FILLER_261_1408 ();
 FILLCELL_X4 FILLER_261_1416 ();
 FILLCELL_X8 FILLER_261_1437 ();
 FILLCELL_X8 FILLER_261_1452 ();
 FILLCELL_X2 FILLER_261_1460 ();
 FILLCELL_X1 FILLER_261_1462 ();
 FILLCELL_X2 FILLER_261_1480 ();
 FILLCELL_X1 FILLER_261_1482 ();
 FILLCELL_X16 FILLER_261_1500 ();
 FILLCELL_X8 FILLER_261_1516 ();
 FILLCELL_X2 FILLER_261_1524 ();
 FILLCELL_X32 FILLER_261_1533 ();
 FILLCELL_X32 FILLER_261_1565 ();
 FILLCELL_X16 FILLER_261_1597 ();
 FILLCELL_X8 FILLER_261_1613 ();
 FILLCELL_X1 FILLER_261_1621 ();
 FILLCELL_X16 FILLER_261_1629 ();
 FILLCELL_X2 FILLER_261_1645 ();
 FILLCELL_X8 FILLER_261_1671 ();
 FILLCELL_X4 FILLER_261_1679 ();
 FILLCELL_X2 FILLER_261_1683 ();
 FILLCELL_X16 FILLER_261_1709 ();
 FILLCELL_X4 FILLER_261_1725 ();
 FILLCELL_X2 FILLER_261_1729 ();
 FILLCELL_X2 FILLER_261_1751 ();
 FILLCELL_X1 FILLER_261_1753 ();
 FILLCELL_X32 FILLER_261_1767 ();
 FILLCELL_X4 FILLER_261_1799 ();
 FILLCELL_X2 FILLER_261_1803 ();
 FILLCELL_X16 FILLER_261_1810 ();
 FILLCELL_X8 FILLER_261_1826 ();
 FILLCELL_X8 FILLER_261_1844 ();
 FILLCELL_X16 FILLER_261_1863 ();
 FILLCELL_X4 FILLER_261_1879 ();
 FILLCELL_X1 FILLER_261_1883 ();
 FILLCELL_X32 FILLER_261_1920 ();
 FILLCELL_X32 FILLER_261_1952 ();
 FILLCELL_X8 FILLER_261_1984 ();
 FILLCELL_X2 FILLER_261_1992 ();
 FILLCELL_X32 FILLER_261_2001 ();
 FILLCELL_X4 FILLER_261_2033 ();
 FILLCELL_X2 FILLER_261_2037 ();
 FILLCELL_X32 FILLER_261_2046 ();
 FILLCELL_X2 FILLER_261_2078 ();
 FILLCELL_X1 FILLER_261_2080 ();
 FILLCELL_X1 FILLER_261_2098 ();
 FILLCELL_X32 FILLER_261_2116 ();
 FILLCELL_X16 FILLER_261_2148 ();
 FILLCELL_X4 FILLER_261_2164 ();
 FILLCELL_X4 FILLER_261_2175 ();
 FILLCELL_X2 FILLER_261_2186 ();
 FILLCELL_X16 FILLER_261_2229 ();
 FILLCELL_X8 FILLER_261_2245 ();
 FILLCELL_X4 FILLER_261_2253 ();
 FILLCELL_X1 FILLER_261_2257 ();
 FILLCELL_X32 FILLER_261_2265 ();
 FILLCELL_X32 FILLER_261_2297 ();
 FILLCELL_X32 FILLER_261_2329 ();
 FILLCELL_X32 FILLER_261_2361 ();
 FILLCELL_X32 FILLER_261_2393 ();
 FILLCELL_X32 FILLER_261_2425 ();
 FILLCELL_X32 FILLER_261_2457 ();
 FILLCELL_X32 FILLER_261_2489 ();
 FILLCELL_X4 FILLER_261_2521 ();
 FILLCELL_X1 FILLER_261_2525 ();
 FILLCELL_X32 FILLER_261_2527 ();
 FILLCELL_X32 FILLER_261_2559 ();
 FILLCELL_X32 FILLER_261_2591 ();
 FILLCELL_X32 FILLER_261_2623 ();
 FILLCELL_X32 FILLER_261_2655 ();
 FILLCELL_X32 FILLER_261_2687 ();
 FILLCELL_X32 FILLER_261_2719 ();
 FILLCELL_X32 FILLER_261_2751 ();
 FILLCELL_X32 FILLER_261_2783 ();
 FILLCELL_X32 FILLER_261_2815 ();
 FILLCELL_X32 FILLER_261_2847 ();
 FILLCELL_X32 FILLER_261_2879 ();
 FILLCELL_X32 FILLER_261_2911 ();
 FILLCELL_X32 FILLER_261_2943 ();
 FILLCELL_X32 FILLER_261_2975 ();
 FILLCELL_X32 FILLER_261_3007 ();
 FILLCELL_X32 FILLER_261_3039 ();
 FILLCELL_X32 FILLER_261_3071 ();
 FILLCELL_X32 FILLER_261_3103 ();
 FILLCELL_X32 FILLER_261_3135 ();
 FILLCELL_X32 FILLER_261_3167 ();
 FILLCELL_X32 FILLER_261_3199 ();
 FILLCELL_X32 FILLER_261_3231 ();
 FILLCELL_X32 FILLER_261_3263 ();
 FILLCELL_X32 FILLER_261_3295 ();
 FILLCELL_X32 FILLER_261_3327 ();
 FILLCELL_X32 FILLER_261_3359 ();
 FILLCELL_X32 FILLER_261_3391 ();
 FILLCELL_X32 FILLER_261_3423 ();
 FILLCELL_X32 FILLER_261_3455 ();
 FILLCELL_X32 FILLER_261_3487 ();
 FILLCELL_X32 FILLER_261_3519 ();
 FILLCELL_X32 FILLER_261_3551 ();
 FILLCELL_X32 FILLER_261_3583 ();
 FILLCELL_X32 FILLER_261_3615 ();
 FILLCELL_X32 FILLER_261_3647 ();
 FILLCELL_X32 FILLER_261_3679 ();
 FILLCELL_X4 FILLER_261_3711 ();
 FILLCELL_X1 FILLER_261_3715 ();
 FILLCELL_X8 FILLER_261_3719 ();
 FILLCELL_X2 FILLER_261_3727 ();
 FILLCELL_X4 FILLER_261_3732 ();
 FILLCELL_X2 FILLER_261_3736 ();
 FILLCELL_X32 FILLER_262_1 ();
 FILLCELL_X32 FILLER_262_33 ();
 FILLCELL_X32 FILLER_262_65 ();
 FILLCELL_X32 FILLER_262_97 ();
 FILLCELL_X32 FILLER_262_129 ();
 FILLCELL_X32 FILLER_262_161 ();
 FILLCELL_X32 FILLER_262_193 ();
 FILLCELL_X32 FILLER_262_225 ();
 FILLCELL_X32 FILLER_262_257 ();
 FILLCELL_X32 FILLER_262_289 ();
 FILLCELL_X32 FILLER_262_321 ();
 FILLCELL_X32 FILLER_262_353 ();
 FILLCELL_X32 FILLER_262_385 ();
 FILLCELL_X32 FILLER_262_417 ();
 FILLCELL_X32 FILLER_262_449 ();
 FILLCELL_X32 FILLER_262_481 ();
 FILLCELL_X32 FILLER_262_513 ();
 FILLCELL_X32 FILLER_262_545 ();
 FILLCELL_X32 FILLER_262_577 ();
 FILLCELL_X16 FILLER_262_609 ();
 FILLCELL_X4 FILLER_262_625 ();
 FILLCELL_X2 FILLER_262_629 ();
 FILLCELL_X32 FILLER_262_632 ();
 FILLCELL_X32 FILLER_262_664 ();
 FILLCELL_X32 FILLER_262_696 ();
 FILLCELL_X32 FILLER_262_728 ();
 FILLCELL_X32 FILLER_262_760 ();
 FILLCELL_X32 FILLER_262_792 ();
 FILLCELL_X32 FILLER_262_824 ();
 FILLCELL_X32 FILLER_262_856 ();
 FILLCELL_X32 FILLER_262_888 ();
 FILLCELL_X32 FILLER_262_920 ();
 FILLCELL_X32 FILLER_262_952 ();
 FILLCELL_X32 FILLER_262_984 ();
 FILLCELL_X32 FILLER_262_1016 ();
 FILLCELL_X32 FILLER_262_1048 ();
 FILLCELL_X32 FILLER_262_1080 ();
 FILLCELL_X32 FILLER_262_1112 ();
 FILLCELL_X32 FILLER_262_1144 ();
 FILLCELL_X32 FILLER_262_1176 ();
 FILLCELL_X32 FILLER_262_1208 ();
 FILLCELL_X32 FILLER_262_1240 ();
 FILLCELL_X32 FILLER_262_1272 ();
 FILLCELL_X32 FILLER_262_1304 ();
 FILLCELL_X32 FILLER_262_1336 ();
 FILLCELL_X32 FILLER_262_1368 ();
 FILLCELL_X32 FILLER_262_1400 ();
 FILLCELL_X16 FILLER_262_1439 ();
 FILLCELL_X2 FILLER_262_1455 ();
 FILLCELL_X32 FILLER_262_1464 ();
 FILLCELL_X16 FILLER_262_1496 ();
 FILLCELL_X1 FILLER_262_1536 ();
 FILLCELL_X16 FILLER_262_1568 ();
 FILLCELL_X8 FILLER_262_1584 ();
 FILLCELL_X4 FILLER_262_1592 ();
 FILLCELL_X2 FILLER_262_1596 ();
 FILLCELL_X1 FILLER_262_1598 ();
 FILLCELL_X32 FILLER_262_1606 ();
 FILLCELL_X32 FILLER_262_1638 ();
 FILLCELL_X16 FILLER_262_1670 ();
 FILLCELL_X8 FILLER_262_1686 ();
 FILLCELL_X4 FILLER_262_1694 ();
 FILLCELL_X2 FILLER_262_1698 ();
 FILLCELL_X16 FILLER_262_1707 ();
 FILLCELL_X8 FILLER_262_1723 ();
 FILLCELL_X1 FILLER_262_1731 ();
 FILLCELL_X2 FILLER_262_1749 ();
 FILLCELL_X1 FILLER_262_1751 ();
 FILLCELL_X4 FILLER_262_1771 ();
 FILLCELL_X1 FILLER_262_1775 ();
 FILLCELL_X32 FILLER_262_1778 ();
 FILLCELL_X2 FILLER_262_1810 ();
 FILLCELL_X1 FILLER_262_1821 ();
 FILLCELL_X8 FILLER_262_1832 ();
 FILLCELL_X4 FILLER_262_1840 ();
 FILLCELL_X1 FILLER_262_1844 ();
 FILLCELL_X1 FILLER_262_1847 ();
 FILLCELL_X8 FILLER_262_1873 ();
 FILLCELL_X1 FILLER_262_1881 ();
 FILLCELL_X2 FILLER_262_1888 ();
 FILLCELL_X2 FILLER_262_1892 ();
 FILLCELL_X4 FILLER_262_1900 ();
 FILLCELL_X2 FILLER_262_1909 ();
 FILLCELL_X1 FILLER_262_1920 ();
 FILLCELL_X32 FILLER_262_1927 ();
 FILLCELL_X8 FILLER_262_1959 ();
 FILLCELL_X2 FILLER_262_1967 ();
 FILLCELL_X1 FILLER_262_1969 ();
 FILLCELL_X2 FILLER_262_1977 ();
 FILLCELL_X1 FILLER_262_1979 ();
 FILLCELL_X4 FILLER_262_1987 ();
 FILLCELL_X2 FILLER_262_1991 ();
 FILLCELL_X32 FILLER_262_1997 ();
 FILLCELL_X4 FILLER_262_2029 ();
 FILLCELL_X2 FILLER_262_2033 ();
 FILLCELL_X8 FILLER_262_2059 ();
 FILLCELL_X4 FILLER_262_2067 ();
 FILLCELL_X2 FILLER_262_2071 ();
 FILLCELL_X2 FILLER_262_2080 ();
 FILLCELL_X1 FILLER_262_2082 ();
 FILLCELL_X32 FILLER_262_2100 ();
 FILLCELL_X8 FILLER_262_2132 ();
 FILLCELL_X2 FILLER_262_2140 ();
 FILLCELL_X1 FILLER_262_2142 ();
 FILLCELL_X8 FILLER_262_2150 ();
 FILLCELL_X4 FILLER_262_2158 ();
 FILLCELL_X2 FILLER_262_2162 ();
 FILLCELL_X1 FILLER_262_2164 ();
 FILLCELL_X32 FILLER_262_2182 ();
 FILLCELL_X32 FILLER_262_2214 ();
 FILLCELL_X8 FILLER_262_2246 ();
 FILLCELL_X1 FILLER_262_2254 ();
 FILLCELL_X32 FILLER_262_2272 ();
 FILLCELL_X4 FILLER_262_2304 ();
 FILLCELL_X1 FILLER_262_2308 ();
 FILLCELL_X32 FILLER_262_2313 ();
 FILLCELL_X32 FILLER_262_2345 ();
 FILLCELL_X32 FILLER_262_2377 ();
 FILLCELL_X32 FILLER_262_2409 ();
 FILLCELL_X32 FILLER_262_2441 ();
 FILLCELL_X32 FILLER_262_2473 ();
 FILLCELL_X32 FILLER_262_2505 ();
 FILLCELL_X32 FILLER_262_2537 ();
 FILLCELL_X32 FILLER_262_2569 ();
 FILLCELL_X32 FILLER_262_2601 ();
 FILLCELL_X32 FILLER_262_2633 ();
 FILLCELL_X32 FILLER_262_2665 ();
 FILLCELL_X32 FILLER_262_2697 ();
 FILLCELL_X32 FILLER_262_2729 ();
 FILLCELL_X32 FILLER_262_2761 ();
 FILLCELL_X32 FILLER_262_2793 ();
 FILLCELL_X32 FILLER_262_2825 ();
 FILLCELL_X32 FILLER_262_2857 ();
 FILLCELL_X32 FILLER_262_2889 ();
 FILLCELL_X32 FILLER_262_2921 ();
 FILLCELL_X32 FILLER_262_2953 ();
 FILLCELL_X32 FILLER_262_2985 ();
 FILLCELL_X32 FILLER_262_3017 ();
 FILLCELL_X32 FILLER_262_3049 ();
 FILLCELL_X32 FILLER_262_3081 ();
 FILLCELL_X32 FILLER_262_3113 ();
 FILLCELL_X8 FILLER_262_3145 ();
 FILLCELL_X4 FILLER_262_3153 ();
 FILLCELL_X32 FILLER_262_3158 ();
 FILLCELL_X32 FILLER_262_3190 ();
 FILLCELL_X32 FILLER_262_3222 ();
 FILLCELL_X32 FILLER_262_3254 ();
 FILLCELL_X32 FILLER_262_3286 ();
 FILLCELL_X32 FILLER_262_3318 ();
 FILLCELL_X32 FILLER_262_3350 ();
 FILLCELL_X32 FILLER_262_3382 ();
 FILLCELL_X32 FILLER_262_3414 ();
 FILLCELL_X32 FILLER_262_3446 ();
 FILLCELL_X32 FILLER_262_3478 ();
 FILLCELL_X32 FILLER_262_3510 ();
 FILLCELL_X32 FILLER_262_3542 ();
 FILLCELL_X32 FILLER_262_3574 ();
 FILLCELL_X32 FILLER_262_3606 ();
 FILLCELL_X32 FILLER_262_3638 ();
 FILLCELL_X32 FILLER_262_3670 ();
 FILLCELL_X32 FILLER_262_3702 ();
 FILLCELL_X4 FILLER_262_3734 ();
 FILLCELL_X32 FILLER_263_1 ();
 FILLCELL_X32 FILLER_263_33 ();
 FILLCELL_X32 FILLER_263_65 ();
 FILLCELL_X32 FILLER_263_97 ();
 FILLCELL_X32 FILLER_263_129 ();
 FILLCELL_X32 FILLER_263_161 ();
 FILLCELL_X32 FILLER_263_193 ();
 FILLCELL_X32 FILLER_263_225 ();
 FILLCELL_X32 FILLER_263_257 ();
 FILLCELL_X32 FILLER_263_289 ();
 FILLCELL_X32 FILLER_263_321 ();
 FILLCELL_X32 FILLER_263_353 ();
 FILLCELL_X32 FILLER_263_385 ();
 FILLCELL_X32 FILLER_263_417 ();
 FILLCELL_X32 FILLER_263_449 ();
 FILLCELL_X32 FILLER_263_481 ();
 FILLCELL_X32 FILLER_263_513 ();
 FILLCELL_X32 FILLER_263_545 ();
 FILLCELL_X32 FILLER_263_577 ();
 FILLCELL_X32 FILLER_263_609 ();
 FILLCELL_X32 FILLER_263_641 ();
 FILLCELL_X32 FILLER_263_673 ();
 FILLCELL_X32 FILLER_263_705 ();
 FILLCELL_X32 FILLER_263_737 ();
 FILLCELL_X32 FILLER_263_769 ();
 FILLCELL_X32 FILLER_263_801 ();
 FILLCELL_X32 FILLER_263_833 ();
 FILLCELL_X32 FILLER_263_865 ();
 FILLCELL_X32 FILLER_263_897 ();
 FILLCELL_X32 FILLER_263_929 ();
 FILLCELL_X32 FILLER_263_961 ();
 FILLCELL_X32 FILLER_263_993 ();
 FILLCELL_X32 FILLER_263_1025 ();
 FILLCELL_X32 FILLER_263_1057 ();
 FILLCELL_X32 FILLER_263_1089 ();
 FILLCELL_X32 FILLER_263_1121 ();
 FILLCELL_X32 FILLER_263_1153 ();
 FILLCELL_X32 FILLER_263_1185 ();
 FILLCELL_X32 FILLER_263_1217 ();
 FILLCELL_X8 FILLER_263_1249 ();
 FILLCELL_X4 FILLER_263_1257 ();
 FILLCELL_X2 FILLER_263_1261 ();
 FILLCELL_X32 FILLER_263_1264 ();
 FILLCELL_X32 FILLER_263_1296 ();
 FILLCELL_X32 FILLER_263_1328 ();
 FILLCELL_X32 FILLER_263_1360 ();
 FILLCELL_X16 FILLER_263_1392 ();
 FILLCELL_X8 FILLER_263_1408 ();
 FILLCELL_X1 FILLER_263_1416 ();
 FILLCELL_X8 FILLER_263_1434 ();
 FILLCELL_X4 FILLER_263_1442 ();
 FILLCELL_X2 FILLER_263_1446 ();
 FILLCELL_X1 FILLER_263_1448 ();
 FILLCELL_X4 FILLER_263_1473 ();
 FILLCELL_X2 FILLER_263_1477 ();
 FILLCELL_X1 FILLER_263_1479 ();
 FILLCELL_X32 FILLER_263_1487 ();
 FILLCELL_X32 FILLER_263_1519 ();
 FILLCELL_X8 FILLER_263_1551 ();
 FILLCELL_X2 FILLER_263_1559 ();
 FILLCELL_X8 FILLER_263_1585 ();
 FILLCELL_X1 FILLER_263_1593 ();
 FILLCELL_X8 FILLER_263_1611 ();
 FILLCELL_X4 FILLER_263_1619 ();
 FILLCELL_X1 FILLER_263_1623 ();
 FILLCELL_X4 FILLER_263_1631 ();
 FILLCELL_X2 FILLER_263_1635 ();
 FILLCELL_X1 FILLER_263_1637 ();
 FILLCELL_X32 FILLER_263_1645 ();
 FILLCELL_X8 FILLER_263_1677 ();
 FILLCELL_X4 FILLER_263_1685 ();
 FILLCELL_X1 FILLER_263_1689 ();
 FILLCELL_X32 FILLER_263_1707 ();
 FILLCELL_X8 FILLER_263_1739 ();
 FILLCELL_X1 FILLER_263_1747 ();
 FILLCELL_X1 FILLER_263_1753 ();
 FILLCELL_X16 FILLER_263_1759 ();
 FILLCELL_X4 FILLER_263_1784 ();
 FILLCELL_X2 FILLER_263_1788 ();
 FILLCELL_X16 FILLER_263_1818 ();
 FILLCELL_X8 FILLER_263_1834 ();
 FILLCELL_X1 FILLER_263_1842 ();
 FILLCELL_X16 FILLER_263_1864 ();
 FILLCELL_X4 FILLER_263_1880 ();
 FILLCELL_X4 FILLER_263_1889 ();
 FILLCELL_X8 FILLER_263_1904 ();
 FILLCELL_X32 FILLER_263_1916 ();
 FILLCELL_X8 FILLER_263_1948 ();
 FILLCELL_X4 FILLER_263_1956 ();
 FILLCELL_X16 FILLER_263_1994 ();
 FILLCELL_X2 FILLER_263_2010 ();
 FILLCELL_X1 FILLER_263_2012 ();
 FILLCELL_X32 FILLER_263_2024 ();
 FILLCELL_X2 FILLER_263_2056 ();
 FILLCELL_X1 FILLER_263_2058 ();
 FILLCELL_X8 FILLER_263_2076 ();
 FILLCELL_X4 FILLER_263_2084 ();
 FILLCELL_X2 FILLER_263_2088 ();
 FILLCELL_X32 FILLER_263_2097 ();
 FILLCELL_X8 FILLER_263_2129 ();
 FILLCELL_X1 FILLER_263_2137 ();
 FILLCELL_X32 FILLER_263_2155 ();
 FILLCELL_X32 FILLER_263_2187 ();
 FILLCELL_X32 FILLER_263_2219 ();
 FILLCELL_X32 FILLER_263_2251 ();
 FILLCELL_X4 FILLER_263_2283 ();
 FILLCELL_X2 FILLER_263_2287 ();
 FILLCELL_X1 FILLER_263_2289 ();
 FILLCELL_X2 FILLER_263_2297 ();
 FILLCELL_X1 FILLER_263_2299 ();
 FILLCELL_X2 FILLER_263_2307 ();
 FILLCELL_X32 FILLER_263_2333 ();
 FILLCELL_X32 FILLER_263_2365 ();
 FILLCELL_X32 FILLER_263_2397 ();
 FILLCELL_X32 FILLER_263_2429 ();
 FILLCELL_X32 FILLER_263_2461 ();
 FILLCELL_X32 FILLER_263_2493 ();
 FILLCELL_X1 FILLER_263_2525 ();
 FILLCELL_X32 FILLER_263_2527 ();
 FILLCELL_X32 FILLER_263_2559 ();
 FILLCELL_X32 FILLER_263_2591 ();
 FILLCELL_X32 FILLER_263_2623 ();
 FILLCELL_X32 FILLER_263_2655 ();
 FILLCELL_X32 FILLER_263_2687 ();
 FILLCELL_X32 FILLER_263_2719 ();
 FILLCELL_X32 FILLER_263_2751 ();
 FILLCELL_X32 FILLER_263_2783 ();
 FILLCELL_X32 FILLER_263_2815 ();
 FILLCELL_X32 FILLER_263_2847 ();
 FILLCELL_X32 FILLER_263_2879 ();
 FILLCELL_X32 FILLER_263_2911 ();
 FILLCELL_X32 FILLER_263_2943 ();
 FILLCELL_X32 FILLER_263_2975 ();
 FILLCELL_X32 FILLER_263_3007 ();
 FILLCELL_X32 FILLER_263_3039 ();
 FILLCELL_X32 FILLER_263_3071 ();
 FILLCELL_X32 FILLER_263_3103 ();
 FILLCELL_X32 FILLER_263_3135 ();
 FILLCELL_X32 FILLER_263_3167 ();
 FILLCELL_X32 FILLER_263_3199 ();
 FILLCELL_X32 FILLER_263_3231 ();
 FILLCELL_X32 FILLER_263_3263 ();
 FILLCELL_X32 FILLER_263_3295 ();
 FILLCELL_X32 FILLER_263_3327 ();
 FILLCELL_X32 FILLER_263_3359 ();
 FILLCELL_X32 FILLER_263_3391 ();
 FILLCELL_X32 FILLER_263_3423 ();
 FILLCELL_X32 FILLER_263_3455 ();
 FILLCELL_X32 FILLER_263_3487 ();
 FILLCELL_X32 FILLER_263_3519 ();
 FILLCELL_X32 FILLER_263_3551 ();
 FILLCELL_X32 FILLER_263_3583 ();
 FILLCELL_X32 FILLER_263_3615 ();
 FILLCELL_X32 FILLER_263_3647 ();
 FILLCELL_X16 FILLER_263_3679 ();
 FILLCELL_X4 FILLER_263_3695 ();
 FILLCELL_X1 FILLER_263_3699 ();
 FILLCELL_X32 FILLER_263_3703 ();
 FILLCELL_X2 FILLER_263_3735 ();
 FILLCELL_X1 FILLER_263_3737 ();
 FILLCELL_X32 FILLER_264_1 ();
 FILLCELL_X32 FILLER_264_33 ();
 FILLCELL_X32 FILLER_264_65 ();
 FILLCELL_X32 FILLER_264_97 ();
 FILLCELL_X32 FILLER_264_129 ();
 FILLCELL_X32 FILLER_264_161 ();
 FILLCELL_X32 FILLER_264_193 ();
 FILLCELL_X32 FILLER_264_225 ();
 FILLCELL_X32 FILLER_264_257 ();
 FILLCELL_X32 FILLER_264_289 ();
 FILLCELL_X32 FILLER_264_321 ();
 FILLCELL_X32 FILLER_264_353 ();
 FILLCELL_X32 FILLER_264_385 ();
 FILLCELL_X32 FILLER_264_417 ();
 FILLCELL_X32 FILLER_264_449 ();
 FILLCELL_X32 FILLER_264_481 ();
 FILLCELL_X32 FILLER_264_513 ();
 FILLCELL_X32 FILLER_264_545 ();
 FILLCELL_X32 FILLER_264_577 ();
 FILLCELL_X16 FILLER_264_609 ();
 FILLCELL_X4 FILLER_264_625 ();
 FILLCELL_X2 FILLER_264_629 ();
 FILLCELL_X32 FILLER_264_632 ();
 FILLCELL_X32 FILLER_264_664 ();
 FILLCELL_X32 FILLER_264_696 ();
 FILLCELL_X32 FILLER_264_728 ();
 FILLCELL_X32 FILLER_264_760 ();
 FILLCELL_X32 FILLER_264_792 ();
 FILLCELL_X32 FILLER_264_824 ();
 FILLCELL_X32 FILLER_264_856 ();
 FILLCELL_X32 FILLER_264_888 ();
 FILLCELL_X32 FILLER_264_920 ();
 FILLCELL_X32 FILLER_264_952 ();
 FILLCELL_X32 FILLER_264_984 ();
 FILLCELL_X32 FILLER_264_1016 ();
 FILLCELL_X32 FILLER_264_1048 ();
 FILLCELL_X32 FILLER_264_1080 ();
 FILLCELL_X32 FILLER_264_1112 ();
 FILLCELL_X32 FILLER_264_1144 ();
 FILLCELL_X32 FILLER_264_1176 ();
 FILLCELL_X32 FILLER_264_1208 ();
 FILLCELL_X32 FILLER_264_1240 ();
 FILLCELL_X32 FILLER_264_1272 ();
 FILLCELL_X32 FILLER_264_1304 ();
 FILLCELL_X32 FILLER_264_1336 ();
 FILLCELL_X32 FILLER_264_1368 ();
 FILLCELL_X16 FILLER_264_1400 ();
 FILLCELL_X8 FILLER_264_1416 ();
 FILLCELL_X4 FILLER_264_1424 ();
 FILLCELL_X1 FILLER_264_1428 ();
 FILLCELL_X16 FILLER_264_1443 ();
 FILLCELL_X8 FILLER_264_1459 ();
 FILLCELL_X2 FILLER_264_1467 ();
 FILLCELL_X1 FILLER_264_1476 ();
 FILLCELL_X16 FILLER_264_1501 ();
 FILLCELL_X8 FILLER_264_1517 ();
 FILLCELL_X1 FILLER_264_1525 ();
 FILLCELL_X1 FILLER_264_1534 ();
 FILLCELL_X32 FILLER_264_1559 ();
 FILLCELL_X4 FILLER_264_1591 ();
 FILLCELL_X2 FILLER_264_1595 ();
 FILLCELL_X1 FILLER_264_1597 ();
 FILLCELL_X8 FILLER_264_1605 ();
 FILLCELL_X4 FILLER_264_1613 ();
 FILLCELL_X2 FILLER_264_1617 ();
 FILLCELL_X1 FILLER_264_1619 ();
 FILLCELL_X4 FILLER_264_1637 ();
 FILLCELL_X2 FILLER_264_1641 ();
 FILLCELL_X16 FILLER_264_1674 ();
 FILLCELL_X2 FILLER_264_1690 ();
 FILLCELL_X1 FILLER_264_1692 ();
 FILLCELL_X1 FILLER_264_1700 ();
 FILLCELL_X2 FILLER_264_1715 ();
 FILLCELL_X1 FILLER_264_1717 ();
 FILLCELL_X4 FILLER_264_1725 ();
 FILLCELL_X2 FILLER_264_1729 ();
 FILLCELL_X1 FILLER_264_1731 ();
 FILLCELL_X4 FILLER_264_1736 ();
 FILLCELL_X2 FILLER_264_1754 ();
 FILLCELL_X4 FILLER_264_1761 ();
 FILLCELL_X4 FILLER_264_1785 ();
 FILLCELL_X2 FILLER_264_1789 ();
 FILLCELL_X1 FILLER_264_1791 ();
 FILLCELL_X32 FILLER_264_1802 ();
 FILLCELL_X8 FILLER_264_1834 ();
 FILLCELL_X2 FILLER_264_1842 ();
 FILLCELL_X1 FILLER_264_1844 ();
 FILLCELL_X32 FILLER_264_1849 ();
 FILLCELL_X4 FILLER_264_1881 ();
 FILLCELL_X1 FILLER_264_1885 ();
 FILLCELL_X1 FILLER_264_1893 ();
 FILLCELL_X16 FILLER_264_1895 ();
 FILLCELL_X2 FILLER_264_1911 ();
 FILLCELL_X32 FILLER_264_1916 ();
 FILLCELL_X32 FILLER_264_1948 ();
 FILLCELL_X16 FILLER_264_1980 ();
 FILLCELL_X8 FILLER_264_1996 ();
 FILLCELL_X4 FILLER_264_2004 ();
 FILLCELL_X2 FILLER_264_2008 ();
 FILLCELL_X4 FILLER_264_2017 ();
 FILLCELL_X2 FILLER_264_2021 ();
 FILLCELL_X1 FILLER_264_2023 ();
 FILLCELL_X8 FILLER_264_2029 ();
 FILLCELL_X4 FILLER_264_2037 ();
 FILLCELL_X16 FILLER_264_2058 ();
 FILLCELL_X8 FILLER_264_2074 ();
 FILLCELL_X4 FILLER_264_2082 ();
 FILLCELL_X1 FILLER_264_2086 ();
 FILLCELL_X16 FILLER_264_2094 ();
 FILLCELL_X4 FILLER_264_2110 ();
 FILLCELL_X32 FILLER_264_2128 ();
 FILLCELL_X32 FILLER_264_2160 ();
 FILLCELL_X4 FILLER_264_2192 ();
 FILLCELL_X2 FILLER_264_2196 ();
 FILLCELL_X1 FILLER_264_2198 ();
 FILLCELL_X8 FILLER_264_2213 ();
 FILLCELL_X2 FILLER_264_2221 ();
 FILLCELL_X1 FILLER_264_2223 ();
 FILLCELL_X32 FILLER_264_2231 ();
 FILLCELL_X16 FILLER_264_2263 ();
 FILLCELL_X4 FILLER_264_2279 ();
 FILLCELL_X2 FILLER_264_2283 ();
 FILLCELL_X1 FILLER_264_2285 ();
 FILLCELL_X32 FILLER_264_2303 ();
 FILLCELL_X32 FILLER_264_2335 ();
 FILLCELL_X32 FILLER_264_2367 ();
 FILLCELL_X32 FILLER_264_2399 ();
 FILLCELL_X32 FILLER_264_2431 ();
 FILLCELL_X32 FILLER_264_2463 ();
 FILLCELL_X32 FILLER_264_2495 ();
 FILLCELL_X32 FILLER_264_2527 ();
 FILLCELL_X32 FILLER_264_2559 ();
 FILLCELL_X32 FILLER_264_2591 ();
 FILLCELL_X32 FILLER_264_2623 ();
 FILLCELL_X32 FILLER_264_2655 ();
 FILLCELL_X32 FILLER_264_2687 ();
 FILLCELL_X32 FILLER_264_2719 ();
 FILLCELL_X32 FILLER_264_2751 ();
 FILLCELL_X32 FILLER_264_2783 ();
 FILLCELL_X32 FILLER_264_2815 ();
 FILLCELL_X32 FILLER_264_2847 ();
 FILLCELL_X32 FILLER_264_2879 ();
 FILLCELL_X32 FILLER_264_2911 ();
 FILLCELL_X32 FILLER_264_2943 ();
 FILLCELL_X32 FILLER_264_2975 ();
 FILLCELL_X32 FILLER_264_3007 ();
 FILLCELL_X32 FILLER_264_3039 ();
 FILLCELL_X32 FILLER_264_3071 ();
 FILLCELL_X32 FILLER_264_3103 ();
 FILLCELL_X16 FILLER_264_3135 ();
 FILLCELL_X4 FILLER_264_3151 ();
 FILLCELL_X2 FILLER_264_3155 ();
 FILLCELL_X32 FILLER_264_3158 ();
 FILLCELL_X32 FILLER_264_3190 ();
 FILLCELL_X32 FILLER_264_3222 ();
 FILLCELL_X32 FILLER_264_3254 ();
 FILLCELL_X32 FILLER_264_3286 ();
 FILLCELL_X32 FILLER_264_3318 ();
 FILLCELL_X32 FILLER_264_3350 ();
 FILLCELL_X32 FILLER_264_3382 ();
 FILLCELL_X32 FILLER_264_3414 ();
 FILLCELL_X32 FILLER_264_3446 ();
 FILLCELL_X32 FILLER_264_3478 ();
 FILLCELL_X32 FILLER_264_3510 ();
 FILLCELL_X32 FILLER_264_3542 ();
 FILLCELL_X32 FILLER_264_3574 ();
 FILLCELL_X32 FILLER_264_3606 ();
 FILLCELL_X32 FILLER_264_3638 ();
 FILLCELL_X32 FILLER_264_3670 ();
 FILLCELL_X32 FILLER_264_3702 ();
 FILLCELL_X4 FILLER_264_3734 ();
 FILLCELL_X32 FILLER_265_1 ();
 FILLCELL_X32 FILLER_265_33 ();
 FILLCELL_X32 FILLER_265_65 ();
 FILLCELL_X32 FILLER_265_97 ();
 FILLCELL_X32 FILLER_265_129 ();
 FILLCELL_X32 FILLER_265_161 ();
 FILLCELL_X32 FILLER_265_193 ();
 FILLCELL_X32 FILLER_265_225 ();
 FILLCELL_X32 FILLER_265_257 ();
 FILLCELL_X32 FILLER_265_289 ();
 FILLCELL_X32 FILLER_265_321 ();
 FILLCELL_X32 FILLER_265_353 ();
 FILLCELL_X32 FILLER_265_385 ();
 FILLCELL_X32 FILLER_265_417 ();
 FILLCELL_X32 FILLER_265_449 ();
 FILLCELL_X32 FILLER_265_481 ();
 FILLCELL_X32 FILLER_265_513 ();
 FILLCELL_X32 FILLER_265_545 ();
 FILLCELL_X32 FILLER_265_577 ();
 FILLCELL_X32 FILLER_265_609 ();
 FILLCELL_X32 FILLER_265_641 ();
 FILLCELL_X32 FILLER_265_673 ();
 FILLCELL_X32 FILLER_265_705 ();
 FILLCELL_X32 FILLER_265_737 ();
 FILLCELL_X32 FILLER_265_769 ();
 FILLCELL_X32 FILLER_265_801 ();
 FILLCELL_X32 FILLER_265_833 ();
 FILLCELL_X32 FILLER_265_865 ();
 FILLCELL_X32 FILLER_265_897 ();
 FILLCELL_X32 FILLER_265_929 ();
 FILLCELL_X32 FILLER_265_961 ();
 FILLCELL_X32 FILLER_265_993 ();
 FILLCELL_X32 FILLER_265_1025 ();
 FILLCELL_X32 FILLER_265_1057 ();
 FILLCELL_X32 FILLER_265_1089 ();
 FILLCELL_X32 FILLER_265_1121 ();
 FILLCELL_X32 FILLER_265_1153 ();
 FILLCELL_X32 FILLER_265_1185 ();
 FILLCELL_X32 FILLER_265_1217 ();
 FILLCELL_X8 FILLER_265_1249 ();
 FILLCELL_X4 FILLER_265_1257 ();
 FILLCELL_X2 FILLER_265_1261 ();
 FILLCELL_X32 FILLER_265_1264 ();
 FILLCELL_X32 FILLER_265_1296 ();
 FILLCELL_X32 FILLER_265_1328 ();
 FILLCELL_X32 FILLER_265_1360 ();
 FILLCELL_X16 FILLER_265_1392 ();
 FILLCELL_X8 FILLER_265_1408 ();
 FILLCELL_X4 FILLER_265_1416 ();
 FILLCELL_X1 FILLER_265_1420 ();
 FILLCELL_X32 FILLER_265_1438 ();
 FILLCELL_X1 FILLER_265_1470 ();
 FILLCELL_X16 FILLER_265_1474 ();
 FILLCELL_X2 FILLER_265_1490 ();
 FILLCELL_X32 FILLER_265_1495 ();
 FILLCELL_X16 FILLER_265_1527 ();
 FILLCELL_X8 FILLER_265_1543 ();
 FILLCELL_X1 FILLER_265_1551 ();
 FILLCELL_X32 FILLER_265_1559 ();
 FILLCELL_X32 FILLER_265_1591 ();
 FILLCELL_X8 FILLER_265_1623 ();
 FILLCELL_X32 FILLER_265_1634 ();
 FILLCELL_X32 FILLER_265_1666 ();
 FILLCELL_X16 FILLER_265_1698 ();
 FILLCELL_X8 FILLER_265_1714 ();
 FILLCELL_X4 FILLER_265_1722 ();
 FILLCELL_X2 FILLER_265_1726 ();
 FILLCELL_X1 FILLER_265_1728 ();
 FILLCELL_X2 FILLER_265_1752 ();
 FILLCELL_X4 FILLER_265_1763 ();
 FILLCELL_X2 FILLER_265_1767 ();
 FILLCELL_X2 FILLER_265_1790 ();
 FILLCELL_X8 FILLER_265_1811 ();
 FILLCELL_X4 FILLER_265_1819 ();
 FILLCELL_X1 FILLER_265_1823 ();
 FILLCELL_X4 FILLER_265_1838 ();
 FILLCELL_X2 FILLER_265_1842 ();
 FILLCELL_X1 FILLER_265_1844 ();
 FILLCELL_X16 FILLER_265_1855 ();
 FILLCELL_X8 FILLER_265_1871 ();
 FILLCELL_X4 FILLER_265_1879 ();
 FILLCELL_X1 FILLER_265_1883 ();
 FILLCELL_X32 FILLER_265_1897 ();
 FILLCELL_X32 FILLER_265_1929 ();
 FILLCELL_X32 FILLER_265_1961 ();
 FILLCELL_X4 FILLER_265_1993 ();
 FILLCELL_X2 FILLER_265_1997 ();
 FILLCELL_X1 FILLER_265_1999 ();
 FILLCELL_X16 FILLER_265_2017 ();
 FILLCELL_X8 FILLER_265_2033 ();
 FILLCELL_X4 FILLER_265_2041 ();
 FILLCELL_X8 FILLER_265_2052 ();
 FILLCELL_X4 FILLER_265_2060 ();
 FILLCELL_X2 FILLER_265_2064 ();
 FILLCELL_X1 FILLER_265_2066 ();
 FILLCELL_X4 FILLER_265_2074 ();
 FILLCELL_X8 FILLER_265_2099 ();
 FILLCELL_X2 FILLER_265_2107 ();
 FILLCELL_X1 FILLER_265_2109 ();
 FILLCELL_X4 FILLER_265_2127 ();
 FILLCELL_X2 FILLER_265_2131 ();
 FILLCELL_X1 FILLER_265_2133 ();
 FILLCELL_X2 FILLER_265_2158 ();
 FILLCELL_X16 FILLER_265_2174 ();
 FILLCELL_X4 FILLER_265_2190 ();
 FILLCELL_X2 FILLER_265_2194 ();
 FILLCELL_X8 FILLER_265_2213 ();
 FILLCELL_X4 FILLER_265_2221 ();
 FILLCELL_X8 FILLER_265_2242 ();
 FILLCELL_X2 FILLER_265_2250 ();
 FILLCELL_X1 FILLER_265_2260 ();
 FILLCELL_X32 FILLER_265_2278 ();
 FILLCELL_X32 FILLER_265_2310 ();
 FILLCELL_X32 FILLER_265_2342 ();
 FILLCELL_X32 FILLER_265_2374 ();
 FILLCELL_X32 FILLER_265_2406 ();
 FILLCELL_X32 FILLER_265_2438 ();
 FILLCELL_X32 FILLER_265_2470 ();
 FILLCELL_X16 FILLER_265_2502 ();
 FILLCELL_X8 FILLER_265_2518 ();
 FILLCELL_X32 FILLER_265_2527 ();
 FILLCELL_X32 FILLER_265_2559 ();
 FILLCELL_X32 FILLER_265_2591 ();
 FILLCELL_X32 FILLER_265_2623 ();
 FILLCELL_X32 FILLER_265_2655 ();
 FILLCELL_X32 FILLER_265_2687 ();
 FILLCELL_X32 FILLER_265_2719 ();
 FILLCELL_X32 FILLER_265_2751 ();
 FILLCELL_X32 FILLER_265_2783 ();
 FILLCELL_X32 FILLER_265_2815 ();
 FILLCELL_X32 FILLER_265_2847 ();
 FILLCELL_X32 FILLER_265_2879 ();
 FILLCELL_X32 FILLER_265_2911 ();
 FILLCELL_X32 FILLER_265_2943 ();
 FILLCELL_X32 FILLER_265_2975 ();
 FILLCELL_X32 FILLER_265_3007 ();
 FILLCELL_X32 FILLER_265_3039 ();
 FILLCELL_X32 FILLER_265_3071 ();
 FILLCELL_X32 FILLER_265_3103 ();
 FILLCELL_X32 FILLER_265_3135 ();
 FILLCELL_X32 FILLER_265_3167 ();
 FILLCELL_X32 FILLER_265_3199 ();
 FILLCELL_X32 FILLER_265_3231 ();
 FILLCELL_X32 FILLER_265_3263 ();
 FILLCELL_X32 FILLER_265_3295 ();
 FILLCELL_X32 FILLER_265_3327 ();
 FILLCELL_X32 FILLER_265_3359 ();
 FILLCELL_X32 FILLER_265_3391 ();
 FILLCELL_X32 FILLER_265_3423 ();
 FILLCELL_X32 FILLER_265_3455 ();
 FILLCELL_X32 FILLER_265_3487 ();
 FILLCELL_X32 FILLER_265_3519 ();
 FILLCELL_X32 FILLER_265_3551 ();
 FILLCELL_X32 FILLER_265_3583 ();
 FILLCELL_X32 FILLER_265_3615 ();
 FILLCELL_X32 FILLER_265_3647 ();
 FILLCELL_X32 FILLER_265_3679 ();
 FILLCELL_X16 FILLER_265_3711 ();
 FILLCELL_X8 FILLER_265_3727 ();
 FILLCELL_X2 FILLER_265_3735 ();
 FILLCELL_X1 FILLER_265_3737 ();
 FILLCELL_X32 FILLER_266_1 ();
 FILLCELL_X32 FILLER_266_33 ();
 FILLCELL_X32 FILLER_266_65 ();
 FILLCELL_X32 FILLER_266_97 ();
 FILLCELL_X32 FILLER_266_129 ();
 FILLCELL_X32 FILLER_266_161 ();
 FILLCELL_X32 FILLER_266_193 ();
 FILLCELL_X32 FILLER_266_225 ();
 FILLCELL_X32 FILLER_266_257 ();
 FILLCELL_X32 FILLER_266_289 ();
 FILLCELL_X32 FILLER_266_321 ();
 FILLCELL_X32 FILLER_266_353 ();
 FILLCELL_X32 FILLER_266_385 ();
 FILLCELL_X32 FILLER_266_417 ();
 FILLCELL_X32 FILLER_266_449 ();
 FILLCELL_X32 FILLER_266_481 ();
 FILLCELL_X32 FILLER_266_513 ();
 FILLCELL_X32 FILLER_266_545 ();
 FILLCELL_X32 FILLER_266_577 ();
 FILLCELL_X16 FILLER_266_609 ();
 FILLCELL_X4 FILLER_266_625 ();
 FILLCELL_X2 FILLER_266_629 ();
 FILLCELL_X32 FILLER_266_632 ();
 FILLCELL_X32 FILLER_266_664 ();
 FILLCELL_X32 FILLER_266_696 ();
 FILLCELL_X32 FILLER_266_728 ();
 FILLCELL_X32 FILLER_266_760 ();
 FILLCELL_X32 FILLER_266_792 ();
 FILLCELL_X32 FILLER_266_824 ();
 FILLCELL_X32 FILLER_266_856 ();
 FILLCELL_X32 FILLER_266_888 ();
 FILLCELL_X32 FILLER_266_920 ();
 FILLCELL_X32 FILLER_266_952 ();
 FILLCELL_X32 FILLER_266_984 ();
 FILLCELL_X32 FILLER_266_1016 ();
 FILLCELL_X32 FILLER_266_1048 ();
 FILLCELL_X32 FILLER_266_1080 ();
 FILLCELL_X32 FILLER_266_1112 ();
 FILLCELL_X32 FILLER_266_1144 ();
 FILLCELL_X32 FILLER_266_1176 ();
 FILLCELL_X32 FILLER_266_1208 ();
 FILLCELL_X32 FILLER_266_1240 ();
 FILLCELL_X32 FILLER_266_1272 ();
 FILLCELL_X32 FILLER_266_1304 ();
 FILLCELL_X32 FILLER_266_1336 ();
 FILLCELL_X32 FILLER_266_1368 ();
 FILLCELL_X32 FILLER_266_1400 ();
 FILLCELL_X16 FILLER_266_1432 ();
 FILLCELL_X8 FILLER_266_1448 ();
 FILLCELL_X4 FILLER_266_1456 ();
 FILLCELL_X2 FILLER_266_1460 ();
 FILLCELL_X4 FILLER_266_1474 ();
 FILLCELL_X2 FILLER_266_1478 ();
 FILLCELL_X1 FILLER_266_1480 ();
 FILLCELL_X2 FILLER_266_1484 ();
 FILLCELL_X8 FILLER_266_1489 ();
 FILLCELL_X2 FILLER_266_1497 ();
 FILLCELL_X1 FILLER_266_1499 ();
 FILLCELL_X16 FILLER_266_1505 ();
 FILLCELL_X2 FILLER_266_1521 ();
 FILLCELL_X1 FILLER_266_1523 ();
 FILLCELL_X8 FILLER_266_1530 ();
 FILLCELL_X2 FILLER_266_1538 ();
 FILLCELL_X2 FILLER_266_1564 ();
 FILLCELL_X1 FILLER_266_1566 ();
 FILLCELL_X2 FILLER_266_1570 ();
 FILLCELL_X1 FILLER_266_1572 ();
 FILLCELL_X32 FILLER_266_1582 ();
 FILLCELL_X32 FILLER_266_1614 ();
 FILLCELL_X4 FILLER_266_1646 ();
 FILLCELL_X2 FILLER_266_1650 ();
 FILLCELL_X4 FILLER_266_1655 ();
 FILLCELL_X1 FILLER_266_1659 ();
 FILLCELL_X32 FILLER_266_1663 ();
 FILLCELL_X8 FILLER_266_1702 ();
 FILLCELL_X1 FILLER_266_1710 ();
 FILLCELL_X16 FILLER_266_1714 ();
 FILLCELL_X8 FILLER_266_1730 ();
 FILLCELL_X1 FILLER_266_1738 ();
 FILLCELL_X8 FILLER_266_1744 ();
 FILLCELL_X4 FILLER_266_1752 ();
 FILLCELL_X2 FILLER_266_1756 ();
 FILLCELL_X8 FILLER_266_1772 ();
 FILLCELL_X4 FILLER_266_1780 ();
 FILLCELL_X4 FILLER_266_1793 ();
 FILLCELL_X2 FILLER_266_1797 ();
 FILLCELL_X16 FILLER_266_1803 ();
 FILLCELL_X4 FILLER_266_1819 ();
 FILLCELL_X2 FILLER_266_1823 ();
 FILLCELL_X1 FILLER_266_1825 ();
 FILLCELL_X32 FILLER_266_1833 ();
 FILLCELL_X16 FILLER_266_1865 ();
 FILLCELL_X8 FILLER_266_1881 ();
 FILLCELL_X4 FILLER_266_1889 ();
 FILLCELL_X1 FILLER_266_1893 ();
 FILLCELL_X32 FILLER_266_1895 ();
 FILLCELL_X32 FILLER_266_1927 ();
 FILLCELL_X16 FILLER_266_1959 ();
 FILLCELL_X8 FILLER_266_1975 ();
 FILLCELL_X2 FILLER_266_1983 ();
 FILLCELL_X32 FILLER_266_1992 ();
 FILLCELL_X16 FILLER_266_2024 ();
 FILLCELL_X8 FILLER_266_2040 ();
 FILLCELL_X4 FILLER_266_2048 ();
 FILLCELL_X2 FILLER_266_2052 ();
 FILLCELL_X1 FILLER_266_2054 ();
 FILLCELL_X32 FILLER_266_2072 ();
 FILLCELL_X32 FILLER_266_2104 ();
 FILLCELL_X16 FILLER_266_2136 ();
 FILLCELL_X8 FILLER_266_2152 ();
 FILLCELL_X4 FILLER_266_2160 ();
 FILLCELL_X2 FILLER_266_2164 ();
 FILLCELL_X32 FILLER_266_2183 ();
 FILLCELL_X16 FILLER_266_2215 ();
 FILLCELL_X4 FILLER_266_2231 ();
 FILLCELL_X2 FILLER_266_2235 ();
 FILLCELL_X1 FILLER_266_2237 ();
 FILLCELL_X8 FILLER_266_2252 ();
 FILLCELL_X4 FILLER_266_2260 ();
 FILLCELL_X1 FILLER_266_2264 ();
 FILLCELL_X8 FILLER_266_2279 ();
 FILLCELL_X4 FILLER_266_2287 ();
 FILLCELL_X1 FILLER_266_2291 ();
 FILLCELL_X32 FILLER_266_2313 ();
 FILLCELL_X4 FILLER_266_2345 ();
 FILLCELL_X1 FILLER_266_2349 ();
 FILLCELL_X32 FILLER_266_2354 ();
 FILLCELL_X32 FILLER_266_2386 ();
 FILLCELL_X32 FILLER_266_2418 ();
 FILLCELL_X32 FILLER_266_2450 ();
 FILLCELL_X32 FILLER_266_2482 ();
 FILLCELL_X32 FILLER_266_2514 ();
 FILLCELL_X32 FILLER_266_2546 ();
 FILLCELL_X32 FILLER_266_2578 ();
 FILLCELL_X32 FILLER_266_2610 ();
 FILLCELL_X32 FILLER_266_2642 ();
 FILLCELL_X32 FILLER_266_2674 ();
 FILLCELL_X32 FILLER_266_2706 ();
 FILLCELL_X32 FILLER_266_2738 ();
 FILLCELL_X32 FILLER_266_2770 ();
 FILLCELL_X32 FILLER_266_2802 ();
 FILLCELL_X32 FILLER_266_2834 ();
 FILLCELL_X32 FILLER_266_2866 ();
 FILLCELL_X32 FILLER_266_2898 ();
 FILLCELL_X32 FILLER_266_2930 ();
 FILLCELL_X32 FILLER_266_2962 ();
 FILLCELL_X32 FILLER_266_2994 ();
 FILLCELL_X32 FILLER_266_3026 ();
 FILLCELL_X32 FILLER_266_3058 ();
 FILLCELL_X32 FILLER_266_3090 ();
 FILLCELL_X32 FILLER_266_3122 ();
 FILLCELL_X2 FILLER_266_3154 ();
 FILLCELL_X1 FILLER_266_3156 ();
 FILLCELL_X32 FILLER_266_3158 ();
 FILLCELL_X32 FILLER_266_3190 ();
 FILLCELL_X32 FILLER_266_3222 ();
 FILLCELL_X32 FILLER_266_3254 ();
 FILLCELL_X32 FILLER_266_3286 ();
 FILLCELL_X32 FILLER_266_3318 ();
 FILLCELL_X32 FILLER_266_3350 ();
 FILLCELL_X32 FILLER_266_3382 ();
 FILLCELL_X32 FILLER_266_3414 ();
 FILLCELL_X32 FILLER_266_3446 ();
 FILLCELL_X32 FILLER_266_3478 ();
 FILLCELL_X32 FILLER_266_3510 ();
 FILLCELL_X32 FILLER_266_3542 ();
 FILLCELL_X32 FILLER_266_3574 ();
 FILLCELL_X32 FILLER_266_3606 ();
 FILLCELL_X32 FILLER_266_3638 ();
 FILLCELL_X32 FILLER_266_3670 ();
 FILLCELL_X32 FILLER_266_3702 ();
 FILLCELL_X4 FILLER_266_3734 ();
 FILLCELL_X32 FILLER_267_1 ();
 FILLCELL_X32 FILLER_267_33 ();
 FILLCELL_X32 FILLER_267_65 ();
 FILLCELL_X32 FILLER_267_97 ();
 FILLCELL_X32 FILLER_267_129 ();
 FILLCELL_X32 FILLER_267_161 ();
 FILLCELL_X32 FILLER_267_193 ();
 FILLCELL_X32 FILLER_267_225 ();
 FILLCELL_X32 FILLER_267_257 ();
 FILLCELL_X32 FILLER_267_289 ();
 FILLCELL_X32 FILLER_267_321 ();
 FILLCELL_X32 FILLER_267_353 ();
 FILLCELL_X32 FILLER_267_385 ();
 FILLCELL_X32 FILLER_267_417 ();
 FILLCELL_X32 FILLER_267_449 ();
 FILLCELL_X32 FILLER_267_481 ();
 FILLCELL_X32 FILLER_267_513 ();
 FILLCELL_X32 FILLER_267_545 ();
 FILLCELL_X32 FILLER_267_577 ();
 FILLCELL_X32 FILLER_267_609 ();
 FILLCELL_X32 FILLER_267_641 ();
 FILLCELL_X32 FILLER_267_673 ();
 FILLCELL_X32 FILLER_267_705 ();
 FILLCELL_X32 FILLER_267_737 ();
 FILLCELL_X32 FILLER_267_769 ();
 FILLCELL_X32 FILLER_267_801 ();
 FILLCELL_X32 FILLER_267_833 ();
 FILLCELL_X32 FILLER_267_865 ();
 FILLCELL_X32 FILLER_267_897 ();
 FILLCELL_X32 FILLER_267_929 ();
 FILLCELL_X32 FILLER_267_961 ();
 FILLCELL_X32 FILLER_267_993 ();
 FILLCELL_X32 FILLER_267_1025 ();
 FILLCELL_X32 FILLER_267_1057 ();
 FILLCELL_X32 FILLER_267_1089 ();
 FILLCELL_X32 FILLER_267_1121 ();
 FILLCELL_X32 FILLER_267_1153 ();
 FILLCELL_X32 FILLER_267_1185 ();
 FILLCELL_X32 FILLER_267_1217 ();
 FILLCELL_X8 FILLER_267_1249 ();
 FILLCELL_X4 FILLER_267_1257 ();
 FILLCELL_X2 FILLER_267_1261 ();
 FILLCELL_X32 FILLER_267_1264 ();
 FILLCELL_X32 FILLER_267_1296 ();
 FILLCELL_X32 FILLER_267_1328 ();
 FILLCELL_X32 FILLER_267_1360 ();
 FILLCELL_X16 FILLER_267_1392 ();
 FILLCELL_X4 FILLER_267_1408 ();
 FILLCELL_X1 FILLER_267_1412 ();
 FILLCELL_X32 FILLER_267_1420 ();
 FILLCELL_X4 FILLER_267_1452 ();
 FILLCELL_X2 FILLER_267_1456 ();
 FILLCELL_X1 FILLER_267_1458 ();
 FILLCELL_X8 FILLER_267_1473 ();
 FILLCELL_X4 FILLER_267_1481 ();
 FILLCELL_X1 FILLER_267_1485 ();
 FILLCELL_X16 FILLER_267_1493 ();
 FILLCELL_X8 FILLER_267_1509 ();
 FILLCELL_X4 FILLER_267_1517 ();
 FILLCELL_X2 FILLER_267_1521 ();
 FILLCELL_X1 FILLER_267_1523 ();
 FILLCELL_X32 FILLER_267_1531 ();
 FILLCELL_X16 FILLER_267_1563 ();
 FILLCELL_X8 FILLER_267_1579 ();
 FILLCELL_X8 FILLER_267_1612 ();
 FILLCELL_X2 FILLER_267_1620 ();
 FILLCELL_X2 FILLER_267_1632 ();
 FILLCELL_X32 FILLER_267_1645 ();
 FILLCELL_X4 FILLER_267_1677 ();
 FILLCELL_X1 FILLER_267_1681 ();
 FILLCELL_X1 FILLER_267_1706 ();
 FILLCELL_X16 FILLER_267_1718 ();
 FILLCELL_X8 FILLER_267_1734 ();
 FILLCELL_X2 FILLER_267_1742 ();
 FILLCELL_X32 FILLER_267_1757 ();
 FILLCELL_X4 FILLER_267_1789 ();
 FILLCELL_X2 FILLER_267_1793 ();
 FILLCELL_X1 FILLER_267_1795 ();
 FILLCELL_X16 FILLER_267_1803 ();
 FILLCELL_X8 FILLER_267_1819 ();
 FILLCELL_X4 FILLER_267_1827 ();
 FILLCELL_X2 FILLER_267_1831 ();
 FILLCELL_X32 FILLER_267_1850 ();
 FILLCELL_X32 FILLER_267_1882 ();
 FILLCELL_X32 FILLER_267_1914 ();
 FILLCELL_X16 FILLER_267_1946 ();
 FILLCELL_X8 FILLER_267_1962 ();
 FILLCELL_X1 FILLER_267_1970 ();
 FILLCELL_X8 FILLER_267_1995 ();
 FILLCELL_X2 FILLER_267_2003 ();
 FILLCELL_X1 FILLER_267_2005 ();
 FILLCELL_X32 FILLER_267_2013 ();
 FILLCELL_X8 FILLER_267_2045 ();
 FILLCELL_X16 FILLER_267_2057 ();
 FILLCELL_X2 FILLER_267_2073 ();
 FILLCELL_X32 FILLER_267_2089 ();
 FILLCELL_X2 FILLER_267_2121 ();
 FILLCELL_X32 FILLER_267_2127 ();
 FILLCELL_X2 FILLER_267_2159 ();
 FILLCELL_X2 FILLER_267_2176 ();
 FILLCELL_X1 FILLER_267_2178 ();
 FILLCELL_X32 FILLER_267_2183 ();
 FILLCELL_X16 FILLER_267_2215 ();
 FILLCELL_X4 FILLER_267_2231 ();
 FILLCELL_X32 FILLER_267_2252 ();
 FILLCELL_X4 FILLER_267_2284 ();
 FILLCELL_X2 FILLER_267_2305 ();
 FILLCELL_X1 FILLER_267_2307 ();
 FILLCELL_X32 FILLER_267_2325 ();
 FILLCELL_X32 FILLER_267_2357 ();
 FILLCELL_X32 FILLER_267_2389 ();
 FILLCELL_X32 FILLER_267_2421 ();
 FILLCELL_X32 FILLER_267_2453 ();
 FILLCELL_X32 FILLER_267_2485 ();
 FILLCELL_X8 FILLER_267_2517 ();
 FILLCELL_X1 FILLER_267_2525 ();
 FILLCELL_X32 FILLER_267_2527 ();
 FILLCELL_X32 FILLER_267_2559 ();
 FILLCELL_X32 FILLER_267_2591 ();
 FILLCELL_X32 FILLER_267_2623 ();
 FILLCELL_X32 FILLER_267_2655 ();
 FILLCELL_X32 FILLER_267_2687 ();
 FILLCELL_X32 FILLER_267_2719 ();
 FILLCELL_X32 FILLER_267_2751 ();
 FILLCELL_X32 FILLER_267_2783 ();
 FILLCELL_X32 FILLER_267_2815 ();
 FILLCELL_X32 FILLER_267_2847 ();
 FILLCELL_X32 FILLER_267_2879 ();
 FILLCELL_X32 FILLER_267_2911 ();
 FILLCELL_X32 FILLER_267_2943 ();
 FILLCELL_X32 FILLER_267_2975 ();
 FILLCELL_X32 FILLER_267_3007 ();
 FILLCELL_X32 FILLER_267_3039 ();
 FILLCELL_X32 FILLER_267_3071 ();
 FILLCELL_X32 FILLER_267_3103 ();
 FILLCELL_X32 FILLER_267_3135 ();
 FILLCELL_X32 FILLER_267_3167 ();
 FILLCELL_X32 FILLER_267_3199 ();
 FILLCELL_X32 FILLER_267_3231 ();
 FILLCELL_X32 FILLER_267_3263 ();
 FILLCELL_X32 FILLER_267_3295 ();
 FILLCELL_X32 FILLER_267_3327 ();
 FILLCELL_X32 FILLER_267_3359 ();
 FILLCELL_X32 FILLER_267_3391 ();
 FILLCELL_X32 FILLER_267_3423 ();
 FILLCELL_X32 FILLER_267_3455 ();
 FILLCELL_X32 FILLER_267_3487 ();
 FILLCELL_X32 FILLER_267_3519 ();
 FILLCELL_X32 FILLER_267_3551 ();
 FILLCELL_X32 FILLER_267_3583 ();
 FILLCELL_X32 FILLER_267_3615 ();
 FILLCELL_X32 FILLER_267_3647 ();
 FILLCELL_X32 FILLER_267_3679 ();
 FILLCELL_X16 FILLER_267_3711 ();
 FILLCELL_X8 FILLER_267_3727 ();
 FILLCELL_X2 FILLER_267_3735 ();
 FILLCELL_X1 FILLER_267_3737 ();
 FILLCELL_X32 FILLER_268_1 ();
 FILLCELL_X32 FILLER_268_33 ();
 FILLCELL_X32 FILLER_268_65 ();
 FILLCELL_X32 FILLER_268_97 ();
 FILLCELL_X32 FILLER_268_129 ();
 FILLCELL_X32 FILLER_268_161 ();
 FILLCELL_X32 FILLER_268_193 ();
 FILLCELL_X32 FILLER_268_225 ();
 FILLCELL_X32 FILLER_268_257 ();
 FILLCELL_X32 FILLER_268_289 ();
 FILLCELL_X32 FILLER_268_321 ();
 FILLCELL_X32 FILLER_268_353 ();
 FILLCELL_X32 FILLER_268_385 ();
 FILLCELL_X32 FILLER_268_417 ();
 FILLCELL_X32 FILLER_268_449 ();
 FILLCELL_X32 FILLER_268_481 ();
 FILLCELL_X32 FILLER_268_513 ();
 FILLCELL_X32 FILLER_268_545 ();
 FILLCELL_X32 FILLER_268_577 ();
 FILLCELL_X16 FILLER_268_609 ();
 FILLCELL_X4 FILLER_268_625 ();
 FILLCELL_X2 FILLER_268_629 ();
 FILLCELL_X32 FILLER_268_632 ();
 FILLCELL_X32 FILLER_268_664 ();
 FILLCELL_X32 FILLER_268_696 ();
 FILLCELL_X32 FILLER_268_728 ();
 FILLCELL_X32 FILLER_268_760 ();
 FILLCELL_X32 FILLER_268_792 ();
 FILLCELL_X32 FILLER_268_824 ();
 FILLCELL_X32 FILLER_268_856 ();
 FILLCELL_X32 FILLER_268_888 ();
 FILLCELL_X32 FILLER_268_920 ();
 FILLCELL_X32 FILLER_268_952 ();
 FILLCELL_X32 FILLER_268_984 ();
 FILLCELL_X32 FILLER_268_1016 ();
 FILLCELL_X32 FILLER_268_1048 ();
 FILLCELL_X32 FILLER_268_1080 ();
 FILLCELL_X32 FILLER_268_1112 ();
 FILLCELL_X32 FILLER_268_1144 ();
 FILLCELL_X32 FILLER_268_1176 ();
 FILLCELL_X32 FILLER_268_1208 ();
 FILLCELL_X32 FILLER_268_1240 ();
 FILLCELL_X32 FILLER_268_1272 ();
 FILLCELL_X32 FILLER_268_1304 ();
 FILLCELL_X32 FILLER_268_1336 ();
 FILLCELL_X32 FILLER_268_1368 ();
 FILLCELL_X2 FILLER_268_1400 ();
 FILLCELL_X8 FILLER_268_1419 ();
 FILLCELL_X2 FILLER_268_1427 ();
 FILLCELL_X8 FILLER_268_1436 ();
 FILLCELL_X2 FILLER_268_1444 ();
 FILLCELL_X8 FILLER_268_1452 ();
 FILLCELL_X2 FILLER_268_1460 ();
 FILLCELL_X1 FILLER_268_1462 ();
 FILLCELL_X32 FILLER_268_1473 ();
 FILLCELL_X16 FILLER_268_1505 ();
 FILLCELL_X4 FILLER_268_1521 ();
 FILLCELL_X1 FILLER_268_1525 ();
 FILLCELL_X32 FILLER_268_1529 ();
 FILLCELL_X8 FILLER_268_1561 ();
 FILLCELL_X2 FILLER_268_1569 ();
 FILLCELL_X1 FILLER_268_1571 ();
 FILLCELL_X1 FILLER_268_1597 ();
 FILLCELL_X4 FILLER_268_1609 ();
 FILLCELL_X1 FILLER_268_1613 ();
 FILLCELL_X16 FILLER_268_1625 ();
 FILLCELL_X2 FILLER_268_1641 ();
 FILLCELL_X8 FILLER_268_1646 ();
 FILLCELL_X2 FILLER_268_1654 ();
 FILLCELL_X1 FILLER_268_1679 ();
 FILLCELL_X16 FILLER_268_1683 ();
 FILLCELL_X8 FILLER_268_1699 ();
 FILLCELL_X1 FILLER_268_1707 ();
 FILLCELL_X8 FILLER_268_1718 ();
 FILLCELL_X8 FILLER_268_1735 ();
 FILLCELL_X1 FILLER_268_1743 ();
 FILLCELL_X8 FILLER_268_1757 ();
 FILLCELL_X2 FILLER_268_1765 ();
 FILLCELL_X2 FILLER_268_1780 ();
 FILLCELL_X2 FILLER_268_1795 ();
 FILLCELL_X32 FILLER_268_1800 ();
 FILLCELL_X32 FILLER_268_1832 ();
 FILLCELL_X16 FILLER_268_1864 ();
 FILLCELL_X8 FILLER_268_1880 ();
 FILLCELL_X4 FILLER_268_1888 ();
 FILLCELL_X2 FILLER_268_1892 ();
 FILLCELL_X32 FILLER_268_1895 ();
 FILLCELL_X32 FILLER_268_1927 ();
 FILLCELL_X32 FILLER_268_1959 ();
 FILLCELL_X8 FILLER_268_1991 ();
 FILLCELL_X4 FILLER_268_1999 ();
 FILLCELL_X8 FILLER_268_2020 ();
 FILLCELL_X2 FILLER_268_2028 ();
 FILLCELL_X1 FILLER_268_2030 ();
 FILLCELL_X4 FILLER_268_2045 ();
 FILLCELL_X1 FILLER_268_2049 ();
 FILLCELL_X16 FILLER_268_2057 ();
 FILLCELL_X16 FILLER_268_2090 ();
 FILLCELL_X8 FILLER_268_2106 ();
 FILLCELL_X4 FILLER_268_2114 ();
 FILLCELL_X8 FILLER_268_2132 ();
 FILLCELL_X4 FILLER_268_2147 ();
 FILLCELL_X4 FILLER_268_2158 ();
 FILLCELL_X2 FILLER_268_2162 ();
 FILLCELL_X1 FILLER_268_2164 ();
 FILLCELL_X16 FILLER_268_2182 ();
 FILLCELL_X4 FILLER_268_2198 ();
 FILLCELL_X1 FILLER_268_2202 ();
 FILLCELL_X4 FILLER_268_2210 ();
 FILLCELL_X32 FILLER_268_2221 ();
 FILLCELL_X8 FILLER_268_2253 ();
 FILLCELL_X4 FILLER_268_2261 ();
 FILLCELL_X2 FILLER_268_2265 ();
 FILLCELL_X1 FILLER_268_2267 ();
 FILLCELL_X16 FILLER_268_2275 ();
 FILLCELL_X4 FILLER_268_2291 ();
 FILLCELL_X1 FILLER_268_2295 ();
 FILLCELL_X32 FILLER_268_2300 ();
 FILLCELL_X8 FILLER_268_2332 ();
 FILLCELL_X4 FILLER_268_2340 ();
 FILLCELL_X32 FILLER_268_2348 ();
 FILLCELL_X32 FILLER_268_2380 ();
 FILLCELL_X32 FILLER_268_2412 ();
 FILLCELL_X32 FILLER_268_2444 ();
 FILLCELL_X32 FILLER_268_2476 ();
 FILLCELL_X32 FILLER_268_2508 ();
 FILLCELL_X32 FILLER_268_2540 ();
 FILLCELL_X32 FILLER_268_2572 ();
 FILLCELL_X32 FILLER_268_2604 ();
 FILLCELL_X32 FILLER_268_2636 ();
 FILLCELL_X32 FILLER_268_2668 ();
 FILLCELL_X32 FILLER_268_2700 ();
 FILLCELL_X32 FILLER_268_2732 ();
 FILLCELL_X32 FILLER_268_2764 ();
 FILLCELL_X32 FILLER_268_2796 ();
 FILLCELL_X32 FILLER_268_2828 ();
 FILLCELL_X32 FILLER_268_2860 ();
 FILLCELL_X32 FILLER_268_2892 ();
 FILLCELL_X32 FILLER_268_2924 ();
 FILLCELL_X32 FILLER_268_2956 ();
 FILLCELL_X32 FILLER_268_2988 ();
 FILLCELL_X32 FILLER_268_3020 ();
 FILLCELL_X32 FILLER_268_3052 ();
 FILLCELL_X32 FILLER_268_3084 ();
 FILLCELL_X32 FILLER_268_3116 ();
 FILLCELL_X8 FILLER_268_3148 ();
 FILLCELL_X1 FILLER_268_3156 ();
 FILLCELL_X32 FILLER_268_3158 ();
 FILLCELL_X32 FILLER_268_3190 ();
 FILLCELL_X32 FILLER_268_3222 ();
 FILLCELL_X32 FILLER_268_3254 ();
 FILLCELL_X32 FILLER_268_3286 ();
 FILLCELL_X32 FILLER_268_3318 ();
 FILLCELL_X32 FILLER_268_3350 ();
 FILLCELL_X32 FILLER_268_3382 ();
 FILLCELL_X32 FILLER_268_3414 ();
 FILLCELL_X32 FILLER_268_3446 ();
 FILLCELL_X32 FILLER_268_3478 ();
 FILLCELL_X32 FILLER_268_3510 ();
 FILLCELL_X32 FILLER_268_3542 ();
 FILLCELL_X32 FILLER_268_3574 ();
 FILLCELL_X32 FILLER_268_3606 ();
 FILLCELL_X32 FILLER_268_3638 ();
 FILLCELL_X32 FILLER_268_3670 ();
 FILLCELL_X1 FILLER_268_3702 ();
 FILLCELL_X32 FILLER_268_3706 ();
 FILLCELL_X32 FILLER_269_1 ();
 FILLCELL_X32 FILLER_269_33 ();
 FILLCELL_X32 FILLER_269_65 ();
 FILLCELL_X32 FILLER_269_97 ();
 FILLCELL_X32 FILLER_269_129 ();
 FILLCELL_X32 FILLER_269_161 ();
 FILLCELL_X32 FILLER_269_193 ();
 FILLCELL_X32 FILLER_269_225 ();
 FILLCELL_X32 FILLER_269_257 ();
 FILLCELL_X32 FILLER_269_289 ();
 FILLCELL_X32 FILLER_269_321 ();
 FILLCELL_X32 FILLER_269_353 ();
 FILLCELL_X32 FILLER_269_385 ();
 FILLCELL_X32 FILLER_269_417 ();
 FILLCELL_X32 FILLER_269_449 ();
 FILLCELL_X32 FILLER_269_481 ();
 FILLCELL_X32 FILLER_269_513 ();
 FILLCELL_X32 FILLER_269_545 ();
 FILLCELL_X32 FILLER_269_577 ();
 FILLCELL_X32 FILLER_269_609 ();
 FILLCELL_X32 FILLER_269_641 ();
 FILLCELL_X32 FILLER_269_673 ();
 FILLCELL_X32 FILLER_269_705 ();
 FILLCELL_X32 FILLER_269_737 ();
 FILLCELL_X32 FILLER_269_769 ();
 FILLCELL_X32 FILLER_269_801 ();
 FILLCELL_X32 FILLER_269_833 ();
 FILLCELL_X32 FILLER_269_865 ();
 FILLCELL_X32 FILLER_269_897 ();
 FILLCELL_X32 FILLER_269_929 ();
 FILLCELL_X32 FILLER_269_961 ();
 FILLCELL_X32 FILLER_269_993 ();
 FILLCELL_X32 FILLER_269_1025 ();
 FILLCELL_X32 FILLER_269_1057 ();
 FILLCELL_X32 FILLER_269_1089 ();
 FILLCELL_X32 FILLER_269_1121 ();
 FILLCELL_X32 FILLER_269_1153 ();
 FILLCELL_X32 FILLER_269_1185 ();
 FILLCELL_X32 FILLER_269_1217 ();
 FILLCELL_X8 FILLER_269_1249 ();
 FILLCELL_X4 FILLER_269_1257 ();
 FILLCELL_X2 FILLER_269_1261 ();
 FILLCELL_X32 FILLER_269_1264 ();
 FILLCELL_X32 FILLER_269_1296 ();
 FILLCELL_X32 FILLER_269_1328 ();
 FILLCELL_X32 FILLER_269_1360 ();
 FILLCELL_X32 FILLER_269_1392 ();
 FILLCELL_X8 FILLER_269_1424 ();
 FILLCELL_X4 FILLER_269_1432 ();
 FILLCELL_X2 FILLER_269_1436 ();
 FILLCELL_X8 FILLER_269_1449 ();
 FILLCELL_X2 FILLER_269_1457 ();
 FILLCELL_X1 FILLER_269_1459 ();
 FILLCELL_X16 FILLER_269_1463 ();
 FILLCELL_X8 FILLER_269_1479 ();
 FILLCELL_X4 FILLER_269_1487 ();
 FILLCELL_X2 FILLER_269_1491 ();
 FILLCELL_X8 FILLER_269_1517 ();
 FILLCELL_X2 FILLER_269_1525 ();
 FILLCELL_X1 FILLER_269_1527 ();
 FILLCELL_X16 FILLER_269_1531 ();
 FILLCELL_X4 FILLER_269_1547 ();
 FILLCELL_X8 FILLER_269_1558 ();
 FILLCELL_X1 FILLER_269_1566 ();
 FILLCELL_X2 FILLER_269_1570 ();
 FILLCELL_X1 FILLER_269_1572 ();
 FILLCELL_X16 FILLER_269_1582 ();
 FILLCELL_X8 FILLER_269_1598 ();
 FILLCELL_X2 FILLER_269_1606 ();
 FILLCELL_X8 FILLER_269_1611 ();
 FILLCELL_X4 FILLER_269_1619 ();
 FILLCELL_X2 FILLER_269_1623 ();
 FILLCELL_X16 FILLER_269_1628 ();
 FILLCELL_X8 FILLER_269_1644 ();
 FILLCELL_X4 FILLER_269_1652 ();
 FILLCELL_X2 FILLER_269_1659 ();
 FILLCELL_X32 FILLER_269_1664 ();
 FILLCELL_X4 FILLER_269_1696 ();
 FILLCELL_X2 FILLER_269_1700 ();
 FILLCELL_X8 FILLER_269_1710 ();
 FILLCELL_X2 FILLER_269_1718 ();
 FILLCELL_X2 FILLER_269_1723 ();
 FILLCELL_X1 FILLER_269_1725 ();
 FILLCELL_X32 FILLER_269_1735 ();
 FILLCELL_X16 FILLER_269_1767 ();
 FILLCELL_X8 FILLER_269_1783 ();
 FILLCELL_X4 FILLER_269_1791 ();
 FILLCELL_X4 FILLER_269_1799 ();
 FILLCELL_X2 FILLER_269_1803 ();
 FILLCELL_X1 FILLER_269_1805 ();
 FILLCELL_X8 FILLER_269_1809 ();
 FILLCELL_X4 FILLER_269_1817 ();
 FILLCELL_X32 FILLER_269_1846 ();
 FILLCELL_X32 FILLER_269_1878 ();
 FILLCELL_X32 FILLER_269_1910 ();
 FILLCELL_X32 FILLER_269_1942 ();
 FILLCELL_X4 FILLER_269_1974 ();
 FILLCELL_X2 FILLER_269_1978 ();
 FILLCELL_X16 FILLER_269_1987 ();
 FILLCELL_X8 FILLER_269_2003 ();
 FILLCELL_X2 FILLER_269_2011 ();
 FILLCELL_X8 FILLER_269_2020 ();
 FILLCELL_X4 FILLER_269_2028 ();
 FILLCELL_X32 FILLER_269_2064 ();
 FILLCELL_X16 FILLER_269_2096 ();
 FILLCELL_X1 FILLER_269_2112 ();
 FILLCELL_X8 FILLER_269_2130 ();
 FILLCELL_X4 FILLER_269_2138 ();
 FILLCELL_X2 FILLER_269_2142 ();
 FILLCELL_X32 FILLER_269_2161 ();
 FILLCELL_X8 FILLER_269_2193 ();
 FILLCELL_X1 FILLER_269_2218 ();
 FILLCELL_X16 FILLER_269_2226 ();
 FILLCELL_X1 FILLER_269_2242 ();
 FILLCELL_X8 FILLER_269_2250 ();
 FILLCELL_X4 FILLER_269_2258 ();
 FILLCELL_X2 FILLER_269_2262 ();
 FILLCELL_X1 FILLER_269_2264 ();
 FILLCELL_X8 FILLER_269_2282 ();
 FILLCELL_X4 FILLER_269_2290 ();
 FILLCELL_X2 FILLER_269_2294 ();
 FILLCELL_X1 FILLER_269_2296 ();
 FILLCELL_X32 FILLER_269_2301 ();
 FILLCELL_X32 FILLER_269_2333 ();
 FILLCELL_X32 FILLER_269_2365 ();
 FILLCELL_X32 FILLER_269_2397 ();
 FILLCELL_X32 FILLER_269_2429 ();
 FILLCELL_X32 FILLER_269_2461 ();
 FILLCELL_X32 FILLER_269_2493 ();
 FILLCELL_X1 FILLER_269_2525 ();
 FILLCELL_X32 FILLER_269_2527 ();
 FILLCELL_X32 FILLER_269_2559 ();
 FILLCELL_X32 FILLER_269_2591 ();
 FILLCELL_X32 FILLER_269_2623 ();
 FILLCELL_X32 FILLER_269_2655 ();
 FILLCELL_X32 FILLER_269_2687 ();
 FILLCELL_X32 FILLER_269_2719 ();
 FILLCELL_X32 FILLER_269_2751 ();
 FILLCELL_X32 FILLER_269_2783 ();
 FILLCELL_X32 FILLER_269_2815 ();
 FILLCELL_X32 FILLER_269_2847 ();
 FILLCELL_X32 FILLER_269_2879 ();
 FILLCELL_X32 FILLER_269_2911 ();
 FILLCELL_X32 FILLER_269_2943 ();
 FILLCELL_X32 FILLER_269_2975 ();
 FILLCELL_X32 FILLER_269_3007 ();
 FILLCELL_X32 FILLER_269_3039 ();
 FILLCELL_X32 FILLER_269_3071 ();
 FILLCELL_X32 FILLER_269_3103 ();
 FILLCELL_X32 FILLER_269_3135 ();
 FILLCELL_X32 FILLER_269_3167 ();
 FILLCELL_X32 FILLER_269_3199 ();
 FILLCELL_X32 FILLER_269_3231 ();
 FILLCELL_X32 FILLER_269_3263 ();
 FILLCELL_X32 FILLER_269_3295 ();
 FILLCELL_X32 FILLER_269_3327 ();
 FILLCELL_X32 FILLER_269_3359 ();
 FILLCELL_X32 FILLER_269_3391 ();
 FILLCELL_X32 FILLER_269_3423 ();
 FILLCELL_X32 FILLER_269_3455 ();
 FILLCELL_X32 FILLER_269_3487 ();
 FILLCELL_X32 FILLER_269_3519 ();
 FILLCELL_X32 FILLER_269_3551 ();
 FILLCELL_X32 FILLER_269_3583 ();
 FILLCELL_X32 FILLER_269_3615 ();
 FILLCELL_X32 FILLER_269_3647 ();
 FILLCELL_X32 FILLER_269_3679 ();
 FILLCELL_X16 FILLER_269_3711 ();
 FILLCELL_X8 FILLER_269_3727 ();
 FILLCELL_X2 FILLER_269_3735 ();
 FILLCELL_X1 FILLER_269_3737 ();
 FILLCELL_X32 FILLER_270_1 ();
 FILLCELL_X32 FILLER_270_33 ();
 FILLCELL_X32 FILLER_270_65 ();
 FILLCELL_X32 FILLER_270_97 ();
 FILLCELL_X32 FILLER_270_129 ();
 FILLCELL_X32 FILLER_270_161 ();
 FILLCELL_X32 FILLER_270_193 ();
 FILLCELL_X32 FILLER_270_225 ();
 FILLCELL_X32 FILLER_270_257 ();
 FILLCELL_X32 FILLER_270_289 ();
 FILLCELL_X32 FILLER_270_321 ();
 FILLCELL_X32 FILLER_270_353 ();
 FILLCELL_X32 FILLER_270_385 ();
 FILLCELL_X32 FILLER_270_417 ();
 FILLCELL_X32 FILLER_270_449 ();
 FILLCELL_X32 FILLER_270_481 ();
 FILLCELL_X32 FILLER_270_513 ();
 FILLCELL_X32 FILLER_270_545 ();
 FILLCELL_X32 FILLER_270_577 ();
 FILLCELL_X16 FILLER_270_609 ();
 FILLCELL_X4 FILLER_270_625 ();
 FILLCELL_X2 FILLER_270_629 ();
 FILLCELL_X32 FILLER_270_632 ();
 FILLCELL_X32 FILLER_270_664 ();
 FILLCELL_X32 FILLER_270_696 ();
 FILLCELL_X32 FILLER_270_728 ();
 FILLCELL_X32 FILLER_270_760 ();
 FILLCELL_X32 FILLER_270_792 ();
 FILLCELL_X32 FILLER_270_824 ();
 FILLCELL_X32 FILLER_270_856 ();
 FILLCELL_X32 FILLER_270_888 ();
 FILLCELL_X32 FILLER_270_920 ();
 FILLCELL_X32 FILLER_270_952 ();
 FILLCELL_X32 FILLER_270_984 ();
 FILLCELL_X32 FILLER_270_1016 ();
 FILLCELL_X32 FILLER_270_1048 ();
 FILLCELL_X32 FILLER_270_1080 ();
 FILLCELL_X32 FILLER_270_1112 ();
 FILLCELL_X32 FILLER_270_1144 ();
 FILLCELL_X32 FILLER_270_1176 ();
 FILLCELL_X32 FILLER_270_1208 ();
 FILLCELL_X32 FILLER_270_1240 ();
 FILLCELL_X32 FILLER_270_1272 ();
 FILLCELL_X32 FILLER_270_1304 ();
 FILLCELL_X32 FILLER_270_1336 ();
 FILLCELL_X32 FILLER_270_1368 ();
 FILLCELL_X16 FILLER_270_1400 ();
 FILLCELL_X2 FILLER_270_1416 ();
 FILLCELL_X1 FILLER_270_1418 ();
 FILLCELL_X8 FILLER_270_1426 ();
 FILLCELL_X4 FILLER_270_1461 ();
 FILLCELL_X1 FILLER_270_1465 ();
 FILLCELL_X4 FILLER_270_1472 ();
 FILLCELL_X1 FILLER_270_1476 ();
 FILLCELL_X8 FILLER_270_1480 ();
 FILLCELL_X1 FILLER_270_1488 ();
 FILLCELL_X16 FILLER_270_1494 ();
 FILLCELL_X4 FILLER_270_1510 ();
 FILLCELL_X2 FILLER_270_1514 ();
 FILLCELL_X1 FILLER_270_1516 ();
 FILLCELL_X16 FILLER_270_1520 ();
 FILLCELL_X8 FILLER_270_1536 ();
 FILLCELL_X16 FILLER_270_1551 ();
 FILLCELL_X8 FILLER_270_1567 ();
 FILLCELL_X1 FILLER_270_1575 ();
 FILLCELL_X1 FILLER_270_1599 ();
 FILLCELL_X4 FILLER_270_1603 ();
 FILLCELL_X1 FILLER_270_1607 ();
 FILLCELL_X4 FILLER_270_1615 ();
 FILLCELL_X2 FILLER_270_1619 ();
 FILLCELL_X4 FILLER_270_1624 ();
 FILLCELL_X1 FILLER_270_1628 ();
 FILLCELL_X32 FILLER_270_1647 ();
 FILLCELL_X1 FILLER_270_1679 ();
 FILLCELL_X4 FILLER_270_1687 ();
 FILLCELL_X1 FILLER_270_1691 ();
 FILLCELL_X2 FILLER_270_1702 ();
 FILLCELL_X1 FILLER_270_1707 ();
 FILLCELL_X4 FILLER_270_1715 ();
 FILLCELL_X2 FILLER_270_1719 ();
 FILLCELL_X4 FILLER_270_1734 ();
 FILLCELL_X2 FILLER_270_1738 ();
 FILLCELL_X1 FILLER_270_1740 ();
 FILLCELL_X16 FILLER_270_1754 ();
 FILLCELL_X8 FILLER_270_1770 ();
 FILLCELL_X8 FILLER_270_1787 ();
 FILLCELL_X2 FILLER_270_1808 ();
 FILLCELL_X4 FILLER_270_1813 ();
 FILLCELL_X32 FILLER_270_1827 ();
 FILLCELL_X32 FILLER_270_1859 ();
 FILLCELL_X2 FILLER_270_1891 ();
 FILLCELL_X1 FILLER_270_1893 ();
 FILLCELL_X4 FILLER_270_1895 ();
 FILLCELL_X32 FILLER_270_1907 ();
 FILLCELL_X32 FILLER_270_1939 ();
 FILLCELL_X4 FILLER_270_1971 ();
 FILLCELL_X1 FILLER_270_1975 ();
 FILLCELL_X32 FILLER_270_1993 ();
 FILLCELL_X8 FILLER_270_2025 ();
 FILLCELL_X4 FILLER_270_2033 ();
 FILLCELL_X1 FILLER_270_2037 ();
 FILLCELL_X32 FILLER_270_2055 ();
 FILLCELL_X32 FILLER_270_2087 ();
 FILLCELL_X32 FILLER_270_2119 ();
 FILLCELL_X32 FILLER_270_2151 ();
 FILLCELL_X16 FILLER_270_2183 ();
 FILLCELL_X4 FILLER_270_2199 ();
 FILLCELL_X2 FILLER_270_2203 ();
 FILLCELL_X1 FILLER_270_2205 ();
 FILLCELL_X32 FILLER_270_2223 ();
 FILLCELL_X32 FILLER_270_2263 ();
 FILLCELL_X32 FILLER_270_2295 ();
 FILLCELL_X32 FILLER_270_2327 ();
 FILLCELL_X32 FILLER_270_2359 ();
 FILLCELL_X32 FILLER_270_2391 ();
 FILLCELL_X32 FILLER_270_2423 ();
 FILLCELL_X32 FILLER_270_2455 ();
 FILLCELL_X32 FILLER_270_2487 ();
 FILLCELL_X32 FILLER_270_2519 ();
 FILLCELL_X32 FILLER_270_2551 ();
 FILLCELL_X32 FILLER_270_2583 ();
 FILLCELL_X32 FILLER_270_2615 ();
 FILLCELL_X32 FILLER_270_2647 ();
 FILLCELL_X32 FILLER_270_2679 ();
 FILLCELL_X32 FILLER_270_2711 ();
 FILLCELL_X32 FILLER_270_2743 ();
 FILLCELL_X32 FILLER_270_2775 ();
 FILLCELL_X32 FILLER_270_2807 ();
 FILLCELL_X32 FILLER_270_2839 ();
 FILLCELL_X32 FILLER_270_2871 ();
 FILLCELL_X32 FILLER_270_2903 ();
 FILLCELL_X32 FILLER_270_2935 ();
 FILLCELL_X32 FILLER_270_2967 ();
 FILLCELL_X32 FILLER_270_2999 ();
 FILLCELL_X32 FILLER_270_3031 ();
 FILLCELL_X32 FILLER_270_3063 ();
 FILLCELL_X32 FILLER_270_3095 ();
 FILLCELL_X16 FILLER_270_3127 ();
 FILLCELL_X8 FILLER_270_3143 ();
 FILLCELL_X4 FILLER_270_3151 ();
 FILLCELL_X2 FILLER_270_3155 ();
 FILLCELL_X32 FILLER_270_3158 ();
 FILLCELL_X32 FILLER_270_3190 ();
 FILLCELL_X32 FILLER_270_3222 ();
 FILLCELL_X32 FILLER_270_3254 ();
 FILLCELL_X32 FILLER_270_3286 ();
 FILLCELL_X32 FILLER_270_3318 ();
 FILLCELL_X32 FILLER_270_3350 ();
 FILLCELL_X32 FILLER_270_3382 ();
 FILLCELL_X32 FILLER_270_3414 ();
 FILLCELL_X32 FILLER_270_3446 ();
 FILLCELL_X32 FILLER_270_3478 ();
 FILLCELL_X32 FILLER_270_3510 ();
 FILLCELL_X32 FILLER_270_3542 ();
 FILLCELL_X32 FILLER_270_3574 ();
 FILLCELL_X32 FILLER_270_3606 ();
 FILLCELL_X32 FILLER_270_3638 ();
 FILLCELL_X32 FILLER_270_3670 ();
 FILLCELL_X32 FILLER_270_3702 ();
 FILLCELL_X4 FILLER_270_3734 ();
 FILLCELL_X32 FILLER_271_1 ();
 FILLCELL_X32 FILLER_271_33 ();
 FILLCELL_X32 FILLER_271_65 ();
 FILLCELL_X32 FILLER_271_97 ();
 FILLCELL_X32 FILLER_271_129 ();
 FILLCELL_X32 FILLER_271_161 ();
 FILLCELL_X32 FILLER_271_193 ();
 FILLCELL_X32 FILLER_271_225 ();
 FILLCELL_X32 FILLER_271_257 ();
 FILLCELL_X32 FILLER_271_289 ();
 FILLCELL_X32 FILLER_271_321 ();
 FILLCELL_X32 FILLER_271_353 ();
 FILLCELL_X32 FILLER_271_385 ();
 FILLCELL_X32 FILLER_271_417 ();
 FILLCELL_X32 FILLER_271_449 ();
 FILLCELL_X32 FILLER_271_481 ();
 FILLCELL_X32 FILLER_271_513 ();
 FILLCELL_X32 FILLER_271_545 ();
 FILLCELL_X32 FILLER_271_577 ();
 FILLCELL_X32 FILLER_271_609 ();
 FILLCELL_X32 FILLER_271_641 ();
 FILLCELL_X32 FILLER_271_673 ();
 FILLCELL_X32 FILLER_271_705 ();
 FILLCELL_X32 FILLER_271_737 ();
 FILLCELL_X32 FILLER_271_769 ();
 FILLCELL_X32 FILLER_271_801 ();
 FILLCELL_X32 FILLER_271_833 ();
 FILLCELL_X32 FILLER_271_865 ();
 FILLCELL_X32 FILLER_271_897 ();
 FILLCELL_X32 FILLER_271_929 ();
 FILLCELL_X32 FILLER_271_961 ();
 FILLCELL_X32 FILLER_271_993 ();
 FILLCELL_X32 FILLER_271_1025 ();
 FILLCELL_X32 FILLER_271_1057 ();
 FILLCELL_X32 FILLER_271_1089 ();
 FILLCELL_X32 FILLER_271_1121 ();
 FILLCELL_X32 FILLER_271_1153 ();
 FILLCELL_X32 FILLER_271_1185 ();
 FILLCELL_X32 FILLER_271_1217 ();
 FILLCELL_X8 FILLER_271_1249 ();
 FILLCELL_X4 FILLER_271_1257 ();
 FILLCELL_X2 FILLER_271_1261 ();
 FILLCELL_X32 FILLER_271_1264 ();
 FILLCELL_X32 FILLER_271_1296 ();
 FILLCELL_X32 FILLER_271_1328 ();
 FILLCELL_X32 FILLER_271_1360 ();
 FILLCELL_X16 FILLER_271_1392 ();
 FILLCELL_X4 FILLER_271_1408 ();
 FILLCELL_X1 FILLER_271_1412 ();
 FILLCELL_X8 FILLER_271_1430 ();
 FILLCELL_X4 FILLER_271_1438 ();
 FILLCELL_X1 FILLER_271_1442 ();
 FILLCELL_X32 FILLER_271_1450 ();
 FILLCELL_X8 FILLER_271_1482 ();
 FILLCELL_X2 FILLER_271_1490 ();
 FILLCELL_X1 FILLER_271_1499 ();
 FILLCELL_X4 FILLER_271_1517 ();
 FILLCELL_X2 FILLER_271_1521 ();
 FILLCELL_X4 FILLER_271_1530 ();
 FILLCELL_X2 FILLER_271_1541 ();
 FILLCELL_X1 FILLER_271_1543 ();
 FILLCELL_X16 FILLER_271_1561 ();
 FILLCELL_X1 FILLER_271_1577 ();
 FILLCELL_X2 FILLER_271_1581 ();
 FILLCELL_X2 FILLER_271_1586 ();
 FILLCELL_X2 FILLER_271_1591 ();
 FILLCELL_X8 FILLER_271_1596 ();
 FILLCELL_X4 FILLER_271_1604 ();
 FILLCELL_X2 FILLER_271_1608 ();
 FILLCELL_X8 FILLER_271_1613 ();
 FILLCELL_X2 FILLER_271_1621 ();
 FILLCELL_X2 FILLER_271_1651 ();
 FILLCELL_X1 FILLER_271_1653 ();
 FILLCELL_X4 FILLER_271_1657 ();
 FILLCELL_X2 FILLER_271_1661 ();
 FILLCELL_X2 FILLER_271_1670 ();
 FILLCELL_X2 FILLER_271_1682 ();
 FILLCELL_X1 FILLER_271_1684 ();
 FILLCELL_X2 FILLER_271_1688 ();
 FILLCELL_X16 FILLER_271_1693 ();
 FILLCELL_X8 FILLER_271_1712 ();
 FILLCELL_X1 FILLER_271_1720 ();
 FILLCELL_X16 FILLER_271_1724 ();
 FILLCELL_X1 FILLER_271_1740 ();
 FILLCELL_X32 FILLER_271_1767 ();
 FILLCELL_X1 FILLER_271_1799 ();
 FILLCELL_X4 FILLER_271_1804 ();
 FILLCELL_X32 FILLER_271_1837 ();
 FILLCELL_X32 FILLER_271_1869 ();
 FILLCELL_X32 FILLER_271_1901 ();
 FILLCELL_X32 FILLER_271_1933 ();
 FILLCELL_X32 FILLER_271_1965 ();
 FILLCELL_X8 FILLER_271_1997 ();
 FILLCELL_X4 FILLER_271_2005 ();
 FILLCELL_X1 FILLER_271_2009 ();
 FILLCELL_X32 FILLER_271_2017 ();
 FILLCELL_X16 FILLER_271_2049 ();
 FILLCELL_X8 FILLER_271_2065 ();
 FILLCELL_X4 FILLER_271_2073 ();
 FILLCELL_X2 FILLER_271_2077 ();
 FILLCELL_X8 FILLER_271_2086 ();
 FILLCELL_X1 FILLER_271_2094 ();
 FILLCELL_X32 FILLER_271_2102 ();
 FILLCELL_X16 FILLER_271_2134 ();
 FILLCELL_X4 FILLER_271_2150 ();
 FILLCELL_X1 FILLER_271_2154 ();
 FILLCELL_X4 FILLER_271_2179 ();
 FILLCELL_X2 FILLER_271_2183 ();
 FILLCELL_X32 FILLER_271_2192 ();
 FILLCELL_X16 FILLER_271_2224 ();
 FILLCELL_X4 FILLER_271_2240 ();
 FILLCELL_X1 FILLER_271_2244 ();
 FILLCELL_X32 FILLER_271_2262 ();
 FILLCELL_X32 FILLER_271_2294 ();
 FILLCELL_X32 FILLER_271_2326 ();
 FILLCELL_X32 FILLER_271_2358 ();
 FILLCELL_X32 FILLER_271_2390 ();
 FILLCELL_X32 FILLER_271_2422 ();
 FILLCELL_X32 FILLER_271_2454 ();
 FILLCELL_X32 FILLER_271_2486 ();
 FILLCELL_X8 FILLER_271_2518 ();
 FILLCELL_X32 FILLER_271_2527 ();
 FILLCELL_X32 FILLER_271_2559 ();
 FILLCELL_X32 FILLER_271_2591 ();
 FILLCELL_X32 FILLER_271_2623 ();
 FILLCELL_X32 FILLER_271_2655 ();
 FILLCELL_X32 FILLER_271_2687 ();
 FILLCELL_X32 FILLER_271_2719 ();
 FILLCELL_X32 FILLER_271_2751 ();
 FILLCELL_X32 FILLER_271_2783 ();
 FILLCELL_X32 FILLER_271_2815 ();
 FILLCELL_X32 FILLER_271_2847 ();
 FILLCELL_X32 FILLER_271_2879 ();
 FILLCELL_X32 FILLER_271_2911 ();
 FILLCELL_X32 FILLER_271_2943 ();
 FILLCELL_X32 FILLER_271_2975 ();
 FILLCELL_X32 FILLER_271_3007 ();
 FILLCELL_X32 FILLER_271_3039 ();
 FILLCELL_X32 FILLER_271_3071 ();
 FILLCELL_X32 FILLER_271_3103 ();
 FILLCELL_X32 FILLER_271_3135 ();
 FILLCELL_X32 FILLER_271_3167 ();
 FILLCELL_X32 FILLER_271_3199 ();
 FILLCELL_X32 FILLER_271_3231 ();
 FILLCELL_X32 FILLER_271_3263 ();
 FILLCELL_X32 FILLER_271_3295 ();
 FILLCELL_X32 FILLER_271_3327 ();
 FILLCELL_X32 FILLER_271_3359 ();
 FILLCELL_X32 FILLER_271_3391 ();
 FILLCELL_X32 FILLER_271_3423 ();
 FILLCELL_X32 FILLER_271_3455 ();
 FILLCELL_X32 FILLER_271_3487 ();
 FILLCELL_X32 FILLER_271_3519 ();
 FILLCELL_X32 FILLER_271_3551 ();
 FILLCELL_X32 FILLER_271_3583 ();
 FILLCELL_X32 FILLER_271_3615 ();
 FILLCELL_X32 FILLER_271_3647 ();
 FILLCELL_X32 FILLER_271_3679 ();
 FILLCELL_X16 FILLER_271_3711 ();
 FILLCELL_X8 FILLER_271_3727 ();
 FILLCELL_X2 FILLER_271_3735 ();
 FILLCELL_X1 FILLER_271_3737 ();
 FILLCELL_X32 FILLER_272_1 ();
 FILLCELL_X32 FILLER_272_33 ();
 FILLCELL_X32 FILLER_272_65 ();
 FILLCELL_X32 FILLER_272_97 ();
 FILLCELL_X32 FILLER_272_129 ();
 FILLCELL_X32 FILLER_272_161 ();
 FILLCELL_X32 FILLER_272_193 ();
 FILLCELL_X32 FILLER_272_225 ();
 FILLCELL_X32 FILLER_272_257 ();
 FILLCELL_X32 FILLER_272_289 ();
 FILLCELL_X32 FILLER_272_321 ();
 FILLCELL_X32 FILLER_272_353 ();
 FILLCELL_X32 FILLER_272_385 ();
 FILLCELL_X32 FILLER_272_417 ();
 FILLCELL_X32 FILLER_272_449 ();
 FILLCELL_X32 FILLER_272_481 ();
 FILLCELL_X32 FILLER_272_513 ();
 FILLCELL_X32 FILLER_272_545 ();
 FILLCELL_X32 FILLER_272_577 ();
 FILLCELL_X16 FILLER_272_609 ();
 FILLCELL_X4 FILLER_272_625 ();
 FILLCELL_X2 FILLER_272_629 ();
 FILLCELL_X32 FILLER_272_632 ();
 FILLCELL_X32 FILLER_272_664 ();
 FILLCELL_X32 FILLER_272_696 ();
 FILLCELL_X32 FILLER_272_728 ();
 FILLCELL_X32 FILLER_272_760 ();
 FILLCELL_X32 FILLER_272_792 ();
 FILLCELL_X32 FILLER_272_824 ();
 FILLCELL_X32 FILLER_272_856 ();
 FILLCELL_X32 FILLER_272_888 ();
 FILLCELL_X32 FILLER_272_920 ();
 FILLCELL_X32 FILLER_272_952 ();
 FILLCELL_X32 FILLER_272_984 ();
 FILLCELL_X32 FILLER_272_1016 ();
 FILLCELL_X32 FILLER_272_1048 ();
 FILLCELL_X32 FILLER_272_1080 ();
 FILLCELL_X32 FILLER_272_1112 ();
 FILLCELL_X32 FILLER_272_1144 ();
 FILLCELL_X32 FILLER_272_1176 ();
 FILLCELL_X32 FILLER_272_1208 ();
 FILLCELL_X32 FILLER_272_1240 ();
 FILLCELL_X32 FILLER_272_1272 ();
 FILLCELL_X32 FILLER_272_1304 ();
 FILLCELL_X32 FILLER_272_1336 ();
 FILLCELL_X32 FILLER_272_1368 ();
 FILLCELL_X32 FILLER_272_1400 ();
 FILLCELL_X8 FILLER_272_1432 ();
 FILLCELL_X4 FILLER_272_1440 ();
 FILLCELL_X1 FILLER_272_1444 ();
 FILLCELL_X32 FILLER_272_1462 ();
 FILLCELL_X16 FILLER_272_1494 ();
 FILLCELL_X8 FILLER_272_1510 ();
 FILLCELL_X2 FILLER_272_1518 ();
 FILLCELL_X1 FILLER_272_1520 ();
 FILLCELL_X32 FILLER_272_1538 ();
 FILLCELL_X32 FILLER_272_1570 ();
 FILLCELL_X16 FILLER_272_1602 ();
 FILLCELL_X8 FILLER_272_1618 ();
 FILLCELL_X4 FILLER_272_1626 ();
 FILLCELL_X2 FILLER_272_1630 ();
 FILLCELL_X8 FILLER_272_1646 ();
 FILLCELL_X4 FILLER_272_1654 ();
 FILLCELL_X32 FILLER_272_1675 ();
 FILLCELL_X32 FILLER_272_1707 ();
 FILLCELL_X4 FILLER_272_1739 ();
 FILLCELL_X8 FILLER_272_1769 ();
 FILLCELL_X8 FILLER_272_1790 ();
 FILLCELL_X4 FILLER_272_1798 ();
 FILLCELL_X32 FILLER_272_1815 ();
 FILLCELL_X32 FILLER_272_1847 ();
 FILLCELL_X8 FILLER_272_1879 ();
 FILLCELL_X4 FILLER_272_1887 ();
 FILLCELL_X2 FILLER_272_1891 ();
 FILLCELL_X1 FILLER_272_1893 ();
 FILLCELL_X32 FILLER_272_1895 ();
 FILLCELL_X32 FILLER_272_1927 ();
 FILLCELL_X32 FILLER_272_1959 ();
 FILLCELL_X8 FILLER_272_1991 ();
 FILLCELL_X4 FILLER_272_1999 ();
 FILLCELL_X4 FILLER_272_2020 ();
 FILLCELL_X1 FILLER_272_2024 ();
 FILLCELL_X8 FILLER_272_2049 ();
 FILLCELL_X1 FILLER_272_2057 ();
 FILLCELL_X8 FILLER_272_2065 ();
 FILLCELL_X4 FILLER_272_2073 ();
 FILLCELL_X2 FILLER_272_2077 ();
 FILLCELL_X1 FILLER_272_2079 ();
 FILLCELL_X16 FILLER_272_2097 ();
 FILLCELL_X2 FILLER_272_2121 ();
 FILLCELL_X4 FILLER_272_2161 ();
 FILLCELL_X2 FILLER_272_2165 ();
 FILLCELL_X1 FILLER_272_2167 ();
 FILLCELL_X2 FILLER_272_2175 ();
 FILLCELL_X1 FILLER_272_2177 ();
 FILLCELL_X32 FILLER_272_2195 ();
 FILLCELL_X32 FILLER_272_2227 ();
 FILLCELL_X32 FILLER_272_2259 ();
 FILLCELL_X32 FILLER_272_2291 ();
 FILLCELL_X32 FILLER_272_2323 ();
 FILLCELL_X32 FILLER_272_2355 ();
 FILLCELL_X32 FILLER_272_2387 ();
 FILLCELL_X32 FILLER_272_2419 ();
 FILLCELL_X32 FILLER_272_2451 ();
 FILLCELL_X32 FILLER_272_2483 ();
 FILLCELL_X32 FILLER_272_2515 ();
 FILLCELL_X32 FILLER_272_2547 ();
 FILLCELL_X32 FILLER_272_2579 ();
 FILLCELL_X32 FILLER_272_2611 ();
 FILLCELL_X32 FILLER_272_2643 ();
 FILLCELL_X32 FILLER_272_2675 ();
 FILLCELL_X32 FILLER_272_2707 ();
 FILLCELL_X32 FILLER_272_2739 ();
 FILLCELL_X32 FILLER_272_2771 ();
 FILLCELL_X32 FILLER_272_2803 ();
 FILLCELL_X32 FILLER_272_2835 ();
 FILLCELL_X32 FILLER_272_2867 ();
 FILLCELL_X32 FILLER_272_2899 ();
 FILLCELL_X32 FILLER_272_2931 ();
 FILLCELL_X32 FILLER_272_2963 ();
 FILLCELL_X32 FILLER_272_2995 ();
 FILLCELL_X32 FILLER_272_3027 ();
 FILLCELL_X32 FILLER_272_3059 ();
 FILLCELL_X32 FILLER_272_3091 ();
 FILLCELL_X32 FILLER_272_3123 ();
 FILLCELL_X2 FILLER_272_3155 ();
 FILLCELL_X32 FILLER_272_3158 ();
 FILLCELL_X32 FILLER_272_3190 ();
 FILLCELL_X32 FILLER_272_3222 ();
 FILLCELL_X32 FILLER_272_3254 ();
 FILLCELL_X32 FILLER_272_3286 ();
 FILLCELL_X32 FILLER_272_3318 ();
 FILLCELL_X32 FILLER_272_3350 ();
 FILLCELL_X32 FILLER_272_3382 ();
 FILLCELL_X32 FILLER_272_3414 ();
 FILLCELL_X32 FILLER_272_3446 ();
 FILLCELL_X32 FILLER_272_3478 ();
 FILLCELL_X32 FILLER_272_3510 ();
 FILLCELL_X32 FILLER_272_3542 ();
 FILLCELL_X32 FILLER_272_3574 ();
 FILLCELL_X32 FILLER_272_3606 ();
 FILLCELL_X32 FILLER_272_3638 ();
 FILLCELL_X32 FILLER_272_3670 ();
 FILLCELL_X32 FILLER_272_3702 ();
 FILLCELL_X4 FILLER_272_3734 ();
 FILLCELL_X32 FILLER_273_1 ();
 FILLCELL_X32 FILLER_273_33 ();
 FILLCELL_X32 FILLER_273_65 ();
 FILLCELL_X32 FILLER_273_97 ();
 FILLCELL_X32 FILLER_273_129 ();
 FILLCELL_X32 FILLER_273_161 ();
 FILLCELL_X32 FILLER_273_193 ();
 FILLCELL_X32 FILLER_273_225 ();
 FILLCELL_X32 FILLER_273_257 ();
 FILLCELL_X32 FILLER_273_289 ();
 FILLCELL_X32 FILLER_273_321 ();
 FILLCELL_X32 FILLER_273_353 ();
 FILLCELL_X32 FILLER_273_385 ();
 FILLCELL_X32 FILLER_273_417 ();
 FILLCELL_X32 FILLER_273_449 ();
 FILLCELL_X32 FILLER_273_481 ();
 FILLCELL_X32 FILLER_273_513 ();
 FILLCELL_X32 FILLER_273_545 ();
 FILLCELL_X32 FILLER_273_577 ();
 FILLCELL_X32 FILLER_273_609 ();
 FILLCELL_X32 FILLER_273_641 ();
 FILLCELL_X32 FILLER_273_673 ();
 FILLCELL_X32 FILLER_273_705 ();
 FILLCELL_X32 FILLER_273_737 ();
 FILLCELL_X32 FILLER_273_769 ();
 FILLCELL_X32 FILLER_273_801 ();
 FILLCELL_X32 FILLER_273_833 ();
 FILLCELL_X32 FILLER_273_865 ();
 FILLCELL_X32 FILLER_273_897 ();
 FILLCELL_X32 FILLER_273_929 ();
 FILLCELL_X32 FILLER_273_961 ();
 FILLCELL_X32 FILLER_273_993 ();
 FILLCELL_X32 FILLER_273_1025 ();
 FILLCELL_X32 FILLER_273_1057 ();
 FILLCELL_X32 FILLER_273_1089 ();
 FILLCELL_X32 FILLER_273_1121 ();
 FILLCELL_X32 FILLER_273_1153 ();
 FILLCELL_X32 FILLER_273_1185 ();
 FILLCELL_X32 FILLER_273_1217 ();
 FILLCELL_X8 FILLER_273_1249 ();
 FILLCELL_X4 FILLER_273_1257 ();
 FILLCELL_X2 FILLER_273_1261 ();
 FILLCELL_X32 FILLER_273_1264 ();
 FILLCELL_X32 FILLER_273_1296 ();
 FILLCELL_X32 FILLER_273_1328 ();
 FILLCELL_X8 FILLER_273_1360 ();
 FILLCELL_X4 FILLER_273_1368 ();
 FILLCELL_X16 FILLER_273_1376 ();
 FILLCELL_X2 FILLER_273_1392 ();
 FILLCELL_X1 FILLER_273_1394 ();
 FILLCELL_X16 FILLER_273_1399 ();
 FILLCELL_X2 FILLER_273_1415 ();
 FILLCELL_X16 FILLER_273_1431 ();
 FILLCELL_X16 FILLER_273_1458 ();
 FILLCELL_X8 FILLER_273_1474 ();
 FILLCELL_X4 FILLER_273_1482 ();
 FILLCELL_X32 FILLER_273_1510 ();
 FILLCELL_X8 FILLER_273_1542 ();
 FILLCELL_X32 FILLER_273_1557 ();
 FILLCELL_X16 FILLER_273_1589 ();
 FILLCELL_X4 FILLER_273_1605 ();
 FILLCELL_X1 FILLER_273_1609 ();
 FILLCELL_X32 FILLER_273_1617 ();
 FILLCELL_X32 FILLER_273_1649 ();
 FILLCELL_X8 FILLER_273_1681 ();
 FILLCELL_X4 FILLER_273_1689 ();
 FILLCELL_X2 FILLER_273_1693 ();
 FILLCELL_X8 FILLER_273_1709 ();
 FILLCELL_X1 FILLER_273_1717 ();
 FILLCELL_X32 FILLER_273_1725 ();
 FILLCELL_X32 FILLER_273_1757 ();
 FILLCELL_X32 FILLER_273_1789 ();
 FILLCELL_X32 FILLER_273_1821 ();
 FILLCELL_X32 FILLER_273_1853 ();
 FILLCELL_X32 FILLER_273_1885 ();
 FILLCELL_X32 FILLER_273_1917 ();
 FILLCELL_X32 FILLER_273_1949 ();
 FILLCELL_X32 FILLER_273_1981 ();
 FILLCELL_X32 FILLER_273_2013 ();
 FILLCELL_X16 FILLER_273_2069 ();
 FILLCELL_X4 FILLER_273_2085 ();
 FILLCELL_X1 FILLER_273_2089 ();
 FILLCELL_X16 FILLER_273_2097 ();
 FILLCELL_X2 FILLER_273_2113 ();
 FILLCELL_X32 FILLER_273_2132 ();
 FILLCELL_X32 FILLER_273_2164 ();
 FILLCELL_X32 FILLER_273_2196 ();
 FILLCELL_X32 FILLER_273_2228 ();
 FILLCELL_X32 FILLER_273_2260 ();
 FILLCELL_X32 FILLER_273_2292 ();
 FILLCELL_X32 FILLER_273_2324 ();
 FILLCELL_X32 FILLER_273_2356 ();
 FILLCELL_X32 FILLER_273_2388 ();
 FILLCELL_X32 FILLER_273_2420 ();
 FILLCELL_X32 FILLER_273_2452 ();
 FILLCELL_X32 FILLER_273_2484 ();
 FILLCELL_X8 FILLER_273_2516 ();
 FILLCELL_X2 FILLER_273_2524 ();
 FILLCELL_X32 FILLER_273_2527 ();
 FILLCELL_X32 FILLER_273_2559 ();
 FILLCELL_X32 FILLER_273_2591 ();
 FILLCELL_X32 FILLER_273_2623 ();
 FILLCELL_X32 FILLER_273_2655 ();
 FILLCELL_X32 FILLER_273_2687 ();
 FILLCELL_X32 FILLER_273_2719 ();
 FILLCELL_X32 FILLER_273_2751 ();
 FILLCELL_X32 FILLER_273_2783 ();
 FILLCELL_X32 FILLER_273_2815 ();
 FILLCELL_X32 FILLER_273_2847 ();
 FILLCELL_X32 FILLER_273_2879 ();
 FILLCELL_X32 FILLER_273_2911 ();
 FILLCELL_X32 FILLER_273_2943 ();
 FILLCELL_X32 FILLER_273_2975 ();
 FILLCELL_X32 FILLER_273_3007 ();
 FILLCELL_X32 FILLER_273_3039 ();
 FILLCELL_X32 FILLER_273_3071 ();
 FILLCELL_X32 FILLER_273_3103 ();
 FILLCELL_X32 FILLER_273_3135 ();
 FILLCELL_X32 FILLER_273_3167 ();
 FILLCELL_X32 FILLER_273_3199 ();
 FILLCELL_X32 FILLER_273_3231 ();
 FILLCELL_X32 FILLER_273_3263 ();
 FILLCELL_X32 FILLER_273_3295 ();
 FILLCELL_X32 FILLER_273_3327 ();
 FILLCELL_X32 FILLER_273_3359 ();
 FILLCELL_X32 FILLER_273_3391 ();
 FILLCELL_X32 FILLER_273_3423 ();
 FILLCELL_X32 FILLER_273_3455 ();
 FILLCELL_X32 FILLER_273_3487 ();
 FILLCELL_X32 FILLER_273_3519 ();
 FILLCELL_X32 FILLER_273_3551 ();
 FILLCELL_X32 FILLER_273_3583 ();
 FILLCELL_X32 FILLER_273_3615 ();
 FILLCELL_X32 FILLER_273_3647 ();
 FILLCELL_X32 FILLER_273_3679 ();
 FILLCELL_X16 FILLER_273_3711 ();
 FILLCELL_X8 FILLER_273_3727 ();
 FILLCELL_X2 FILLER_273_3735 ();
 FILLCELL_X1 FILLER_273_3737 ();
 FILLCELL_X32 FILLER_274_1 ();
 FILLCELL_X32 FILLER_274_33 ();
 FILLCELL_X32 FILLER_274_65 ();
 FILLCELL_X32 FILLER_274_97 ();
 FILLCELL_X32 FILLER_274_129 ();
 FILLCELL_X32 FILLER_274_161 ();
 FILLCELL_X32 FILLER_274_193 ();
 FILLCELL_X32 FILLER_274_225 ();
 FILLCELL_X32 FILLER_274_257 ();
 FILLCELL_X32 FILLER_274_289 ();
 FILLCELL_X32 FILLER_274_321 ();
 FILLCELL_X32 FILLER_274_353 ();
 FILLCELL_X32 FILLER_274_385 ();
 FILLCELL_X32 FILLER_274_417 ();
 FILLCELL_X32 FILLER_274_449 ();
 FILLCELL_X32 FILLER_274_481 ();
 FILLCELL_X32 FILLER_274_513 ();
 FILLCELL_X32 FILLER_274_545 ();
 FILLCELL_X32 FILLER_274_577 ();
 FILLCELL_X16 FILLER_274_609 ();
 FILLCELL_X4 FILLER_274_625 ();
 FILLCELL_X2 FILLER_274_629 ();
 FILLCELL_X32 FILLER_274_632 ();
 FILLCELL_X32 FILLER_274_664 ();
 FILLCELL_X32 FILLER_274_696 ();
 FILLCELL_X32 FILLER_274_728 ();
 FILLCELL_X32 FILLER_274_760 ();
 FILLCELL_X32 FILLER_274_792 ();
 FILLCELL_X32 FILLER_274_824 ();
 FILLCELL_X32 FILLER_274_856 ();
 FILLCELL_X32 FILLER_274_888 ();
 FILLCELL_X32 FILLER_274_920 ();
 FILLCELL_X32 FILLER_274_952 ();
 FILLCELL_X32 FILLER_274_984 ();
 FILLCELL_X32 FILLER_274_1016 ();
 FILLCELL_X32 FILLER_274_1048 ();
 FILLCELL_X32 FILLER_274_1080 ();
 FILLCELL_X32 FILLER_274_1112 ();
 FILLCELL_X32 FILLER_274_1144 ();
 FILLCELL_X32 FILLER_274_1176 ();
 FILLCELL_X32 FILLER_274_1208 ();
 FILLCELL_X32 FILLER_274_1240 ();
 FILLCELL_X32 FILLER_274_1272 ();
 FILLCELL_X32 FILLER_274_1304 ();
 FILLCELL_X32 FILLER_274_1336 ();
 FILLCELL_X32 FILLER_274_1368 ();
 FILLCELL_X8 FILLER_274_1400 ();
 FILLCELL_X4 FILLER_274_1408 ();
 FILLCELL_X1 FILLER_274_1412 ();
 FILLCELL_X32 FILLER_274_1430 ();
 FILLCELL_X16 FILLER_274_1462 ();
 FILLCELL_X4 FILLER_274_1478 ();
 FILLCELL_X16 FILLER_274_1489 ();
 FILLCELL_X1 FILLER_274_1505 ();
 FILLCELL_X16 FILLER_274_1513 ();
 FILLCELL_X8 FILLER_274_1529 ();
 FILLCELL_X4 FILLER_274_1537 ();
 FILLCELL_X2 FILLER_274_1541 ();
 FILLCELL_X1 FILLER_274_1543 ();
 FILLCELL_X8 FILLER_274_1551 ();
 FILLCELL_X2 FILLER_274_1559 ();
 FILLCELL_X1 FILLER_274_1561 ();
 FILLCELL_X4 FILLER_274_1569 ();
 FILLCELL_X1 FILLER_274_1573 ();
 FILLCELL_X16 FILLER_274_1581 ();
 FILLCELL_X8 FILLER_274_1597 ();
 FILLCELL_X2 FILLER_274_1605 ();
 FILLCELL_X16 FILLER_274_1624 ();
 FILLCELL_X2 FILLER_274_1640 ();
 FILLCELL_X16 FILLER_274_1649 ();
 FILLCELL_X4 FILLER_274_1665 ();
 FILLCELL_X1 FILLER_274_1669 ();
 FILLCELL_X16 FILLER_274_1677 ();
 FILLCELL_X4 FILLER_274_1693 ();
 FILLCELL_X1 FILLER_274_1697 ();
 FILLCELL_X2 FILLER_274_1715 ();
 FILLCELL_X32 FILLER_274_1734 ();
 FILLCELL_X32 FILLER_274_1766 ();
 FILLCELL_X32 FILLER_274_1798 ();
 FILLCELL_X32 FILLER_274_1830 ();
 FILLCELL_X32 FILLER_274_1862 ();
 FILLCELL_X32 FILLER_274_1895 ();
 FILLCELL_X32 FILLER_274_1927 ();
 FILLCELL_X32 FILLER_274_1959 ();
 FILLCELL_X32 FILLER_274_1991 ();
 FILLCELL_X32 FILLER_274_2023 ();
 FILLCELL_X32 FILLER_274_2055 ();
 FILLCELL_X4 FILLER_274_2087 ();
 FILLCELL_X32 FILLER_274_2108 ();
 FILLCELL_X32 FILLER_274_2140 ();
 FILLCELL_X32 FILLER_274_2172 ();
 FILLCELL_X32 FILLER_274_2204 ();
 FILLCELL_X32 FILLER_274_2236 ();
 FILLCELL_X32 FILLER_274_2268 ();
 FILLCELL_X32 FILLER_274_2300 ();
 FILLCELL_X32 FILLER_274_2332 ();
 FILLCELL_X32 FILLER_274_2364 ();
 FILLCELL_X32 FILLER_274_2396 ();
 FILLCELL_X32 FILLER_274_2428 ();
 FILLCELL_X32 FILLER_274_2460 ();
 FILLCELL_X32 FILLER_274_2492 ();
 FILLCELL_X32 FILLER_274_2524 ();
 FILLCELL_X32 FILLER_274_2556 ();
 FILLCELL_X32 FILLER_274_2588 ();
 FILLCELL_X32 FILLER_274_2620 ();
 FILLCELL_X32 FILLER_274_2652 ();
 FILLCELL_X32 FILLER_274_2684 ();
 FILLCELL_X32 FILLER_274_2716 ();
 FILLCELL_X32 FILLER_274_2748 ();
 FILLCELL_X32 FILLER_274_2780 ();
 FILLCELL_X32 FILLER_274_2812 ();
 FILLCELL_X32 FILLER_274_2844 ();
 FILLCELL_X32 FILLER_274_2876 ();
 FILLCELL_X32 FILLER_274_2908 ();
 FILLCELL_X32 FILLER_274_2940 ();
 FILLCELL_X32 FILLER_274_2972 ();
 FILLCELL_X32 FILLER_274_3004 ();
 FILLCELL_X32 FILLER_274_3036 ();
 FILLCELL_X32 FILLER_274_3068 ();
 FILLCELL_X32 FILLER_274_3100 ();
 FILLCELL_X16 FILLER_274_3132 ();
 FILLCELL_X8 FILLER_274_3148 ();
 FILLCELL_X1 FILLER_274_3156 ();
 FILLCELL_X32 FILLER_274_3158 ();
 FILLCELL_X32 FILLER_274_3190 ();
 FILLCELL_X32 FILLER_274_3222 ();
 FILLCELL_X32 FILLER_274_3254 ();
 FILLCELL_X32 FILLER_274_3286 ();
 FILLCELL_X32 FILLER_274_3318 ();
 FILLCELL_X32 FILLER_274_3350 ();
 FILLCELL_X32 FILLER_274_3382 ();
 FILLCELL_X32 FILLER_274_3414 ();
 FILLCELL_X32 FILLER_274_3446 ();
 FILLCELL_X32 FILLER_274_3478 ();
 FILLCELL_X32 FILLER_274_3510 ();
 FILLCELL_X32 FILLER_274_3542 ();
 FILLCELL_X32 FILLER_274_3574 ();
 FILLCELL_X32 FILLER_274_3606 ();
 FILLCELL_X32 FILLER_274_3638 ();
 FILLCELL_X32 FILLER_274_3670 ();
 FILLCELL_X32 FILLER_274_3702 ();
 FILLCELL_X4 FILLER_274_3734 ();
 FILLCELL_X32 FILLER_275_1 ();
 FILLCELL_X32 FILLER_275_33 ();
 FILLCELL_X32 FILLER_275_65 ();
 FILLCELL_X32 FILLER_275_97 ();
 FILLCELL_X32 FILLER_275_129 ();
 FILLCELL_X32 FILLER_275_161 ();
 FILLCELL_X32 FILLER_275_193 ();
 FILLCELL_X32 FILLER_275_225 ();
 FILLCELL_X32 FILLER_275_257 ();
 FILLCELL_X32 FILLER_275_289 ();
 FILLCELL_X32 FILLER_275_321 ();
 FILLCELL_X32 FILLER_275_353 ();
 FILLCELL_X32 FILLER_275_385 ();
 FILLCELL_X32 FILLER_275_417 ();
 FILLCELL_X32 FILLER_275_449 ();
 FILLCELL_X32 FILLER_275_481 ();
 FILLCELL_X32 FILLER_275_513 ();
 FILLCELL_X32 FILLER_275_545 ();
 FILLCELL_X32 FILLER_275_577 ();
 FILLCELL_X32 FILLER_275_609 ();
 FILLCELL_X32 FILLER_275_641 ();
 FILLCELL_X32 FILLER_275_673 ();
 FILLCELL_X32 FILLER_275_705 ();
 FILLCELL_X32 FILLER_275_737 ();
 FILLCELL_X32 FILLER_275_769 ();
 FILLCELL_X32 FILLER_275_801 ();
 FILLCELL_X32 FILLER_275_833 ();
 FILLCELL_X32 FILLER_275_865 ();
 FILLCELL_X32 FILLER_275_897 ();
 FILLCELL_X32 FILLER_275_929 ();
 FILLCELL_X32 FILLER_275_961 ();
 FILLCELL_X32 FILLER_275_993 ();
 FILLCELL_X32 FILLER_275_1025 ();
 FILLCELL_X32 FILLER_275_1057 ();
 FILLCELL_X32 FILLER_275_1089 ();
 FILLCELL_X32 FILLER_275_1121 ();
 FILLCELL_X32 FILLER_275_1153 ();
 FILLCELL_X32 FILLER_275_1185 ();
 FILLCELL_X32 FILLER_275_1217 ();
 FILLCELL_X8 FILLER_275_1249 ();
 FILLCELL_X4 FILLER_275_1257 ();
 FILLCELL_X2 FILLER_275_1261 ();
 FILLCELL_X32 FILLER_275_1264 ();
 FILLCELL_X32 FILLER_275_1296 ();
 FILLCELL_X32 FILLER_275_1328 ();
 FILLCELL_X32 FILLER_275_1360 ();
 FILLCELL_X16 FILLER_275_1392 ();
 FILLCELL_X2 FILLER_275_1408 ();
 FILLCELL_X16 FILLER_275_1434 ();
 FILLCELL_X4 FILLER_275_1450 ();
 FILLCELL_X16 FILLER_275_1461 ();
 FILLCELL_X2 FILLER_275_1477 ();
 FILLCELL_X8 FILLER_275_1486 ();
 FILLCELL_X4 FILLER_275_1494 ();
 FILLCELL_X1 FILLER_275_1498 ();
 FILLCELL_X8 FILLER_275_1523 ();
 FILLCELL_X4 FILLER_275_1531 ();
 FILLCELL_X1 FILLER_275_1535 ();
 FILLCELL_X4 FILLER_275_1553 ();
 FILLCELL_X2 FILLER_275_1557 ();
 FILLCELL_X16 FILLER_275_1600 ();
 FILLCELL_X2 FILLER_275_1616 ();
 FILLCELL_X8 FILLER_275_1625 ();
 FILLCELL_X4 FILLER_275_1633 ();
 FILLCELL_X2 FILLER_275_1637 ();
 FILLCELL_X1 FILLER_275_1639 ();
 FILLCELL_X8 FILLER_275_1657 ();
 FILLCELL_X2 FILLER_275_1665 ();
 FILLCELL_X1 FILLER_275_1667 ();
 FILLCELL_X16 FILLER_275_1685 ();
 FILLCELL_X4 FILLER_275_1701 ();
 FILLCELL_X2 FILLER_275_1705 ();
 FILLCELL_X1 FILLER_275_1707 ();
 FILLCELL_X32 FILLER_275_1713 ();
 FILLCELL_X32 FILLER_275_1745 ();
 FILLCELL_X16 FILLER_275_1777 ();
 FILLCELL_X1 FILLER_275_1793 ();
 FILLCELL_X32 FILLER_275_1798 ();
 FILLCELL_X32 FILLER_275_1830 ();
 FILLCELL_X32 FILLER_275_1862 ();
 FILLCELL_X32 FILLER_275_1894 ();
 FILLCELL_X32 FILLER_275_1926 ();
 FILLCELL_X32 FILLER_275_1958 ();
 FILLCELL_X32 FILLER_275_1990 ();
 FILLCELL_X32 FILLER_275_2022 ();
 FILLCELL_X32 FILLER_275_2054 ();
 FILLCELL_X32 FILLER_275_2086 ();
 FILLCELL_X32 FILLER_275_2118 ();
 FILLCELL_X32 FILLER_275_2150 ();
 FILLCELL_X32 FILLER_275_2182 ();
 FILLCELL_X32 FILLER_275_2214 ();
 FILLCELL_X32 FILLER_275_2246 ();
 FILLCELL_X32 FILLER_275_2278 ();
 FILLCELL_X32 FILLER_275_2310 ();
 FILLCELL_X32 FILLER_275_2342 ();
 FILLCELL_X32 FILLER_275_2374 ();
 FILLCELL_X32 FILLER_275_2406 ();
 FILLCELL_X32 FILLER_275_2438 ();
 FILLCELL_X32 FILLER_275_2470 ();
 FILLCELL_X16 FILLER_275_2502 ();
 FILLCELL_X8 FILLER_275_2518 ();
 FILLCELL_X32 FILLER_275_2527 ();
 FILLCELL_X32 FILLER_275_2559 ();
 FILLCELL_X32 FILLER_275_2591 ();
 FILLCELL_X32 FILLER_275_2623 ();
 FILLCELL_X32 FILLER_275_2655 ();
 FILLCELL_X32 FILLER_275_2687 ();
 FILLCELL_X32 FILLER_275_2719 ();
 FILLCELL_X32 FILLER_275_2751 ();
 FILLCELL_X32 FILLER_275_2783 ();
 FILLCELL_X32 FILLER_275_2815 ();
 FILLCELL_X32 FILLER_275_2847 ();
 FILLCELL_X32 FILLER_275_2879 ();
 FILLCELL_X32 FILLER_275_2911 ();
 FILLCELL_X32 FILLER_275_2943 ();
 FILLCELL_X32 FILLER_275_2975 ();
 FILLCELL_X32 FILLER_275_3007 ();
 FILLCELL_X32 FILLER_275_3039 ();
 FILLCELL_X32 FILLER_275_3071 ();
 FILLCELL_X32 FILLER_275_3103 ();
 FILLCELL_X32 FILLER_275_3135 ();
 FILLCELL_X32 FILLER_275_3167 ();
 FILLCELL_X32 FILLER_275_3199 ();
 FILLCELL_X32 FILLER_275_3231 ();
 FILLCELL_X32 FILLER_275_3263 ();
 FILLCELL_X32 FILLER_275_3295 ();
 FILLCELL_X32 FILLER_275_3327 ();
 FILLCELL_X32 FILLER_275_3359 ();
 FILLCELL_X32 FILLER_275_3391 ();
 FILLCELL_X32 FILLER_275_3423 ();
 FILLCELL_X32 FILLER_275_3455 ();
 FILLCELL_X32 FILLER_275_3487 ();
 FILLCELL_X32 FILLER_275_3519 ();
 FILLCELL_X32 FILLER_275_3551 ();
 FILLCELL_X32 FILLER_275_3583 ();
 FILLCELL_X32 FILLER_275_3615 ();
 FILLCELL_X32 FILLER_275_3647 ();
 FILLCELL_X32 FILLER_275_3679 ();
 FILLCELL_X16 FILLER_275_3711 ();
 FILLCELL_X8 FILLER_275_3727 ();
 FILLCELL_X2 FILLER_275_3735 ();
 FILLCELL_X1 FILLER_275_3737 ();
 FILLCELL_X32 FILLER_276_1 ();
 FILLCELL_X32 FILLER_276_33 ();
 FILLCELL_X32 FILLER_276_65 ();
 FILLCELL_X32 FILLER_276_97 ();
 FILLCELL_X32 FILLER_276_129 ();
 FILLCELL_X32 FILLER_276_161 ();
 FILLCELL_X32 FILLER_276_193 ();
 FILLCELL_X32 FILLER_276_225 ();
 FILLCELL_X32 FILLER_276_257 ();
 FILLCELL_X32 FILLER_276_289 ();
 FILLCELL_X32 FILLER_276_321 ();
 FILLCELL_X32 FILLER_276_353 ();
 FILLCELL_X32 FILLER_276_385 ();
 FILLCELL_X32 FILLER_276_417 ();
 FILLCELL_X32 FILLER_276_449 ();
 FILLCELL_X32 FILLER_276_481 ();
 FILLCELL_X32 FILLER_276_513 ();
 FILLCELL_X32 FILLER_276_545 ();
 FILLCELL_X32 FILLER_276_577 ();
 FILLCELL_X16 FILLER_276_609 ();
 FILLCELL_X4 FILLER_276_625 ();
 FILLCELL_X2 FILLER_276_629 ();
 FILLCELL_X32 FILLER_276_632 ();
 FILLCELL_X32 FILLER_276_664 ();
 FILLCELL_X32 FILLER_276_696 ();
 FILLCELL_X32 FILLER_276_728 ();
 FILLCELL_X32 FILLER_276_760 ();
 FILLCELL_X32 FILLER_276_792 ();
 FILLCELL_X32 FILLER_276_824 ();
 FILLCELL_X32 FILLER_276_856 ();
 FILLCELL_X32 FILLER_276_888 ();
 FILLCELL_X32 FILLER_276_920 ();
 FILLCELL_X32 FILLER_276_952 ();
 FILLCELL_X32 FILLER_276_984 ();
 FILLCELL_X32 FILLER_276_1016 ();
 FILLCELL_X32 FILLER_276_1048 ();
 FILLCELL_X32 FILLER_276_1080 ();
 FILLCELL_X32 FILLER_276_1112 ();
 FILLCELL_X32 FILLER_276_1144 ();
 FILLCELL_X32 FILLER_276_1176 ();
 FILLCELL_X32 FILLER_276_1208 ();
 FILLCELL_X32 FILLER_276_1240 ();
 FILLCELL_X32 FILLER_276_1272 ();
 FILLCELL_X32 FILLER_276_1304 ();
 FILLCELL_X32 FILLER_276_1336 ();
 FILLCELL_X32 FILLER_276_1368 ();
 FILLCELL_X32 FILLER_276_1400 ();
 FILLCELL_X4 FILLER_276_1432 ();
 FILLCELL_X1 FILLER_276_1436 ();
 FILLCELL_X8 FILLER_276_1444 ();
 FILLCELL_X2 FILLER_276_1452 ();
 FILLCELL_X16 FILLER_276_1461 ();
 FILLCELL_X1 FILLER_276_1477 ();
 FILLCELL_X32 FILLER_276_1495 ();
 FILLCELL_X16 FILLER_276_1527 ();
 FILLCELL_X4 FILLER_276_1543 ();
 FILLCELL_X1 FILLER_276_1547 ();
 FILLCELL_X4 FILLER_276_1555 ();
 FILLCELL_X4 FILLER_276_1566 ();
 FILLCELL_X1 FILLER_276_1570 ();
 FILLCELL_X16 FILLER_276_1579 ();
 FILLCELL_X2 FILLER_276_1595 ();
 FILLCELL_X32 FILLER_276_1621 ();
 FILLCELL_X32 FILLER_276_1653 ();
 FILLCELL_X16 FILLER_276_1685 ();
 FILLCELL_X1 FILLER_276_1701 ();
 FILLCELL_X8 FILLER_276_1728 ();
 FILLCELL_X4 FILLER_276_1736 ();
 FILLCELL_X2 FILLER_276_1740 ();
 FILLCELL_X32 FILLER_276_1766 ();
 FILLCELL_X32 FILLER_276_1798 ();
 FILLCELL_X32 FILLER_276_1830 ();
 FILLCELL_X32 FILLER_276_1862 ();
 FILLCELL_X32 FILLER_276_1895 ();
 FILLCELL_X32 FILLER_276_1927 ();
 FILLCELL_X32 FILLER_276_1959 ();
 FILLCELL_X32 FILLER_276_1991 ();
 FILLCELL_X32 FILLER_276_2023 ();
 FILLCELL_X32 FILLER_276_2055 ();
 FILLCELL_X32 FILLER_276_2087 ();
 FILLCELL_X32 FILLER_276_2119 ();
 FILLCELL_X32 FILLER_276_2151 ();
 FILLCELL_X32 FILLER_276_2183 ();
 FILLCELL_X32 FILLER_276_2215 ();
 FILLCELL_X32 FILLER_276_2247 ();
 FILLCELL_X32 FILLER_276_2279 ();
 FILLCELL_X32 FILLER_276_2311 ();
 FILLCELL_X32 FILLER_276_2343 ();
 FILLCELL_X32 FILLER_276_2375 ();
 FILLCELL_X32 FILLER_276_2407 ();
 FILLCELL_X32 FILLER_276_2439 ();
 FILLCELL_X32 FILLER_276_2471 ();
 FILLCELL_X32 FILLER_276_2503 ();
 FILLCELL_X32 FILLER_276_2535 ();
 FILLCELL_X32 FILLER_276_2567 ();
 FILLCELL_X32 FILLER_276_2599 ();
 FILLCELL_X32 FILLER_276_2631 ();
 FILLCELL_X32 FILLER_276_2663 ();
 FILLCELL_X32 FILLER_276_2695 ();
 FILLCELL_X32 FILLER_276_2727 ();
 FILLCELL_X32 FILLER_276_2759 ();
 FILLCELL_X32 FILLER_276_2791 ();
 FILLCELL_X32 FILLER_276_2823 ();
 FILLCELL_X32 FILLER_276_2855 ();
 FILLCELL_X32 FILLER_276_2887 ();
 FILLCELL_X32 FILLER_276_2919 ();
 FILLCELL_X32 FILLER_276_2951 ();
 FILLCELL_X32 FILLER_276_2983 ();
 FILLCELL_X32 FILLER_276_3015 ();
 FILLCELL_X32 FILLER_276_3047 ();
 FILLCELL_X32 FILLER_276_3079 ();
 FILLCELL_X32 FILLER_276_3111 ();
 FILLCELL_X8 FILLER_276_3143 ();
 FILLCELL_X4 FILLER_276_3151 ();
 FILLCELL_X2 FILLER_276_3155 ();
 FILLCELL_X32 FILLER_276_3158 ();
 FILLCELL_X32 FILLER_276_3190 ();
 FILLCELL_X32 FILLER_276_3222 ();
 FILLCELL_X32 FILLER_276_3254 ();
 FILLCELL_X32 FILLER_276_3286 ();
 FILLCELL_X32 FILLER_276_3318 ();
 FILLCELL_X32 FILLER_276_3350 ();
 FILLCELL_X32 FILLER_276_3382 ();
 FILLCELL_X32 FILLER_276_3414 ();
 FILLCELL_X32 FILLER_276_3446 ();
 FILLCELL_X32 FILLER_276_3478 ();
 FILLCELL_X32 FILLER_276_3510 ();
 FILLCELL_X32 FILLER_276_3542 ();
 FILLCELL_X32 FILLER_276_3574 ();
 FILLCELL_X32 FILLER_276_3606 ();
 FILLCELL_X32 FILLER_276_3638 ();
 FILLCELL_X32 FILLER_276_3670 ();
 FILLCELL_X32 FILLER_276_3702 ();
 FILLCELL_X4 FILLER_276_3734 ();
 FILLCELL_X32 FILLER_277_1 ();
 FILLCELL_X32 FILLER_277_33 ();
 FILLCELL_X32 FILLER_277_65 ();
 FILLCELL_X32 FILLER_277_97 ();
 FILLCELL_X32 FILLER_277_129 ();
 FILLCELL_X32 FILLER_277_161 ();
 FILLCELL_X32 FILLER_277_193 ();
 FILLCELL_X32 FILLER_277_225 ();
 FILLCELL_X32 FILLER_277_257 ();
 FILLCELL_X32 FILLER_277_289 ();
 FILLCELL_X32 FILLER_277_321 ();
 FILLCELL_X32 FILLER_277_353 ();
 FILLCELL_X32 FILLER_277_385 ();
 FILLCELL_X32 FILLER_277_417 ();
 FILLCELL_X32 FILLER_277_449 ();
 FILLCELL_X32 FILLER_277_481 ();
 FILLCELL_X32 FILLER_277_513 ();
 FILLCELL_X32 FILLER_277_545 ();
 FILLCELL_X32 FILLER_277_577 ();
 FILLCELL_X32 FILLER_277_609 ();
 FILLCELL_X32 FILLER_277_641 ();
 FILLCELL_X32 FILLER_277_673 ();
 FILLCELL_X32 FILLER_277_705 ();
 FILLCELL_X32 FILLER_277_737 ();
 FILLCELL_X32 FILLER_277_769 ();
 FILLCELL_X32 FILLER_277_801 ();
 FILLCELL_X32 FILLER_277_833 ();
 FILLCELL_X32 FILLER_277_865 ();
 FILLCELL_X32 FILLER_277_897 ();
 FILLCELL_X32 FILLER_277_929 ();
 FILLCELL_X32 FILLER_277_961 ();
 FILLCELL_X32 FILLER_277_993 ();
 FILLCELL_X32 FILLER_277_1025 ();
 FILLCELL_X32 FILLER_277_1057 ();
 FILLCELL_X32 FILLER_277_1089 ();
 FILLCELL_X32 FILLER_277_1121 ();
 FILLCELL_X32 FILLER_277_1153 ();
 FILLCELL_X32 FILLER_277_1185 ();
 FILLCELL_X32 FILLER_277_1217 ();
 FILLCELL_X8 FILLER_277_1249 ();
 FILLCELL_X4 FILLER_277_1257 ();
 FILLCELL_X2 FILLER_277_1261 ();
 FILLCELL_X32 FILLER_277_1264 ();
 FILLCELL_X32 FILLER_277_1296 ();
 FILLCELL_X32 FILLER_277_1328 ();
 FILLCELL_X32 FILLER_277_1360 ();
 FILLCELL_X32 FILLER_277_1392 ();
 FILLCELL_X8 FILLER_277_1441 ();
 FILLCELL_X2 FILLER_277_1449 ();
 FILLCELL_X32 FILLER_277_1468 ();
 FILLCELL_X32 FILLER_277_1500 ();
 FILLCELL_X8 FILLER_277_1532 ();
 FILLCELL_X1 FILLER_277_1540 ();
 FILLCELL_X2 FILLER_277_1558 ();
 FILLCELL_X1 FILLER_277_1560 ();
 FILLCELL_X16 FILLER_277_1568 ();
 FILLCELL_X4 FILLER_277_1584 ();
 FILLCELL_X32 FILLER_277_1595 ();
 FILLCELL_X32 FILLER_277_1627 ();
 FILLCELL_X32 FILLER_277_1659 ();
 FILLCELL_X8 FILLER_277_1691 ();
 FILLCELL_X4 FILLER_277_1699 ();
 FILLCELL_X2 FILLER_277_1710 ();
 FILLCELL_X1 FILLER_277_1719 ();
 FILLCELL_X32 FILLER_277_1724 ();
 FILLCELL_X32 FILLER_277_1756 ();
 FILLCELL_X32 FILLER_277_1788 ();
 FILLCELL_X32 FILLER_277_1820 ();
 FILLCELL_X32 FILLER_277_1852 ();
 FILLCELL_X32 FILLER_277_1884 ();
 FILLCELL_X32 FILLER_277_1916 ();
 FILLCELL_X32 FILLER_277_1948 ();
 FILLCELL_X32 FILLER_277_1980 ();
 FILLCELL_X32 FILLER_277_2012 ();
 FILLCELL_X32 FILLER_277_2044 ();
 FILLCELL_X32 FILLER_277_2076 ();
 FILLCELL_X32 FILLER_277_2108 ();
 FILLCELL_X32 FILLER_277_2140 ();
 FILLCELL_X32 FILLER_277_2172 ();
 FILLCELL_X32 FILLER_277_2204 ();
 FILLCELL_X32 FILLER_277_2236 ();
 FILLCELL_X32 FILLER_277_2268 ();
 FILLCELL_X32 FILLER_277_2300 ();
 FILLCELL_X32 FILLER_277_2332 ();
 FILLCELL_X32 FILLER_277_2364 ();
 FILLCELL_X32 FILLER_277_2396 ();
 FILLCELL_X32 FILLER_277_2428 ();
 FILLCELL_X32 FILLER_277_2460 ();
 FILLCELL_X32 FILLER_277_2492 ();
 FILLCELL_X2 FILLER_277_2524 ();
 FILLCELL_X32 FILLER_277_2527 ();
 FILLCELL_X32 FILLER_277_2559 ();
 FILLCELL_X32 FILLER_277_2591 ();
 FILLCELL_X32 FILLER_277_2623 ();
 FILLCELL_X32 FILLER_277_2655 ();
 FILLCELL_X32 FILLER_277_2687 ();
 FILLCELL_X32 FILLER_277_2719 ();
 FILLCELL_X32 FILLER_277_2751 ();
 FILLCELL_X32 FILLER_277_2783 ();
 FILLCELL_X32 FILLER_277_2815 ();
 FILLCELL_X32 FILLER_277_2847 ();
 FILLCELL_X32 FILLER_277_2879 ();
 FILLCELL_X32 FILLER_277_2911 ();
 FILLCELL_X32 FILLER_277_2943 ();
 FILLCELL_X32 FILLER_277_2975 ();
 FILLCELL_X32 FILLER_277_3007 ();
 FILLCELL_X32 FILLER_277_3039 ();
 FILLCELL_X32 FILLER_277_3071 ();
 FILLCELL_X32 FILLER_277_3103 ();
 FILLCELL_X32 FILLER_277_3135 ();
 FILLCELL_X32 FILLER_277_3167 ();
 FILLCELL_X32 FILLER_277_3199 ();
 FILLCELL_X32 FILLER_277_3231 ();
 FILLCELL_X32 FILLER_277_3263 ();
 FILLCELL_X32 FILLER_277_3295 ();
 FILLCELL_X32 FILLER_277_3327 ();
 FILLCELL_X32 FILLER_277_3359 ();
 FILLCELL_X32 FILLER_277_3391 ();
 FILLCELL_X32 FILLER_277_3423 ();
 FILLCELL_X32 FILLER_277_3455 ();
 FILLCELL_X32 FILLER_277_3487 ();
 FILLCELL_X32 FILLER_277_3519 ();
 FILLCELL_X32 FILLER_277_3551 ();
 FILLCELL_X32 FILLER_277_3583 ();
 FILLCELL_X32 FILLER_277_3615 ();
 FILLCELL_X32 FILLER_277_3647 ();
 FILLCELL_X32 FILLER_277_3679 ();
 FILLCELL_X16 FILLER_277_3711 ();
 FILLCELL_X8 FILLER_277_3727 ();
 FILLCELL_X2 FILLER_277_3735 ();
 FILLCELL_X1 FILLER_277_3737 ();
 FILLCELL_X32 FILLER_278_1 ();
 FILLCELL_X32 FILLER_278_33 ();
 FILLCELL_X32 FILLER_278_65 ();
 FILLCELL_X32 FILLER_278_97 ();
 FILLCELL_X32 FILLER_278_129 ();
 FILLCELL_X32 FILLER_278_161 ();
 FILLCELL_X32 FILLER_278_193 ();
 FILLCELL_X32 FILLER_278_225 ();
 FILLCELL_X32 FILLER_278_257 ();
 FILLCELL_X32 FILLER_278_289 ();
 FILLCELL_X32 FILLER_278_321 ();
 FILLCELL_X32 FILLER_278_353 ();
 FILLCELL_X32 FILLER_278_385 ();
 FILLCELL_X32 FILLER_278_417 ();
 FILLCELL_X32 FILLER_278_449 ();
 FILLCELL_X32 FILLER_278_481 ();
 FILLCELL_X32 FILLER_278_513 ();
 FILLCELL_X32 FILLER_278_545 ();
 FILLCELL_X32 FILLER_278_577 ();
 FILLCELL_X16 FILLER_278_609 ();
 FILLCELL_X4 FILLER_278_625 ();
 FILLCELL_X2 FILLER_278_629 ();
 FILLCELL_X32 FILLER_278_632 ();
 FILLCELL_X32 FILLER_278_664 ();
 FILLCELL_X32 FILLER_278_696 ();
 FILLCELL_X32 FILLER_278_728 ();
 FILLCELL_X32 FILLER_278_760 ();
 FILLCELL_X32 FILLER_278_792 ();
 FILLCELL_X32 FILLER_278_824 ();
 FILLCELL_X32 FILLER_278_856 ();
 FILLCELL_X32 FILLER_278_888 ();
 FILLCELL_X32 FILLER_278_920 ();
 FILLCELL_X32 FILLER_278_952 ();
 FILLCELL_X32 FILLER_278_984 ();
 FILLCELL_X32 FILLER_278_1016 ();
 FILLCELL_X32 FILLER_278_1048 ();
 FILLCELL_X32 FILLER_278_1080 ();
 FILLCELL_X32 FILLER_278_1112 ();
 FILLCELL_X32 FILLER_278_1144 ();
 FILLCELL_X32 FILLER_278_1176 ();
 FILLCELL_X32 FILLER_278_1208 ();
 FILLCELL_X32 FILLER_278_1240 ();
 FILLCELL_X32 FILLER_278_1272 ();
 FILLCELL_X32 FILLER_278_1304 ();
 FILLCELL_X32 FILLER_278_1336 ();
 FILLCELL_X32 FILLER_278_1368 ();
 FILLCELL_X8 FILLER_278_1400 ();
 FILLCELL_X1 FILLER_278_1408 ();
 FILLCELL_X32 FILLER_278_1426 ();
 FILLCELL_X8 FILLER_278_1458 ();
 FILLCELL_X4 FILLER_278_1466 ();
 FILLCELL_X1 FILLER_278_1470 ();
 FILLCELL_X4 FILLER_278_1475 ();
 FILLCELL_X1 FILLER_278_1479 ();
 FILLCELL_X2 FILLER_278_1487 ();
 FILLCELL_X1 FILLER_278_1489 ();
 FILLCELL_X32 FILLER_278_1521 ();
 FILLCELL_X8 FILLER_278_1570 ();
 FILLCELL_X4 FILLER_278_1578 ();
 FILLCELL_X2 FILLER_278_1582 ();
 FILLCELL_X1 FILLER_278_1584 ();
 FILLCELL_X32 FILLER_278_1602 ();
 FILLCELL_X16 FILLER_278_1634 ();
 FILLCELL_X8 FILLER_278_1650 ();
 FILLCELL_X2 FILLER_278_1658 ();
 FILLCELL_X1 FILLER_278_1660 ();
 FILLCELL_X16 FILLER_278_1678 ();
 FILLCELL_X4 FILLER_278_1694 ();
 FILLCELL_X1 FILLER_278_1698 ();
 FILLCELL_X16 FILLER_278_1716 ();
 FILLCELL_X2 FILLER_278_1732 ();
 FILLCELL_X1 FILLER_278_1734 ();
 FILLCELL_X32 FILLER_278_1759 ();
 FILLCELL_X32 FILLER_278_1791 ();
 FILLCELL_X32 FILLER_278_1823 ();
 FILLCELL_X32 FILLER_278_1855 ();
 FILLCELL_X4 FILLER_278_1887 ();
 FILLCELL_X2 FILLER_278_1891 ();
 FILLCELL_X1 FILLER_278_1893 ();
 FILLCELL_X32 FILLER_278_1895 ();
 FILLCELL_X32 FILLER_278_1927 ();
 FILLCELL_X32 FILLER_278_1959 ();
 FILLCELL_X32 FILLER_278_1991 ();
 FILLCELL_X32 FILLER_278_2023 ();
 FILLCELL_X32 FILLER_278_2055 ();
 FILLCELL_X32 FILLER_278_2087 ();
 FILLCELL_X32 FILLER_278_2119 ();
 FILLCELL_X32 FILLER_278_2151 ();
 FILLCELL_X32 FILLER_278_2183 ();
 FILLCELL_X32 FILLER_278_2215 ();
 FILLCELL_X32 FILLER_278_2247 ();
 FILLCELL_X32 FILLER_278_2279 ();
 FILLCELL_X32 FILLER_278_2311 ();
 FILLCELL_X32 FILLER_278_2343 ();
 FILLCELL_X32 FILLER_278_2375 ();
 FILLCELL_X32 FILLER_278_2407 ();
 FILLCELL_X32 FILLER_278_2439 ();
 FILLCELL_X32 FILLER_278_2471 ();
 FILLCELL_X32 FILLER_278_2503 ();
 FILLCELL_X32 FILLER_278_2535 ();
 FILLCELL_X32 FILLER_278_2567 ();
 FILLCELL_X32 FILLER_278_2599 ();
 FILLCELL_X32 FILLER_278_2631 ();
 FILLCELL_X32 FILLER_278_2663 ();
 FILLCELL_X32 FILLER_278_2695 ();
 FILLCELL_X32 FILLER_278_2727 ();
 FILLCELL_X32 FILLER_278_2759 ();
 FILLCELL_X32 FILLER_278_2791 ();
 FILLCELL_X32 FILLER_278_2823 ();
 FILLCELL_X32 FILLER_278_2855 ();
 FILLCELL_X32 FILLER_278_2887 ();
 FILLCELL_X32 FILLER_278_2919 ();
 FILLCELL_X32 FILLER_278_2951 ();
 FILLCELL_X32 FILLER_278_2983 ();
 FILLCELL_X32 FILLER_278_3015 ();
 FILLCELL_X32 FILLER_278_3047 ();
 FILLCELL_X32 FILLER_278_3079 ();
 FILLCELL_X32 FILLER_278_3111 ();
 FILLCELL_X8 FILLER_278_3143 ();
 FILLCELL_X4 FILLER_278_3151 ();
 FILLCELL_X2 FILLER_278_3155 ();
 FILLCELL_X32 FILLER_278_3158 ();
 FILLCELL_X32 FILLER_278_3190 ();
 FILLCELL_X32 FILLER_278_3222 ();
 FILLCELL_X32 FILLER_278_3254 ();
 FILLCELL_X32 FILLER_278_3286 ();
 FILLCELL_X32 FILLER_278_3318 ();
 FILLCELL_X32 FILLER_278_3350 ();
 FILLCELL_X32 FILLER_278_3382 ();
 FILLCELL_X32 FILLER_278_3414 ();
 FILLCELL_X32 FILLER_278_3446 ();
 FILLCELL_X32 FILLER_278_3478 ();
 FILLCELL_X32 FILLER_278_3510 ();
 FILLCELL_X32 FILLER_278_3542 ();
 FILLCELL_X32 FILLER_278_3574 ();
 FILLCELL_X32 FILLER_278_3606 ();
 FILLCELL_X32 FILLER_278_3638 ();
 FILLCELL_X32 FILLER_278_3670 ();
 FILLCELL_X32 FILLER_278_3702 ();
 FILLCELL_X4 FILLER_278_3734 ();
 FILLCELL_X32 FILLER_279_1 ();
 FILLCELL_X32 FILLER_279_33 ();
 FILLCELL_X32 FILLER_279_65 ();
 FILLCELL_X32 FILLER_279_97 ();
 FILLCELL_X32 FILLER_279_129 ();
 FILLCELL_X32 FILLER_279_161 ();
 FILLCELL_X32 FILLER_279_193 ();
 FILLCELL_X32 FILLER_279_225 ();
 FILLCELL_X32 FILLER_279_257 ();
 FILLCELL_X32 FILLER_279_289 ();
 FILLCELL_X32 FILLER_279_321 ();
 FILLCELL_X32 FILLER_279_353 ();
 FILLCELL_X32 FILLER_279_385 ();
 FILLCELL_X32 FILLER_279_417 ();
 FILLCELL_X32 FILLER_279_449 ();
 FILLCELL_X32 FILLER_279_481 ();
 FILLCELL_X32 FILLER_279_513 ();
 FILLCELL_X32 FILLER_279_545 ();
 FILLCELL_X32 FILLER_279_577 ();
 FILLCELL_X32 FILLER_279_609 ();
 FILLCELL_X32 FILLER_279_641 ();
 FILLCELL_X32 FILLER_279_673 ();
 FILLCELL_X32 FILLER_279_705 ();
 FILLCELL_X32 FILLER_279_737 ();
 FILLCELL_X32 FILLER_279_769 ();
 FILLCELL_X32 FILLER_279_801 ();
 FILLCELL_X32 FILLER_279_833 ();
 FILLCELL_X32 FILLER_279_865 ();
 FILLCELL_X32 FILLER_279_897 ();
 FILLCELL_X32 FILLER_279_929 ();
 FILLCELL_X32 FILLER_279_961 ();
 FILLCELL_X32 FILLER_279_993 ();
 FILLCELL_X32 FILLER_279_1025 ();
 FILLCELL_X32 FILLER_279_1057 ();
 FILLCELL_X32 FILLER_279_1089 ();
 FILLCELL_X32 FILLER_279_1121 ();
 FILLCELL_X32 FILLER_279_1153 ();
 FILLCELL_X32 FILLER_279_1185 ();
 FILLCELL_X32 FILLER_279_1217 ();
 FILLCELL_X8 FILLER_279_1249 ();
 FILLCELL_X4 FILLER_279_1257 ();
 FILLCELL_X2 FILLER_279_1261 ();
 FILLCELL_X32 FILLER_279_1264 ();
 FILLCELL_X32 FILLER_279_1296 ();
 FILLCELL_X32 FILLER_279_1328 ();
 FILLCELL_X32 FILLER_279_1360 ();
 FILLCELL_X16 FILLER_279_1392 ();
 FILLCELL_X4 FILLER_279_1408 ();
 FILLCELL_X1 FILLER_279_1412 ();
 FILLCELL_X4 FILLER_279_1420 ();
 FILLCELL_X2 FILLER_279_1424 ();
 FILLCELL_X1 FILLER_279_1426 ();
 FILLCELL_X16 FILLER_279_1434 ();
 FILLCELL_X2 FILLER_279_1450 ();
 FILLCELL_X1 FILLER_279_1452 ();
 FILLCELL_X2 FILLER_279_1460 ();
 FILLCELL_X1 FILLER_279_1462 ();
 FILLCELL_X4 FILLER_279_1470 ();
 FILLCELL_X2 FILLER_279_1474 ();
 FILLCELL_X16 FILLER_279_1481 ();
 FILLCELL_X4 FILLER_279_1497 ();
 FILLCELL_X32 FILLER_279_1518 ();
 FILLCELL_X32 FILLER_279_1550 ();
 FILLCELL_X8 FILLER_279_1582 ();
 FILLCELL_X2 FILLER_279_1590 ();
 FILLCELL_X1 FILLER_279_1592 ();
 FILLCELL_X8 FILLER_279_1600 ();
 FILLCELL_X4 FILLER_279_1608 ();
 FILLCELL_X1 FILLER_279_1612 ();
 FILLCELL_X16 FILLER_279_1630 ();
 FILLCELL_X8 FILLER_279_1660 ();
 FILLCELL_X4 FILLER_279_1668 ();
 FILLCELL_X16 FILLER_279_1686 ();
 FILLCELL_X4 FILLER_279_1702 ();
 FILLCELL_X1 FILLER_279_1706 ();
 FILLCELL_X16 FILLER_279_1714 ();
 FILLCELL_X8 FILLER_279_1730 ();
 FILLCELL_X2 FILLER_279_1738 ();
 FILLCELL_X1 FILLER_279_1740 ();
 FILLCELL_X32 FILLER_279_1748 ();
 FILLCELL_X32 FILLER_279_1780 ();
 FILLCELL_X32 FILLER_279_1812 ();
 FILLCELL_X32 FILLER_279_1844 ();
 FILLCELL_X32 FILLER_279_1876 ();
 FILLCELL_X32 FILLER_279_1908 ();
 FILLCELL_X32 FILLER_279_1940 ();
 FILLCELL_X32 FILLER_279_1972 ();
 FILLCELL_X32 FILLER_279_2004 ();
 FILLCELL_X32 FILLER_279_2036 ();
 FILLCELL_X32 FILLER_279_2068 ();
 FILLCELL_X32 FILLER_279_2100 ();
 FILLCELL_X32 FILLER_279_2132 ();
 FILLCELL_X32 FILLER_279_2164 ();
 FILLCELL_X32 FILLER_279_2196 ();
 FILLCELL_X32 FILLER_279_2228 ();
 FILLCELL_X32 FILLER_279_2260 ();
 FILLCELL_X32 FILLER_279_2292 ();
 FILLCELL_X32 FILLER_279_2324 ();
 FILLCELL_X32 FILLER_279_2356 ();
 FILLCELL_X32 FILLER_279_2388 ();
 FILLCELL_X32 FILLER_279_2420 ();
 FILLCELL_X32 FILLER_279_2452 ();
 FILLCELL_X32 FILLER_279_2484 ();
 FILLCELL_X8 FILLER_279_2516 ();
 FILLCELL_X2 FILLER_279_2524 ();
 FILLCELL_X32 FILLER_279_2527 ();
 FILLCELL_X32 FILLER_279_2559 ();
 FILLCELL_X32 FILLER_279_2591 ();
 FILLCELL_X32 FILLER_279_2623 ();
 FILLCELL_X32 FILLER_279_2655 ();
 FILLCELL_X32 FILLER_279_2687 ();
 FILLCELL_X32 FILLER_279_2719 ();
 FILLCELL_X32 FILLER_279_2751 ();
 FILLCELL_X32 FILLER_279_2783 ();
 FILLCELL_X32 FILLER_279_2815 ();
 FILLCELL_X32 FILLER_279_2847 ();
 FILLCELL_X32 FILLER_279_2879 ();
 FILLCELL_X32 FILLER_279_2911 ();
 FILLCELL_X32 FILLER_279_2943 ();
 FILLCELL_X32 FILLER_279_2975 ();
 FILLCELL_X32 FILLER_279_3007 ();
 FILLCELL_X32 FILLER_279_3039 ();
 FILLCELL_X32 FILLER_279_3071 ();
 FILLCELL_X32 FILLER_279_3103 ();
 FILLCELL_X32 FILLER_279_3135 ();
 FILLCELL_X32 FILLER_279_3167 ();
 FILLCELL_X32 FILLER_279_3199 ();
 FILLCELL_X32 FILLER_279_3231 ();
 FILLCELL_X32 FILLER_279_3263 ();
 FILLCELL_X32 FILLER_279_3295 ();
 FILLCELL_X32 FILLER_279_3327 ();
 FILLCELL_X32 FILLER_279_3359 ();
 FILLCELL_X32 FILLER_279_3391 ();
 FILLCELL_X32 FILLER_279_3423 ();
 FILLCELL_X32 FILLER_279_3455 ();
 FILLCELL_X32 FILLER_279_3487 ();
 FILLCELL_X32 FILLER_279_3519 ();
 FILLCELL_X32 FILLER_279_3551 ();
 FILLCELL_X32 FILLER_279_3583 ();
 FILLCELL_X32 FILLER_279_3615 ();
 FILLCELL_X32 FILLER_279_3647 ();
 FILLCELL_X32 FILLER_279_3679 ();
 FILLCELL_X16 FILLER_279_3711 ();
 FILLCELL_X8 FILLER_279_3727 ();
 FILLCELL_X2 FILLER_279_3735 ();
 FILLCELL_X1 FILLER_279_3737 ();
 FILLCELL_X32 FILLER_280_1 ();
 FILLCELL_X32 FILLER_280_33 ();
 FILLCELL_X32 FILLER_280_65 ();
 FILLCELL_X32 FILLER_280_97 ();
 FILLCELL_X32 FILLER_280_129 ();
 FILLCELL_X32 FILLER_280_161 ();
 FILLCELL_X32 FILLER_280_193 ();
 FILLCELL_X32 FILLER_280_225 ();
 FILLCELL_X32 FILLER_280_257 ();
 FILLCELL_X32 FILLER_280_289 ();
 FILLCELL_X32 FILLER_280_321 ();
 FILLCELL_X32 FILLER_280_353 ();
 FILLCELL_X32 FILLER_280_385 ();
 FILLCELL_X32 FILLER_280_417 ();
 FILLCELL_X32 FILLER_280_449 ();
 FILLCELL_X32 FILLER_280_481 ();
 FILLCELL_X32 FILLER_280_513 ();
 FILLCELL_X32 FILLER_280_545 ();
 FILLCELL_X32 FILLER_280_577 ();
 FILLCELL_X16 FILLER_280_609 ();
 FILLCELL_X4 FILLER_280_625 ();
 FILLCELL_X2 FILLER_280_629 ();
 FILLCELL_X32 FILLER_280_632 ();
 FILLCELL_X32 FILLER_280_664 ();
 FILLCELL_X32 FILLER_280_696 ();
 FILLCELL_X32 FILLER_280_728 ();
 FILLCELL_X32 FILLER_280_760 ();
 FILLCELL_X32 FILLER_280_792 ();
 FILLCELL_X32 FILLER_280_824 ();
 FILLCELL_X32 FILLER_280_856 ();
 FILLCELL_X32 FILLER_280_888 ();
 FILLCELL_X32 FILLER_280_920 ();
 FILLCELL_X32 FILLER_280_952 ();
 FILLCELL_X32 FILLER_280_984 ();
 FILLCELL_X32 FILLER_280_1016 ();
 FILLCELL_X32 FILLER_280_1048 ();
 FILLCELL_X32 FILLER_280_1080 ();
 FILLCELL_X32 FILLER_280_1112 ();
 FILLCELL_X32 FILLER_280_1144 ();
 FILLCELL_X32 FILLER_280_1176 ();
 FILLCELL_X32 FILLER_280_1208 ();
 FILLCELL_X32 FILLER_280_1240 ();
 FILLCELL_X32 FILLER_280_1272 ();
 FILLCELL_X32 FILLER_280_1304 ();
 FILLCELL_X32 FILLER_280_1336 ();
 FILLCELL_X32 FILLER_280_1368 ();
 FILLCELL_X8 FILLER_280_1400 ();
 FILLCELL_X4 FILLER_280_1408 ();
 FILLCELL_X8 FILLER_280_1436 ();
 FILLCELL_X4 FILLER_280_1444 ();
 FILLCELL_X32 FILLER_280_1465 ();
 FILLCELL_X32 FILLER_280_1497 ();
 FILLCELL_X16 FILLER_280_1529 ();
 FILLCELL_X8 FILLER_280_1545 ();
 FILLCELL_X2 FILLER_280_1553 ();
 FILLCELL_X1 FILLER_280_1555 ();
 FILLCELL_X16 FILLER_280_1587 ();
 FILLCELL_X8 FILLER_280_1603 ();
 FILLCELL_X4 FILLER_280_1611 ();
 FILLCELL_X2 FILLER_280_1615 ();
 FILLCELL_X2 FILLER_280_1624 ();
 FILLCELL_X1 FILLER_280_1626 ();
 FILLCELL_X8 FILLER_280_1634 ();
 FILLCELL_X4 FILLER_280_1642 ();
 FILLCELL_X2 FILLER_280_1646 ();
 FILLCELL_X8 FILLER_280_1665 ();
 FILLCELL_X2 FILLER_280_1673 ();
 FILLCELL_X16 FILLER_280_1682 ();
 FILLCELL_X4 FILLER_280_1698 ();
 FILLCELL_X2 FILLER_280_1702 ();
 FILLCELL_X32 FILLER_280_1728 ();
 FILLCELL_X32 FILLER_280_1760 ();
 FILLCELL_X32 FILLER_280_1792 ();
 FILLCELL_X32 FILLER_280_1824 ();
 FILLCELL_X32 FILLER_280_1856 ();
 FILLCELL_X4 FILLER_280_1888 ();
 FILLCELL_X2 FILLER_280_1892 ();
 FILLCELL_X32 FILLER_280_1895 ();
 FILLCELL_X32 FILLER_280_1927 ();
 FILLCELL_X32 FILLER_280_1959 ();
 FILLCELL_X32 FILLER_280_1991 ();
 FILLCELL_X32 FILLER_280_2023 ();
 FILLCELL_X32 FILLER_280_2055 ();
 FILLCELL_X32 FILLER_280_2087 ();
 FILLCELL_X32 FILLER_280_2119 ();
 FILLCELL_X32 FILLER_280_2151 ();
 FILLCELL_X32 FILLER_280_2183 ();
 FILLCELL_X32 FILLER_280_2215 ();
 FILLCELL_X32 FILLER_280_2247 ();
 FILLCELL_X32 FILLER_280_2279 ();
 FILLCELL_X32 FILLER_280_2311 ();
 FILLCELL_X32 FILLER_280_2343 ();
 FILLCELL_X32 FILLER_280_2375 ();
 FILLCELL_X32 FILLER_280_2407 ();
 FILLCELL_X32 FILLER_280_2439 ();
 FILLCELL_X32 FILLER_280_2471 ();
 FILLCELL_X32 FILLER_280_2503 ();
 FILLCELL_X32 FILLER_280_2535 ();
 FILLCELL_X32 FILLER_280_2567 ();
 FILLCELL_X32 FILLER_280_2599 ();
 FILLCELL_X32 FILLER_280_2631 ();
 FILLCELL_X32 FILLER_280_2663 ();
 FILLCELL_X32 FILLER_280_2695 ();
 FILLCELL_X32 FILLER_280_2727 ();
 FILLCELL_X32 FILLER_280_2759 ();
 FILLCELL_X32 FILLER_280_2791 ();
 FILLCELL_X32 FILLER_280_2823 ();
 FILLCELL_X32 FILLER_280_2855 ();
 FILLCELL_X32 FILLER_280_2887 ();
 FILLCELL_X32 FILLER_280_2919 ();
 FILLCELL_X32 FILLER_280_2951 ();
 FILLCELL_X32 FILLER_280_2983 ();
 FILLCELL_X32 FILLER_280_3015 ();
 FILLCELL_X32 FILLER_280_3047 ();
 FILLCELL_X32 FILLER_280_3079 ();
 FILLCELL_X32 FILLER_280_3111 ();
 FILLCELL_X8 FILLER_280_3143 ();
 FILLCELL_X4 FILLER_280_3151 ();
 FILLCELL_X2 FILLER_280_3155 ();
 FILLCELL_X32 FILLER_280_3158 ();
 FILLCELL_X32 FILLER_280_3190 ();
 FILLCELL_X32 FILLER_280_3222 ();
 FILLCELL_X32 FILLER_280_3254 ();
 FILLCELL_X32 FILLER_280_3286 ();
 FILLCELL_X32 FILLER_280_3318 ();
 FILLCELL_X32 FILLER_280_3350 ();
 FILLCELL_X32 FILLER_280_3382 ();
 FILLCELL_X32 FILLER_280_3414 ();
 FILLCELL_X32 FILLER_280_3446 ();
 FILLCELL_X32 FILLER_280_3478 ();
 FILLCELL_X32 FILLER_280_3510 ();
 FILLCELL_X32 FILLER_280_3542 ();
 FILLCELL_X32 FILLER_280_3574 ();
 FILLCELL_X32 FILLER_280_3606 ();
 FILLCELL_X32 FILLER_280_3638 ();
 FILLCELL_X32 FILLER_280_3670 ();
 FILLCELL_X32 FILLER_280_3702 ();
 FILLCELL_X4 FILLER_280_3734 ();
 FILLCELL_X32 FILLER_281_1 ();
 FILLCELL_X32 FILLER_281_33 ();
 FILLCELL_X32 FILLER_281_65 ();
 FILLCELL_X32 FILLER_281_97 ();
 FILLCELL_X32 FILLER_281_129 ();
 FILLCELL_X32 FILLER_281_161 ();
 FILLCELL_X32 FILLER_281_193 ();
 FILLCELL_X32 FILLER_281_225 ();
 FILLCELL_X32 FILLER_281_257 ();
 FILLCELL_X32 FILLER_281_289 ();
 FILLCELL_X32 FILLER_281_321 ();
 FILLCELL_X32 FILLER_281_353 ();
 FILLCELL_X32 FILLER_281_385 ();
 FILLCELL_X32 FILLER_281_417 ();
 FILLCELL_X32 FILLER_281_449 ();
 FILLCELL_X32 FILLER_281_481 ();
 FILLCELL_X32 FILLER_281_513 ();
 FILLCELL_X32 FILLER_281_545 ();
 FILLCELL_X32 FILLER_281_577 ();
 FILLCELL_X32 FILLER_281_609 ();
 FILLCELL_X32 FILLER_281_641 ();
 FILLCELL_X32 FILLER_281_673 ();
 FILLCELL_X32 FILLER_281_705 ();
 FILLCELL_X32 FILLER_281_737 ();
 FILLCELL_X32 FILLER_281_769 ();
 FILLCELL_X32 FILLER_281_801 ();
 FILLCELL_X32 FILLER_281_833 ();
 FILLCELL_X32 FILLER_281_865 ();
 FILLCELL_X32 FILLER_281_897 ();
 FILLCELL_X32 FILLER_281_929 ();
 FILLCELL_X32 FILLER_281_961 ();
 FILLCELL_X32 FILLER_281_993 ();
 FILLCELL_X32 FILLER_281_1025 ();
 FILLCELL_X32 FILLER_281_1057 ();
 FILLCELL_X32 FILLER_281_1089 ();
 FILLCELL_X32 FILLER_281_1121 ();
 FILLCELL_X32 FILLER_281_1153 ();
 FILLCELL_X32 FILLER_281_1185 ();
 FILLCELL_X32 FILLER_281_1217 ();
 FILLCELL_X8 FILLER_281_1249 ();
 FILLCELL_X4 FILLER_281_1257 ();
 FILLCELL_X2 FILLER_281_1261 ();
 FILLCELL_X32 FILLER_281_1264 ();
 FILLCELL_X32 FILLER_281_1296 ();
 FILLCELL_X32 FILLER_281_1328 ();
 FILLCELL_X32 FILLER_281_1360 ();
 FILLCELL_X32 FILLER_281_1392 ();
 FILLCELL_X32 FILLER_281_1424 ();
 FILLCELL_X32 FILLER_281_1456 ();
 FILLCELL_X16 FILLER_281_1488 ();
 FILLCELL_X8 FILLER_281_1504 ();
 FILLCELL_X32 FILLER_281_1536 ();
 FILLCELL_X4 FILLER_281_1568 ();
 FILLCELL_X2 FILLER_281_1572 ();
 FILLCELL_X1 FILLER_281_1574 ();
 FILLCELL_X32 FILLER_281_1589 ();
 FILLCELL_X8 FILLER_281_1621 ();
 FILLCELL_X4 FILLER_281_1629 ();
 FILLCELL_X2 FILLER_281_1633 ();
 FILLCELL_X32 FILLER_281_1639 ();
 FILLCELL_X32 FILLER_281_1671 ();
 FILLCELL_X32 FILLER_281_1703 ();
 FILLCELL_X8 FILLER_281_1735 ();
 FILLCELL_X1 FILLER_281_1743 ();
 FILLCELL_X32 FILLER_281_1751 ();
 FILLCELL_X32 FILLER_281_1783 ();
 FILLCELL_X32 FILLER_281_1815 ();
 FILLCELL_X32 FILLER_281_1847 ();
 FILLCELL_X32 FILLER_281_1879 ();
 FILLCELL_X32 FILLER_281_1911 ();
 FILLCELL_X32 FILLER_281_1943 ();
 FILLCELL_X32 FILLER_281_1975 ();
 FILLCELL_X32 FILLER_281_2007 ();
 FILLCELL_X32 FILLER_281_2039 ();
 FILLCELL_X32 FILLER_281_2071 ();
 FILLCELL_X32 FILLER_281_2103 ();
 FILLCELL_X32 FILLER_281_2135 ();
 FILLCELL_X32 FILLER_281_2167 ();
 FILLCELL_X32 FILLER_281_2199 ();
 FILLCELL_X32 FILLER_281_2231 ();
 FILLCELL_X32 FILLER_281_2263 ();
 FILLCELL_X32 FILLER_281_2295 ();
 FILLCELL_X32 FILLER_281_2327 ();
 FILLCELL_X32 FILLER_281_2359 ();
 FILLCELL_X32 FILLER_281_2391 ();
 FILLCELL_X32 FILLER_281_2423 ();
 FILLCELL_X32 FILLER_281_2455 ();
 FILLCELL_X32 FILLER_281_2487 ();
 FILLCELL_X4 FILLER_281_2519 ();
 FILLCELL_X2 FILLER_281_2523 ();
 FILLCELL_X1 FILLER_281_2525 ();
 FILLCELL_X32 FILLER_281_2527 ();
 FILLCELL_X32 FILLER_281_2559 ();
 FILLCELL_X32 FILLER_281_2591 ();
 FILLCELL_X32 FILLER_281_2623 ();
 FILLCELL_X32 FILLER_281_2655 ();
 FILLCELL_X32 FILLER_281_2687 ();
 FILLCELL_X32 FILLER_281_2719 ();
 FILLCELL_X32 FILLER_281_2751 ();
 FILLCELL_X32 FILLER_281_2783 ();
 FILLCELL_X32 FILLER_281_2815 ();
 FILLCELL_X32 FILLER_281_2847 ();
 FILLCELL_X32 FILLER_281_2879 ();
 FILLCELL_X32 FILLER_281_2911 ();
 FILLCELL_X32 FILLER_281_2943 ();
 FILLCELL_X32 FILLER_281_2975 ();
 FILLCELL_X32 FILLER_281_3007 ();
 FILLCELL_X32 FILLER_281_3039 ();
 FILLCELL_X32 FILLER_281_3071 ();
 FILLCELL_X32 FILLER_281_3103 ();
 FILLCELL_X32 FILLER_281_3135 ();
 FILLCELL_X32 FILLER_281_3167 ();
 FILLCELL_X32 FILLER_281_3199 ();
 FILLCELL_X32 FILLER_281_3231 ();
 FILLCELL_X32 FILLER_281_3263 ();
 FILLCELL_X32 FILLER_281_3295 ();
 FILLCELL_X32 FILLER_281_3327 ();
 FILLCELL_X32 FILLER_281_3359 ();
 FILLCELL_X32 FILLER_281_3391 ();
 FILLCELL_X32 FILLER_281_3423 ();
 FILLCELL_X32 FILLER_281_3455 ();
 FILLCELL_X32 FILLER_281_3487 ();
 FILLCELL_X32 FILLER_281_3519 ();
 FILLCELL_X32 FILLER_281_3551 ();
 FILLCELL_X32 FILLER_281_3583 ();
 FILLCELL_X32 FILLER_281_3615 ();
 FILLCELL_X32 FILLER_281_3647 ();
 FILLCELL_X32 FILLER_281_3679 ();
 FILLCELL_X16 FILLER_281_3711 ();
 FILLCELL_X8 FILLER_281_3727 ();
 FILLCELL_X2 FILLER_281_3735 ();
 FILLCELL_X1 FILLER_281_3737 ();
 FILLCELL_X32 FILLER_282_1 ();
 FILLCELL_X32 FILLER_282_33 ();
 FILLCELL_X32 FILLER_282_65 ();
 FILLCELL_X32 FILLER_282_97 ();
 FILLCELL_X32 FILLER_282_129 ();
 FILLCELL_X32 FILLER_282_161 ();
 FILLCELL_X32 FILLER_282_193 ();
 FILLCELL_X32 FILLER_282_225 ();
 FILLCELL_X32 FILLER_282_257 ();
 FILLCELL_X32 FILLER_282_289 ();
 FILLCELL_X32 FILLER_282_321 ();
 FILLCELL_X32 FILLER_282_353 ();
 FILLCELL_X32 FILLER_282_385 ();
 FILLCELL_X32 FILLER_282_417 ();
 FILLCELL_X32 FILLER_282_449 ();
 FILLCELL_X32 FILLER_282_481 ();
 FILLCELL_X32 FILLER_282_513 ();
 FILLCELL_X32 FILLER_282_545 ();
 FILLCELL_X32 FILLER_282_577 ();
 FILLCELL_X16 FILLER_282_609 ();
 FILLCELL_X4 FILLER_282_625 ();
 FILLCELL_X2 FILLER_282_629 ();
 FILLCELL_X32 FILLER_282_632 ();
 FILLCELL_X32 FILLER_282_664 ();
 FILLCELL_X32 FILLER_282_696 ();
 FILLCELL_X32 FILLER_282_728 ();
 FILLCELL_X32 FILLER_282_760 ();
 FILLCELL_X32 FILLER_282_792 ();
 FILLCELL_X32 FILLER_282_824 ();
 FILLCELL_X32 FILLER_282_856 ();
 FILLCELL_X32 FILLER_282_888 ();
 FILLCELL_X32 FILLER_282_920 ();
 FILLCELL_X32 FILLER_282_952 ();
 FILLCELL_X32 FILLER_282_984 ();
 FILLCELL_X32 FILLER_282_1016 ();
 FILLCELL_X32 FILLER_282_1048 ();
 FILLCELL_X32 FILLER_282_1080 ();
 FILLCELL_X32 FILLER_282_1112 ();
 FILLCELL_X32 FILLER_282_1144 ();
 FILLCELL_X32 FILLER_282_1176 ();
 FILLCELL_X32 FILLER_282_1208 ();
 FILLCELL_X32 FILLER_282_1240 ();
 FILLCELL_X32 FILLER_282_1272 ();
 FILLCELL_X32 FILLER_282_1304 ();
 FILLCELL_X32 FILLER_282_1336 ();
 FILLCELL_X16 FILLER_282_1368 ();
 FILLCELL_X8 FILLER_282_1384 ();
 FILLCELL_X2 FILLER_282_1392 ();
 FILLCELL_X1 FILLER_282_1394 ();
 FILLCELL_X16 FILLER_282_1399 ();
 FILLCELL_X16 FILLER_282_1432 ();
 FILLCELL_X8 FILLER_282_1448 ();
 FILLCELL_X1 FILLER_282_1456 ();
 FILLCELL_X8 FILLER_282_1464 ();
 FILLCELL_X4 FILLER_282_1472 ();
 FILLCELL_X2 FILLER_282_1476 ();
 FILLCELL_X1 FILLER_282_1478 ();
 FILLCELL_X4 FILLER_282_1486 ();
 FILLCELL_X4 FILLER_282_1494 ();
 FILLCELL_X8 FILLER_282_1505 ();
 FILLCELL_X1 FILLER_282_1513 ();
 FILLCELL_X32 FILLER_282_1521 ();
 FILLCELL_X16 FILLER_282_1553 ();
 FILLCELL_X4 FILLER_282_1569 ();
 FILLCELL_X4 FILLER_282_1590 ();
 FILLCELL_X2 FILLER_282_1594 ();
 FILLCELL_X16 FILLER_282_1603 ();
 FILLCELL_X4 FILLER_282_1619 ();
 FILLCELL_X1 FILLER_282_1623 ();
 FILLCELL_X8 FILLER_282_1631 ();
 FILLCELL_X4 FILLER_282_1639 ();
 FILLCELL_X2 FILLER_282_1643 ();
 FILLCELL_X8 FILLER_282_1652 ();
 FILLCELL_X1 FILLER_282_1660 ();
 FILLCELL_X4 FILLER_282_1665 ();
 FILLCELL_X4 FILLER_282_1676 ();
 FILLCELL_X2 FILLER_282_1680 ();
 FILLCELL_X32 FILLER_282_1706 ();
 FILLCELL_X4 FILLER_282_1738 ();
 FILLCELL_X2 FILLER_282_1742 ();
 FILLCELL_X32 FILLER_282_1761 ();
 FILLCELL_X32 FILLER_282_1793 ();
 FILLCELL_X32 FILLER_282_1825 ();
 FILLCELL_X32 FILLER_282_1857 ();
 FILLCELL_X4 FILLER_282_1889 ();
 FILLCELL_X1 FILLER_282_1893 ();
 FILLCELL_X32 FILLER_282_1895 ();
 FILLCELL_X32 FILLER_282_1927 ();
 FILLCELL_X32 FILLER_282_1959 ();
 FILLCELL_X32 FILLER_282_1991 ();
 FILLCELL_X32 FILLER_282_2023 ();
 FILLCELL_X32 FILLER_282_2055 ();
 FILLCELL_X32 FILLER_282_2087 ();
 FILLCELL_X32 FILLER_282_2119 ();
 FILLCELL_X32 FILLER_282_2151 ();
 FILLCELL_X32 FILLER_282_2183 ();
 FILLCELL_X32 FILLER_282_2215 ();
 FILLCELL_X32 FILLER_282_2247 ();
 FILLCELL_X32 FILLER_282_2279 ();
 FILLCELL_X32 FILLER_282_2311 ();
 FILLCELL_X32 FILLER_282_2343 ();
 FILLCELL_X32 FILLER_282_2375 ();
 FILLCELL_X32 FILLER_282_2407 ();
 FILLCELL_X32 FILLER_282_2439 ();
 FILLCELL_X32 FILLER_282_2471 ();
 FILLCELL_X32 FILLER_282_2503 ();
 FILLCELL_X32 FILLER_282_2535 ();
 FILLCELL_X32 FILLER_282_2567 ();
 FILLCELL_X32 FILLER_282_2599 ();
 FILLCELL_X32 FILLER_282_2631 ();
 FILLCELL_X32 FILLER_282_2663 ();
 FILLCELL_X32 FILLER_282_2695 ();
 FILLCELL_X32 FILLER_282_2727 ();
 FILLCELL_X32 FILLER_282_2759 ();
 FILLCELL_X32 FILLER_282_2791 ();
 FILLCELL_X32 FILLER_282_2823 ();
 FILLCELL_X32 FILLER_282_2855 ();
 FILLCELL_X32 FILLER_282_2887 ();
 FILLCELL_X32 FILLER_282_2919 ();
 FILLCELL_X32 FILLER_282_2951 ();
 FILLCELL_X32 FILLER_282_2983 ();
 FILLCELL_X32 FILLER_282_3015 ();
 FILLCELL_X32 FILLER_282_3047 ();
 FILLCELL_X32 FILLER_282_3079 ();
 FILLCELL_X32 FILLER_282_3111 ();
 FILLCELL_X8 FILLER_282_3143 ();
 FILLCELL_X4 FILLER_282_3151 ();
 FILLCELL_X2 FILLER_282_3155 ();
 FILLCELL_X32 FILLER_282_3158 ();
 FILLCELL_X32 FILLER_282_3190 ();
 FILLCELL_X32 FILLER_282_3222 ();
 FILLCELL_X32 FILLER_282_3254 ();
 FILLCELL_X32 FILLER_282_3286 ();
 FILLCELL_X32 FILLER_282_3318 ();
 FILLCELL_X32 FILLER_282_3350 ();
 FILLCELL_X32 FILLER_282_3382 ();
 FILLCELL_X32 FILLER_282_3414 ();
 FILLCELL_X32 FILLER_282_3446 ();
 FILLCELL_X32 FILLER_282_3478 ();
 FILLCELL_X32 FILLER_282_3510 ();
 FILLCELL_X32 FILLER_282_3542 ();
 FILLCELL_X32 FILLER_282_3574 ();
 FILLCELL_X32 FILLER_282_3606 ();
 FILLCELL_X32 FILLER_282_3638 ();
 FILLCELL_X32 FILLER_282_3670 ();
 FILLCELL_X32 FILLER_282_3702 ();
 FILLCELL_X4 FILLER_282_3734 ();
 FILLCELL_X32 FILLER_283_1 ();
 FILLCELL_X32 FILLER_283_33 ();
 FILLCELL_X32 FILLER_283_65 ();
 FILLCELL_X32 FILLER_283_97 ();
 FILLCELL_X32 FILLER_283_129 ();
 FILLCELL_X32 FILLER_283_161 ();
 FILLCELL_X32 FILLER_283_193 ();
 FILLCELL_X32 FILLER_283_225 ();
 FILLCELL_X32 FILLER_283_257 ();
 FILLCELL_X32 FILLER_283_289 ();
 FILLCELL_X32 FILLER_283_321 ();
 FILLCELL_X32 FILLER_283_353 ();
 FILLCELL_X32 FILLER_283_385 ();
 FILLCELL_X32 FILLER_283_417 ();
 FILLCELL_X32 FILLER_283_449 ();
 FILLCELL_X32 FILLER_283_481 ();
 FILLCELL_X32 FILLER_283_513 ();
 FILLCELL_X32 FILLER_283_545 ();
 FILLCELL_X32 FILLER_283_577 ();
 FILLCELL_X32 FILLER_283_609 ();
 FILLCELL_X32 FILLER_283_641 ();
 FILLCELL_X32 FILLER_283_673 ();
 FILLCELL_X32 FILLER_283_705 ();
 FILLCELL_X32 FILLER_283_737 ();
 FILLCELL_X32 FILLER_283_769 ();
 FILLCELL_X32 FILLER_283_801 ();
 FILLCELL_X32 FILLER_283_833 ();
 FILLCELL_X32 FILLER_283_865 ();
 FILLCELL_X32 FILLER_283_897 ();
 FILLCELL_X32 FILLER_283_929 ();
 FILLCELL_X32 FILLER_283_961 ();
 FILLCELL_X32 FILLER_283_993 ();
 FILLCELL_X32 FILLER_283_1025 ();
 FILLCELL_X32 FILLER_283_1057 ();
 FILLCELL_X32 FILLER_283_1089 ();
 FILLCELL_X32 FILLER_283_1121 ();
 FILLCELL_X32 FILLER_283_1153 ();
 FILLCELL_X32 FILLER_283_1185 ();
 FILLCELL_X32 FILLER_283_1217 ();
 FILLCELL_X8 FILLER_283_1249 ();
 FILLCELL_X4 FILLER_283_1257 ();
 FILLCELL_X2 FILLER_283_1261 ();
 FILLCELL_X32 FILLER_283_1264 ();
 FILLCELL_X32 FILLER_283_1296 ();
 FILLCELL_X32 FILLER_283_1328 ();
 FILLCELL_X16 FILLER_283_1360 ();
 FILLCELL_X8 FILLER_283_1376 ();
 FILLCELL_X2 FILLER_283_1384 ();
 FILLCELL_X1 FILLER_283_1386 ();
 FILLCELL_X16 FILLER_283_1391 ();
 FILLCELL_X4 FILLER_283_1407 ();
 FILLCELL_X2 FILLER_283_1411 ();
 FILLCELL_X1 FILLER_283_1413 ();
 FILLCELL_X8 FILLER_283_1421 ();
 FILLCELL_X4 FILLER_283_1429 ();
 FILLCELL_X2 FILLER_283_1433 ();
 FILLCELL_X8 FILLER_283_1442 ();
 FILLCELL_X2 FILLER_283_1450 ();
 FILLCELL_X8 FILLER_283_1469 ();
 FILLCELL_X1 FILLER_283_1477 ();
 FILLCELL_X4 FILLER_283_1495 ();
 FILLCELL_X32 FILLER_283_1516 ();
 FILLCELL_X8 FILLER_283_1548 ();
 FILLCELL_X1 FILLER_283_1556 ();
 FILLCELL_X8 FILLER_283_1561 ();
 FILLCELL_X4 FILLER_283_1569 ();
 FILLCELL_X2 FILLER_283_1573 ();
 FILLCELL_X1 FILLER_283_1575 ();
 FILLCELL_X8 FILLER_283_1583 ();
 FILLCELL_X1 FILLER_283_1591 ();
 FILLCELL_X4 FILLER_283_1616 ();
 FILLCELL_X4 FILLER_283_1637 ();
 FILLCELL_X1 FILLER_283_1641 ();
 FILLCELL_X4 FILLER_283_1659 ();
 FILLCELL_X2 FILLER_283_1663 ();
 FILLCELL_X8 FILLER_283_1682 ();
 FILLCELL_X4 FILLER_283_1690 ();
 FILLCELL_X1 FILLER_283_1694 ();
 FILLCELL_X8 FILLER_283_1709 ();
 FILLCELL_X1 FILLER_283_1717 ();
 FILLCELL_X4 FILLER_283_1725 ();
 FILLCELL_X2 FILLER_283_1729 ();
 FILLCELL_X1 FILLER_283_1731 ();
 FILLCELL_X32 FILLER_283_1739 ();
 FILLCELL_X32 FILLER_283_1771 ();
 FILLCELL_X32 FILLER_283_1803 ();
 FILLCELL_X32 FILLER_283_1835 ();
 FILLCELL_X32 FILLER_283_1867 ();
 FILLCELL_X32 FILLER_283_1899 ();
 FILLCELL_X32 FILLER_283_1931 ();
 FILLCELL_X32 FILLER_283_1963 ();
 FILLCELL_X32 FILLER_283_1995 ();
 FILLCELL_X32 FILLER_283_2027 ();
 FILLCELL_X32 FILLER_283_2059 ();
 FILLCELL_X32 FILLER_283_2091 ();
 FILLCELL_X32 FILLER_283_2123 ();
 FILLCELL_X32 FILLER_283_2155 ();
 FILLCELL_X32 FILLER_283_2187 ();
 FILLCELL_X32 FILLER_283_2219 ();
 FILLCELL_X32 FILLER_283_2251 ();
 FILLCELL_X32 FILLER_283_2283 ();
 FILLCELL_X32 FILLER_283_2315 ();
 FILLCELL_X32 FILLER_283_2347 ();
 FILLCELL_X32 FILLER_283_2379 ();
 FILLCELL_X32 FILLER_283_2411 ();
 FILLCELL_X32 FILLER_283_2443 ();
 FILLCELL_X32 FILLER_283_2475 ();
 FILLCELL_X16 FILLER_283_2507 ();
 FILLCELL_X2 FILLER_283_2523 ();
 FILLCELL_X1 FILLER_283_2525 ();
 FILLCELL_X32 FILLER_283_2527 ();
 FILLCELL_X32 FILLER_283_2559 ();
 FILLCELL_X32 FILLER_283_2591 ();
 FILLCELL_X32 FILLER_283_2623 ();
 FILLCELL_X32 FILLER_283_2655 ();
 FILLCELL_X32 FILLER_283_2687 ();
 FILLCELL_X32 FILLER_283_2719 ();
 FILLCELL_X32 FILLER_283_2751 ();
 FILLCELL_X32 FILLER_283_2783 ();
 FILLCELL_X32 FILLER_283_2815 ();
 FILLCELL_X32 FILLER_283_2847 ();
 FILLCELL_X32 FILLER_283_2879 ();
 FILLCELL_X32 FILLER_283_2911 ();
 FILLCELL_X32 FILLER_283_2943 ();
 FILLCELL_X32 FILLER_283_2975 ();
 FILLCELL_X32 FILLER_283_3007 ();
 FILLCELL_X32 FILLER_283_3039 ();
 FILLCELL_X32 FILLER_283_3071 ();
 FILLCELL_X32 FILLER_283_3103 ();
 FILLCELL_X32 FILLER_283_3135 ();
 FILLCELL_X32 FILLER_283_3167 ();
 FILLCELL_X32 FILLER_283_3199 ();
 FILLCELL_X32 FILLER_283_3231 ();
 FILLCELL_X32 FILLER_283_3263 ();
 FILLCELL_X32 FILLER_283_3295 ();
 FILLCELL_X32 FILLER_283_3327 ();
 FILLCELL_X32 FILLER_283_3359 ();
 FILLCELL_X32 FILLER_283_3391 ();
 FILLCELL_X32 FILLER_283_3423 ();
 FILLCELL_X32 FILLER_283_3455 ();
 FILLCELL_X32 FILLER_283_3487 ();
 FILLCELL_X32 FILLER_283_3519 ();
 FILLCELL_X32 FILLER_283_3551 ();
 FILLCELL_X32 FILLER_283_3583 ();
 FILLCELL_X32 FILLER_283_3615 ();
 FILLCELL_X32 FILLER_283_3647 ();
 FILLCELL_X32 FILLER_283_3679 ();
 FILLCELL_X16 FILLER_283_3711 ();
 FILLCELL_X8 FILLER_283_3727 ();
 FILLCELL_X2 FILLER_283_3735 ();
 FILLCELL_X1 FILLER_283_3737 ();
 FILLCELL_X32 FILLER_284_1 ();
 FILLCELL_X32 FILLER_284_33 ();
 FILLCELL_X32 FILLER_284_65 ();
 FILLCELL_X32 FILLER_284_97 ();
 FILLCELL_X32 FILLER_284_129 ();
 FILLCELL_X32 FILLER_284_161 ();
 FILLCELL_X32 FILLER_284_193 ();
 FILLCELL_X32 FILLER_284_225 ();
 FILLCELL_X32 FILLER_284_257 ();
 FILLCELL_X32 FILLER_284_289 ();
 FILLCELL_X32 FILLER_284_321 ();
 FILLCELL_X32 FILLER_284_353 ();
 FILLCELL_X32 FILLER_284_385 ();
 FILLCELL_X32 FILLER_284_417 ();
 FILLCELL_X32 FILLER_284_449 ();
 FILLCELL_X32 FILLER_284_481 ();
 FILLCELL_X32 FILLER_284_513 ();
 FILLCELL_X32 FILLER_284_545 ();
 FILLCELL_X32 FILLER_284_577 ();
 FILLCELL_X16 FILLER_284_609 ();
 FILLCELL_X4 FILLER_284_625 ();
 FILLCELL_X2 FILLER_284_629 ();
 FILLCELL_X32 FILLER_284_632 ();
 FILLCELL_X32 FILLER_284_664 ();
 FILLCELL_X32 FILLER_284_696 ();
 FILLCELL_X32 FILLER_284_728 ();
 FILLCELL_X32 FILLER_284_760 ();
 FILLCELL_X32 FILLER_284_792 ();
 FILLCELL_X32 FILLER_284_824 ();
 FILLCELL_X32 FILLER_284_856 ();
 FILLCELL_X32 FILLER_284_888 ();
 FILLCELL_X32 FILLER_284_920 ();
 FILLCELL_X32 FILLER_284_952 ();
 FILLCELL_X32 FILLER_284_984 ();
 FILLCELL_X32 FILLER_284_1016 ();
 FILLCELL_X32 FILLER_284_1048 ();
 FILLCELL_X32 FILLER_284_1080 ();
 FILLCELL_X32 FILLER_284_1112 ();
 FILLCELL_X32 FILLER_284_1144 ();
 FILLCELL_X32 FILLER_284_1176 ();
 FILLCELL_X32 FILLER_284_1208 ();
 FILLCELL_X32 FILLER_284_1240 ();
 FILLCELL_X32 FILLER_284_1272 ();
 FILLCELL_X32 FILLER_284_1304 ();
 FILLCELL_X32 FILLER_284_1336 ();
 FILLCELL_X32 FILLER_284_1368 ();
 FILLCELL_X16 FILLER_284_1400 ();
 FILLCELL_X32 FILLER_284_1440 ();
 FILLCELL_X32 FILLER_284_1472 ();
 FILLCELL_X32 FILLER_284_1504 ();
 FILLCELL_X32 FILLER_284_1536 ();
 FILLCELL_X8 FILLER_284_1585 ();
 FILLCELL_X32 FILLER_284_1600 ();
 FILLCELL_X32 FILLER_284_1632 ();
 FILLCELL_X16 FILLER_284_1664 ();
 FILLCELL_X32 FILLER_284_1688 ();
 FILLCELL_X8 FILLER_284_1720 ();
 FILLCELL_X32 FILLER_284_1745 ();
 FILLCELL_X32 FILLER_284_1777 ();
 FILLCELL_X32 FILLER_284_1809 ();
 FILLCELL_X32 FILLER_284_1841 ();
 FILLCELL_X16 FILLER_284_1873 ();
 FILLCELL_X4 FILLER_284_1889 ();
 FILLCELL_X1 FILLER_284_1893 ();
 FILLCELL_X32 FILLER_284_1895 ();
 FILLCELL_X32 FILLER_284_1927 ();
 FILLCELL_X32 FILLER_284_1959 ();
 FILLCELL_X32 FILLER_284_1991 ();
 FILLCELL_X32 FILLER_284_2023 ();
 FILLCELL_X32 FILLER_284_2055 ();
 FILLCELL_X32 FILLER_284_2087 ();
 FILLCELL_X32 FILLER_284_2119 ();
 FILLCELL_X32 FILLER_284_2151 ();
 FILLCELL_X32 FILLER_284_2183 ();
 FILLCELL_X32 FILLER_284_2215 ();
 FILLCELL_X32 FILLER_284_2247 ();
 FILLCELL_X32 FILLER_284_2279 ();
 FILLCELL_X32 FILLER_284_2311 ();
 FILLCELL_X32 FILLER_284_2343 ();
 FILLCELL_X32 FILLER_284_2375 ();
 FILLCELL_X32 FILLER_284_2407 ();
 FILLCELL_X32 FILLER_284_2439 ();
 FILLCELL_X32 FILLER_284_2471 ();
 FILLCELL_X32 FILLER_284_2503 ();
 FILLCELL_X32 FILLER_284_2535 ();
 FILLCELL_X32 FILLER_284_2567 ();
 FILLCELL_X32 FILLER_284_2599 ();
 FILLCELL_X32 FILLER_284_2631 ();
 FILLCELL_X32 FILLER_284_2663 ();
 FILLCELL_X32 FILLER_284_2695 ();
 FILLCELL_X32 FILLER_284_2727 ();
 FILLCELL_X32 FILLER_284_2759 ();
 FILLCELL_X32 FILLER_284_2791 ();
 FILLCELL_X32 FILLER_284_2823 ();
 FILLCELL_X32 FILLER_284_2855 ();
 FILLCELL_X32 FILLER_284_2887 ();
 FILLCELL_X32 FILLER_284_2919 ();
 FILLCELL_X32 FILLER_284_2951 ();
 FILLCELL_X32 FILLER_284_2983 ();
 FILLCELL_X32 FILLER_284_3015 ();
 FILLCELL_X32 FILLER_284_3047 ();
 FILLCELL_X32 FILLER_284_3079 ();
 FILLCELL_X32 FILLER_284_3111 ();
 FILLCELL_X8 FILLER_284_3143 ();
 FILLCELL_X4 FILLER_284_3151 ();
 FILLCELL_X2 FILLER_284_3155 ();
 FILLCELL_X32 FILLER_284_3158 ();
 FILLCELL_X32 FILLER_284_3190 ();
 FILLCELL_X32 FILLER_284_3222 ();
 FILLCELL_X32 FILLER_284_3254 ();
 FILLCELL_X32 FILLER_284_3286 ();
 FILLCELL_X32 FILLER_284_3318 ();
 FILLCELL_X32 FILLER_284_3350 ();
 FILLCELL_X32 FILLER_284_3382 ();
 FILLCELL_X32 FILLER_284_3414 ();
 FILLCELL_X32 FILLER_284_3446 ();
 FILLCELL_X32 FILLER_284_3478 ();
 FILLCELL_X32 FILLER_284_3510 ();
 FILLCELL_X32 FILLER_284_3542 ();
 FILLCELL_X32 FILLER_284_3574 ();
 FILLCELL_X32 FILLER_284_3606 ();
 FILLCELL_X32 FILLER_284_3638 ();
 FILLCELL_X32 FILLER_284_3670 ();
 FILLCELL_X32 FILLER_284_3702 ();
 FILLCELL_X4 FILLER_284_3734 ();
 FILLCELL_X32 FILLER_285_1 ();
 FILLCELL_X32 FILLER_285_33 ();
 FILLCELL_X32 FILLER_285_65 ();
 FILLCELL_X32 FILLER_285_97 ();
 FILLCELL_X32 FILLER_285_129 ();
 FILLCELL_X32 FILLER_285_161 ();
 FILLCELL_X32 FILLER_285_193 ();
 FILLCELL_X32 FILLER_285_225 ();
 FILLCELL_X32 FILLER_285_257 ();
 FILLCELL_X32 FILLER_285_289 ();
 FILLCELL_X32 FILLER_285_321 ();
 FILLCELL_X32 FILLER_285_353 ();
 FILLCELL_X32 FILLER_285_385 ();
 FILLCELL_X32 FILLER_285_417 ();
 FILLCELL_X32 FILLER_285_449 ();
 FILLCELL_X32 FILLER_285_481 ();
 FILLCELL_X32 FILLER_285_513 ();
 FILLCELL_X32 FILLER_285_545 ();
 FILLCELL_X32 FILLER_285_577 ();
 FILLCELL_X32 FILLER_285_609 ();
 FILLCELL_X32 FILLER_285_641 ();
 FILLCELL_X32 FILLER_285_673 ();
 FILLCELL_X32 FILLER_285_705 ();
 FILLCELL_X32 FILLER_285_737 ();
 FILLCELL_X32 FILLER_285_769 ();
 FILLCELL_X32 FILLER_285_801 ();
 FILLCELL_X32 FILLER_285_833 ();
 FILLCELL_X32 FILLER_285_865 ();
 FILLCELL_X32 FILLER_285_897 ();
 FILLCELL_X32 FILLER_285_929 ();
 FILLCELL_X32 FILLER_285_961 ();
 FILLCELL_X32 FILLER_285_993 ();
 FILLCELL_X32 FILLER_285_1025 ();
 FILLCELL_X32 FILLER_285_1057 ();
 FILLCELL_X32 FILLER_285_1089 ();
 FILLCELL_X32 FILLER_285_1121 ();
 FILLCELL_X32 FILLER_285_1153 ();
 FILLCELL_X32 FILLER_285_1185 ();
 FILLCELL_X32 FILLER_285_1217 ();
 FILLCELL_X8 FILLER_285_1249 ();
 FILLCELL_X4 FILLER_285_1257 ();
 FILLCELL_X2 FILLER_285_1261 ();
 FILLCELL_X32 FILLER_285_1264 ();
 FILLCELL_X32 FILLER_285_1296 ();
 FILLCELL_X32 FILLER_285_1328 ();
 FILLCELL_X32 FILLER_285_1360 ();
 FILLCELL_X32 FILLER_285_1392 ();
 FILLCELL_X32 FILLER_285_1424 ();
 FILLCELL_X4 FILLER_285_1456 ();
 FILLCELL_X2 FILLER_285_1460 ();
 FILLCELL_X32 FILLER_285_1469 ();
 FILLCELL_X8 FILLER_285_1501 ();
 FILLCELL_X4 FILLER_285_1509 ();
 FILLCELL_X2 FILLER_285_1513 ();
 FILLCELL_X1 FILLER_285_1515 ();
 FILLCELL_X1 FILLER_285_1523 ();
 FILLCELL_X1 FILLER_285_1531 ();
 FILLCELL_X16 FILLER_285_1556 ();
 FILLCELL_X8 FILLER_285_1572 ();
 FILLCELL_X2 FILLER_285_1580 ();
 FILLCELL_X1 FILLER_285_1582 ();
 FILLCELL_X32 FILLER_285_1590 ();
 FILLCELL_X32 FILLER_285_1622 ();
 FILLCELL_X32 FILLER_285_1654 ();
 FILLCELL_X4 FILLER_285_1686 ();
 FILLCELL_X1 FILLER_285_1690 ();
 FILLCELL_X8 FILLER_285_1698 ();
 FILLCELL_X2 FILLER_285_1714 ();
 FILLCELL_X32 FILLER_285_1723 ();
 FILLCELL_X32 FILLER_285_1755 ();
 FILLCELL_X32 FILLER_285_1787 ();
 FILLCELL_X32 FILLER_285_1819 ();
 FILLCELL_X32 FILLER_285_1851 ();
 FILLCELL_X32 FILLER_285_1883 ();
 FILLCELL_X32 FILLER_285_1915 ();
 FILLCELL_X32 FILLER_285_1947 ();
 FILLCELL_X32 FILLER_285_1979 ();
 FILLCELL_X32 FILLER_285_2011 ();
 FILLCELL_X32 FILLER_285_2043 ();
 FILLCELL_X32 FILLER_285_2075 ();
 FILLCELL_X32 FILLER_285_2107 ();
 FILLCELL_X32 FILLER_285_2139 ();
 FILLCELL_X32 FILLER_285_2171 ();
 FILLCELL_X32 FILLER_285_2203 ();
 FILLCELL_X32 FILLER_285_2235 ();
 FILLCELL_X32 FILLER_285_2267 ();
 FILLCELL_X32 FILLER_285_2299 ();
 FILLCELL_X32 FILLER_285_2331 ();
 FILLCELL_X32 FILLER_285_2363 ();
 FILLCELL_X32 FILLER_285_2395 ();
 FILLCELL_X32 FILLER_285_2427 ();
 FILLCELL_X32 FILLER_285_2459 ();
 FILLCELL_X32 FILLER_285_2491 ();
 FILLCELL_X2 FILLER_285_2523 ();
 FILLCELL_X1 FILLER_285_2525 ();
 FILLCELL_X32 FILLER_285_2527 ();
 FILLCELL_X32 FILLER_285_2559 ();
 FILLCELL_X32 FILLER_285_2591 ();
 FILLCELL_X32 FILLER_285_2623 ();
 FILLCELL_X32 FILLER_285_2655 ();
 FILLCELL_X32 FILLER_285_2687 ();
 FILLCELL_X32 FILLER_285_2719 ();
 FILLCELL_X32 FILLER_285_2751 ();
 FILLCELL_X32 FILLER_285_2783 ();
 FILLCELL_X32 FILLER_285_2815 ();
 FILLCELL_X32 FILLER_285_2847 ();
 FILLCELL_X32 FILLER_285_2879 ();
 FILLCELL_X32 FILLER_285_2911 ();
 FILLCELL_X32 FILLER_285_2943 ();
 FILLCELL_X32 FILLER_285_2975 ();
 FILLCELL_X32 FILLER_285_3007 ();
 FILLCELL_X32 FILLER_285_3039 ();
 FILLCELL_X32 FILLER_285_3071 ();
 FILLCELL_X32 FILLER_285_3103 ();
 FILLCELL_X32 FILLER_285_3135 ();
 FILLCELL_X32 FILLER_285_3167 ();
 FILLCELL_X32 FILLER_285_3199 ();
 FILLCELL_X32 FILLER_285_3231 ();
 FILLCELL_X32 FILLER_285_3263 ();
 FILLCELL_X32 FILLER_285_3295 ();
 FILLCELL_X32 FILLER_285_3327 ();
 FILLCELL_X32 FILLER_285_3359 ();
 FILLCELL_X32 FILLER_285_3391 ();
 FILLCELL_X32 FILLER_285_3423 ();
 FILLCELL_X32 FILLER_285_3455 ();
 FILLCELL_X32 FILLER_285_3487 ();
 FILLCELL_X32 FILLER_285_3519 ();
 FILLCELL_X32 FILLER_285_3551 ();
 FILLCELL_X32 FILLER_285_3583 ();
 FILLCELL_X32 FILLER_285_3615 ();
 FILLCELL_X32 FILLER_285_3647 ();
 FILLCELL_X32 FILLER_285_3679 ();
 FILLCELL_X16 FILLER_285_3711 ();
 FILLCELL_X8 FILLER_285_3727 ();
 FILLCELL_X2 FILLER_285_3735 ();
 FILLCELL_X1 FILLER_285_3737 ();
 FILLCELL_X32 FILLER_286_1 ();
 FILLCELL_X32 FILLER_286_33 ();
 FILLCELL_X32 FILLER_286_65 ();
 FILLCELL_X32 FILLER_286_97 ();
 FILLCELL_X32 FILLER_286_129 ();
 FILLCELL_X32 FILLER_286_161 ();
 FILLCELL_X32 FILLER_286_193 ();
 FILLCELL_X32 FILLER_286_225 ();
 FILLCELL_X32 FILLER_286_257 ();
 FILLCELL_X32 FILLER_286_289 ();
 FILLCELL_X32 FILLER_286_321 ();
 FILLCELL_X32 FILLER_286_353 ();
 FILLCELL_X32 FILLER_286_385 ();
 FILLCELL_X32 FILLER_286_417 ();
 FILLCELL_X32 FILLER_286_449 ();
 FILLCELL_X32 FILLER_286_481 ();
 FILLCELL_X32 FILLER_286_513 ();
 FILLCELL_X32 FILLER_286_545 ();
 FILLCELL_X32 FILLER_286_577 ();
 FILLCELL_X16 FILLER_286_609 ();
 FILLCELL_X4 FILLER_286_625 ();
 FILLCELL_X2 FILLER_286_629 ();
 FILLCELL_X32 FILLER_286_632 ();
 FILLCELL_X32 FILLER_286_664 ();
 FILLCELL_X32 FILLER_286_696 ();
 FILLCELL_X32 FILLER_286_728 ();
 FILLCELL_X32 FILLER_286_760 ();
 FILLCELL_X32 FILLER_286_792 ();
 FILLCELL_X32 FILLER_286_824 ();
 FILLCELL_X32 FILLER_286_856 ();
 FILLCELL_X32 FILLER_286_888 ();
 FILLCELL_X32 FILLER_286_920 ();
 FILLCELL_X32 FILLER_286_952 ();
 FILLCELL_X32 FILLER_286_984 ();
 FILLCELL_X32 FILLER_286_1016 ();
 FILLCELL_X32 FILLER_286_1048 ();
 FILLCELL_X32 FILLER_286_1080 ();
 FILLCELL_X32 FILLER_286_1112 ();
 FILLCELL_X32 FILLER_286_1144 ();
 FILLCELL_X32 FILLER_286_1176 ();
 FILLCELL_X32 FILLER_286_1208 ();
 FILLCELL_X32 FILLER_286_1240 ();
 FILLCELL_X32 FILLER_286_1272 ();
 FILLCELL_X32 FILLER_286_1304 ();
 FILLCELL_X32 FILLER_286_1336 ();
 FILLCELL_X32 FILLER_286_1368 ();
 FILLCELL_X32 FILLER_286_1400 ();
 FILLCELL_X16 FILLER_286_1432 ();
 FILLCELL_X16 FILLER_286_1472 ();
 FILLCELL_X4 FILLER_286_1488 ();
 FILLCELL_X8 FILLER_286_1499 ();
 FILLCELL_X2 FILLER_286_1507 ();
 FILLCELL_X1 FILLER_286_1509 ();
 FILLCELL_X32 FILLER_286_1527 ();
 FILLCELL_X16 FILLER_286_1559 ();
 FILLCELL_X4 FILLER_286_1575 ();
 FILLCELL_X1 FILLER_286_1579 ();
 FILLCELL_X4 FILLER_286_1597 ();
 FILLCELL_X2 FILLER_286_1601 ();
 FILLCELL_X1 FILLER_286_1603 ();
 FILLCELL_X8 FILLER_286_1611 ();
 FILLCELL_X1 FILLER_286_1619 ();
 FILLCELL_X16 FILLER_286_1634 ();
 FILLCELL_X2 FILLER_286_1657 ();
 FILLCELL_X2 FILLER_286_1666 ();
 FILLCELL_X8 FILLER_286_1675 ();
 FILLCELL_X4 FILLER_286_1683 ();
 FILLCELL_X2 FILLER_286_1687 ();
 FILLCELL_X1 FILLER_286_1689 ();
 FILLCELL_X8 FILLER_286_1707 ();
 FILLCELL_X32 FILLER_286_1735 ();
 FILLCELL_X32 FILLER_286_1767 ();
 FILLCELL_X32 FILLER_286_1799 ();
 FILLCELL_X32 FILLER_286_1831 ();
 FILLCELL_X16 FILLER_286_1863 ();
 FILLCELL_X8 FILLER_286_1879 ();
 FILLCELL_X4 FILLER_286_1887 ();
 FILLCELL_X2 FILLER_286_1891 ();
 FILLCELL_X1 FILLER_286_1893 ();
 FILLCELL_X32 FILLER_286_1895 ();
 FILLCELL_X32 FILLER_286_1927 ();
 FILLCELL_X32 FILLER_286_1959 ();
 FILLCELL_X32 FILLER_286_1991 ();
 FILLCELL_X32 FILLER_286_2023 ();
 FILLCELL_X32 FILLER_286_2055 ();
 FILLCELL_X32 FILLER_286_2087 ();
 FILLCELL_X32 FILLER_286_2119 ();
 FILLCELL_X32 FILLER_286_2151 ();
 FILLCELL_X32 FILLER_286_2183 ();
 FILLCELL_X32 FILLER_286_2215 ();
 FILLCELL_X32 FILLER_286_2247 ();
 FILLCELL_X32 FILLER_286_2279 ();
 FILLCELL_X32 FILLER_286_2311 ();
 FILLCELL_X32 FILLER_286_2343 ();
 FILLCELL_X32 FILLER_286_2375 ();
 FILLCELL_X32 FILLER_286_2407 ();
 FILLCELL_X32 FILLER_286_2439 ();
 FILLCELL_X32 FILLER_286_2471 ();
 FILLCELL_X32 FILLER_286_2503 ();
 FILLCELL_X32 FILLER_286_2535 ();
 FILLCELL_X32 FILLER_286_2567 ();
 FILLCELL_X32 FILLER_286_2599 ();
 FILLCELL_X32 FILLER_286_2631 ();
 FILLCELL_X32 FILLER_286_2663 ();
 FILLCELL_X32 FILLER_286_2695 ();
 FILLCELL_X32 FILLER_286_2727 ();
 FILLCELL_X32 FILLER_286_2759 ();
 FILLCELL_X32 FILLER_286_2791 ();
 FILLCELL_X32 FILLER_286_2823 ();
 FILLCELL_X32 FILLER_286_2855 ();
 FILLCELL_X32 FILLER_286_2887 ();
 FILLCELL_X32 FILLER_286_2919 ();
 FILLCELL_X32 FILLER_286_2951 ();
 FILLCELL_X32 FILLER_286_2983 ();
 FILLCELL_X32 FILLER_286_3015 ();
 FILLCELL_X32 FILLER_286_3047 ();
 FILLCELL_X32 FILLER_286_3079 ();
 FILLCELL_X32 FILLER_286_3111 ();
 FILLCELL_X8 FILLER_286_3143 ();
 FILLCELL_X4 FILLER_286_3151 ();
 FILLCELL_X2 FILLER_286_3155 ();
 FILLCELL_X32 FILLER_286_3158 ();
 FILLCELL_X32 FILLER_286_3190 ();
 FILLCELL_X32 FILLER_286_3222 ();
 FILLCELL_X32 FILLER_286_3254 ();
 FILLCELL_X32 FILLER_286_3286 ();
 FILLCELL_X32 FILLER_286_3318 ();
 FILLCELL_X32 FILLER_286_3350 ();
 FILLCELL_X32 FILLER_286_3382 ();
 FILLCELL_X32 FILLER_286_3414 ();
 FILLCELL_X32 FILLER_286_3446 ();
 FILLCELL_X32 FILLER_286_3478 ();
 FILLCELL_X32 FILLER_286_3510 ();
 FILLCELL_X32 FILLER_286_3542 ();
 FILLCELL_X32 FILLER_286_3574 ();
 FILLCELL_X32 FILLER_286_3606 ();
 FILLCELL_X32 FILLER_286_3638 ();
 FILLCELL_X32 FILLER_286_3670 ();
 FILLCELL_X32 FILLER_286_3702 ();
 FILLCELL_X4 FILLER_286_3734 ();
 FILLCELL_X32 FILLER_287_1 ();
 FILLCELL_X32 FILLER_287_33 ();
 FILLCELL_X32 FILLER_287_65 ();
 FILLCELL_X32 FILLER_287_97 ();
 FILLCELL_X32 FILLER_287_129 ();
 FILLCELL_X32 FILLER_287_161 ();
 FILLCELL_X32 FILLER_287_193 ();
 FILLCELL_X32 FILLER_287_225 ();
 FILLCELL_X32 FILLER_287_257 ();
 FILLCELL_X32 FILLER_287_289 ();
 FILLCELL_X32 FILLER_287_321 ();
 FILLCELL_X32 FILLER_287_353 ();
 FILLCELL_X32 FILLER_287_385 ();
 FILLCELL_X32 FILLER_287_417 ();
 FILLCELL_X32 FILLER_287_449 ();
 FILLCELL_X32 FILLER_287_481 ();
 FILLCELL_X32 FILLER_287_513 ();
 FILLCELL_X32 FILLER_287_545 ();
 FILLCELL_X32 FILLER_287_577 ();
 FILLCELL_X32 FILLER_287_609 ();
 FILLCELL_X32 FILLER_287_641 ();
 FILLCELL_X32 FILLER_287_673 ();
 FILLCELL_X32 FILLER_287_705 ();
 FILLCELL_X32 FILLER_287_737 ();
 FILLCELL_X32 FILLER_287_769 ();
 FILLCELL_X32 FILLER_287_801 ();
 FILLCELL_X32 FILLER_287_833 ();
 FILLCELL_X32 FILLER_287_865 ();
 FILLCELL_X32 FILLER_287_897 ();
 FILLCELL_X32 FILLER_287_929 ();
 FILLCELL_X32 FILLER_287_961 ();
 FILLCELL_X32 FILLER_287_993 ();
 FILLCELL_X32 FILLER_287_1025 ();
 FILLCELL_X32 FILLER_287_1057 ();
 FILLCELL_X32 FILLER_287_1089 ();
 FILLCELL_X32 FILLER_287_1121 ();
 FILLCELL_X32 FILLER_287_1153 ();
 FILLCELL_X32 FILLER_287_1185 ();
 FILLCELL_X32 FILLER_287_1217 ();
 FILLCELL_X8 FILLER_287_1249 ();
 FILLCELL_X4 FILLER_287_1257 ();
 FILLCELL_X2 FILLER_287_1261 ();
 FILLCELL_X32 FILLER_287_1264 ();
 FILLCELL_X32 FILLER_287_1296 ();
 FILLCELL_X32 FILLER_287_1328 ();
 FILLCELL_X32 FILLER_287_1360 ();
 FILLCELL_X32 FILLER_287_1392 ();
 FILLCELL_X16 FILLER_287_1424 ();
 FILLCELL_X8 FILLER_287_1440 ();
 FILLCELL_X4 FILLER_287_1448 ();
 FILLCELL_X1 FILLER_287_1459 ();
 FILLCELL_X32 FILLER_287_1467 ();
 FILLCELL_X2 FILLER_287_1499 ();
 FILLCELL_X1 FILLER_287_1501 ();
 FILLCELL_X32 FILLER_287_1519 ();
 FILLCELL_X32 FILLER_287_1551 ();
 FILLCELL_X16 FILLER_287_1583 ();
 FILLCELL_X1 FILLER_287_1599 ();
 FILLCELL_X8 FILLER_287_1617 ();
 FILLCELL_X2 FILLER_287_1642 ();
 FILLCELL_X8 FILLER_287_1661 ();
 FILLCELL_X1 FILLER_287_1669 ();
 FILLCELL_X32 FILLER_287_1687 ();
 FILLCELL_X32 FILLER_287_1719 ();
 FILLCELL_X32 FILLER_287_1751 ();
 FILLCELL_X32 FILLER_287_1783 ();
 FILLCELL_X32 FILLER_287_1815 ();
 FILLCELL_X32 FILLER_287_1847 ();
 FILLCELL_X32 FILLER_287_1879 ();
 FILLCELL_X32 FILLER_287_1911 ();
 FILLCELL_X32 FILLER_287_1943 ();
 FILLCELL_X32 FILLER_287_1975 ();
 FILLCELL_X32 FILLER_287_2007 ();
 FILLCELL_X32 FILLER_287_2039 ();
 FILLCELL_X32 FILLER_287_2071 ();
 FILLCELL_X32 FILLER_287_2103 ();
 FILLCELL_X32 FILLER_287_2135 ();
 FILLCELL_X32 FILLER_287_2167 ();
 FILLCELL_X32 FILLER_287_2199 ();
 FILLCELL_X32 FILLER_287_2231 ();
 FILLCELL_X32 FILLER_287_2263 ();
 FILLCELL_X32 FILLER_287_2295 ();
 FILLCELL_X32 FILLER_287_2327 ();
 FILLCELL_X32 FILLER_287_2359 ();
 FILLCELL_X32 FILLER_287_2391 ();
 FILLCELL_X32 FILLER_287_2423 ();
 FILLCELL_X32 FILLER_287_2455 ();
 FILLCELL_X32 FILLER_287_2487 ();
 FILLCELL_X4 FILLER_287_2519 ();
 FILLCELL_X2 FILLER_287_2523 ();
 FILLCELL_X1 FILLER_287_2525 ();
 FILLCELL_X32 FILLER_287_2527 ();
 FILLCELL_X32 FILLER_287_2559 ();
 FILLCELL_X32 FILLER_287_2591 ();
 FILLCELL_X32 FILLER_287_2623 ();
 FILLCELL_X32 FILLER_287_2655 ();
 FILLCELL_X32 FILLER_287_2687 ();
 FILLCELL_X32 FILLER_287_2719 ();
 FILLCELL_X32 FILLER_287_2751 ();
 FILLCELL_X32 FILLER_287_2783 ();
 FILLCELL_X32 FILLER_287_2815 ();
 FILLCELL_X32 FILLER_287_2847 ();
 FILLCELL_X32 FILLER_287_2879 ();
 FILLCELL_X32 FILLER_287_2911 ();
 FILLCELL_X32 FILLER_287_2943 ();
 FILLCELL_X32 FILLER_287_2975 ();
 FILLCELL_X32 FILLER_287_3007 ();
 FILLCELL_X32 FILLER_287_3039 ();
 FILLCELL_X32 FILLER_287_3071 ();
 FILLCELL_X32 FILLER_287_3103 ();
 FILLCELL_X32 FILLER_287_3135 ();
 FILLCELL_X32 FILLER_287_3167 ();
 FILLCELL_X32 FILLER_287_3199 ();
 FILLCELL_X32 FILLER_287_3231 ();
 FILLCELL_X32 FILLER_287_3263 ();
 FILLCELL_X32 FILLER_287_3295 ();
 FILLCELL_X32 FILLER_287_3327 ();
 FILLCELL_X32 FILLER_287_3359 ();
 FILLCELL_X32 FILLER_287_3391 ();
 FILLCELL_X32 FILLER_287_3423 ();
 FILLCELL_X32 FILLER_287_3455 ();
 FILLCELL_X32 FILLER_287_3487 ();
 FILLCELL_X32 FILLER_287_3519 ();
 FILLCELL_X32 FILLER_287_3551 ();
 FILLCELL_X32 FILLER_287_3583 ();
 FILLCELL_X32 FILLER_287_3615 ();
 FILLCELL_X32 FILLER_287_3647 ();
 FILLCELL_X32 FILLER_287_3679 ();
 FILLCELL_X16 FILLER_287_3711 ();
 FILLCELL_X8 FILLER_287_3727 ();
 FILLCELL_X2 FILLER_287_3735 ();
 FILLCELL_X1 FILLER_287_3737 ();
 FILLCELL_X32 FILLER_288_1 ();
 FILLCELL_X32 FILLER_288_33 ();
 FILLCELL_X32 FILLER_288_65 ();
 FILLCELL_X32 FILLER_288_97 ();
 FILLCELL_X32 FILLER_288_129 ();
 FILLCELL_X32 FILLER_288_161 ();
 FILLCELL_X32 FILLER_288_193 ();
 FILLCELL_X32 FILLER_288_225 ();
 FILLCELL_X32 FILLER_288_257 ();
 FILLCELL_X32 FILLER_288_289 ();
 FILLCELL_X32 FILLER_288_321 ();
 FILLCELL_X32 FILLER_288_353 ();
 FILLCELL_X32 FILLER_288_385 ();
 FILLCELL_X32 FILLER_288_417 ();
 FILLCELL_X32 FILLER_288_449 ();
 FILLCELL_X32 FILLER_288_481 ();
 FILLCELL_X32 FILLER_288_513 ();
 FILLCELL_X32 FILLER_288_545 ();
 FILLCELL_X32 FILLER_288_577 ();
 FILLCELL_X16 FILLER_288_609 ();
 FILLCELL_X4 FILLER_288_625 ();
 FILLCELL_X2 FILLER_288_629 ();
 FILLCELL_X32 FILLER_288_632 ();
 FILLCELL_X32 FILLER_288_664 ();
 FILLCELL_X32 FILLER_288_696 ();
 FILLCELL_X32 FILLER_288_728 ();
 FILLCELL_X32 FILLER_288_760 ();
 FILLCELL_X32 FILLER_288_792 ();
 FILLCELL_X32 FILLER_288_824 ();
 FILLCELL_X32 FILLER_288_856 ();
 FILLCELL_X32 FILLER_288_888 ();
 FILLCELL_X32 FILLER_288_920 ();
 FILLCELL_X32 FILLER_288_952 ();
 FILLCELL_X32 FILLER_288_984 ();
 FILLCELL_X32 FILLER_288_1016 ();
 FILLCELL_X32 FILLER_288_1048 ();
 FILLCELL_X32 FILLER_288_1080 ();
 FILLCELL_X32 FILLER_288_1112 ();
 FILLCELL_X32 FILLER_288_1144 ();
 FILLCELL_X32 FILLER_288_1176 ();
 FILLCELL_X32 FILLER_288_1208 ();
 FILLCELL_X32 FILLER_288_1240 ();
 FILLCELL_X32 FILLER_288_1272 ();
 FILLCELL_X32 FILLER_288_1304 ();
 FILLCELL_X32 FILLER_288_1336 ();
 FILLCELL_X32 FILLER_288_1368 ();
 FILLCELL_X32 FILLER_288_1400 ();
 FILLCELL_X16 FILLER_288_1432 ();
 FILLCELL_X8 FILLER_288_1448 ();
 FILLCELL_X4 FILLER_288_1456 ();
 FILLCELL_X1 FILLER_288_1460 ();
 FILLCELL_X32 FILLER_288_1478 ();
 FILLCELL_X4 FILLER_288_1510 ();
 FILLCELL_X2 FILLER_288_1514 ();
 FILLCELL_X8 FILLER_288_1530 ();
 FILLCELL_X2 FILLER_288_1538 ();
 FILLCELL_X32 FILLER_288_1547 ();
 FILLCELL_X32 FILLER_288_1579 ();
 FILLCELL_X32 FILLER_288_1611 ();
 FILLCELL_X32 FILLER_288_1643 ();
 FILLCELL_X32 FILLER_288_1675 ();
 FILLCELL_X32 FILLER_288_1707 ();
 FILLCELL_X32 FILLER_288_1739 ();
 FILLCELL_X32 FILLER_288_1771 ();
 FILLCELL_X32 FILLER_288_1803 ();
 FILLCELL_X32 FILLER_288_1835 ();
 FILLCELL_X16 FILLER_288_1867 ();
 FILLCELL_X8 FILLER_288_1883 ();
 FILLCELL_X2 FILLER_288_1891 ();
 FILLCELL_X1 FILLER_288_1893 ();
 FILLCELL_X32 FILLER_288_1895 ();
 FILLCELL_X32 FILLER_288_1927 ();
 FILLCELL_X32 FILLER_288_1959 ();
 FILLCELL_X32 FILLER_288_1991 ();
 FILLCELL_X32 FILLER_288_2023 ();
 FILLCELL_X32 FILLER_288_2055 ();
 FILLCELL_X32 FILLER_288_2087 ();
 FILLCELL_X32 FILLER_288_2119 ();
 FILLCELL_X32 FILLER_288_2151 ();
 FILLCELL_X32 FILLER_288_2183 ();
 FILLCELL_X32 FILLER_288_2215 ();
 FILLCELL_X32 FILLER_288_2247 ();
 FILLCELL_X32 FILLER_288_2279 ();
 FILLCELL_X32 FILLER_288_2311 ();
 FILLCELL_X32 FILLER_288_2343 ();
 FILLCELL_X32 FILLER_288_2375 ();
 FILLCELL_X32 FILLER_288_2407 ();
 FILLCELL_X32 FILLER_288_2439 ();
 FILLCELL_X32 FILLER_288_2471 ();
 FILLCELL_X32 FILLER_288_2503 ();
 FILLCELL_X32 FILLER_288_2535 ();
 FILLCELL_X32 FILLER_288_2567 ();
 FILLCELL_X32 FILLER_288_2599 ();
 FILLCELL_X32 FILLER_288_2631 ();
 FILLCELL_X32 FILLER_288_2663 ();
 FILLCELL_X32 FILLER_288_2695 ();
 FILLCELL_X32 FILLER_288_2727 ();
 FILLCELL_X32 FILLER_288_2759 ();
 FILLCELL_X32 FILLER_288_2791 ();
 FILLCELL_X32 FILLER_288_2823 ();
 FILLCELL_X32 FILLER_288_2855 ();
 FILLCELL_X32 FILLER_288_2887 ();
 FILLCELL_X32 FILLER_288_2919 ();
 FILLCELL_X32 FILLER_288_2951 ();
 FILLCELL_X32 FILLER_288_2983 ();
 FILLCELL_X32 FILLER_288_3015 ();
 FILLCELL_X32 FILLER_288_3047 ();
 FILLCELL_X32 FILLER_288_3079 ();
 FILLCELL_X32 FILLER_288_3111 ();
 FILLCELL_X8 FILLER_288_3143 ();
 FILLCELL_X4 FILLER_288_3151 ();
 FILLCELL_X2 FILLER_288_3155 ();
 FILLCELL_X32 FILLER_288_3158 ();
 FILLCELL_X32 FILLER_288_3190 ();
 FILLCELL_X32 FILLER_288_3222 ();
 FILLCELL_X32 FILLER_288_3254 ();
 FILLCELL_X32 FILLER_288_3286 ();
 FILLCELL_X32 FILLER_288_3318 ();
 FILLCELL_X32 FILLER_288_3350 ();
 FILLCELL_X32 FILLER_288_3382 ();
 FILLCELL_X32 FILLER_288_3414 ();
 FILLCELL_X32 FILLER_288_3446 ();
 FILLCELL_X32 FILLER_288_3478 ();
 FILLCELL_X32 FILLER_288_3510 ();
 FILLCELL_X32 FILLER_288_3542 ();
 FILLCELL_X32 FILLER_288_3574 ();
 FILLCELL_X32 FILLER_288_3606 ();
 FILLCELL_X32 FILLER_288_3638 ();
 FILLCELL_X32 FILLER_288_3670 ();
 FILLCELL_X32 FILLER_288_3702 ();
 FILLCELL_X4 FILLER_288_3734 ();
 FILLCELL_X32 FILLER_289_1 ();
 FILLCELL_X32 FILLER_289_33 ();
 FILLCELL_X32 FILLER_289_65 ();
 FILLCELL_X32 FILLER_289_97 ();
 FILLCELL_X32 FILLER_289_129 ();
 FILLCELL_X32 FILLER_289_161 ();
 FILLCELL_X32 FILLER_289_193 ();
 FILLCELL_X32 FILLER_289_225 ();
 FILLCELL_X32 FILLER_289_257 ();
 FILLCELL_X32 FILLER_289_289 ();
 FILLCELL_X32 FILLER_289_321 ();
 FILLCELL_X32 FILLER_289_353 ();
 FILLCELL_X32 FILLER_289_385 ();
 FILLCELL_X32 FILLER_289_417 ();
 FILLCELL_X32 FILLER_289_449 ();
 FILLCELL_X32 FILLER_289_481 ();
 FILLCELL_X32 FILLER_289_513 ();
 FILLCELL_X32 FILLER_289_545 ();
 FILLCELL_X32 FILLER_289_577 ();
 FILLCELL_X32 FILLER_289_609 ();
 FILLCELL_X32 FILLER_289_641 ();
 FILLCELL_X32 FILLER_289_673 ();
 FILLCELL_X32 FILLER_289_705 ();
 FILLCELL_X32 FILLER_289_737 ();
 FILLCELL_X32 FILLER_289_769 ();
 FILLCELL_X32 FILLER_289_801 ();
 FILLCELL_X32 FILLER_289_833 ();
 FILLCELL_X32 FILLER_289_865 ();
 FILLCELL_X32 FILLER_289_897 ();
 FILLCELL_X32 FILLER_289_929 ();
 FILLCELL_X32 FILLER_289_961 ();
 FILLCELL_X32 FILLER_289_993 ();
 FILLCELL_X32 FILLER_289_1025 ();
 FILLCELL_X32 FILLER_289_1057 ();
 FILLCELL_X32 FILLER_289_1089 ();
 FILLCELL_X32 FILLER_289_1121 ();
 FILLCELL_X32 FILLER_289_1153 ();
 FILLCELL_X32 FILLER_289_1185 ();
 FILLCELL_X32 FILLER_289_1217 ();
 FILLCELL_X8 FILLER_289_1249 ();
 FILLCELL_X4 FILLER_289_1257 ();
 FILLCELL_X2 FILLER_289_1261 ();
 FILLCELL_X32 FILLER_289_1264 ();
 FILLCELL_X32 FILLER_289_1296 ();
 FILLCELL_X32 FILLER_289_1328 ();
 FILLCELL_X32 FILLER_289_1360 ();
 FILLCELL_X32 FILLER_289_1392 ();
 FILLCELL_X32 FILLER_289_1424 ();
 FILLCELL_X32 FILLER_289_1456 ();
 FILLCELL_X16 FILLER_289_1488 ();
 FILLCELL_X4 FILLER_289_1504 ();
 FILLCELL_X1 FILLER_289_1508 ();
 FILLCELL_X8 FILLER_289_1526 ();
 FILLCELL_X4 FILLER_289_1534 ();
 FILLCELL_X1 FILLER_289_1538 ();
 FILLCELL_X8 FILLER_289_1556 ();
 FILLCELL_X4 FILLER_289_1564 ();
 FILLCELL_X2 FILLER_289_1568 ();
 FILLCELL_X1 FILLER_289_1570 ();
 FILLCELL_X4 FILLER_289_1579 ();
 FILLCELL_X1 FILLER_289_1583 ();
 FILLCELL_X8 FILLER_289_1588 ();
 FILLCELL_X4 FILLER_289_1596 ();
 FILLCELL_X2 FILLER_289_1600 ();
 FILLCELL_X32 FILLER_289_1619 ();
 FILLCELL_X32 FILLER_289_1675 ();
 FILLCELL_X32 FILLER_289_1707 ();
 FILLCELL_X32 FILLER_289_1739 ();
 FILLCELL_X16 FILLER_289_1771 ();
 FILLCELL_X8 FILLER_289_1787 ();
 FILLCELL_X32 FILLER_289_1799 ();
 FILLCELL_X32 FILLER_289_1831 ();
 FILLCELL_X32 FILLER_289_1863 ();
 FILLCELL_X32 FILLER_289_1895 ();
 FILLCELL_X32 FILLER_289_1927 ();
 FILLCELL_X32 FILLER_289_1959 ();
 FILLCELL_X32 FILLER_289_1991 ();
 FILLCELL_X32 FILLER_289_2023 ();
 FILLCELL_X32 FILLER_289_2055 ();
 FILLCELL_X32 FILLER_289_2087 ();
 FILLCELL_X32 FILLER_289_2119 ();
 FILLCELL_X32 FILLER_289_2151 ();
 FILLCELL_X32 FILLER_289_2183 ();
 FILLCELL_X32 FILLER_289_2215 ();
 FILLCELL_X32 FILLER_289_2247 ();
 FILLCELL_X32 FILLER_289_2279 ();
 FILLCELL_X32 FILLER_289_2311 ();
 FILLCELL_X32 FILLER_289_2343 ();
 FILLCELL_X32 FILLER_289_2375 ();
 FILLCELL_X32 FILLER_289_2407 ();
 FILLCELL_X32 FILLER_289_2439 ();
 FILLCELL_X32 FILLER_289_2471 ();
 FILLCELL_X16 FILLER_289_2503 ();
 FILLCELL_X4 FILLER_289_2519 ();
 FILLCELL_X2 FILLER_289_2523 ();
 FILLCELL_X1 FILLER_289_2525 ();
 FILLCELL_X32 FILLER_289_2527 ();
 FILLCELL_X32 FILLER_289_2559 ();
 FILLCELL_X32 FILLER_289_2591 ();
 FILLCELL_X32 FILLER_289_2623 ();
 FILLCELL_X32 FILLER_289_2655 ();
 FILLCELL_X32 FILLER_289_2687 ();
 FILLCELL_X32 FILLER_289_2719 ();
 FILLCELL_X32 FILLER_289_2751 ();
 FILLCELL_X32 FILLER_289_2783 ();
 FILLCELL_X32 FILLER_289_2815 ();
 FILLCELL_X32 FILLER_289_2847 ();
 FILLCELL_X32 FILLER_289_2879 ();
 FILLCELL_X32 FILLER_289_2911 ();
 FILLCELL_X32 FILLER_289_2943 ();
 FILLCELL_X32 FILLER_289_2975 ();
 FILLCELL_X32 FILLER_289_3007 ();
 FILLCELL_X32 FILLER_289_3039 ();
 FILLCELL_X32 FILLER_289_3071 ();
 FILLCELL_X32 FILLER_289_3103 ();
 FILLCELL_X32 FILLER_289_3135 ();
 FILLCELL_X32 FILLER_289_3167 ();
 FILLCELL_X32 FILLER_289_3199 ();
 FILLCELL_X32 FILLER_289_3231 ();
 FILLCELL_X32 FILLER_289_3263 ();
 FILLCELL_X32 FILLER_289_3295 ();
 FILLCELL_X32 FILLER_289_3327 ();
 FILLCELL_X32 FILLER_289_3359 ();
 FILLCELL_X32 FILLER_289_3391 ();
 FILLCELL_X32 FILLER_289_3423 ();
 FILLCELL_X32 FILLER_289_3455 ();
 FILLCELL_X32 FILLER_289_3487 ();
 FILLCELL_X32 FILLER_289_3519 ();
 FILLCELL_X32 FILLER_289_3551 ();
 FILLCELL_X32 FILLER_289_3583 ();
 FILLCELL_X32 FILLER_289_3615 ();
 FILLCELL_X32 FILLER_289_3647 ();
 FILLCELL_X32 FILLER_289_3679 ();
 FILLCELL_X16 FILLER_289_3711 ();
 FILLCELL_X8 FILLER_289_3727 ();
 FILLCELL_X2 FILLER_289_3735 ();
 FILLCELL_X1 FILLER_289_3737 ();
 FILLCELL_X32 FILLER_290_1 ();
 FILLCELL_X32 FILLER_290_33 ();
 FILLCELL_X32 FILLER_290_65 ();
 FILLCELL_X32 FILLER_290_97 ();
 FILLCELL_X32 FILLER_290_129 ();
 FILLCELL_X32 FILLER_290_161 ();
 FILLCELL_X32 FILLER_290_193 ();
 FILLCELL_X32 FILLER_290_225 ();
 FILLCELL_X32 FILLER_290_257 ();
 FILLCELL_X32 FILLER_290_289 ();
 FILLCELL_X32 FILLER_290_321 ();
 FILLCELL_X32 FILLER_290_353 ();
 FILLCELL_X32 FILLER_290_385 ();
 FILLCELL_X32 FILLER_290_417 ();
 FILLCELL_X32 FILLER_290_449 ();
 FILLCELL_X32 FILLER_290_481 ();
 FILLCELL_X32 FILLER_290_513 ();
 FILLCELL_X32 FILLER_290_545 ();
 FILLCELL_X32 FILLER_290_577 ();
 FILLCELL_X16 FILLER_290_609 ();
 FILLCELL_X4 FILLER_290_625 ();
 FILLCELL_X2 FILLER_290_629 ();
 FILLCELL_X32 FILLER_290_632 ();
 FILLCELL_X32 FILLER_290_664 ();
 FILLCELL_X32 FILLER_290_696 ();
 FILLCELL_X32 FILLER_290_728 ();
 FILLCELL_X32 FILLER_290_760 ();
 FILLCELL_X32 FILLER_290_792 ();
 FILLCELL_X32 FILLER_290_824 ();
 FILLCELL_X32 FILLER_290_856 ();
 FILLCELL_X32 FILLER_290_888 ();
 FILLCELL_X32 FILLER_290_920 ();
 FILLCELL_X32 FILLER_290_952 ();
 FILLCELL_X32 FILLER_290_984 ();
 FILLCELL_X32 FILLER_290_1016 ();
 FILLCELL_X32 FILLER_290_1048 ();
 FILLCELL_X32 FILLER_290_1080 ();
 FILLCELL_X32 FILLER_290_1112 ();
 FILLCELL_X32 FILLER_290_1144 ();
 FILLCELL_X32 FILLER_290_1176 ();
 FILLCELL_X32 FILLER_290_1208 ();
 FILLCELL_X32 FILLER_290_1240 ();
 FILLCELL_X32 FILLER_290_1272 ();
 FILLCELL_X32 FILLER_290_1304 ();
 FILLCELL_X32 FILLER_290_1336 ();
 FILLCELL_X32 FILLER_290_1368 ();
 FILLCELL_X32 FILLER_290_1400 ();
 FILLCELL_X32 FILLER_290_1432 ();
 FILLCELL_X32 FILLER_290_1464 ();
 FILLCELL_X32 FILLER_290_1496 ();
 FILLCELL_X32 FILLER_290_1528 ();
 FILLCELL_X32 FILLER_290_1560 ();
 FILLCELL_X8 FILLER_290_1592 ();
 FILLCELL_X4 FILLER_290_1600 ();
 FILLCELL_X4 FILLER_290_1611 ();
 FILLCELL_X2 FILLER_290_1615 ();
 FILLCELL_X16 FILLER_290_1624 ();
 FILLCELL_X4 FILLER_290_1640 ();
 FILLCELL_X2 FILLER_290_1644 ();
 FILLCELL_X1 FILLER_290_1646 ();
 FILLCELL_X2 FILLER_290_1654 ();
 FILLCELL_X1 FILLER_290_1656 ();
 FILLCELL_X32 FILLER_290_1664 ();
 FILLCELL_X32 FILLER_290_1696 ();
 FILLCELL_X32 FILLER_290_1728 ();
 FILLCELL_X32 FILLER_290_1760 ();
 FILLCELL_X32 FILLER_290_1792 ();
 FILLCELL_X32 FILLER_290_1824 ();
 FILLCELL_X32 FILLER_290_1856 ();
 FILLCELL_X4 FILLER_290_1888 ();
 FILLCELL_X2 FILLER_290_1892 ();
 FILLCELL_X32 FILLER_290_1895 ();
 FILLCELL_X32 FILLER_290_1927 ();
 FILLCELL_X32 FILLER_290_1959 ();
 FILLCELL_X32 FILLER_290_1991 ();
 FILLCELL_X32 FILLER_290_2023 ();
 FILLCELL_X32 FILLER_290_2055 ();
 FILLCELL_X32 FILLER_290_2087 ();
 FILLCELL_X32 FILLER_290_2119 ();
 FILLCELL_X32 FILLER_290_2151 ();
 FILLCELL_X32 FILLER_290_2183 ();
 FILLCELL_X32 FILLER_290_2215 ();
 FILLCELL_X32 FILLER_290_2247 ();
 FILLCELL_X32 FILLER_290_2279 ();
 FILLCELL_X32 FILLER_290_2311 ();
 FILLCELL_X32 FILLER_290_2343 ();
 FILLCELL_X32 FILLER_290_2375 ();
 FILLCELL_X32 FILLER_290_2407 ();
 FILLCELL_X32 FILLER_290_2439 ();
 FILLCELL_X32 FILLER_290_2471 ();
 FILLCELL_X32 FILLER_290_2503 ();
 FILLCELL_X32 FILLER_290_2535 ();
 FILLCELL_X32 FILLER_290_2567 ();
 FILLCELL_X32 FILLER_290_2599 ();
 FILLCELL_X32 FILLER_290_2631 ();
 FILLCELL_X32 FILLER_290_2663 ();
 FILLCELL_X32 FILLER_290_2695 ();
 FILLCELL_X32 FILLER_290_2727 ();
 FILLCELL_X32 FILLER_290_2759 ();
 FILLCELL_X32 FILLER_290_2791 ();
 FILLCELL_X32 FILLER_290_2823 ();
 FILLCELL_X32 FILLER_290_2855 ();
 FILLCELL_X32 FILLER_290_2887 ();
 FILLCELL_X32 FILLER_290_2919 ();
 FILLCELL_X32 FILLER_290_2951 ();
 FILLCELL_X32 FILLER_290_2983 ();
 FILLCELL_X32 FILLER_290_3015 ();
 FILLCELL_X32 FILLER_290_3047 ();
 FILLCELL_X32 FILLER_290_3079 ();
 FILLCELL_X32 FILLER_290_3111 ();
 FILLCELL_X8 FILLER_290_3143 ();
 FILLCELL_X4 FILLER_290_3151 ();
 FILLCELL_X2 FILLER_290_3155 ();
 FILLCELL_X32 FILLER_290_3158 ();
 FILLCELL_X32 FILLER_290_3190 ();
 FILLCELL_X32 FILLER_290_3222 ();
 FILLCELL_X32 FILLER_290_3254 ();
 FILLCELL_X32 FILLER_290_3286 ();
 FILLCELL_X32 FILLER_290_3318 ();
 FILLCELL_X32 FILLER_290_3350 ();
 FILLCELL_X32 FILLER_290_3382 ();
 FILLCELL_X32 FILLER_290_3414 ();
 FILLCELL_X32 FILLER_290_3446 ();
 FILLCELL_X32 FILLER_290_3478 ();
 FILLCELL_X32 FILLER_290_3510 ();
 FILLCELL_X32 FILLER_290_3542 ();
 FILLCELL_X32 FILLER_290_3574 ();
 FILLCELL_X32 FILLER_290_3606 ();
 FILLCELL_X32 FILLER_290_3638 ();
 FILLCELL_X32 FILLER_290_3670 ();
 FILLCELL_X32 FILLER_290_3702 ();
 FILLCELL_X4 FILLER_290_3734 ();
 FILLCELL_X32 FILLER_291_1 ();
 FILLCELL_X32 FILLER_291_33 ();
 FILLCELL_X32 FILLER_291_65 ();
 FILLCELL_X32 FILLER_291_97 ();
 FILLCELL_X32 FILLER_291_129 ();
 FILLCELL_X32 FILLER_291_161 ();
 FILLCELL_X32 FILLER_291_193 ();
 FILLCELL_X32 FILLER_291_225 ();
 FILLCELL_X32 FILLER_291_257 ();
 FILLCELL_X32 FILLER_291_289 ();
 FILLCELL_X32 FILLER_291_321 ();
 FILLCELL_X32 FILLER_291_353 ();
 FILLCELL_X32 FILLER_291_385 ();
 FILLCELL_X32 FILLER_291_417 ();
 FILLCELL_X32 FILLER_291_449 ();
 FILLCELL_X32 FILLER_291_481 ();
 FILLCELL_X32 FILLER_291_513 ();
 FILLCELL_X32 FILLER_291_545 ();
 FILLCELL_X32 FILLER_291_577 ();
 FILLCELL_X32 FILLER_291_609 ();
 FILLCELL_X32 FILLER_291_641 ();
 FILLCELL_X32 FILLER_291_673 ();
 FILLCELL_X32 FILLER_291_705 ();
 FILLCELL_X32 FILLER_291_737 ();
 FILLCELL_X32 FILLER_291_769 ();
 FILLCELL_X32 FILLER_291_801 ();
 FILLCELL_X32 FILLER_291_833 ();
 FILLCELL_X32 FILLER_291_865 ();
 FILLCELL_X32 FILLER_291_897 ();
 FILLCELL_X32 FILLER_291_929 ();
 FILLCELL_X32 FILLER_291_961 ();
 FILLCELL_X32 FILLER_291_993 ();
 FILLCELL_X32 FILLER_291_1025 ();
 FILLCELL_X32 FILLER_291_1057 ();
 FILLCELL_X32 FILLER_291_1089 ();
 FILLCELL_X32 FILLER_291_1121 ();
 FILLCELL_X32 FILLER_291_1153 ();
 FILLCELL_X32 FILLER_291_1185 ();
 FILLCELL_X32 FILLER_291_1217 ();
 FILLCELL_X8 FILLER_291_1249 ();
 FILLCELL_X4 FILLER_291_1257 ();
 FILLCELL_X2 FILLER_291_1261 ();
 FILLCELL_X32 FILLER_291_1264 ();
 FILLCELL_X32 FILLER_291_1296 ();
 FILLCELL_X32 FILLER_291_1328 ();
 FILLCELL_X32 FILLER_291_1360 ();
 FILLCELL_X32 FILLER_291_1392 ();
 FILLCELL_X32 FILLER_291_1424 ();
 FILLCELL_X32 FILLER_291_1456 ();
 FILLCELL_X32 FILLER_291_1488 ();
 FILLCELL_X32 FILLER_291_1520 ();
 FILLCELL_X32 FILLER_291_1552 ();
 FILLCELL_X16 FILLER_291_1584 ();
 FILLCELL_X8 FILLER_291_1600 ();
 FILLCELL_X1 FILLER_291_1608 ();
 FILLCELL_X8 FILLER_291_1633 ();
 FILLCELL_X32 FILLER_291_1658 ();
 FILLCELL_X32 FILLER_291_1690 ();
 FILLCELL_X32 FILLER_291_1722 ();
 FILLCELL_X32 FILLER_291_1754 ();
 FILLCELL_X32 FILLER_291_1786 ();
 FILLCELL_X32 FILLER_291_1818 ();
 FILLCELL_X32 FILLER_291_1850 ();
 FILLCELL_X32 FILLER_291_1882 ();
 FILLCELL_X32 FILLER_291_1914 ();
 FILLCELL_X32 FILLER_291_1946 ();
 FILLCELL_X32 FILLER_291_1978 ();
 FILLCELL_X32 FILLER_291_2010 ();
 FILLCELL_X32 FILLER_291_2042 ();
 FILLCELL_X32 FILLER_291_2074 ();
 FILLCELL_X32 FILLER_291_2106 ();
 FILLCELL_X32 FILLER_291_2138 ();
 FILLCELL_X32 FILLER_291_2170 ();
 FILLCELL_X32 FILLER_291_2202 ();
 FILLCELL_X32 FILLER_291_2234 ();
 FILLCELL_X32 FILLER_291_2266 ();
 FILLCELL_X32 FILLER_291_2298 ();
 FILLCELL_X32 FILLER_291_2330 ();
 FILLCELL_X32 FILLER_291_2362 ();
 FILLCELL_X32 FILLER_291_2394 ();
 FILLCELL_X32 FILLER_291_2426 ();
 FILLCELL_X32 FILLER_291_2458 ();
 FILLCELL_X32 FILLER_291_2490 ();
 FILLCELL_X4 FILLER_291_2522 ();
 FILLCELL_X32 FILLER_291_2527 ();
 FILLCELL_X32 FILLER_291_2559 ();
 FILLCELL_X32 FILLER_291_2591 ();
 FILLCELL_X32 FILLER_291_2623 ();
 FILLCELL_X32 FILLER_291_2655 ();
 FILLCELL_X32 FILLER_291_2687 ();
 FILLCELL_X32 FILLER_291_2719 ();
 FILLCELL_X32 FILLER_291_2751 ();
 FILLCELL_X32 FILLER_291_2783 ();
 FILLCELL_X32 FILLER_291_2815 ();
 FILLCELL_X32 FILLER_291_2847 ();
 FILLCELL_X32 FILLER_291_2879 ();
 FILLCELL_X32 FILLER_291_2911 ();
 FILLCELL_X32 FILLER_291_2943 ();
 FILLCELL_X32 FILLER_291_2975 ();
 FILLCELL_X32 FILLER_291_3007 ();
 FILLCELL_X32 FILLER_291_3039 ();
 FILLCELL_X32 FILLER_291_3071 ();
 FILLCELL_X32 FILLER_291_3103 ();
 FILLCELL_X32 FILLER_291_3135 ();
 FILLCELL_X32 FILLER_291_3167 ();
 FILLCELL_X32 FILLER_291_3199 ();
 FILLCELL_X32 FILLER_291_3231 ();
 FILLCELL_X32 FILLER_291_3263 ();
 FILLCELL_X32 FILLER_291_3295 ();
 FILLCELL_X32 FILLER_291_3327 ();
 FILLCELL_X32 FILLER_291_3359 ();
 FILLCELL_X32 FILLER_291_3391 ();
 FILLCELL_X32 FILLER_291_3423 ();
 FILLCELL_X32 FILLER_291_3455 ();
 FILLCELL_X32 FILLER_291_3487 ();
 FILLCELL_X32 FILLER_291_3519 ();
 FILLCELL_X32 FILLER_291_3551 ();
 FILLCELL_X32 FILLER_291_3583 ();
 FILLCELL_X32 FILLER_291_3615 ();
 FILLCELL_X32 FILLER_291_3647 ();
 FILLCELL_X32 FILLER_291_3679 ();
 FILLCELL_X16 FILLER_291_3711 ();
 FILLCELL_X8 FILLER_291_3727 ();
 FILLCELL_X2 FILLER_291_3735 ();
 FILLCELL_X1 FILLER_291_3737 ();
 FILLCELL_X32 FILLER_292_1 ();
 FILLCELL_X32 FILLER_292_33 ();
 FILLCELL_X32 FILLER_292_65 ();
 FILLCELL_X32 FILLER_292_97 ();
 FILLCELL_X32 FILLER_292_129 ();
 FILLCELL_X32 FILLER_292_161 ();
 FILLCELL_X32 FILLER_292_193 ();
 FILLCELL_X32 FILLER_292_225 ();
 FILLCELL_X32 FILLER_292_257 ();
 FILLCELL_X32 FILLER_292_289 ();
 FILLCELL_X32 FILLER_292_321 ();
 FILLCELL_X32 FILLER_292_353 ();
 FILLCELL_X32 FILLER_292_385 ();
 FILLCELL_X32 FILLER_292_417 ();
 FILLCELL_X32 FILLER_292_449 ();
 FILLCELL_X32 FILLER_292_481 ();
 FILLCELL_X32 FILLER_292_513 ();
 FILLCELL_X32 FILLER_292_545 ();
 FILLCELL_X32 FILLER_292_577 ();
 FILLCELL_X16 FILLER_292_609 ();
 FILLCELL_X4 FILLER_292_625 ();
 FILLCELL_X2 FILLER_292_629 ();
 FILLCELL_X32 FILLER_292_632 ();
 FILLCELL_X32 FILLER_292_664 ();
 FILLCELL_X32 FILLER_292_696 ();
 FILLCELL_X32 FILLER_292_728 ();
 FILLCELL_X32 FILLER_292_760 ();
 FILLCELL_X32 FILLER_292_792 ();
 FILLCELL_X32 FILLER_292_824 ();
 FILLCELL_X32 FILLER_292_856 ();
 FILLCELL_X32 FILLER_292_888 ();
 FILLCELL_X32 FILLER_292_920 ();
 FILLCELL_X32 FILLER_292_952 ();
 FILLCELL_X32 FILLER_292_984 ();
 FILLCELL_X32 FILLER_292_1016 ();
 FILLCELL_X32 FILLER_292_1048 ();
 FILLCELL_X32 FILLER_292_1080 ();
 FILLCELL_X32 FILLER_292_1112 ();
 FILLCELL_X32 FILLER_292_1144 ();
 FILLCELL_X32 FILLER_292_1176 ();
 FILLCELL_X32 FILLER_292_1208 ();
 FILLCELL_X32 FILLER_292_1240 ();
 FILLCELL_X32 FILLER_292_1272 ();
 FILLCELL_X32 FILLER_292_1304 ();
 FILLCELL_X32 FILLER_292_1336 ();
 FILLCELL_X32 FILLER_292_1368 ();
 FILLCELL_X32 FILLER_292_1400 ();
 FILLCELL_X32 FILLER_292_1432 ();
 FILLCELL_X32 FILLER_292_1464 ();
 FILLCELL_X32 FILLER_292_1496 ();
 FILLCELL_X32 FILLER_292_1528 ();
 FILLCELL_X32 FILLER_292_1560 ();
 FILLCELL_X32 FILLER_292_1592 ();
 FILLCELL_X32 FILLER_292_1624 ();
 FILLCELL_X32 FILLER_292_1656 ();
 FILLCELL_X32 FILLER_292_1688 ();
 FILLCELL_X32 FILLER_292_1720 ();
 FILLCELL_X32 FILLER_292_1752 ();
 FILLCELL_X32 FILLER_292_1784 ();
 FILLCELL_X32 FILLER_292_1816 ();
 FILLCELL_X32 FILLER_292_1848 ();
 FILLCELL_X8 FILLER_292_1880 ();
 FILLCELL_X4 FILLER_292_1888 ();
 FILLCELL_X2 FILLER_292_1892 ();
 FILLCELL_X32 FILLER_292_1895 ();
 FILLCELL_X32 FILLER_292_1927 ();
 FILLCELL_X32 FILLER_292_1959 ();
 FILLCELL_X32 FILLER_292_1991 ();
 FILLCELL_X32 FILLER_292_2023 ();
 FILLCELL_X32 FILLER_292_2055 ();
 FILLCELL_X32 FILLER_292_2087 ();
 FILLCELL_X32 FILLER_292_2119 ();
 FILLCELL_X32 FILLER_292_2151 ();
 FILLCELL_X32 FILLER_292_2183 ();
 FILLCELL_X32 FILLER_292_2215 ();
 FILLCELL_X32 FILLER_292_2247 ();
 FILLCELL_X32 FILLER_292_2279 ();
 FILLCELL_X32 FILLER_292_2311 ();
 FILLCELL_X32 FILLER_292_2343 ();
 FILLCELL_X32 FILLER_292_2375 ();
 FILLCELL_X32 FILLER_292_2407 ();
 FILLCELL_X32 FILLER_292_2439 ();
 FILLCELL_X32 FILLER_292_2471 ();
 FILLCELL_X32 FILLER_292_2503 ();
 FILLCELL_X32 FILLER_292_2535 ();
 FILLCELL_X32 FILLER_292_2567 ();
 FILLCELL_X32 FILLER_292_2599 ();
 FILLCELL_X32 FILLER_292_2631 ();
 FILLCELL_X32 FILLER_292_2663 ();
 FILLCELL_X32 FILLER_292_2695 ();
 FILLCELL_X32 FILLER_292_2727 ();
 FILLCELL_X32 FILLER_292_2759 ();
 FILLCELL_X32 FILLER_292_2791 ();
 FILLCELL_X32 FILLER_292_2823 ();
 FILLCELL_X32 FILLER_292_2855 ();
 FILLCELL_X32 FILLER_292_2887 ();
 FILLCELL_X32 FILLER_292_2919 ();
 FILLCELL_X32 FILLER_292_2951 ();
 FILLCELL_X32 FILLER_292_2983 ();
 FILLCELL_X32 FILLER_292_3015 ();
 FILLCELL_X32 FILLER_292_3047 ();
 FILLCELL_X32 FILLER_292_3079 ();
 FILLCELL_X32 FILLER_292_3111 ();
 FILLCELL_X8 FILLER_292_3143 ();
 FILLCELL_X4 FILLER_292_3151 ();
 FILLCELL_X2 FILLER_292_3155 ();
 FILLCELL_X32 FILLER_292_3158 ();
 FILLCELL_X32 FILLER_292_3190 ();
 FILLCELL_X32 FILLER_292_3222 ();
 FILLCELL_X32 FILLER_292_3254 ();
 FILLCELL_X32 FILLER_292_3286 ();
 FILLCELL_X32 FILLER_292_3318 ();
 FILLCELL_X32 FILLER_292_3350 ();
 FILLCELL_X32 FILLER_292_3382 ();
 FILLCELL_X32 FILLER_292_3414 ();
 FILLCELL_X32 FILLER_292_3446 ();
 FILLCELL_X32 FILLER_292_3478 ();
 FILLCELL_X32 FILLER_292_3510 ();
 FILLCELL_X32 FILLER_292_3542 ();
 FILLCELL_X32 FILLER_292_3574 ();
 FILLCELL_X32 FILLER_292_3606 ();
 FILLCELL_X32 FILLER_292_3638 ();
 FILLCELL_X32 FILLER_292_3670 ();
 FILLCELL_X32 FILLER_292_3702 ();
 FILLCELL_X4 FILLER_292_3734 ();
 FILLCELL_X32 FILLER_293_1 ();
 FILLCELL_X32 FILLER_293_33 ();
 FILLCELL_X32 FILLER_293_65 ();
 FILLCELL_X32 FILLER_293_97 ();
 FILLCELL_X32 FILLER_293_129 ();
 FILLCELL_X32 FILLER_293_161 ();
 FILLCELL_X32 FILLER_293_193 ();
 FILLCELL_X32 FILLER_293_225 ();
 FILLCELL_X32 FILLER_293_257 ();
 FILLCELL_X32 FILLER_293_289 ();
 FILLCELL_X32 FILLER_293_321 ();
 FILLCELL_X32 FILLER_293_353 ();
 FILLCELL_X32 FILLER_293_385 ();
 FILLCELL_X32 FILLER_293_417 ();
 FILLCELL_X32 FILLER_293_449 ();
 FILLCELL_X32 FILLER_293_481 ();
 FILLCELL_X32 FILLER_293_513 ();
 FILLCELL_X32 FILLER_293_545 ();
 FILLCELL_X32 FILLER_293_577 ();
 FILLCELL_X32 FILLER_293_609 ();
 FILLCELL_X32 FILLER_293_641 ();
 FILLCELL_X32 FILLER_293_673 ();
 FILLCELL_X32 FILLER_293_705 ();
 FILLCELL_X32 FILLER_293_737 ();
 FILLCELL_X32 FILLER_293_769 ();
 FILLCELL_X32 FILLER_293_801 ();
 FILLCELL_X32 FILLER_293_833 ();
 FILLCELL_X32 FILLER_293_865 ();
 FILLCELL_X32 FILLER_293_897 ();
 FILLCELL_X32 FILLER_293_929 ();
 FILLCELL_X32 FILLER_293_961 ();
 FILLCELL_X32 FILLER_293_993 ();
 FILLCELL_X32 FILLER_293_1025 ();
 FILLCELL_X32 FILLER_293_1057 ();
 FILLCELL_X32 FILLER_293_1089 ();
 FILLCELL_X32 FILLER_293_1121 ();
 FILLCELL_X32 FILLER_293_1153 ();
 FILLCELL_X32 FILLER_293_1185 ();
 FILLCELL_X32 FILLER_293_1217 ();
 FILLCELL_X8 FILLER_293_1249 ();
 FILLCELL_X4 FILLER_293_1257 ();
 FILLCELL_X2 FILLER_293_1261 ();
 FILLCELL_X32 FILLER_293_1264 ();
 FILLCELL_X32 FILLER_293_1296 ();
 FILLCELL_X32 FILLER_293_1328 ();
 FILLCELL_X32 FILLER_293_1360 ();
 FILLCELL_X32 FILLER_293_1392 ();
 FILLCELL_X32 FILLER_293_1424 ();
 FILLCELL_X32 FILLER_293_1456 ();
 FILLCELL_X32 FILLER_293_1488 ();
 FILLCELL_X32 FILLER_293_1520 ();
 FILLCELL_X32 FILLER_293_1552 ();
 FILLCELL_X32 FILLER_293_1584 ();
 FILLCELL_X32 FILLER_293_1616 ();
 FILLCELL_X8 FILLER_293_1648 ();
 FILLCELL_X4 FILLER_293_1656 ();
 FILLCELL_X2 FILLER_293_1660 ();
 FILLCELL_X16 FILLER_293_1666 ();
 FILLCELL_X8 FILLER_293_1682 ();
 FILLCELL_X2 FILLER_293_1690 ();
 FILLCELL_X32 FILLER_293_1696 ();
 FILLCELL_X32 FILLER_293_1728 ();
 FILLCELL_X32 FILLER_293_1760 ();
 FILLCELL_X32 FILLER_293_1792 ();
 FILLCELL_X32 FILLER_293_1824 ();
 FILLCELL_X32 FILLER_293_1856 ();
 FILLCELL_X32 FILLER_293_1888 ();
 FILLCELL_X32 FILLER_293_1920 ();
 FILLCELL_X32 FILLER_293_1952 ();
 FILLCELL_X32 FILLER_293_1984 ();
 FILLCELL_X32 FILLER_293_2016 ();
 FILLCELL_X32 FILLER_293_2048 ();
 FILLCELL_X32 FILLER_293_2080 ();
 FILLCELL_X32 FILLER_293_2112 ();
 FILLCELL_X32 FILLER_293_2144 ();
 FILLCELL_X32 FILLER_293_2176 ();
 FILLCELL_X32 FILLER_293_2208 ();
 FILLCELL_X32 FILLER_293_2240 ();
 FILLCELL_X32 FILLER_293_2272 ();
 FILLCELL_X32 FILLER_293_2304 ();
 FILLCELL_X32 FILLER_293_2336 ();
 FILLCELL_X32 FILLER_293_2368 ();
 FILLCELL_X32 FILLER_293_2400 ();
 FILLCELL_X32 FILLER_293_2432 ();
 FILLCELL_X32 FILLER_293_2464 ();
 FILLCELL_X16 FILLER_293_2496 ();
 FILLCELL_X8 FILLER_293_2512 ();
 FILLCELL_X4 FILLER_293_2520 ();
 FILLCELL_X2 FILLER_293_2524 ();
 FILLCELL_X32 FILLER_293_2527 ();
 FILLCELL_X32 FILLER_293_2559 ();
 FILLCELL_X32 FILLER_293_2591 ();
 FILLCELL_X32 FILLER_293_2623 ();
 FILLCELL_X32 FILLER_293_2655 ();
 FILLCELL_X32 FILLER_293_2687 ();
 FILLCELL_X32 FILLER_293_2719 ();
 FILLCELL_X32 FILLER_293_2751 ();
 FILLCELL_X32 FILLER_293_2783 ();
 FILLCELL_X32 FILLER_293_2815 ();
 FILLCELL_X32 FILLER_293_2847 ();
 FILLCELL_X32 FILLER_293_2879 ();
 FILLCELL_X32 FILLER_293_2911 ();
 FILLCELL_X32 FILLER_293_2943 ();
 FILLCELL_X32 FILLER_293_2975 ();
 FILLCELL_X32 FILLER_293_3007 ();
 FILLCELL_X32 FILLER_293_3039 ();
 FILLCELL_X32 FILLER_293_3071 ();
 FILLCELL_X32 FILLER_293_3103 ();
 FILLCELL_X32 FILLER_293_3135 ();
 FILLCELL_X32 FILLER_293_3167 ();
 FILLCELL_X32 FILLER_293_3199 ();
 FILLCELL_X32 FILLER_293_3231 ();
 FILLCELL_X32 FILLER_293_3263 ();
 FILLCELL_X32 FILLER_293_3295 ();
 FILLCELL_X32 FILLER_293_3327 ();
 FILLCELL_X32 FILLER_293_3359 ();
 FILLCELL_X32 FILLER_293_3391 ();
 FILLCELL_X32 FILLER_293_3423 ();
 FILLCELL_X32 FILLER_293_3455 ();
 FILLCELL_X32 FILLER_293_3487 ();
 FILLCELL_X32 FILLER_293_3519 ();
 FILLCELL_X32 FILLER_293_3551 ();
 FILLCELL_X32 FILLER_293_3583 ();
 FILLCELL_X32 FILLER_293_3615 ();
 FILLCELL_X32 FILLER_293_3647 ();
 FILLCELL_X32 FILLER_293_3679 ();
 FILLCELL_X16 FILLER_293_3711 ();
 FILLCELL_X8 FILLER_293_3727 ();
 FILLCELL_X2 FILLER_293_3735 ();
 FILLCELL_X1 FILLER_293_3737 ();
 FILLCELL_X32 FILLER_294_1 ();
 FILLCELL_X32 FILLER_294_33 ();
 FILLCELL_X32 FILLER_294_65 ();
 FILLCELL_X32 FILLER_294_97 ();
 FILLCELL_X32 FILLER_294_129 ();
 FILLCELL_X32 FILLER_294_161 ();
 FILLCELL_X32 FILLER_294_193 ();
 FILLCELL_X32 FILLER_294_225 ();
 FILLCELL_X32 FILLER_294_257 ();
 FILLCELL_X32 FILLER_294_289 ();
 FILLCELL_X32 FILLER_294_321 ();
 FILLCELL_X32 FILLER_294_353 ();
 FILLCELL_X32 FILLER_294_385 ();
 FILLCELL_X32 FILLER_294_417 ();
 FILLCELL_X32 FILLER_294_449 ();
 FILLCELL_X32 FILLER_294_481 ();
 FILLCELL_X32 FILLER_294_513 ();
 FILLCELL_X32 FILLER_294_545 ();
 FILLCELL_X32 FILLER_294_577 ();
 FILLCELL_X16 FILLER_294_609 ();
 FILLCELL_X4 FILLER_294_625 ();
 FILLCELL_X2 FILLER_294_629 ();
 FILLCELL_X32 FILLER_294_632 ();
 FILLCELL_X32 FILLER_294_664 ();
 FILLCELL_X32 FILLER_294_696 ();
 FILLCELL_X32 FILLER_294_728 ();
 FILLCELL_X32 FILLER_294_760 ();
 FILLCELL_X32 FILLER_294_792 ();
 FILLCELL_X32 FILLER_294_824 ();
 FILLCELL_X32 FILLER_294_856 ();
 FILLCELL_X32 FILLER_294_888 ();
 FILLCELL_X32 FILLER_294_920 ();
 FILLCELL_X32 FILLER_294_952 ();
 FILLCELL_X32 FILLER_294_984 ();
 FILLCELL_X32 FILLER_294_1016 ();
 FILLCELL_X32 FILLER_294_1048 ();
 FILLCELL_X32 FILLER_294_1080 ();
 FILLCELL_X32 FILLER_294_1112 ();
 FILLCELL_X32 FILLER_294_1144 ();
 FILLCELL_X32 FILLER_294_1176 ();
 FILLCELL_X32 FILLER_294_1208 ();
 FILLCELL_X32 FILLER_294_1240 ();
 FILLCELL_X32 FILLER_294_1272 ();
 FILLCELL_X32 FILLER_294_1304 ();
 FILLCELL_X32 FILLER_294_1336 ();
 FILLCELL_X32 FILLER_294_1368 ();
 FILLCELL_X32 FILLER_294_1400 ();
 FILLCELL_X32 FILLER_294_1432 ();
 FILLCELL_X32 FILLER_294_1464 ();
 FILLCELL_X32 FILLER_294_1496 ();
 FILLCELL_X32 FILLER_294_1528 ();
 FILLCELL_X32 FILLER_294_1560 ();
 FILLCELL_X32 FILLER_294_1592 ();
 FILLCELL_X32 FILLER_294_1624 ();
 FILLCELL_X32 FILLER_294_1656 ();
 FILLCELL_X32 FILLER_294_1688 ();
 FILLCELL_X32 FILLER_294_1720 ();
 FILLCELL_X32 FILLER_294_1752 ();
 FILLCELL_X32 FILLER_294_1784 ();
 FILLCELL_X32 FILLER_294_1816 ();
 FILLCELL_X32 FILLER_294_1848 ();
 FILLCELL_X8 FILLER_294_1880 ();
 FILLCELL_X4 FILLER_294_1888 ();
 FILLCELL_X2 FILLER_294_1892 ();
 FILLCELL_X32 FILLER_294_1895 ();
 FILLCELL_X32 FILLER_294_1927 ();
 FILLCELL_X32 FILLER_294_1959 ();
 FILLCELL_X32 FILLER_294_1991 ();
 FILLCELL_X32 FILLER_294_2023 ();
 FILLCELL_X32 FILLER_294_2055 ();
 FILLCELL_X32 FILLER_294_2087 ();
 FILLCELL_X32 FILLER_294_2119 ();
 FILLCELL_X32 FILLER_294_2151 ();
 FILLCELL_X32 FILLER_294_2183 ();
 FILLCELL_X32 FILLER_294_2215 ();
 FILLCELL_X32 FILLER_294_2247 ();
 FILLCELL_X32 FILLER_294_2279 ();
 FILLCELL_X32 FILLER_294_2311 ();
 FILLCELL_X32 FILLER_294_2343 ();
 FILLCELL_X32 FILLER_294_2375 ();
 FILLCELL_X32 FILLER_294_2407 ();
 FILLCELL_X32 FILLER_294_2439 ();
 FILLCELL_X32 FILLER_294_2471 ();
 FILLCELL_X32 FILLER_294_2503 ();
 FILLCELL_X32 FILLER_294_2535 ();
 FILLCELL_X32 FILLER_294_2567 ();
 FILLCELL_X32 FILLER_294_2599 ();
 FILLCELL_X32 FILLER_294_2631 ();
 FILLCELL_X32 FILLER_294_2663 ();
 FILLCELL_X32 FILLER_294_2695 ();
 FILLCELL_X32 FILLER_294_2727 ();
 FILLCELL_X32 FILLER_294_2759 ();
 FILLCELL_X32 FILLER_294_2791 ();
 FILLCELL_X32 FILLER_294_2823 ();
 FILLCELL_X32 FILLER_294_2855 ();
 FILLCELL_X32 FILLER_294_2887 ();
 FILLCELL_X32 FILLER_294_2919 ();
 FILLCELL_X32 FILLER_294_2951 ();
 FILLCELL_X32 FILLER_294_2983 ();
 FILLCELL_X32 FILLER_294_3015 ();
 FILLCELL_X32 FILLER_294_3047 ();
 FILLCELL_X32 FILLER_294_3079 ();
 FILLCELL_X32 FILLER_294_3111 ();
 FILLCELL_X8 FILLER_294_3143 ();
 FILLCELL_X4 FILLER_294_3151 ();
 FILLCELL_X2 FILLER_294_3155 ();
 FILLCELL_X32 FILLER_294_3158 ();
 FILLCELL_X32 FILLER_294_3190 ();
 FILLCELL_X32 FILLER_294_3222 ();
 FILLCELL_X32 FILLER_294_3254 ();
 FILLCELL_X32 FILLER_294_3286 ();
 FILLCELL_X32 FILLER_294_3318 ();
 FILLCELL_X32 FILLER_294_3350 ();
 FILLCELL_X32 FILLER_294_3382 ();
 FILLCELL_X32 FILLER_294_3414 ();
 FILLCELL_X32 FILLER_294_3446 ();
 FILLCELL_X32 FILLER_294_3478 ();
 FILLCELL_X32 FILLER_294_3510 ();
 FILLCELL_X32 FILLER_294_3542 ();
 FILLCELL_X32 FILLER_294_3574 ();
 FILLCELL_X32 FILLER_294_3606 ();
 FILLCELL_X32 FILLER_294_3638 ();
 FILLCELL_X32 FILLER_294_3670 ();
 FILLCELL_X32 FILLER_294_3702 ();
 FILLCELL_X4 FILLER_294_3734 ();
 FILLCELL_X32 FILLER_295_1 ();
 FILLCELL_X32 FILLER_295_33 ();
 FILLCELL_X32 FILLER_295_65 ();
 FILLCELL_X32 FILLER_295_97 ();
 FILLCELL_X32 FILLER_295_129 ();
 FILLCELL_X32 FILLER_295_161 ();
 FILLCELL_X32 FILLER_295_193 ();
 FILLCELL_X32 FILLER_295_225 ();
 FILLCELL_X32 FILLER_295_257 ();
 FILLCELL_X32 FILLER_295_289 ();
 FILLCELL_X32 FILLER_295_321 ();
 FILLCELL_X32 FILLER_295_353 ();
 FILLCELL_X32 FILLER_295_385 ();
 FILLCELL_X32 FILLER_295_417 ();
 FILLCELL_X32 FILLER_295_449 ();
 FILLCELL_X32 FILLER_295_481 ();
 FILLCELL_X32 FILLER_295_513 ();
 FILLCELL_X32 FILLER_295_545 ();
 FILLCELL_X32 FILLER_295_577 ();
 FILLCELL_X32 FILLER_295_609 ();
 FILLCELL_X32 FILLER_295_641 ();
 FILLCELL_X32 FILLER_295_673 ();
 FILLCELL_X32 FILLER_295_705 ();
 FILLCELL_X32 FILLER_295_737 ();
 FILLCELL_X32 FILLER_295_769 ();
 FILLCELL_X32 FILLER_295_801 ();
 FILLCELL_X32 FILLER_295_833 ();
 FILLCELL_X32 FILLER_295_865 ();
 FILLCELL_X32 FILLER_295_897 ();
 FILLCELL_X32 FILLER_295_929 ();
 FILLCELL_X32 FILLER_295_961 ();
 FILLCELL_X32 FILLER_295_993 ();
 FILLCELL_X32 FILLER_295_1025 ();
 FILLCELL_X32 FILLER_295_1057 ();
 FILLCELL_X32 FILLER_295_1089 ();
 FILLCELL_X32 FILLER_295_1121 ();
 FILLCELL_X32 FILLER_295_1153 ();
 FILLCELL_X32 FILLER_295_1185 ();
 FILLCELL_X32 FILLER_295_1217 ();
 FILLCELL_X8 FILLER_295_1249 ();
 FILLCELL_X4 FILLER_295_1257 ();
 FILLCELL_X2 FILLER_295_1261 ();
 FILLCELL_X32 FILLER_295_1264 ();
 FILLCELL_X32 FILLER_295_1296 ();
 FILLCELL_X32 FILLER_295_1328 ();
 FILLCELL_X32 FILLER_295_1360 ();
 FILLCELL_X32 FILLER_295_1392 ();
 FILLCELL_X32 FILLER_295_1424 ();
 FILLCELL_X32 FILLER_295_1456 ();
 FILLCELL_X32 FILLER_295_1488 ();
 FILLCELL_X32 FILLER_295_1520 ();
 FILLCELL_X32 FILLER_295_1552 ();
 FILLCELL_X32 FILLER_295_1584 ();
 FILLCELL_X32 FILLER_295_1616 ();
 FILLCELL_X32 FILLER_295_1648 ();
 FILLCELL_X32 FILLER_295_1680 ();
 FILLCELL_X32 FILLER_295_1712 ();
 FILLCELL_X32 FILLER_295_1744 ();
 FILLCELL_X32 FILLER_295_1776 ();
 FILLCELL_X32 FILLER_295_1808 ();
 FILLCELL_X32 FILLER_295_1840 ();
 FILLCELL_X32 FILLER_295_1872 ();
 FILLCELL_X32 FILLER_295_1904 ();
 FILLCELL_X32 FILLER_295_1936 ();
 FILLCELL_X32 FILLER_295_1968 ();
 FILLCELL_X32 FILLER_295_2000 ();
 FILLCELL_X32 FILLER_295_2032 ();
 FILLCELL_X32 FILLER_295_2064 ();
 FILLCELL_X32 FILLER_295_2096 ();
 FILLCELL_X32 FILLER_295_2128 ();
 FILLCELL_X32 FILLER_295_2160 ();
 FILLCELL_X32 FILLER_295_2192 ();
 FILLCELL_X32 FILLER_295_2224 ();
 FILLCELL_X32 FILLER_295_2256 ();
 FILLCELL_X32 FILLER_295_2288 ();
 FILLCELL_X32 FILLER_295_2320 ();
 FILLCELL_X32 FILLER_295_2352 ();
 FILLCELL_X32 FILLER_295_2384 ();
 FILLCELL_X32 FILLER_295_2416 ();
 FILLCELL_X32 FILLER_295_2448 ();
 FILLCELL_X32 FILLER_295_2480 ();
 FILLCELL_X8 FILLER_295_2512 ();
 FILLCELL_X4 FILLER_295_2520 ();
 FILLCELL_X2 FILLER_295_2524 ();
 FILLCELL_X32 FILLER_295_2527 ();
 FILLCELL_X32 FILLER_295_2559 ();
 FILLCELL_X32 FILLER_295_2591 ();
 FILLCELL_X32 FILLER_295_2623 ();
 FILLCELL_X32 FILLER_295_2655 ();
 FILLCELL_X32 FILLER_295_2687 ();
 FILLCELL_X32 FILLER_295_2719 ();
 FILLCELL_X32 FILLER_295_2751 ();
 FILLCELL_X32 FILLER_295_2783 ();
 FILLCELL_X32 FILLER_295_2815 ();
 FILLCELL_X32 FILLER_295_2847 ();
 FILLCELL_X32 FILLER_295_2879 ();
 FILLCELL_X32 FILLER_295_2911 ();
 FILLCELL_X32 FILLER_295_2943 ();
 FILLCELL_X32 FILLER_295_2975 ();
 FILLCELL_X32 FILLER_295_3007 ();
 FILLCELL_X32 FILLER_295_3039 ();
 FILLCELL_X32 FILLER_295_3071 ();
 FILLCELL_X32 FILLER_295_3103 ();
 FILLCELL_X32 FILLER_295_3135 ();
 FILLCELL_X32 FILLER_295_3167 ();
 FILLCELL_X32 FILLER_295_3199 ();
 FILLCELL_X32 FILLER_295_3231 ();
 FILLCELL_X32 FILLER_295_3263 ();
 FILLCELL_X32 FILLER_295_3295 ();
 FILLCELL_X32 FILLER_295_3327 ();
 FILLCELL_X32 FILLER_295_3359 ();
 FILLCELL_X32 FILLER_295_3391 ();
 FILLCELL_X32 FILLER_295_3423 ();
 FILLCELL_X32 FILLER_295_3455 ();
 FILLCELL_X32 FILLER_295_3487 ();
 FILLCELL_X32 FILLER_295_3519 ();
 FILLCELL_X32 FILLER_295_3551 ();
 FILLCELL_X32 FILLER_295_3583 ();
 FILLCELL_X32 FILLER_295_3615 ();
 FILLCELL_X32 FILLER_295_3647 ();
 FILLCELL_X32 FILLER_295_3679 ();
 FILLCELL_X16 FILLER_295_3711 ();
 FILLCELL_X8 FILLER_295_3727 ();
 FILLCELL_X2 FILLER_295_3735 ();
 FILLCELL_X1 FILLER_295_3737 ();
 FILLCELL_X32 FILLER_296_1 ();
 FILLCELL_X32 FILLER_296_33 ();
 FILLCELL_X32 FILLER_296_65 ();
 FILLCELL_X32 FILLER_296_97 ();
 FILLCELL_X32 FILLER_296_129 ();
 FILLCELL_X32 FILLER_296_161 ();
 FILLCELL_X32 FILLER_296_193 ();
 FILLCELL_X32 FILLER_296_225 ();
 FILLCELL_X32 FILLER_296_257 ();
 FILLCELL_X32 FILLER_296_289 ();
 FILLCELL_X32 FILLER_296_321 ();
 FILLCELL_X32 FILLER_296_353 ();
 FILLCELL_X32 FILLER_296_385 ();
 FILLCELL_X32 FILLER_296_417 ();
 FILLCELL_X32 FILLER_296_449 ();
 FILLCELL_X32 FILLER_296_481 ();
 FILLCELL_X32 FILLER_296_513 ();
 FILLCELL_X32 FILLER_296_545 ();
 FILLCELL_X32 FILLER_296_577 ();
 FILLCELL_X16 FILLER_296_609 ();
 FILLCELL_X4 FILLER_296_625 ();
 FILLCELL_X2 FILLER_296_629 ();
 FILLCELL_X32 FILLER_296_632 ();
 FILLCELL_X32 FILLER_296_664 ();
 FILLCELL_X32 FILLER_296_696 ();
 FILLCELL_X32 FILLER_296_728 ();
 FILLCELL_X32 FILLER_296_760 ();
 FILLCELL_X32 FILLER_296_792 ();
 FILLCELL_X32 FILLER_296_824 ();
 FILLCELL_X32 FILLER_296_856 ();
 FILLCELL_X32 FILLER_296_888 ();
 FILLCELL_X32 FILLER_296_920 ();
 FILLCELL_X32 FILLER_296_952 ();
 FILLCELL_X32 FILLER_296_984 ();
 FILLCELL_X32 FILLER_296_1016 ();
 FILLCELL_X32 FILLER_296_1048 ();
 FILLCELL_X32 FILLER_296_1080 ();
 FILLCELL_X32 FILLER_296_1112 ();
 FILLCELL_X32 FILLER_296_1144 ();
 FILLCELL_X32 FILLER_296_1176 ();
 FILLCELL_X32 FILLER_296_1208 ();
 FILLCELL_X32 FILLER_296_1240 ();
 FILLCELL_X32 FILLER_296_1272 ();
 FILLCELL_X32 FILLER_296_1304 ();
 FILLCELL_X32 FILLER_296_1336 ();
 FILLCELL_X32 FILLER_296_1368 ();
 FILLCELL_X32 FILLER_296_1400 ();
 FILLCELL_X32 FILLER_296_1432 ();
 FILLCELL_X32 FILLER_296_1464 ();
 FILLCELL_X32 FILLER_296_1496 ();
 FILLCELL_X32 FILLER_296_1528 ();
 FILLCELL_X32 FILLER_296_1560 ();
 FILLCELL_X32 FILLER_296_1592 ();
 FILLCELL_X32 FILLER_296_1624 ();
 FILLCELL_X32 FILLER_296_1656 ();
 FILLCELL_X32 FILLER_296_1688 ();
 FILLCELL_X32 FILLER_296_1720 ();
 FILLCELL_X32 FILLER_296_1752 ();
 FILLCELL_X32 FILLER_296_1784 ();
 FILLCELL_X32 FILLER_296_1816 ();
 FILLCELL_X32 FILLER_296_1848 ();
 FILLCELL_X8 FILLER_296_1880 ();
 FILLCELL_X4 FILLER_296_1888 ();
 FILLCELL_X2 FILLER_296_1892 ();
 FILLCELL_X32 FILLER_296_1895 ();
 FILLCELL_X32 FILLER_296_1927 ();
 FILLCELL_X32 FILLER_296_1959 ();
 FILLCELL_X32 FILLER_296_1991 ();
 FILLCELL_X32 FILLER_296_2023 ();
 FILLCELL_X32 FILLER_296_2055 ();
 FILLCELL_X32 FILLER_296_2087 ();
 FILLCELL_X32 FILLER_296_2119 ();
 FILLCELL_X32 FILLER_296_2151 ();
 FILLCELL_X32 FILLER_296_2183 ();
 FILLCELL_X32 FILLER_296_2215 ();
 FILLCELL_X32 FILLER_296_2247 ();
 FILLCELL_X32 FILLER_296_2279 ();
 FILLCELL_X32 FILLER_296_2311 ();
 FILLCELL_X32 FILLER_296_2343 ();
 FILLCELL_X32 FILLER_296_2375 ();
 FILLCELL_X32 FILLER_296_2407 ();
 FILLCELL_X32 FILLER_296_2439 ();
 FILLCELL_X32 FILLER_296_2471 ();
 FILLCELL_X32 FILLER_296_2503 ();
 FILLCELL_X32 FILLER_296_2535 ();
 FILLCELL_X32 FILLER_296_2567 ();
 FILLCELL_X32 FILLER_296_2599 ();
 FILLCELL_X32 FILLER_296_2631 ();
 FILLCELL_X32 FILLER_296_2663 ();
 FILLCELL_X32 FILLER_296_2695 ();
 FILLCELL_X32 FILLER_296_2727 ();
 FILLCELL_X32 FILLER_296_2759 ();
 FILLCELL_X32 FILLER_296_2791 ();
 FILLCELL_X32 FILLER_296_2823 ();
 FILLCELL_X32 FILLER_296_2855 ();
 FILLCELL_X32 FILLER_296_2887 ();
 FILLCELL_X32 FILLER_296_2919 ();
 FILLCELL_X32 FILLER_296_2951 ();
 FILLCELL_X32 FILLER_296_2983 ();
 FILLCELL_X32 FILLER_296_3015 ();
 FILLCELL_X32 FILLER_296_3047 ();
 FILLCELL_X32 FILLER_296_3079 ();
 FILLCELL_X32 FILLER_296_3111 ();
 FILLCELL_X8 FILLER_296_3143 ();
 FILLCELL_X4 FILLER_296_3151 ();
 FILLCELL_X2 FILLER_296_3155 ();
 FILLCELL_X32 FILLER_296_3158 ();
 FILLCELL_X32 FILLER_296_3190 ();
 FILLCELL_X32 FILLER_296_3222 ();
 FILLCELL_X32 FILLER_296_3254 ();
 FILLCELL_X32 FILLER_296_3286 ();
 FILLCELL_X32 FILLER_296_3318 ();
 FILLCELL_X32 FILLER_296_3350 ();
 FILLCELL_X32 FILLER_296_3382 ();
 FILLCELL_X32 FILLER_296_3414 ();
 FILLCELL_X32 FILLER_296_3446 ();
 FILLCELL_X32 FILLER_296_3478 ();
 FILLCELL_X32 FILLER_296_3510 ();
 FILLCELL_X32 FILLER_296_3542 ();
 FILLCELL_X32 FILLER_296_3574 ();
 FILLCELL_X32 FILLER_296_3606 ();
 FILLCELL_X32 FILLER_296_3638 ();
 FILLCELL_X32 FILLER_296_3670 ();
 FILLCELL_X32 FILLER_296_3702 ();
 FILLCELL_X4 FILLER_296_3734 ();
 FILLCELL_X32 FILLER_297_1 ();
 FILLCELL_X32 FILLER_297_33 ();
 FILLCELL_X32 FILLER_297_65 ();
 FILLCELL_X32 FILLER_297_97 ();
 FILLCELL_X32 FILLER_297_129 ();
 FILLCELL_X32 FILLER_297_161 ();
 FILLCELL_X32 FILLER_297_193 ();
 FILLCELL_X32 FILLER_297_225 ();
 FILLCELL_X32 FILLER_297_257 ();
 FILLCELL_X32 FILLER_297_289 ();
 FILLCELL_X32 FILLER_297_321 ();
 FILLCELL_X32 FILLER_297_353 ();
 FILLCELL_X32 FILLER_297_385 ();
 FILLCELL_X32 FILLER_297_417 ();
 FILLCELL_X32 FILLER_297_449 ();
 FILLCELL_X32 FILLER_297_481 ();
 FILLCELL_X32 FILLER_297_513 ();
 FILLCELL_X32 FILLER_297_545 ();
 FILLCELL_X32 FILLER_297_577 ();
 FILLCELL_X32 FILLER_297_609 ();
 FILLCELL_X32 FILLER_297_641 ();
 FILLCELL_X32 FILLER_297_673 ();
 FILLCELL_X32 FILLER_297_705 ();
 FILLCELL_X32 FILLER_297_737 ();
 FILLCELL_X32 FILLER_297_769 ();
 FILLCELL_X32 FILLER_297_801 ();
 FILLCELL_X32 FILLER_297_833 ();
 FILLCELL_X32 FILLER_297_865 ();
 FILLCELL_X32 FILLER_297_897 ();
 FILLCELL_X32 FILLER_297_929 ();
 FILLCELL_X32 FILLER_297_961 ();
 FILLCELL_X32 FILLER_297_993 ();
 FILLCELL_X32 FILLER_297_1025 ();
 FILLCELL_X32 FILLER_297_1057 ();
 FILLCELL_X32 FILLER_297_1089 ();
 FILLCELL_X32 FILLER_297_1121 ();
 FILLCELL_X32 FILLER_297_1153 ();
 FILLCELL_X32 FILLER_297_1185 ();
 FILLCELL_X32 FILLER_297_1217 ();
 FILLCELL_X8 FILLER_297_1249 ();
 FILLCELL_X4 FILLER_297_1257 ();
 FILLCELL_X2 FILLER_297_1261 ();
 FILLCELL_X32 FILLER_297_1264 ();
 FILLCELL_X32 FILLER_297_1296 ();
 FILLCELL_X32 FILLER_297_1328 ();
 FILLCELL_X32 FILLER_297_1360 ();
 FILLCELL_X32 FILLER_297_1392 ();
 FILLCELL_X32 FILLER_297_1424 ();
 FILLCELL_X32 FILLER_297_1456 ();
 FILLCELL_X32 FILLER_297_1488 ();
 FILLCELL_X32 FILLER_297_1520 ();
 FILLCELL_X32 FILLER_297_1552 ();
 FILLCELL_X32 FILLER_297_1584 ();
 FILLCELL_X32 FILLER_297_1616 ();
 FILLCELL_X32 FILLER_297_1648 ();
 FILLCELL_X32 FILLER_297_1680 ();
 FILLCELL_X32 FILLER_297_1712 ();
 FILLCELL_X32 FILLER_297_1744 ();
 FILLCELL_X32 FILLER_297_1776 ();
 FILLCELL_X32 FILLER_297_1808 ();
 FILLCELL_X32 FILLER_297_1840 ();
 FILLCELL_X32 FILLER_297_1872 ();
 FILLCELL_X32 FILLER_297_1904 ();
 FILLCELL_X32 FILLER_297_1936 ();
 FILLCELL_X32 FILLER_297_1968 ();
 FILLCELL_X32 FILLER_297_2000 ();
 FILLCELL_X32 FILLER_297_2032 ();
 FILLCELL_X32 FILLER_297_2064 ();
 FILLCELL_X32 FILLER_297_2096 ();
 FILLCELL_X32 FILLER_297_2128 ();
 FILLCELL_X32 FILLER_297_2160 ();
 FILLCELL_X32 FILLER_297_2192 ();
 FILLCELL_X32 FILLER_297_2224 ();
 FILLCELL_X32 FILLER_297_2256 ();
 FILLCELL_X32 FILLER_297_2288 ();
 FILLCELL_X32 FILLER_297_2320 ();
 FILLCELL_X32 FILLER_297_2352 ();
 FILLCELL_X32 FILLER_297_2384 ();
 FILLCELL_X32 FILLER_297_2416 ();
 FILLCELL_X32 FILLER_297_2448 ();
 FILLCELL_X32 FILLER_297_2480 ();
 FILLCELL_X8 FILLER_297_2512 ();
 FILLCELL_X4 FILLER_297_2520 ();
 FILLCELL_X2 FILLER_297_2524 ();
 FILLCELL_X32 FILLER_297_2527 ();
 FILLCELL_X32 FILLER_297_2559 ();
 FILLCELL_X32 FILLER_297_2591 ();
 FILLCELL_X32 FILLER_297_2623 ();
 FILLCELL_X32 FILLER_297_2655 ();
 FILLCELL_X32 FILLER_297_2687 ();
 FILLCELL_X32 FILLER_297_2719 ();
 FILLCELL_X32 FILLER_297_2751 ();
 FILLCELL_X32 FILLER_297_2783 ();
 FILLCELL_X32 FILLER_297_2815 ();
 FILLCELL_X32 FILLER_297_2847 ();
 FILLCELL_X32 FILLER_297_2879 ();
 FILLCELL_X32 FILLER_297_2911 ();
 FILLCELL_X32 FILLER_297_2943 ();
 FILLCELL_X32 FILLER_297_2975 ();
 FILLCELL_X32 FILLER_297_3007 ();
 FILLCELL_X32 FILLER_297_3039 ();
 FILLCELL_X32 FILLER_297_3071 ();
 FILLCELL_X32 FILLER_297_3103 ();
 FILLCELL_X32 FILLER_297_3135 ();
 FILLCELL_X32 FILLER_297_3167 ();
 FILLCELL_X32 FILLER_297_3199 ();
 FILLCELL_X32 FILLER_297_3231 ();
 FILLCELL_X32 FILLER_297_3263 ();
 FILLCELL_X32 FILLER_297_3295 ();
 FILLCELL_X32 FILLER_297_3327 ();
 FILLCELL_X32 FILLER_297_3359 ();
 FILLCELL_X32 FILLER_297_3391 ();
 FILLCELL_X32 FILLER_297_3423 ();
 FILLCELL_X32 FILLER_297_3455 ();
 FILLCELL_X32 FILLER_297_3487 ();
 FILLCELL_X32 FILLER_297_3519 ();
 FILLCELL_X32 FILLER_297_3551 ();
 FILLCELL_X32 FILLER_297_3583 ();
 FILLCELL_X32 FILLER_297_3615 ();
 FILLCELL_X32 FILLER_297_3647 ();
 FILLCELL_X32 FILLER_297_3679 ();
 FILLCELL_X16 FILLER_297_3711 ();
 FILLCELL_X8 FILLER_297_3727 ();
 FILLCELL_X2 FILLER_297_3735 ();
 FILLCELL_X1 FILLER_297_3737 ();
 FILLCELL_X32 FILLER_298_1 ();
 FILLCELL_X32 FILLER_298_33 ();
 FILLCELL_X32 FILLER_298_65 ();
 FILLCELL_X32 FILLER_298_97 ();
 FILLCELL_X32 FILLER_298_129 ();
 FILLCELL_X32 FILLER_298_161 ();
 FILLCELL_X32 FILLER_298_193 ();
 FILLCELL_X32 FILLER_298_225 ();
 FILLCELL_X32 FILLER_298_257 ();
 FILLCELL_X32 FILLER_298_289 ();
 FILLCELL_X32 FILLER_298_321 ();
 FILLCELL_X32 FILLER_298_353 ();
 FILLCELL_X32 FILLER_298_385 ();
 FILLCELL_X32 FILLER_298_417 ();
 FILLCELL_X32 FILLER_298_449 ();
 FILLCELL_X32 FILLER_298_481 ();
 FILLCELL_X32 FILLER_298_513 ();
 FILLCELL_X32 FILLER_298_545 ();
 FILLCELL_X32 FILLER_298_577 ();
 FILLCELL_X16 FILLER_298_609 ();
 FILLCELL_X4 FILLER_298_625 ();
 FILLCELL_X2 FILLER_298_629 ();
 FILLCELL_X32 FILLER_298_632 ();
 FILLCELL_X32 FILLER_298_664 ();
 FILLCELL_X32 FILLER_298_696 ();
 FILLCELL_X32 FILLER_298_728 ();
 FILLCELL_X32 FILLER_298_760 ();
 FILLCELL_X32 FILLER_298_792 ();
 FILLCELL_X32 FILLER_298_824 ();
 FILLCELL_X32 FILLER_298_856 ();
 FILLCELL_X32 FILLER_298_888 ();
 FILLCELL_X32 FILLER_298_920 ();
 FILLCELL_X32 FILLER_298_952 ();
 FILLCELL_X32 FILLER_298_984 ();
 FILLCELL_X32 FILLER_298_1016 ();
 FILLCELL_X32 FILLER_298_1048 ();
 FILLCELL_X32 FILLER_298_1080 ();
 FILLCELL_X32 FILLER_298_1112 ();
 FILLCELL_X32 FILLER_298_1144 ();
 FILLCELL_X32 FILLER_298_1176 ();
 FILLCELL_X32 FILLER_298_1208 ();
 FILLCELL_X32 FILLER_298_1240 ();
 FILLCELL_X32 FILLER_298_1272 ();
 FILLCELL_X32 FILLER_298_1304 ();
 FILLCELL_X32 FILLER_298_1336 ();
 FILLCELL_X32 FILLER_298_1368 ();
 FILLCELL_X32 FILLER_298_1400 ();
 FILLCELL_X32 FILLER_298_1432 ();
 FILLCELL_X32 FILLER_298_1464 ();
 FILLCELL_X32 FILLER_298_1496 ();
 FILLCELL_X32 FILLER_298_1528 ();
 FILLCELL_X32 FILLER_298_1560 ();
 FILLCELL_X32 FILLER_298_1592 ();
 FILLCELL_X32 FILLER_298_1624 ();
 FILLCELL_X32 FILLER_298_1656 ();
 FILLCELL_X32 FILLER_298_1688 ();
 FILLCELL_X32 FILLER_298_1720 ();
 FILLCELL_X32 FILLER_298_1752 ();
 FILLCELL_X32 FILLER_298_1784 ();
 FILLCELL_X32 FILLER_298_1816 ();
 FILLCELL_X32 FILLER_298_1848 ();
 FILLCELL_X8 FILLER_298_1880 ();
 FILLCELL_X4 FILLER_298_1888 ();
 FILLCELL_X2 FILLER_298_1892 ();
 FILLCELL_X32 FILLER_298_1895 ();
 FILLCELL_X32 FILLER_298_1927 ();
 FILLCELL_X32 FILLER_298_1959 ();
 FILLCELL_X32 FILLER_298_1991 ();
 FILLCELL_X32 FILLER_298_2023 ();
 FILLCELL_X32 FILLER_298_2055 ();
 FILLCELL_X32 FILLER_298_2087 ();
 FILLCELL_X32 FILLER_298_2119 ();
 FILLCELL_X32 FILLER_298_2151 ();
 FILLCELL_X32 FILLER_298_2183 ();
 FILLCELL_X32 FILLER_298_2215 ();
 FILLCELL_X32 FILLER_298_2247 ();
 FILLCELL_X32 FILLER_298_2279 ();
 FILLCELL_X32 FILLER_298_2311 ();
 FILLCELL_X32 FILLER_298_2343 ();
 FILLCELL_X32 FILLER_298_2375 ();
 FILLCELL_X32 FILLER_298_2407 ();
 FILLCELL_X32 FILLER_298_2439 ();
 FILLCELL_X32 FILLER_298_2471 ();
 FILLCELL_X32 FILLER_298_2503 ();
 FILLCELL_X32 FILLER_298_2535 ();
 FILLCELL_X32 FILLER_298_2567 ();
 FILLCELL_X32 FILLER_298_2599 ();
 FILLCELL_X32 FILLER_298_2631 ();
 FILLCELL_X32 FILLER_298_2663 ();
 FILLCELL_X32 FILLER_298_2695 ();
 FILLCELL_X32 FILLER_298_2727 ();
 FILLCELL_X32 FILLER_298_2759 ();
 FILLCELL_X32 FILLER_298_2791 ();
 FILLCELL_X32 FILLER_298_2823 ();
 FILLCELL_X32 FILLER_298_2855 ();
 FILLCELL_X32 FILLER_298_2887 ();
 FILLCELL_X32 FILLER_298_2919 ();
 FILLCELL_X32 FILLER_298_2951 ();
 FILLCELL_X32 FILLER_298_2983 ();
 FILLCELL_X32 FILLER_298_3015 ();
 FILLCELL_X32 FILLER_298_3047 ();
 FILLCELL_X32 FILLER_298_3079 ();
 FILLCELL_X32 FILLER_298_3111 ();
 FILLCELL_X8 FILLER_298_3143 ();
 FILLCELL_X4 FILLER_298_3151 ();
 FILLCELL_X2 FILLER_298_3155 ();
 FILLCELL_X32 FILLER_298_3158 ();
 FILLCELL_X32 FILLER_298_3190 ();
 FILLCELL_X32 FILLER_298_3222 ();
 FILLCELL_X32 FILLER_298_3254 ();
 FILLCELL_X32 FILLER_298_3286 ();
 FILLCELL_X32 FILLER_298_3318 ();
 FILLCELL_X32 FILLER_298_3350 ();
 FILLCELL_X32 FILLER_298_3382 ();
 FILLCELL_X32 FILLER_298_3414 ();
 FILLCELL_X32 FILLER_298_3446 ();
 FILLCELL_X32 FILLER_298_3478 ();
 FILLCELL_X32 FILLER_298_3510 ();
 FILLCELL_X32 FILLER_298_3542 ();
 FILLCELL_X32 FILLER_298_3574 ();
 FILLCELL_X32 FILLER_298_3606 ();
 FILLCELL_X32 FILLER_298_3638 ();
 FILLCELL_X32 FILLER_298_3670 ();
 FILLCELL_X32 FILLER_298_3702 ();
 FILLCELL_X4 FILLER_298_3734 ();
 FILLCELL_X32 FILLER_299_1 ();
 FILLCELL_X32 FILLER_299_33 ();
 FILLCELL_X32 FILLER_299_65 ();
 FILLCELL_X32 FILLER_299_97 ();
 FILLCELL_X32 FILLER_299_129 ();
 FILLCELL_X32 FILLER_299_161 ();
 FILLCELL_X32 FILLER_299_193 ();
 FILLCELL_X32 FILLER_299_225 ();
 FILLCELL_X32 FILLER_299_257 ();
 FILLCELL_X32 FILLER_299_289 ();
 FILLCELL_X32 FILLER_299_321 ();
 FILLCELL_X32 FILLER_299_353 ();
 FILLCELL_X32 FILLER_299_385 ();
 FILLCELL_X32 FILLER_299_417 ();
 FILLCELL_X32 FILLER_299_449 ();
 FILLCELL_X32 FILLER_299_481 ();
 FILLCELL_X32 FILLER_299_513 ();
 FILLCELL_X32 FILLER_299_545 ();
 FILLCELL_X32 FILLER_299_577 ();
 FILLCELL_X32 FILLER_299_609 ();
 FILLCELL_X32 FILLER_299_641 ();
 FILLCELL_X32 FILLER_299_673 ();
 FILLCELL_X32 FILLER_299_705 ();
 FILLCELL_X32 FILLER_299_737 ();
 FILLCELL_X32 FILLER_299_769 ();
 FILLCELL_X32 FILLER_299_801 ();
 FILLCELL_X32 FILLER_299_833 ();
 FILLCELL_X32 FILLER_299_865 ();
 FILLCELL_X32 FILLER_299_897 ();
 FILLCELL_X32 FILLER_299_929 ();
 FILLCELL_X32 FILLER_299_961 ();
 FILLCELL_X32 FILLER_299_993 ();
 FILLCELL_X32 FILLER_299_1025 ();
 FILLCELL_X32 FILLER_299_1057 ();
 FILLCELL_X32 FILLER_299_1089 ();
 FILLCELL_X32 FILLER_299_1121 ();
 FILLCELL_X32 FILLER_299_1153 ();
 FILLCELL_X32 FILLER_299_1185 ();
 FILLCELL_X32 FILLER_299_1217 ();
 FILLCELL_X8 FILLER_299_1249 ();
 FILLCELL_X4 FILLER_299_1257 ();
 FILLCELL_X2 FILLER_299_1261 ();
 FILLCELL_X32 FILLER_299_1264 ();
 FILLCELL_X32 FILLER_299_1296 ();
 FILLCELL_X32 FILLER_299_1328 ();
 FILLCELL_X32 FILLER_299_1360 ();
 FILLCELL_X32 FILLER_299_1392 ();
 FILLCELL_X32 FILLER_299_1424 ();
 FILLCELL_X32 FILLER_299_1456 ();
 FILLCELL_X32 FILLER_299_1488 ();
 FILLCELL_X32 FILLER_299_1520 ();
 FILLCELL_X32 FILLER_299_1552 ();
 FILLCELL_X32 FILLER_299_1584 ();
 FILLCELL_X32 FILLER_299_1616 ();
 FILLCELL_X32 FILLER_299_1648 ();
 FILLCELL_X32 FILLER_299_1680 ();
 FILLCELL_X32 FILLER_299_1712 ();
 FILLCELL_X32 FILLER_299_1744 ();
 FILLCELL_X32 FILLER_299_1776 ();
 FILLCELL_X32 FILLER_299_1808 ();
 FILLCELL_X32 FILLER_299_1840 ();
 FILLCELL_X32 FILLER_299_1872 ();
 FILLCELL_X32 FILLER_299_1904 ();
 FILLCELL_X32 FILLER_299_1936 ();
 FILLCELL_X32 FILLER_299_1968 ();
 FILLCELL_X32 FILLER_299_2000 ();
 FILLCELL_X32 FILLER_299_2032 ();
 FILLCELL_X32 FILLER_299_2064 ();
 FILLCELL_X32 FILLER_299_2096 ();
 FILLCELL_X32 FILLER_299_2128 ();
 FILLCELL_X32 FILLER_299_2160 ();
 FILLCELL_X32 FILLER_299_2192 ();
 FILLCELL_X32 FILLER_299_2224 ();
 FILLCELL_X32 FILLER_299_2256 ();
 FILLCELL_X32 FILLER_299_2288 ();
 FILLCELL_X32 FILLER_299_2320 ();
 FILLCELL_X32 FILLER_299_2352 ();
 FILLCELL_X32 FILLER_299_2384 ();
 FILLCELL_X32 FILLER_299_2416 ();
 FILLCELL_X32 FILLER_299_2448 ();
 FILLCELL_X32 FILLER_299_2480 ();
 FILLCELL_X8 FILLER_299_2512 ();
 FILLCELL_X4 FILLER_299_2520 ();
 FILLCELL_X2 FILLER_299_2524 ();
 FILLCELL_X32 FILLER_299_2527 ();
 FILLCELL_X32 FILLER_299_2559 ();
 FILLCELL_X32 FILLER_299_2591 ();
 FILLCELL_X32 FILLER_299_2623 ();
 FILLCELL_X32 FILLER_299_2655 ();
 FILLCELL_X32 FILLER_299_2687 ();
 FILLCELL_X32 FILLER_299_2719 ();
 FILLCELL_X32 FILLER_299_2751 ();
 FILLCELL_X32 FILLER_299_2783 ();
 FILLCELL_X32 FILLER_299_2815 ();
 FILLCELL_X32 FILLER_299_2847 ();
 FILLCELL_X32 FILLER_299_2879 ();
 FILLCELL_X32 FILLER_299_2911 ();
 FILLCELL_X32 FILLER_299_2943 ();
 FILLCELL_X32 FILLER_299_2975 ();
 FILLCELL_X32 FILLER_299_3007 ();
 FILLCELL_X32 FILLER_299_3039 ();
 FILLCELL_X32 FILLER_299_3071 ();
 FILLCELL_X32 FILLER_299_3103 ();
 FILLCELL_X32 FILLER_299_3135 ();
 FILLCELL_X32 FILLER_299_3167 ();
 FILLCELL_X32 FILLER_299_3199 ();
 FILLCELL_X32 FILLER_299_3231 ();
 FILLCELL_X32 FILLER_299_3263 ();
 FILLCELL_X32 FILLER_299_3295 ();
 FILLCELL_X32 FILLER_299_3327 ();
 FILLCELL_X32 FILLER_299_3359 ();
 FILLCELL_X32 FILLER_299_3391 ();
 FILLCELL_X32 FILLER_299_3423 ();
 FILLCELL_X32 FILLER_299_3455 ();
 FILLCELL_X32 FILLER_299_3487 ();
 FILLCELL_X32 FILLER_299_3519 ();
 FILLCELL_X32 FILLER_299_3551 ();
 FILLCELL_X32 FILLER_299_3583 ();
 FILLCELL_X32 FILLER_299_3615 ();
 FILLCELL_X32 FILLER_299_3647 ();
 FILLCELL_X32 FILLER_299_3679 ();
 FILLCELL_X16 FILLER_299_3711 ();
 FILLCELL_X8 FILLER_299_3727 ();
 FILLCELL_X2 FILLER_299_3735 ();
 FILLCELL_X1 FILLER_299_3737 ();
 FILLCELL_X32 FILLER_300_1 ();
 FILLCELL_X32 FILLER_300_33 ();
 FILLCELL_X32 FILLER_300_65 ();
 FILLCELL_X32 FILLER_300_97 ();
 FILLCELL_X32 FILLER_300_129 ();
 FILLCELL_X32 FILLER_300_161 ();
 FILLCELL_X32 FILLER_300_193 ();
 FILLCELL_X32 FILLER_300_225 ();
 FILLCELL_X32 FILLER_300_257 ();
 FILLCELL_X32 FILLER_300_289 ();
 FILLCELL_X32 FILLER_300_321 ();
 FILLCELL_X32 FILLER_300_353 ();
 FILLCELL_X32 FILLER_300_385 ();
 FILLCELL_X32 FILLER_300_417 ();
 FILLCELL_X32 FILLER_300_449 ();
 FILLCELL_X32 FILLER_300_481 ();
 FILLCELL_X32 FILLER_300_513 ();
 FILLCELL_X32 FILLER_300_545 ();
 FILLCELL_X32 FILLER_300_577 ();
 FILLCELL_X16 FILLER_300_609 ();
 FILLCELL_X4 FILLER_300_625 ();
 FILLCELL_X2 FILLER_300_629 ();
 FILLCELL_X32 FILLER_300_632 ();
 FILLCELL_X32 FILLER_300_664 ();
 FILLCELL_X32 FILLER_300_696 ();
 FILLCELL_X32 FILLER_300_728 ();
 FILLCELL_X32 FILLER_300_760 ();
 FILLCELL_X32 FILLER_300_792 ();
 FILLCELL_X32 FILLER_300_824 ();
 FILLCELL_X32 FILLER_300_856 ();
 FILLCELL_X32 FILLER_300_888 ();
 FILLCELL_X32 FILLER_300_920 ();
 FILLCELL_X32 FILLER_300_952 ();
 FILLCELL_X32 FILLER_300_984 ();
 FILLCELL_X32 FILLER_300_1016 ();
 FILLCELL_X32 FILLER_300_1048 ();
 FILLCELL_X32 FILLER_300_1080 ();
 FILLCELL_X32 FILLER_300_1112 ();
 FILLCELL_X32 FILLER_300_1144 ();
 FILLCELL_X32 FILLER_300_1176 ();
 FILLCELL_X32 FILLER_300_1208 ();
 FILLCELL_X32 FILLER_300_1240 ();
 FILLCELL_X32 FILLER_300_1272 ();
 FILLCELL_X32 FILLER_300_1304 ();
 FILLCELL_X32 FILLER_300_1336 ();
 FILLCELL_X32 FILLER_300_1368 ();
 FILLCELL_X32 FILLER_300_1400 ();
 FILLCELL_X32 FILLER_300_1432 ();
 FILLCELL_X32 FILLER_300_1464 ();
 FILLCELL_X32 FILLER_300_1496 ();
 FILLCELL_X32 FILLER_300_1528 ();
 FILLCELL_X32 FILLER_300_1560 ();
 FILLCELL_X32 FILLER_300_1592 ();
 FILLCELL_X32 FILLER_300_1624 ();
 FILLCELL_X32 FILLER_300_1656 ();
 FILLCELL_X32 FILLER_300_1688 ();
 FILLCELL_X32 FILLER_300_1720 ();
 FILLCELL_X32 FILLER_300_1752 ();
 FILLCELL_X32 FILLER_300_1784 ();
 FILLCELL_X32 FILLER_300_1816 ();
 FILLCELL_X32 FILLER_300_1848 ();
 FILLCELL_X8 FILLER_300_1880 ();
 FILLCELL_X4 FILLER_300_1888 ();
 FILLCELL_X2 FILLER_300_1892 ();
 FILLCELL_X32 FILLER_300_1895 ();
 FILLCELL_X32 FILLER_300_1927 ();
 FILLCELL_X32 FILLER_300_1959 ();
 FILLCELL_X32 FILLER_300_1991 ();
 FILLCELL_X32 FILLER_300_2023 ();
 FILLCELL_X32 FILLER_300_2055 ();
 FILLCELL_X32 FILLER_300_2087 ();
 FILLCELL_X32 FILLER_300_2119 ();
 FILLCELL_X32 FILLER_300_2151 ();
 FILLCELL_X32 FILLER_300_2183 ();
 FILLCELL_X32 FILLER_300_2215 ();
 FILLCELL_X32 FILLER_300_2247 ();
 FILLCELL_X32 FILLER_300_2279 ();
 FILLCELL_X32 FILLER_300_2311 ();
 FILLCELL_X32 FILLER_300_2343 ();
 FILLCELL_X32 FILLER_300_2375 ();
 FILLCELL_X32 FILLER_300_2407 ();
 FILLCELL_X32 FILLER_300_2439 ();
 FILLCELL_X32 FILLER_300_2471 ();
 FILLCELL_X32 FILLER_300_2503 ();
 FILLCELL_X32 FILLER_300_2535 ();
 FILLCELL_X32 FILLER_300_2567 ();
 FILLCELL_X32 FILLER_300_2599 ();
 FILLCELL_X32 FILLER_300_2631 ();
 FILLCELL_X32 FILLER_300_2663 ();
 FILLCELL_X32 FILLER_300_2695 ();
 FILLCELL_X32 FILLER_300_2727 ();
 FILLCELL_X32 FILLER_300_2759 ();
 FILLCELL_X32 FILLER_300_2791 ();
 FILLCELL_X32 FILLER_300_2823 ();
 FILLCELL_X32 FILLER_300_2855 ();
 FILLCELL_X32 FILLER_300_2887 ();
 FILLCELL_X32 FILLER_300_2919 ();
 FILLCELL_X32 FILLER_300_2951 ();
 FILLCELL_X32 FILLER_300_2983 ();
 FILLCELL_X32 FILLER_300_3015 ();
 FILLCELL_X32 FILLER_300_3047 ();
 FILLCELL_X32 FILLER_300_3079 ();
 FILLCELL_X32 FILLER_300_3111 ();
 FILLCELL_X8 FILLER_300_3143 ();
 FILLCELL_X4 FILLER_300_3151 ();
 FILLCELL_X2 FILLER_300_3155 ();
 FILLCELL_X32 FILLER_300_3158 ();
 FILLCELL_X32 FILLER_300_3190 ();
 FILLCELL_X32 FILLER_300_3222 ();
 FILLCELL_X32 FILLER_300_3254 ();
 FILLCELL_X32 FILLER_300_3286 ();
 FILLCELL_X32 FILLER_300_3318 ();
 FILLCELL_X32 FILLER_300_3350 ();
 FILLCELL_X32 FILLER_300_3382 ();
 FILLCELL_X32 FILLER_300_3414 ();
 FILLCELL_X32 FILLER_300_3446 ();
 FILLCELL_X32 FILLER_300_3478 ();
 FILLCELL_X32 FILLER_300_3510 ();
 FILLCELL_X32 FILLER_300_3542 ();
 FILLCELL_X32 FILLER_300_3574 ();
 FILLCELL_X32 FILLER_300_3606 ();
 FILLCELL_X32 FILLER_300_3638 ();
 FILLCELL_X32 FILLER_300_3670 ();
 FILLCELL_X32 FILLER_300_3702 ();
 FILLCELL_X4 FILLER_300_3734 ();
 FILLCELL_X32 FILLER_301_1 ();
 FILLCELL_X32 FILLER_301_33 ();
 FILLCELL_X32 FILLER_301_65 ();
 FILLCELL_X32 FILLER_301_97 ();
 FILLCELL_X32 FILLER_301_129 ();
 FILLCELL_X32 FILLER_301_161 ();
 FILLCELL_X32 FILLER_301_193 ();
 FILLCELL_X32 FILLER_301_225 ();
 FILLCELL_X32 FILLER_301_257 ();
 FILLCELL_X32 FILLER_301_289 ();
 FILLCELL_X32 FILLER_301_321 ();
 FILLCELL_X32 FILLER_301_353 ();
 FILLCELL_X32 FILLER_301_385 ();
 FILLCELL_X32 FILLER_301_417 ();
 FILLCELL_X32 FILLER_301_449 ();
 FILLCELL_X32 FILLER_301_481 ();
 FILLCELL_X32 FILLER_301_513 ();
 FILLCELL_X32 FILLER_301_545 ();
 FILLCELL_X32 FILLER_301_577 ();
 FILLCELL_X32 FILLER_301_609 ();
 FILLCELL_X32 FILLER_301_641 ();
 FILLCELL_X32 FILLER_301_673 ();
 FILLCELL_X32 FILLER_301_705 ();
 FILLCELL_X32 FILLER_301_737 ();
 FILLCELL_X32 FILLER_301_769 ();
 FILLCELL_X32 FILLER_301_801 ();
 FILLCELL_X32 FILLER_301_833 ();
 FILLCELL_X32 FILLER_301_865 ();
 FILLCELL_X32 FILLER_301_897 ();
 FILLCELL_X32 FILLER_301_929 ();
 FILLCELL_X32 FILLER_301_961 ();
 FILLCELL_X32 FILLER_301_993 ();
 FILLCELL_X32 FILLER_301_1025 ();
 FILLCELL_X32 FILLER_301_1057 ();
 FILLCELL_X32 FILLER_301_1089 ();
 FILLCELL_X32 FILLER_301_1121 ();
 FILLCELL_X32 FILLER_301_1153 ();
 FILLCELL_X32 FILLER_301_1185 ();
 FILLCELL_X32 FILLER_301_1217 ();
 FILLCELL_X8 FILLER_301_1249 ();
 FILLCELL_X4 FILLER_301_1257 ();
 FILLCELL_X2 FILLER_301_1261 ();
 FILLCELL_X32 FILLER_301_1264 ();
 FILLCELL_X32 FILLER_301_1296 ();
 FILLCELL_X32 FILLER_301_1328 ();
 FILLCELL_X32 FILLER_301_1360 ();
 FILLCELL_X32 FILLER_301_1392 ();
 FILLCELL_X32 FILLER_301_1424 ();
 FILLCELL_X32 FILLER_301_1456 ();
 FILLCELL_X32 FILLER_301_1488 ();
 FILLCELL_X32 FILLER_301_1520 ();
 FILLCELL_X32 FILLER_301_1552 ();
 FILLCELL_X32 FILLER_301_1584 ();
 FILLCELL_X32 FILLER_301_1616 ();
 FILLCELL_X32 FILLER_301_1648 ();
 FILLCELL_X32 FILLER_301_1680 ();
 FILLCELL_X32 FILLER_301_1712 ();
 FILLCELL_X32 FILLER_301_1744 ();
 FILLCELL_X32 FILLER_301_1776 ();
 FILLCELL_X32 FILLER_301_1808 ();
 FILLCELL_X32 FILLER_301_1840 ();
 FILLCELL_X32 FILLER_301_1872 ();
 FILLCELL_X32 FILLER_301_1904 ();
 FILLCELL_X32 FILLER_301_1936 ();
 FILLCELL_X32 FILLER_301_1968 ();
 FILLCELL_X32 FILLER_301_2000 ();
 FILLCELL_X32 FILLER_301_2032 ();
 FILLCELL_X32 FILLER_301_2064 ();
 FILLCELL_X32 FILLER_301_2096 ();
 FILLCELL_X32 FILLER_301_2128 ();
 FILLCELL_X32 FILLER_301_2160 ();
 FILLCELL_X32 FILLER_301_2192 ();
 FILLCELL_X32 FILLER_301_2224 ();
 FILLCELL_X32 FILLER_301_2256 ();
 FILLCELL_X32 FILLER_301_2288 ();
 FILLCELL_X32 FILLER_301_2320 ();
 FILLCELL_X32 FILLER_301_2352 ();
 FILLCELL_X32 FILLER_301_2384 ();
 FILLCELL_X32 FILLER_301_2416 ();
 FILLCELL_X32 FILLER_301_2448 ();
 FILLCELL_X32 FILLER_301_2480 ();
 FILLCELL_X8 FILLER_301_2512 ();
 FILLCELL_X4 FILLER_301_2520 ();
 FILLCELL_X2 FILLER_301_2524 ();
 FILLCELL_X32 FILLER_301_2527 ();
 FILLCELL_X32 FILLER_301_2559 ();
 FILLCELL_X32 FILLER_301_2591 ();
 FILLCELL_X32 FILLER_301_2623 ();
 FILLCELL_X32 FILLER_301_2655 ();
 FILLCELL_X32 FILLER_301_2687 ();
 FILLCELL_X32 FILLER_301_2719 ();
 FILLCELL_X32 FILLER_301_2751 ();
 FILLCELL_X32 FILLER_301_2783 ();
 FILLCELL_X32 FILLER_301_2815 ();
 FILLCELL_X32 FILLER_301_2847 ();
 FILLCELL_X32 FILLER_301_2879 ();
 FILLCELL_X32 FILLER_301_2911 ();
 FILLCELL_X32 FILLER_301_2943 ();
 FILLCELL_X32 FILLER_301_2975 ();
 FILLCELL_X32 FILLER_301_3007 ();
 FILLCELL_X32 FILLER_301_3039 ();
 FILLCELL_X32 FILLER_301_3071 ();
 FILLCELL_X32 FILLER_301_3103 ();
 FILLCELL_X32 FILLER_301_3135 ();
 FILLCELL_X32 FILLER_301_3167 ();
 FILLCELL_X32 FILLER_301_3199 ();
 FILLCELL_X32 FILLER_301_3231 ();
 FILLCELL_X32 FILLER_301_3263 ();
 FILLCELL_X32 FILLER_301_3295 ();
 FILLCELL_X32 FILLER_301_3327 ();
 FILLCELL_X32 FILLER_301_3359 ();
 FILLCELL_X32 FILLER_301_3391 ();
 FILLCELL_X32 FILLER_301_3423 ();
 FILLCELL_X32 FILLER_301_3455 ();
 FILLCELL_X32 FILLER_301_3487 ();
 FILLCELL_X32 FILLER_301_3519 ();
 FILLCELL_X32 FILLER_301_3551 ();
 FILLCELL_X32 FILLER_301_3583 ();
 FILLCELL_X32 FILLER_301_3615 ();
 FILLCELL_X32 FILLER_301_3647 ();
 FILLCELL_X32 FILLER_301_3679 ();
 FILLCELL_X16 FILLER_301_3711 ();
 FILLCELL_X8 FILLER_301_3727 ();
 FILLCELL_X2 FILLER_301_3735 ();
 FILLCELL_X1 FILLER_301_3737 ();
 FILLCELL_X32 FILLER_302_1 ();
 FILLCELL_X32 FILLER_302_33 ();
 FILLCELL_X32 FILLER_302_65 ();
 FILLCELL_X32 FILLER_302_97 ();
 FILLCELL_X32 FILLER_302_129 ();
 FILLCELL_X32 FILLER_302_161 ();
 FILLCELL_X32 FILLER_302_193 ();
 FILLCELL_X32 FILLER_302_225 ();
 FILLCELL_X32 FILLER_302_257 ();
 FILLCELL_X32 FILLER_302_289 ();
 FILLCELL_X32 FILLER_302_321 ();
 FILLCELL_X32 FILLER_302_353 ();
 FILLCELL_X32 FILLER_302_385 ();
 FILLCELL_X32 FILLER_302_417 ();
 FILLCELL_X32 FILLER_302_449 ();
 FILLCELL_X32 FILLER_302_481 ();
 FILLCELL_X32 FILLER_302_513 ();
 FILLCELL_X32 FILLER_302_545 ();
 FILLCELL_X32 FILLER_302_577 ();
 FILLCELL_X16 FILLER_302_609 ();
 FILLCELL_X4 FILLER_302_625 ();
 FILLCELL_X2 FILLER_302_629 ();
 FILLCELL_X32 FILLER_302_632 ();
 FILLCELL_X32 FILLER_302_664 ();
 FILLCELL_X32 FILLER_302_696 ();
 FILLCELL_X32 FILLER_302_728 ();
 FILLCELL_X32 FILLER_302_760 ();
 FILLCELL_X32 FILLER_302_792 ();
 FILLCELL_X32 FILLER_302_824 ();
 FILLCELL_X32 FILLER_302_856 ();
 FILLCELL_X32 FILLER_302_888 ();
 FILLCELL_X32 FILLER_302_920 ();
 FILLCELL_X32 FILLER_302_952 ();
 FILLCELL_X32 FILLER_302_984 ();
 FILLCELL_X32 FILLER_302_1016 ();
 FILLCELL_X32 FILLER_302_1048 ();
 FILLCELL_X32 FILLER_302_1080 ();
 FILLCELL_X32 FILLER_302_1112 ();
 FILLCELL_X32 FILLER_302_1144 ();
 FILLCELL_X32 FILLER_302_1176 ();
 FILLCELL_X32 FILLER_302_1208 ();
 FILLCELL_X32 FILLER_302_1240 ();
 FILLCELL_X32 FILLER_302_1272 ();
 FILLCELL_X32 FILLER_302_1304 ();
 FILLCELL_X32 FILLER_302_1336 ();
 FILLCELL_X32 FILLER_302_1368 ();
 FILLCELL_X32 FILLER_302_1400 ();
 FILLCELL_X32 FILLER_302_1432 ();
 FILLCELL_X32 FILLER_302_1464 ();
 FILLCELL_X32 FILLER_302_1496 ();
 FILLCELL_X32 FILLER_302_1528 ();
 FILLCELL_X32 FILLER_302_1560 ();
 FILLCELL_X32 FILLER_302_1592 ();
 FILLCELL_X32 FILLER_302_1624 ();
 FILLCELL_X32 FILLER_302_1656 ();
 FILLCELL_X32 FILLER_302_1688 ();
 FILLCELL_X32 FILLER_302_1720 ();
 FILLCELL_X32 FILLER_302_1752 ();
 FILLCELL_X32 FILLER_302_1784 ();
 FILLCELL_X32 FILLER_302_1816 ();
 FILLCELL_X32 FILLER_302_1848 ();
 FILLCELL_X8 FILLER_302_1880 ();
 FILLCELL_X4 FILLER_302_1888 ();
 FILLCELL_X2 FILLER_302_1892 ();
 FILLCELL_X32 FILLER_302_1895 ();
 FILLCELL_X32 FILLER_302_1927 ();
 FILLCELL_X32 FILLER_302_1959 ();
 FILLCELL_X32 FILLER_302_1991 ();
 FILLCELL_X32 FILLER_302_2023 ();
 FILLCELL_X32 FILLER_302_2055 ();
 FILLCELL_X32 FILLER_302_2087 ();
 FILLCELL_X32 FILLER_302_2119 ();
 FILLCELL_X32 FILLER_302_2151 ();
 FILLCELL_X32 FILLER_302_2183 ();
 FILLCELL_X32 FILLER_302_2215 ();
 FILLCELL_X32 FILLER_302_2247 ();
 FILLCELL_X32 FILLER_302_2279 ();
 FILLCELL_X32 FILLER_302_2311 ();
 FILLCELL_X32 FILLER_302_2343 ();
 FILLCELL_X32 FILLER_302_2375 ();
 FILLCELL_X32 FILLER_302_2407 ();
 FILLCELL_X32 FILLER_302_2439 ();
 FILLCELL_X32 FILLER_302_2471 ();
 FILLCELL_X32 FILLER_302_2503 ();
 FILLCELL_X32 FILLER_302_2535 ();
 FILLCELL_X32 FILLER_302_2567 ();
 FILLCELL_X32 FILLER_302_2599 ();
 FILLCELL_X32 FILLER_302_2631 ();
 FILLCELL_X32 FILLER_302_2663 ();
 FILLCELL_X32 FILLER_302_2695 ();
 FILLCELL_X32 FILLER_302_2727 ();
 FILLCELL_X32 FILLER_302_2759 ();
 FILLCELL_X32 FILLER_302_2791 ();
 FILLCELL_X32 FILLER_302_2823 ();
 FILLCELL_X32 FILLER_302_2855 ();
 FILLCELL_X32 FILLER_302_2887 ();
 FILLCELL_X32 FILLER_302_2919 ();
 FILLCELL_X32 FILLER_302_2951 ();
 FILLCELL_X32 FILLER_302_2983 ();
 FILLCELL_X32 FILLER_302_3015 ();
 FILLCELL_X32 FILLER_302_3047 ();
 FILLCELL_X32 FILLER_302_3079 ();
 FILLCELL_X32 FILLER_302_3111 ();
 FILLCELL_X8 FILLER_302_3143 ();
 FILLCELL_X4 FILLER_302_3151 ();
 FILLCELL_X2 FILLER_302_3155 ();
 FILLCELL_X32 FILLER_302_3158 ();
 FILLCELL_X32 FILLER_302_3190 ();
 FILLCELL_X32 FILLER_302_3222 ();
 FILLCELL_X32 FILLER_302_3254 ();
 FILLCELL_X32 FILLER_302_3286 ();
 FILLCELL_X32 FILLER_302_3318 ();
 FILLCELL_X32 FILLER_302_3350 ();
 FILLCELL_X32 FILLER_302_3382 ();
 FILLCELL_X32 FILLER_302_3414 ();
 FILLCELL_X32 FILLER_302_3446 ();
 FILLCELL_X32 FILLER_302_3478 ();
 FILLCELL_X32 FILLER_302_3510 ();
 FILLCELL_X32 FILLER_302_3542 ();
 FILLCELL_X32 FILLER_302_3574 ();
 FILLCELL_X32 FILLER_302_3606 ();
 FILLCELL_X32 FILLER_302_3638 ();
 FILLCELL_X32 FILLER_302_3670 ();
 FILLCELL_X32 FILLER_302_3702 ();
 FILLCELL_X4 FILLER_302_3734 ();
 FILLCELL_X32 FILLER_303_1 ();
 FILLCELL_X32 FILLER_303_33 ();
 FILLCELL_X32 FILLER_303_65 ();
 FILLCELL_X32 FILLER_303_97 ();
 FILLCELL_X32 FILLER_303_129 ();
 FILLCELL_X32 FILLER_303_161 ();
 FILLCELL_X32 FILLER_303_193 ();
 FILLCELL_X32 FILLER_303_225 ();
 FILLCELL_X32 FILLER_303_257 ();
 FILLCELL_X32 FILLER_303_289 ();
 FILLCELL_X32 FILLER_303_321 ();
 FILLCELL_X32 FILLER_303_353 ();
 FILLCELL_X32 FILLER_303_385 ();
 FILLCELL_X32 FILLER_303_417 ();
 FILLCELL_X32 FILLER_303_449 ();
 FILLCELL_X32 FILLER_303_481 ();
 FILLCELL_X32 FILLER_303_513 ();
 FILLCELL_X32 FILLER_303_545 ();
 FILLCELL_X32 FILLER_303_577 ();
 FILLCELL_X32 FILLER_303_609 ();
 FILLCELL_X32 FILLER_303_641 ();
 FILLCELL_X32 FILLER_303_673 ();
 FILLCELL_X32 FILLER_303_705 ();
 FILLCELL_X32 FILLER_303_737 ();
 FILLCELL_X32 FILLER_303_769 ();
 FILLCELL_X32 FILLER_303_801 ();
 FILLCELL_X32 FILLER_303_833 ();
 FILLCELL_X32 FILLER_303_865 ();
 FILLCELL_X32 FILLER_303_897 ();
 FILLCELL_X32 FILLER_303_929 ();
 FILLCELL_X32 FILLER_303_961 ();
 FILLCELL_X32 FILLER_303_993 ();
 FILLCELL_X32 FILLER_303_1025 ();
 FILLCELL_X32 FILLER_303_1057 ();
 FILLCELL_X32 FILLER_303_1089 ();
 FILLCELL_X32 FILLER_303_1121 ();
 FILLCELL_X32 FILLER_303_1153 ();
 FILLCELL_X32 FILLER_303_1185 ();
 FILLCELL_X32 FILLER_303_1217 ();
 FILLCELL_X8 FILLER_303_1249 ();
 FILLCELL_X4 FILLER_303_1257 ();
 FILLCELL_X2 FILLER_303_1261 ();
 FILLCELL_X32 FILLER_303_1264 ();
 FILLCELL_X32 FILLER_303_1296 ();
 FILLCELL_X32 FILLER_303_1328 ();
 FILLCELL_X32 FILLER_303_1360 ();
 FILLCELL_X32 FILLER_303_1392 ();
 FILLCELL_X32 FILLER_303_1424 ();
 FILLCELL_X32 FILLER_303_1456 ();
 FILLCELL_X32 FILLER_303_1488 ();
 FILLCELL_X32 FILLER_303_1520 ();
 FILLCELL_X32 FILLER_303_1552 ();
 FILLCELL_X32 FILLER_303_1584 ();
 FILLCELL_X32 FILLER_303_1616 ();
 FILLCELL_X32 FILLER_303_1648 ();
 FILLCELL_X32 FILLER_303_1680 ();
 FILLCELL_X32 FILLER_303_1712 ();
 FILLCELL_X32 FILLER_303_1744 ();
 FILLCELL_X32 FILLER_303_1776 ();
 FILLCELL_X32 FILLER_303_1808 ();
 FILLCELL_X32 FILLER_303_1840 ();
 FILLCELL_X32 FILLER_303_1872 ();
 FILLCELL_X32 FILLER_303_1904 ();
 FILLCELL_X32 FILLER_303_1936 ();
 FILLCELL_X32 FILLER_303_1968 ();
 FILLCELL_X32 FILLER_303_2000 ();
 FILLCELL_X32 FILLER_303_2032 ();
 FILLCELL_X32 FILLER_303_2064 ();
 FILLCELL_X32 FILLER_303_2096 ();
 FILLCELL_X32 FILLER_303_2128 ();
 FILLCELL_X32 FILLER_303_2160 ();
 FILLCELL_X32 FILLER_303_2192 ();
 FILLCELL_X32 FILLER_303_2224 ();
 FILLCELL_X32 FILLER_303_2256 ();
 FILLCELL_X32 FILLER_303_2288 ();
 FILLCELL_X32 FILLER_303_2320 ();
 FILLCELL_X32 FILLER_303_2352 ();
 FILLCELL_X32 FILLER_303_2384 ();
 FILLCELL_X32 FILLER_303_2416 ();
 FILLCELL_X32 FILLER_303_2448 ();
 FILLCELL_X32 FILLER_303_2480 ();
 FILLCELL_X8 FILLER_303_2512 ();
 FILLCELL_X4 FILLER_303_2520 ();
 FILLCELL_X2 FILLER_303_2524 ();
 FILLCELL_X32 FILLER_303_2527 ();
 FILLCELL_X32 FILLER_303_2559 ();
 FILLCELL_X32 FILLER_303_2591 ();
 FILLCELL_X32 FILLER_303_2623 ();
 FILLCELL_X32 FILLER_303_2655 ();
 FILLCELL_X32 FILLER_303_2687 ();
 FILLCELL_X32 FILLER_303_2719 ();
 FILLCELL_X32 FILLER_303_2751 ();
 FILLCELL_X32 FILLER_303_2783 ();
 FILLCELL_X32 FILLER_303_2815 ();
 FILLCELL_X32 FILLER_303_2847 ();
 FILLCELL_X32 FILLER_303_2879 ();
 FILLCELL_X32 FILLER_303_2911 ();
 FILLCELL_X32 FILLER_303_2943 ();
 FILLCELL_X32 FILLER_303_2975 ();
 FILLCELL_X32 FILLER_303_3007 ();
 FILLCELL_X32 FILLER_303_3039 ();
 FILLCELL_X32 FILLER_303_3071 ();
 FILLCELL_X32 FILLER_303_3103 ();
 FILLCELL_X32 FILLER_303_3135 ();
 FILLCELL_X32 FILLER_303_3167 ();
 FILLCELL_X32 FILLER_303_3199 ();
 FILLCELL_X32 FILLER_303_3231 ();
 FILLCELL_X32 FILLER_303_3263 ();
 FILLCELL_X32 FILLER_303_3295 ();
 FILLCELL_X32 FILLER_303_3327 ();
 FILLCELL_X32 FILLER_303_3359 ();
 FILLCELL_X32 FILLER_303_3391 ();
 FILLCELL_X32 FILLER_303_3423 ();
 FILLCELL_X32 FILLER_303_3455 ();
 FILLCELL_X32 FILLER_303_3487 ();
 FILLCELL_X32 FILLER_303_3519 ();
 FILLCELL_X32 FILLER_303_3551 ();
 FILLCELL_X32 FILLER_303_3583 ();
 FILLCELL_X32 FILLER_303_3615 ();
 FILLCELL_X32 FILLER_303_3647 ();
 FILLCELL_X32 FILLER_303_3679 ();
 FILLCELL_X16 FILLER_303_3711 ();
 FILLCELL_X8 FILLER_303_3727 ();
 FILLCELL_X2 FILLER_303_3735 ();
 FILLCELL_X1 FILLER_303_3737 ();
 FILLCELL_X32 FILLER_304_1 ();
 FILLCELL_X32 FILLER_304_33 ();
 FILLCELL_X32 FILLER_304_65 ();
 FILLCELL_X32 FILLER_304_97 ();
 FILLCELL_X32 FILLER_304_129 ();
 FILLCELL_X32 FILLER_304_161 ();
 FILLCELL_X32 FILLER_304_193 ();
 FILLCELL_X32 FILLER_304_225 ();
 FILLCELL_X32 FILLER_304_257 ();
 FILLCELL_X32 FILLER_304_289 ();
 FILLCELL_X32 FILLER_304_321 ();
 FILLCELL_X32 FILLER_304_353 ();
 FILLCELL_X32 FILLER_304_385 ();
 FILLCELL_X32 FILLER_304_417 ();
 FILLCELL_X32 FILLER_304_449 ();
 FILLCELL_X32 FILLER_304_481 ();
 FILLCELL_X32 FILLER_304_513 ();
 FILLCELL_X32 FILLER_304_545 ();
 FILLCELL_X32 FILLER_304_577 ();
 FILLCELL_X16 FILLER_304_609 ();
 FILLCELL_X4 FILLER_304_625 ();
 FILLCELL_X2 FILLER_304_629 ();
 FILLCELL_X32 FILLER_304_632 ();
 FILLCELL_X32 FILLER_304_664 ();
 FILLCELL_X32 FILLER_304_696 ();
 FILLCELL_X32 FILLER_304_728 ();
 FILLCELL_X32 FILLER_304_760 ();
 FILLCELL_X32 FILLER_304_792 ();
 FILLCELL_X32 FILLER_304_824 ();
 FILLCELL_X32 FILLER_304_856 ();
 FILLCELL_X32 FILLER_304_888 ();
 FILLCELL_X32 FILLER_304_920 ();
 FILLCELL_X32 FILLER_304_952 ();
 FILLCELL_X32 FILLER_304_984 ();
 FILLCELL_X32 FILLER_304_1016 ();
 FILLCELL_X32 FILLER_304_1048 ();
 FILLCELL_X32 FILLER_304_1080 ();
 FILLCELL_X32 FILLER_304_1112 ();
 FILLCELL_X32 FILLER_304_1144 ();
 FILLCELL_X32 FILLER_304_1176 ();
 FILLCELL_X32 FILLER_304_1208 ();
 FILLCELL_X32 FILLER_304_1240 ();
 FILLCELL_X32 FILLER_304_1272 ();
 FILLCELL_X32 FILLER_304_1304 ();
 FILLCELL_X32 FILLER_304_1336 ();
 FILLCELL_X32 FILLER_304_1368 ();
 FILLCELL_X32 FILLER_304_1400 ();
 FILLCELL_X32 FILLER_304_1432 ();
 FILLCELL_X32 FILLER_304_1464 ();
 FILLCELL_X32 FILLER_304_1496 ();
 FILLCELL_X32 FILLER_304_1528 ();
 FILLCELL_X32 FILLER_304_1560 ();
 FILLCELL_X32 FILLER_304_1592 ();
 FILLCELL_X32 FILLER_304_1624 ();
 FILLCELL_X32 FILLER_304_1656 ();
 FILLCELL_X32 FILLER_304_1688 ();
 FILLCELL_X32 FILLER_304_1720 ();
 FILLCELL_X32 FILLER_304_1752 ();
 FILLCELL_X32 FILLER_304_1784 ();
 FILLCELL_X32 FILLER_304_1816 ();
 FILLCELL_X32 FILLER_304_1848 ();
 FILLCELL_X8 FILLER_304_1880 ();
 FILLCELL_X4 FILLER_304_1888 ();
 FILLCELL_X2 FILLER_304_1892 ();
 FILLCELL_X32 FILLER_304_1895 ();
 FILLCELL_X32 FILLER_304_1927 ();
 FILLCELL_X32 FILLER_304_1959 ();
 FILLCELL_X32 FILLER_304_1991 ();
 FILLCELL_X32 FILLER_304_2023 ();
 FILLCELL_X32 FILLER_304_2055 ();
 FILLCELL_X32 FILLER_304_2087 ();
 FILLCELL_X32 FILLER_304_2119 ();
 FILLCELL_X32 FILLER_304_2151 ();
 FILLCELL_X32 FILLER_304_2183 ();
 FILLCELL_X32 FILLER_304_2215 ();
 FILLCELL_X32 FILLER_304_2247 ();
 FILLCELL_X32 FILLER_304_2279 ();
 FILLCELL_X32 FILLER_304_2311 ();
 FILLCELL_X32 FILLER_304_2343 ();
 FILLCELL_X32 FILLER_304_2375 ();
 FILLCELL_X32 FILLER_304_2407 ();
 FILLCELL_X32 FILLER_304_2439 ();
 FILLCELL_X32 FILLER_304_2471 ();
 FILLCELL_X32 FILLER_304_2503 ();
 FILLCELL_X32 FILLER_304_2535 ();
 FILLCELL_X32 FILLER_304_2567 ();
 FILLCELL_X32 FILLER_304_2599 ();
 FILLCELL_X32 FILLER_304_2631 ();
 FILLCELL_X32 FILLER_304_2663 ();
 FILLCELL_X32 FILLER_304_2695 ();
 FILLCELL_X32 FILLER_304_2727 ();
 FILLCELL_X32 FILLER_304_2759 ();
 FILLCELL_X32 FILLER_304_2791 ();
 FILLCELL_X32 FILLER_304_2823 ();
 FILLCELL_X32 FILLER_304_2855 ();
 FILLCELL_X32 FILLER_304_2887 ();
 FILLCELL_X32 FILLER_304_2919 ();
 FILLCELL_X32 FILLER_304_2951 ();
 FILLCELL_X32 FILLER_304_2983 ();
 FILLCELL_X32 FILLER_304_3015 ();
 FILLCELL_X32 FILLER_304_3047 ();
 FILLCELL_X32 FILLER_304_3079 ();
 FILLCELL_X32 FILLER_304_3111 ();
 FILLCELL_X8 FILLER_304_3143 ();
 FILLCELL_X4 FILLER_304_3151 ();
 FILLCELL_X2 FILLER_304_3155 ();
 FILLCELL_X32 FILLER_304_3158 ();
 FILLCELL_X32 FILLER_304_3190 ();
 FILLCELL_X32 FILLER_304_3222 ();
 FILLCELL_X32 FILLER_304_3254 ();
 FILLCELL_X32 FILLER_304_3286 ();
 FILLCELL_X32 FILLER_304_3318 ();
 FILLCELL_X32 FILLER_304_3350 ();
 FILLCELL_X32 FILLER_304_3382 ();
 FILLCELL_X32 FILLER_304_3414 ();
 FILLCELL_X32 FILLER_304_3446 ();
 FILLCELL_X32 FILLER_304_3478 ();
 FILLCELL_X32 FILLER_304_3510 ();
 FILLCELL_X32 FILLER_304_3542 ();
 FILLCELL_X32 FILLER_304_3574 ();
 FILLCELL_X32 FILLER_304_3606 ();
 FILLCELL_X32 FILLER_304_3638 ();
 FILLCELL_X32 FILLER_304_3670 ();
 FILLCELL_X32 FILLER_304_3702 ();
 FILLCELL_X4 FILLER_304_3734 ();
 FILLCELL_X32 FILLER_305_1 ();
 FILLCELL_X32 FILLER_305_33 ();
 FILLCELL_X32 FILLER_305_65 ();
 FILLCELL_X32 FILLER_305_97 ();
 FILLCELL_X32 FILLER_305_129 ();
 FILLCELL_X32 FILLER_305_161 ();
 FILLCELL_X32 FILLER_305_193 ();
 FILLCELL_X32 FILLER_305_225 ();
 FILLCELL_X32 FILLER_305_257 ();
 FILLCELL_X32 FILLER_305_289 ();
 FILLCELL_X32 FILLER_305_321 ();
 FILLCELL_X32 FILLER_305_353 ();
 FILLCELL_X32 FILLER_305_385 ();
 FILLCELL_X32 FILLER_305_417 ();
 FILLCELL_X32 FILLER_305_449 ();
 FILLCELL_X32 FILLER_305_481 ();
 FILLCELL_X32 FILLER_305_513 ();
 FILLCELL_X32 FILLER_305_545 ();
 FILLCELL_X32 FILLER_305_577 ();
 FILLCELL_X32 FILLER_305_609 ();
 FILLCELL_X32 FILLER_305_641 ();
 FILLCELL_X32 FILLER_305_673 ();
 FILLCELL_X32 FILLER_305_705 ();
 FILLCELL_X32 FILLER_305_737 ();
 FILLCELL_X32 FILLER_305_769 ();
 FILLCELL_X32 FILLER_305_801 ();
 FILLCELL_X32 FILLER_305_833 ();
 FILLCELL_X32 FILLER_305_865 ();
 FILLCELL_X32 FILLER_305_897 ();
 FILLCELL_X32 FILLER_305_929 ();
 FILLCELL_X32 FILLER_305_961 ();
 FILLCELL_X32 FILLER_305_993 ();
 FILLCELL_X32 FILLER_305_1025 ();
 FILLCELL_X32 FILLER_305_1057 ();
 FILLCELL_X32 FILLER_305_1089 ();
 FILLCELL_X32 FILLER_305_1121 ();
 FILLCELL_X32 FILLER_305_1153 ();
 FILLCELL_X32 FILLER_305_1185 ();
 FILLCELL_X32 FILLER_305_1217 ();
 FILLCELL_X8 FILLER_305_1249 ();
 FILLCELL_X4 FILLER_305_1257 ();
 FILLCELL_X2 FILLER_305_1261 ();
 FILLCELL_X32 FILLER_305_1264 ();
 FILLCELL_X32 FILLER_305_1296 ();
 FILLCELL_X32 FILLER_305_1328 ();
 FILLCELL_X32 FILLER_305_1360 ();
 FILLCELL_X32 FILLER_305_1392 ();
 FILLCELL_X32 FILLER_305_1424 ();
 FILLCELL_X32 FILLER_305_1456 ();
 FILLCELL_X32 FILLER_305_1488 ();
 FILLCELL_X32 FILLER_305_1520 ();
 FILLCELL_X32 FILLER_305_1552 ();
 FILLCELL_X32 FILLER_305_1584 ();
 FILLCELL_X32 FILLER_305_1616 ();
 FILLCELL_X32 FILLER_305_1648 ();
 FILLCELL_X32 FILLER_305_1680 ();
 FILLCELL_X32 FILLER_305_1712 ();
 FILLCELL_X32 FILLER_305_1744 ();
 FILLCELL_X32 FILLER_305_1776 ();
 FILLCELL_X32 FILLER_305_1808 ();
 FILLCELL_X32 FILLER_305_1840 ();
 FILLCELL_X32 FILLER_305_1872 ();
 FILLCELL_X32 FILLER_305_1904 ();
 FILLCELL_X32 FILLER_305_1936 ();
 FILLCELL_X32 FILLER_305_1968 ();
 FILLCELL_X32 FILLER_305_2000 ();
 FILLCELL_X32 FILLER_305_2032 ();
 FILLCELL_X32 FILLER_305_2064 ();
 FILLCELL_X32 FILLER_305_2096 ();
 FILLCELL_X32 FILLER_305_2128 ();
 FILLCELL_X32 FILLER_305_2160 ();
 FILLCELL_X32 FILLER_305_2192 ();
 FILLCELL_X32 FILLER_305_2224 ();
 FILLCELL_X32 FILLER_305_2256 ();
 FILLCELL_X32 FILLER_305_2288 ();
 FILLCELL_X32 FILLER_305_2320 ();
 FILLCELL_X32 FILLER_305_2352 ();
 FILLCELL_X32 FILLER_305_2384 ();
 FILLCELL_X32 FILLER_305_2416 ();
 FILLCELL_X32 FILLER_305_2448 ();
 FILLCELL_X32 FILLER_305_2480 ();
 FILLCELL_X8 FILLER_305_2512 ();
 FILLCELL_X4 FILLER_305_2520 ();
 FILLCELL_X2 FILLER_305_2524 ();
 FILLCELL_X32 FILLER_305_2527 ();
 FILLCELL_X32 FILLER_305_2559 ();
 FILLCELL_X32 FILLER_305_2591 ();
 FILLCELL_X32 FILLER_305_2623 ();
 FILLCELL_X32 FILLER_305_2655 ();
 FILLCELL_X32 FILLER_305_2687 ();
 FILLCELL_X32 FILLER_305_2719 ();
 FILLCELL_X32 FILLER_305_2751 ();
 FILLCELL_X32 FILLER_305_2783 ();
 FILLCELL_X32 FILLER_305_2815 ();
 FILLCELL_X32 FILLER_305_2847 ();
 FILLCELL_X32 FILLER_305_2879 ();
 FILLCELL_X32 FILLER_305_2911 ();
 FILLCELL_X32 FILLER_305_2943 ();
 FILLCELL_X32 FILLER_305_2975 ();
 FILLCELL_X32 FILLER_305_3007 ();
 FILLCELL_X32 FILLER_305_3039 ();
 FILLCELL_X32 FILLER_305_3071 ();
 FILLCELL_X32 FILLER_305_3103 ();
 FILLCELL_X32 FILLER_305_3135 ();
 FILLCELL_X32 FILLER_305_3167 ();
 FILLCELL_X32 FILLER_305_3199 ();
 FILLCELL_X32 FILLER_305_3231 ();
 FILLCELL_X32 FILLER_305_3263 ();
 FILLCELL_X32 FILLER_305_3295 ();
 FILLCELL_X32 FILLER_305_3327 ();
 FILLCELL_X32 FILLER_305_3359 ();
 FILLCELL_X32 FILLER_305_3391 ();
 FILLCELL_X32 FILLER_305_3423 ();
 FILLCELL_X32 FILLER_305_3455 ();
 FILLCELL_X32 FILLER_305_3487 ();
 FILLCELL_X32 FILLER_305_3519 ();
 FILLCELL_X32 FILLER_305_3551 ();
 FILLCELL_X32 FILLER_305_3583 ();
 FILLCELL_X32 FILLER_305_3615 ();
 FILLCELL_X32 FILLER_305_3647 ();
 FILLCELL_X32 FILLER_305_3679 ();
 FILLCELL_X16 FILLER_305_3711 ();
 FILLCELL_X8 FILLER_305_3727 ();
 FILLCELL_X2 FILLER_305_3735 ();
 FILLCELL_X1 FILLER_305_3737 ();
 FILLCELL_X32 FILLER_306_1 ();
 FILLCELL_X32 FILLER_306_33 ();
 FILLCELL_X32 FILLER_306_65 ();
 FILLCELL_X32 FILLER_306_97 ();
 FILLCELL_X32 FILLER_306_129 ();
 FILLCELL_X32 FILLER_306_161 ();
 FILLCELL_X32 FILLER_306_193 ();
 FILLCELL_X32 FILLER_306_225 ();
 FILLCELL_X32 FILLER_306_257 ();
 FILLCELL_X32 FILLER_306_289 ();
 FILLCELL_X32 FILLER_306_321 ();
 FILLCELL_X32 FILLER_306_353 ();
 FILLCELL_X32 FILLER_306_385 ();
 FILLCELL_X32 FILLER_306_417 ();
 FILLCELL_X32 FILLER_306_449 ();
 FILLCELL_X32 FILLER_306_481 ();
 FILLCELL_X32 FILLER_306_513 ();
 FILLCELL_X32 FILLER_306_545 ();
 FILLCELL_X32 FILLER_306_577 ();
 FILLCELL_X16 FILLER_306_609 ();
 FILLCELL_X4 FILLER_306_625 ();
 FILLCELL_X2 FILLER_306_629 ();
 FILLCELL_X32 FILLER_306_632 ();
 FILLCELL_X32 FILLER_306_664 ();
 FILLCELL_X32 FILLER_306_696 ();
 FILLCELL_X32 FILLER_306_728 ();
 FILLCELL_X32 FILLER_306_760 ();
 FILLCELL_X32 FILLER_306_792 ();
 FILLCELL_X32 FILLER_306_824 ();
 FILLCELL_X32 FILLER_306_856 ();
 FILLCELL_X32 FILLER_306_888 ();
 FILLCELL_X32 FILLER_306_920 ();
 FILLCELL_X32 FILLER_306_952 ();
 FILLCELL_X32 FILLER_306_984 ();
 FILLCELL_X32 FILLER_306_1016 ();
 FILLCELL_X32 FILLER_306_1048 ();
 FILLCELL_X32 FILLER_306_1080 ();
 FILLCELL_X32 FILLER_306_1112 ();
 FILLCELL_X32 FILLER_306_1144 ();
 FILLCELL_X32 FILLER_306_1176 ();
 FILLCELL_X32 FILLER_306_1208 ();
 FILLCELL_X32 FILLER_306_1240 ();
 FILLCELL_X32 FILLER_306_1272 ();
 FILLCELL_X32 FILLER_306_1304 ();
 FILLCELL_X32 FILLER_306_1336 ();
 FILLCELL_X32 FILLER_306_1368 ();
 FILLCELL_X32 FILLER_306_1400 ();
 FILLCELL_X32 FILLER_306_1432 ();
 FILLCELL_X32 FILLER_306_1464 ();
 FILLCELL_X32 FILLER_306_1496 ();
 FILLCELL_X32 FILLER_306_1528 ();
 FILLCELL_X32 FILLER_306_1560 ();
 FILLCELL_X32 FILLER_306_1592 ();
 FILLCELL_X32 FILLER_306_1624 ();
 FILLCELL_X32 FILLER_306_1656 ();
 FILLCELL_X32 FILLER_306_1688 ();
 FILLCELL_X32 FILLER_306_1720 ();
 FILLCELL_X32 FILLER_306_1752 ();
 FILLCELL_X32 FILLER_306_1784 ();
 FILLCELL_X32 FILLER_306_1816 ();
 FILLCELL_X32 FILLER_306_1848 ();
 FILLCELL_X8 FILLER_306_1880 ();
 FILLCELL_X4 FILLER_306_1888 ();
 FILLCELL_X2 FILLER_306_1892 ();
 FILLCELL_X32 FILLER_306_1895 ();
 FILLCELL_X32 FILLER_306_1927 ();
 FILLCELL_X32 FILLER_306_1959 ();
 FILLCELL_X32 FILLER_306_1991 ();
 FILLCELL_X32 FILLER_306_2023 ();
 FILLCELL_X32 FILLER_306_2055 ();
 FILLCELL_X32 FILLER_306_2087 ();
 FILLCELL_X32 FILLER_306_2119 ();
 FILLCELL_X32 FILLER_306_2151 ();
 FILLCELL_X32 FILLER_306_2183 ();
 FILLCELL_X32 FILLER_306_2215 ();
 FILLCELL_X32 FILLER_306_2247 ();
 FILLCELL_X32 FILLER_306_2279 ();
 FILLCELL_X32 FILLER_306_2311 ();
 FILLCELL_X32 FILLER_306_2343 ();
 FILLCELL_X32 FILLER_306_2375 ();
 FILLCELL_X32 FILLER_306_2407 ();
 FILLCELL_X32 FILLER_306_2439 ();
 FILLCELL_X32 FILLER_306_2471 ();
 FILLCELL_X32 FILLER_306_2503 ();
 FILLCELL_X32 FILLER_306_2535 ();
 FILLCELL_X32 FILLER_306_2567 ();
 FILLCELL_X32 FILLER_306_2599 ();
 FILLCELL_X32 FILLER_306_2631 ();
 FILLCELL_X32 FILLER_306_2663 ();
 FILLCELL_X32 FILLER_306_2695 ();
 FILLCELL_X32 FILLER_306_2727 ();
 FILLCELL_X32 FILLER_306_2759 ();
 FILLCELL_X32 FILLER_306_2791 ();
 FILLCELL_X32 FILLER_306_2823 ();
 FILLCELL_X32 FILLER_306_2855 ();
 FILLCELL_X32 FILLER_306_2887 ();
 FILLCELL_X32 FILLER_306_2919 ();
 FILLCELL_X32 FILLER_306_2951 ();
 FILLCELL_X32 FILLER_306_2983 ();
 FILLCELL_X32 FILLER_306_3015 ();
 FILLCELL_X32 FILLER_306_3047 ();
 FILLCELL_X32 FILLER_306_3079 ();
 FILLCELL_X32 FILLER_306_3111 ();
 FILLCELL_X8 FILLER_306_3143 ();
 FILLCELL_X4 FILLER_306_3151 ();
 FILLCELL_X2 FILLER_306_3155 ();
 FILLCELL_X32 FILLER_306_3158 ();
 FILLCELL_X32 FILLER_306_3190 ();
 FILLCELL_X32 FILLER_306_3222 ();
 FILLCELL_X32 FILLER_306_3254 ();
 FILLCELL_X32 FILLER_306_3286 ();
 FILLCELL_X32 FILLER_306_3318 ();
 FILLCELL_X32 FILLER_306_3350 ();
 FILLCELL_X32 FILLER_306_3382 ();
 FILLCELL_X32 FILLER_306_3414 ();
 FILLCELL_X32 FILLER_306_3446 ();
 FILLCELL_X32 FILLER_306_3478 ();
 FILLCELL_X32 FILLER_306_3510 ();
 FILLCELL_X32 FILLER_306_3542 ();
 FILLCELL_X32 FILLER_306_3574 ();
 FILLCELL_X32 FILLER_306_3606 ();
 FILLCELL_X32 FILLER_306_3638 ();
 FILLCELL_X32 FILLER_306_3670 ();
 FILLCELL_X32 FILLER_306_3702 ();
 FILLCELL_X4 FILLER_306_3734 ();
 FILLCELL_X32 FILLER_307_1 ();
 FILLCELL_X32 FILLER_307_33 ();
 FILLCELL_X32 FILLER_307_65 ();
 FILLCELL_X32 FILLER_307_97 ();
 FILLCELL_X32 FILLER_307_129 ();
 FILLCELL_X32 FILLER_307_161 ();
 FILLCELL_X32 FILLER_307_193 ();
 FILLCELL_X32 FILLER_307_225 ();
 FILLCELL_X32 FILLER_307_257 ();
 FILLCELL_X32 FILLER_307_289 ();
 FILLCELL_X32 FILLER_307_321 ();
 FILLCELL_X32 FILLER_307_353 ();
 FILLCELL_X32 FILLER_307_385 ();
 FILLCELL_X32 FILLER_307_417 ();
 FILLCELL_X32 FILLER_307_449 ();
 FILLCELL_X32 FILLER_307_481 ();
 FILLCELL_X32 FILLER_307_513 ();
 FILLCELL_X32 FILLER_307_545 ();
 FILLCELL_X32 FILLER_307_577 ();
 FILLCELL_X32 FILLER_307_609 ();
 FILLCELL_X32 FILLER_307_641 ();
 FILLCELL_X32 FILLER_307_673 ();
 FILLCELL_X32 FILLER_307_705 ();
 FILLCELL_X32 FILLER_307_737 ();
 FILLCELL_X32 FILLER_307_769 ();
 FILLCELL_X32 FILLER_307_801 ();
 FILLCELL_X32 FILLER_307_833 ();
 FILLCELL_X32 FILLER_307_865 ();
 FILLCELL_X32 FILLER_307_897 ();
 FILLCELL_X32 FILLER_307_929 ();
 FILLCELL_X32 FILLER_307_961 ();
 FILLCELL_X32 FILLER_307_993 ();
 FILLCELL_X32 FILLER_307_1025 ();
 FILLCELL_X32 FILLER_307_1057 ();
 FILLCELL_X32 FILLER_307_1089 ();
 FILLCELL_X32 FILLER_307_1121 ();
 FILLCELL_X32 FILLER_307_1153 ();
 FILLCELL_X32 FILLER_307_1185 ();
 FILLCELL_X32 FILLER_307_1217 ();
 FILLCELL_X8 FILLER_307_1249 ();
 FILLCELL_X4 FILLER_307_1257 ();
 FILLCELL_X2 FILLER_307_1261 ();
 FILLCELL_X32 FILLER_307_1264 ();
 FILLCELL_X32 FILLER_307_1296 ();
 FILLCELL_X32 FILLER_307_1328 ();
 FILLCELL_X32 FILLER_307_1360 ();
 FILLCELL_X32 FILLER_307_1392 ();
 FILLCELL_X32 FILLER_307_1424 ();
 FILLCELL_X32 FILLER_307_1456 ();
 FILLCELL_X32 FILLER_307_1488 ();
 FILLCELL_X32 FILLER_307_1520 ();
 FILLCELL_X32 FILLER_307_1552 ();
 FILLCELL_X32 FILLER_307_1584 ();
 FILLCELL_X32 FILLER_307_1616 ();
 FILLCELL_X32 FILLER_307_1648 ();
 FILLCELL_X32 FILLER_307_1680 ();
 FILLCELL_X32 FILLER_307_1712 ();
 FILLCELL_X32 FILLER_307_1744 ();
 FILLCELL_X32 FILLER_307_1776 ();
 FILLCELL_X32 FILLER_307_1808 ();
 FILLCELL_X32 FILLER_307_1840 ();
 FILLCELL_X32 FILLER_307_1872 ();
 FILLCELL_X32 FILLER_307_1904 ();
 FILLCELL_X32 FILLER_307_1936 ();
 FILLCELL_X32 FILLER_307_1968 ();
 FILLCELL_X32 FILLER_307_2000 ();
 FILLCELL_X32 FILLER_307_2032 ();
 FILLCELL_X32 FILLER_307_2064 ();
 FILLCELL_X32 FILLER_307_2096 ();
 FILLCELL_X32 FILLER_307_2128 ();
 FILLCELL_X32 FILLER_307_2160 ();
 FILLCELL_X32 FILLER_307_2192 ();
 FILLCELL_X32 FILLER_307_2224 ();
 FILLCELL_X32 FILLER_307_2256 ();
 FILLCELL_X32 FILLER_307_2288 ();
 FILLCELL_X32 FILLER_307_2320 ();
 FILLCELL_X32 FILLER_307_2352 ();
 FILLCELL_X32 FILLER_307_2384 ();
 FILLCELL_X32 FILLER_307_2416 ();
 FILLCELL_X32 FILLER_307_2448 ();
 FILLCELL_X32 FILLER_307_2480 ();
 FILLCELL_X8 FILLER_307_2512 ();
 FILLCELL_X4 FILLER_307_2520 ();
 FILLCELL_X2 FILLER_307_2524 ();
 FILLCELL_X32 FILLER_307_2527 ();
 FILLCELL_X32 FILLER_307_2559 ();
 FILLCELL_X32 FILLER_307_2591 ();
 FILLCELL_X32 FILLER_307_2623 ();
 FILLCELL_X32 FILLER_307_2655 ();
 FILLCELL_X32 FILLER_307_2687 ();
 FILLCELL_X32 FILLER_307_2719 ();
 FILLCELL_X32 FILLER_307_2751 ();
 FILLCELL_X32 FILLER_307_2783 ();
 FILLCELL_X32 FILLER_307_2815 ();
 FILLCELL_X32 FILLER_307_2847 ();
 FILLCELL_X32 FILLER_307_2879 ();
 FILLCELL_X32 FILLER_307_2911 ();
 FILLCELL_X32 FILLER_307_2943 ();
 FILLCELL_X32 FILLER_307_2975 ();
 FILLCELL_X32 FILLER_307_3007 ();
 FILLCELL_X32 FILLER_307_3039 ();
 FILLCELL_X32 FILLER_307_3071 ();
 FILLCELL_X32 FILLER_307_3103 ();
 FILLCELL_X32 FILLER_307_3135 ();
 FILLCELL_X32 FILLER_307_3167 ();
 FILLCELL_X32 FILLER_307_3199 ();
 FILLCELL_X32 FILLER_307_3231 ();
 FILLCELL_X32 FILLER_307_3263 ();
 FILLCELL_X32 FILLER_307_3295 ();
 FILLCELL_X32 FILLER_307_3327 ();
 FILLCELL_X32 FILLER_307_3359 ();
 FILLCELL_X32 FILLER_307_3391 ();
 FILLCELL_X32 FILLER_307_3423 ();
 FILLCELL_X32 FILLER_307_3455 ();
 FILLCELL_X32 FILLER_307_3487 ();
 FILLCELL_X32 FILLER_307_3519 ();
 FILLCELL_X32 FILLER_307_3551 ();
 FILLCELL_X32 FILLER_307_3583 ();
 FILLCELL_X32 FILLER_307_3615 ();
 FILLCELL_X32 FILLER_307_3647 ();
 FILLCELL_X32 FILLER_307_3679 ();
 FILLCELL_X16 FILLER_307_3711 ();
 FILLCELL_X8 FILLER_307_3727 ();
 FILLCELL_X2 FILLER_307_3735 ();
 FILLCELL_X1 FILLER_307_3737 ();
 FILLCELL_X32 FILLER_308_1 ();
 FILLCELL_X32 FILLER_308_33 ();
 FILLCELL_X32 FILLER_308_65 ();
 FILLCELL_X32 FILLER_308_97 ();
 FILLCELL_X32 FILLER_308_129 ();
 FILLCELL_X32 FILLER_308_161 ();
 FILLCELL_X32 FILLER_308_193 ();
 FILLCELL_X32 FILLER_308_225 ();
 FILLCELL_X32 FILLER_308_257 ();
 FILLCELL_X32 FILLER_308_289 ();
 FILLCELL_X32 FILLER_308_321 ();
 FILLCELL_X32 FILLER_308_353 ();
 FILLCELL_X32 FILLER_308_385 ();
 FILLCELL_X32 FILLER_308_417 ();
 FILLCELL_X32 FILLER_308_449 ();
 FILLCELL_X32 FILLER_308_481 ();
 FILLCELL_X32 FILLER_308_513 ();
 FILLCELL_X32 FILLER_308_545 ();
 FILLCELL_X32 FILLER_308_577 ();
 FILLCELL_X16 FILLER_308_609 ();
 FILLCELL_X4 FILLER_308_625 ();
 FILLCELL_X2 FILLER_308_629 ();
 FILLCELL_X32 FILLER_308_632 ();
 FILLCELL_X32 FILLER_308_664 ();
 FILLCELL_X32 FILLER_308_696 ();
 FILLCELL_X32 FILLER_308_728 ();
 FILLCELL_X32 FILLER_308_760 ();
 FILLCELL_X32 FILLER_308_792 ();
 FILLCELL_X32 FILLER_308_824 ();
 FILLCELL_X32 FILLER_308_856 ();
 FILLCELL_X32 FILLER_308_888 ();
 FILLCELL_X32 FILLER_308_920 ();
 FILLCELL_X32 FILLER_308_952 ();
 FILLCELL_X32 FILLER_308_984 ();
 FILLCELL_X32 FILLER_308_1016 ();
 FILLCELL_X32 FILLER_308_1048 ();
 FILLCELL_X32 FILLER_308_1080 ();
 FILLCELL_X32 FILLER_308_1112 ();
 FILLCELL_X32 FILLER_308_1144 ();
 FILLCELL_X32 FILLER_308_1176 ();
 FILLCELL_X32 FILLER_308_1208 ();
 FILLCELL_X32 FILLER_308_1240 ();
 FILLCELL_X32 FILLER_308_1272 ();
 FILLCELL_X32 FILLER_308_1304 ();
 FILLCELL_X32 FILLER_308_1336 ();
 FILLCELL_X32 FILLER_308_1368 ();
 FILLCELL_X32 FILLER_308_1400 ();
 FILLCELL_X32 FILLER_308_1432 ();
 FILLCELL_X32 FILLER_308_1464 ();
 FILLCELL_X32 FILLER_308_1496 ();
 FILLCELL_X32 FILLER_308_1528 ();
 FILLCELL_X32 FILLER_308_1560 ();
 FILLCELL_X32 FILLER_308_1592 ();
 FILLCELL_X32 FILLER_308_1624 ();
 FILLCELL_X32 FILLER_308_1656 ();
 FILLCELL_X32 FILLER_308_1688 ();
 FILLCELL_X32 FILLER_308_1720 ();
 FILLCELL_X32 FILLER_308_1752 ();
 FILLCELL_X32 FILLER_308_1784 ();
 FILLCELL_X32 FILLER_308_1816 ();
 FILLCELL_X32 FILLER_308_1848 ();
 FILLCELL_X8 FILLER_308_1880 ();
 FILLCELL_X4 FILLER_308_1888 ();
 FILLCELL_X2 FILLER_308_1892 ();
 FILLCELL_X32 FILLER_308_1895 ();
 FILLCELL_X32 FILLER_308_1927 ();
 FILLCELL_X32 FILLER_308_1959 ();
 FILLCELL_X32 FILLER_308_1991 ();
 FILLCELL_X32 FILLER_308_2023 ();
 FILLCELL_X32 FILLER_308_2055 ();
 FILLCELL_X32 FILLER_308_2087 ();
 FILLCELL_X32 FILLER_308_2119 ();
 FILLCELL_X32 FILLER_308_2151 ();
 FILLCELL_X32 FILLER_308_2183 ();
 FILLCELL_X32 FILLER_308_2215 ();
 FILLCELL_X32 FILLER_308_2247 ();
 FILLCELL_X32 FILLER_308_2279 ();
 FILLCELL_X32 FILLER_308_2311 ();
 FILLCELL_X32 FILLER_308_2343 ();
 FILLCELL_X32 FILLER_308_2375 ();
 FILLCELL_X32 FILLER_308_2407 ();
 FILLCELL_X32 FILLER_308_2439 ();
 FILLCELL_X32 FILLER_308_2471 ();
 FILLCELL_X32 FILLER_308_2503 ();
 FILLCELL_X32 FILLER_308_2535 ();
 FILLCELL_X32 FILLER_308_2567 ();
 FILLCELL_X32 FILLER_308_2599 ();
 FILLCELL_X32 FILLER_308_2631 ();
 FILLCELL_X32 FILLER_308_2663 ();
 FILLCELL_X32 FILLER_308_2695 ();
 FILLCELL_X32 FILLER_308_2727 ();
 FILLCELL_X32 FILLER_308_2759 ();
 FILLCELL_X32 FILLER_308_2791 ();
 FILLCELL_X32 FILLER_308_2823 ();
 FILLCELL_X32 FILLER_308_2855 ();
 FILLCELL_X32 FILLER_308_2887 ();
 FILLCELL_X32 FILLER_308_2919 ();
 FILLCELL_X32 FILLER_308_2951 ();
 FILLCELL_X32 FILLER_308_2983 ();
 FILLCELL_X32 FILLER_308_3015 ();
 FILLCELL_X32 FILLER_308_3047 ();
 FILLCELL_X32 FILLER_308_3079 ();
 FILLCELL_X32 FILLER_308_3111 ();
 FILLCELL_X8 FILLER_308_3143 ();
 FILLCELL_X4 FILLER_308_3151 ();
 FILLCELL_X2 FILLER_308_3155 ();
 FILLCELL_X32 FILLER_308_3158 ();
 FILLCELL_X32 FILLER_308_3190 ();
 FILLCELL_X32 FILLER_308_3222 ();
 FILLCELL_X32 FILLER_308_3254 ();
 FILLCELL_X32 FILLER_308_3286 ();
 FILLCELL_X32 FILLER_308_3318 ();
 FILLCELL_X32 FILLER_308_3350 ();
 FILLCELL_X32 FILLER_308_3382 ();
 FILLCELL_X32 FILLER_308_3414 ();
 FILLCELL_X32 FILLER_308_3446 ();
 FILLCELL_X32 FILLER_308_3478 ();
 FILLCELL_X32 FILLER_308_3510 ();
 FILLCELL_X32 FILLER_308_3542 ();
 FILLCELL_X32 FILLER_308_3574 ();
 FILLCELL_X32 FILLER_308_3606 ();
 FILLCELL_X32 FILLER_308_3638 ();
 FILLCELL_X32 FILLER_308_3670 ();
 FILLCELL_X32 FILLER_308_3702 ();
 FILLCELL_X4 FILLER_308_3734 ();
 FILLCELL_X32 FILLER_309_1 ();
 FILLCELL_X32 FILLER_309_33 ();
 FILLCELL_X32 FILLER_309_65 ();
 FILLCELL_X32 FILLER_309_97 ();
 FILLCELL_X32 FILLER_309_129 ();
 FILLCELL_X32 FILLER_309_161 ();
 FILLCELL_X32 FILLER_309_193 ();
 FILLCELL_X32 FILLER_309_225 ();
 FILLCELL_X32 FILLER_309_257 ();
 FILLCELL_X32 FILLER_309_289 ();
 FILLCELL_X32 FILLER_309_321 ();
 FILLCELL_X32 FILLER_309_353 ();
 FILLCELL_X32 FILLER_309_385 ();
 FILLCELL_X32 FILLER_309_417 ();
 FILLCELL_X32 FILLER_309_449 ();
 FILLCELL_X32 FILLER_309_481 ();
 FILLCELL_X32 FILLER_309_513 ();
 FILLCELL_X32 FILLER_309_545 ();
 FILLCELL_X32 FILLER_309_577 ();
 FILLCELL_X32 FILLER_309_609 ();
 FILLCELL_X32 FILLER_309_641 ();
 FILLCELL_X32 FILLER_309_673 ();
 FILLCELL_X32 FILLER_309_705 ();
 FILLCELL_X32 FILLER_309_737 ();
 FILLCELL_X32 FILLER_309_769 ();
 FILLCELL_X32 FILLER_309_801 ();
 FILLCELL_X32 FILLER_309_833 ();
 FILLCELL_X32 FILLER_309_865 ();
 FILLCELL_X32 FILLER_309_897 ();
 FILLCELL_X32 FILLER_309_929 ();
 FILLCELL_X32 FILLER_309_961 ();
 FILLCELL_X32 FILLER_309_993 ();
 FILLCELL_X32 FILLER_309_1025 ();
 FILLCELL_X32 FILLER_309_1057 ();
 FILLCELL_X32 FILLER_309_1089 ();
 FILLCELL_X32 FILLER_309_1121 ();
 FILLCELL_X32 FILLER_309_1153 ();
 FILLCELL_X32 FILLER_309_1185 ();
 FILLCELL_X32 FILLER_309_1217 ();
 FILLCELL_X8 FILLER_309_1249 ();
 FILLCELL_X4 FILLER_309_1257 ();
 FILLCELL_X2 FILLER_309_1261 ();
 FILLCELL_X32 FILLER_309_1264 ();
 FILLCELL_X32 FILLER_309_1296 ();
 FILLCELL_X32 FILLER_309_1328 ();
 FILLCELL_X32 FILLER_309_1360 ();
 FILLCELL_X32 FILLER_309_1392 ();
 FILLCELL_X32 FILLER_309_1424 ();
 FILLCELL_X32 FILLER_309_1456 ();
 FILLCELL_X32 FILLER_309_1488 ();
 FILLCELL_X32 FILLER_309_1520 ();
 FILLCELL_X32 FILLER_309_1552 ();
 FILLCELL_X32 FILLER_309_1584 ();
 FILLCELL_X32 FILLER_309_1616 ();
 FILLCELL_X32 FILLER_309_1648 ();
 FILLCELL_X32 FILLER_309_1680 ();
 FILLCELL_X32 FILLER_309_1712 ();
 FILLCELL_X32 FILLER_309_1744 ();
 FILLCELL_X32 FILLER_309_1776 ();
 FILLCELL_X32 FILLER_309_1808 ();
 FILLCELL_X32 FILLER_309_1840 ();
 FILLCELL_X32 FILLER_309_1872 ();
 FILLCELL_X32 FILLER_309_1904 ();
 FILLCELL_X32 FILLER_309_1936 ();
 FILLCELL_X32 FILLER_309_1968 ();
 FILLCELL_X32 FILLER_309_2000 ();
 FILLCELL_X32 FILLER_309_2032 ();
 FILLCELL_X32 FILLER_309_2064 ();
 FILLCELL_X32 FILLER_309_2096 ();
 FILLCELL_X32 FILLER_309_2128 ();
 FILLCELL_X32 FILLER_309_2160 ();
 FILLCELL_X32 FILLER_309_2192 ();
 FILLCELL_X32 FILLER_309_2224 ();
 FILLCELL_X32 FILLER_309_2256 ();
 FILLCELL_X32 FILLER_309_2288 ();
 FILLCELL_X32 FILLER_309_2320 ();
 FILLCELL_X32 FILLER_309_2352 ();
 FILLCELL_X32 FILLER_309_2384 ();
 FILLCELL_X32 FILLER_309_2416 ();
 FILLCELL_X32 FILLER_309_2448 ();
 FILLCELL_X32 FILLER_309_2480 ();
 FILLCELL_X8 FILLER_309_2512 ();
 FILLCELL_X4 FILLER_309_2520 ();
 FILLCELL_X2 FILLER_309_2524 ();
 FILLCELL_X32 FILLER_309_2527 ();
 FILLCELL_X32 FILLER_309_2559 ();
 FILLCELL_X32 FILLER_309_2591 ();
 FILLCELL_X32 FILLER_309_2623 ();
 FILLCELL_X32 FILLER_309_2655 ();
 FILLCELL_X32 FILLER_309_2687 ();
 FILLCELL_X32 FILLER_309_2719 ();
 FILLCELL_X32 FILLER_309_2751 ();
 FILLCELL_X32 FILLER_309_2783 ();
 FILLCELL_X32 FILLER_309_2815 ();
 FILLCELL_X32 FILLER_309_2847 ();
 FILLCELL_X32 FILLER_309_2879 ();
 FILLCELL_X32 FILLER_309_2911 ();
 FILLCELL_X32 FILLER_309_2943 ();
 FILLCELL_X32 FILLER_309_2975 ();
 FILLCELL_X32 FILLER_309_3007 ();
 FILLCELL_X32 FILLER_309_3039 ();
 FILLCELL_X32 FILLER_309_3071 ();
 FILLCELL_X32 FILLER_309_3103 ();
 FILLCELL_X32 FILLER_309_3135 ();
 FILLCELL_X32 FILLER_309_3167 ();
 FILLCELL_X32 FILLER_309_3199 ();
 FILLCELL_X32 FILLER_309_3231 ();
 FILLCELL_X32 FILLER_309_3263 ();
 FILLCELL_X32 FILLER_309_3295 ();
 FILLCELL_X32 FILLER_309_3327 ();
 FILLCELL_X32 FILLER_309_3359 ();
 FILLCELL_X32 FILLER_309_3391 ();
 FILLCELL_X32 FILLER_309_3423 ();
 FILLCELL_X32 FILLER_309_3455 ();
 FILLCELL_X32 FILLER_309_3487 ();
 FILLCELL_X32 FILLER_309_3519 ();
 FILLCELL_X32 FILLER_309_3551 ();
 FILLCELL_X32 FILLER_309_3583 ();
 FILLCELL_X32 FILLER_309_3615 ();
 FILLCELL_X32 FILLER_309_3647 ();
 FILLCELL_X32 FILLER_309_3679 ();
 FILLCELL_X16 FILLER_309_3711 ();
 FILLCELL_X8 FILLER_309_3727 ();
 FILLCELL_X2 FILLER_309_3735 ();
 FILLCELL_X1 FILLER_309_3737 ();
 FILLCELL_X32 FILLER_310_1 ();
 FILLCELL_X32 FILLER_310_33 ();
 FILLCELL_X32 FILLER_310_65 ();
 FILLCELL_X32 FILLER_310_97 ();
 FILLCELL_X32 FILLER_310_129 ();
 FILLCELL_X32 FILLER_310_161 ();
 FILLCELL_X32 FILLER_310_193 ();
 FILLCELL_X32 FILLER_310_225 ();
 FILLCELL_X32 FILLER_310_257 ();
 FILLCELL_X32 FILLER_310_289 ();
 FILLCELL_X32 FILLER_310_321 ();
 FILLCELL_X32 FILLER_310_353 ();
 FILLCELL_X32 FILLER_310_385 ();
 FILLCELL_X32 FILLER_310_417 ();
 FILLCELL_X32 FILLER_310_449 ();
 FILLCELL_X32 FILLER_310_481 ();
 FILLCELL_X32 FILLER_310_513 ();
 FILLCELL_X32 FILLER_310_545 ();
 FILLCELL_X32 FILLER_310_577 ();
 FILLCELL_X16 FILLER_310_609 ();
 FILLCELL_X4 FILLER_310_625 ();
 FILLCELL_X2 FILLER_310_629 ();
 FILLCELL_X32 FILLER_310_632 ();
 FILLCELL_X32 FILLER_310_664 ();
 FILLCELL_X32 FILLER_310_696 ();
 FILLCELL_X32 FILLER_310_728 ();
 FILLCELL_X32 FILLER_310_760 ();
 FILLCELL_X32 FILLER_310_792 ();
 FILLCELL_X32 FILLER_310_824 ();
 FILLCELL_X32 FILLER_310_856 ();
 FILLCELL_X32 FILLER_310_888 ();
 FILLCELL_X32 FILLER_310_920 ();
 FILLCELL_X32 FILLER_310_952 ();
 FILLCELL_X32 FILLER_310_984 ();
 FILLCELL_X32 FILLER_310_1016 ();
 FILLCELL_X32 FILLER_310_1048 ();
 FILLCELL_X32 FILLER_310_1080 ();
 FILLCELL_X32 FILLER_310_1112 ();
 FILLCELL_X32 FILLER_310_1144 ();
 FILLCELL_X32 FILLER_310_1176 ();
 FILLCELL_X32 FILLER_310_1208 ();
 FILLCELL_X32 FILLER_310_1240 ();
 FILLCELL_X32 FILLER_310_1272 ();
 FILLCELL_X32 FILLER_310_1304 ();
 FILLCELL_X32 FILLER_310_1336 ();
 FILLCELL_X32 FILLER_310_1368 ();
 FILLCELL_X32 FILLER_310_1400 ();
 FILLCELL_X32 FILLER_310_1432 ();
 FILLCELL_X32 FILLER_310_1464 ();
 FILLCELL_X32 FILLER_310_1496 ();
 FILLCELL_X32 FILLER_310_1528 ();
 FILLCELL_X32 FILLER_310_1560 ();
 FILLCELL_X32 FILLER_310_1592 ();
 FILLCELL_X32 FILLER_310_1624 ();
 FILLCELL_X32 FILLER_310_1656 ();
 FILLCELL_X32 FILLER_310_1688 ();
 FILLCELL_X32 FILLER_310_1720 ();
 FILLCELL_X32 FILLER_310_1752 ();
 FILLCELL_X32 FILLER_310_1784 ();
 FILLCELL_X32 FILLER_310_1816 ();
 FILLCELL_X32 FILLER_310_1848 ();
 FILLCELL_X8 FILLER_310_1880 ();
 FILLCELL_X4 FILLER_310_1888 ();
 FILLCELL_X2 FILLER_310_1892 ();
 FILLCELL_X32 FILLER_310_1895 ();
 FILLCELL_X32 FILLER_310_1927 ();
 FILLCELL_X32 FILLER_310_1959 ();
 FILLCELL_X32 FILLER_310_1991 ();
 FILLCELL_X32 FILLER_310_2023 ();
 FILLCELL_X32 FILLER_310_2055 ();
 FILLCELL_X32 FILLER_310_2087 ();
 FILLCELL_X32 FILLER_310_2119 ();
 FILLCELL_X32 FILLER_310_2151 ();
 FILLCELL_X32 FILLER_310_2183 ();
 FILLCELL_X32 FILLER_310_2215 ();
 FILLCELL_X32 FILLER_310_2247 ();
 FILLCELL_X32 FILLER_310_2279 ();
 FILLCELL_X32 FILLER_310_2311 ();
 FILLCELL_X32 FILLER_310_2343 ();
 FILLCELL_X32 FILLER_310_2375 ();
 FILLCELL_X32 FILLER_310_2407 ();
 FILLCELL_X32 FILLER_310_2439 ();
 FILLCELL_X32 FILLER_310_2471 ();
 FILLCELL_X32 FILLER_310_2503 ();
 FILLCELL_X32 FILLER_310_2535 ();
 FILLCELL_X32 FILLER_310_2567 ();
 FILLCELL_X32 FILLER_310_2599 ();
 FILLCELL_X32 FILLER_310_2631 ();
 FILLCELL_X32 FILLER_310_2663 ();
 FILLCELL_X32 FILLER_310_2695 ();
 FILLCELL_X32 FILLER_310_2727 ();
 FILLCELL_X32 FILLER_310_2759 ();
 FILLCELL_X32 FILLER_310_2791 ();
 FILLCELL_X32 FILLER_310_2823 ();
 FILLCELL_X32 FILLER_310_2855 ();
 FILLCELL_X32 FILLER_310_2887 ();
 FILLCELL_X32 FILLER_310_2919 ();
 FILLCELL_X32 FILLER_310_2951 ();
 FILLCELL_X32 FILLER_310_2983 ();
 FILLCELL_X32 FILLER_310_3015 ();
 FILLCELL_X32 FILLER_310_3047 ();
 FILLCELL_X32 FILLER_310_3079 ();
 FILLCELL_X32 FILLER_310_3111 ();
 FILLCELL_X8 FILLER_310_3143 ();
 FILLCELL_X4 FILLER_310_3151 ();
 FILLCELL_X2 FILLER_310_3155 ();
 FILLCELL_X32 FILLER_310_3158 ();
 FILLCELL_X32 FILLER_310_3190 ();
 FILLCELL_X32 FILLER_310_3222 ();
 FILLCELL_X32 FILLER_310_3254 ();
 FILLCELL_X32 FILLER_310_3286 ();
 FILLCELL_X32 FILLER_310_3318 ();
 FILLCELL_X32 FILLER_310_3350 ();
 FILLCELL_X32 FILLER_310_3382 ();
 FILLCELL_X32 FILLER_310_3414 ();
 FILLCELL_X32 FILLER_310_3446 ();
 FILLCELL_X32 FILLER_310_3478 ();
 FILLCELL_X32 FILLER_310_3510 ();
 FILLCELL_X32 FILLER_310_3542 ();
 FILLCELL_X32 FILLER_310_3574 ();
 FILLCELL_X32 FILLER_310_3606 ();
 FILLCELL_X32 FILLER_310_3638 ();
 FILLCELL_X32 FILLER_310_3670 ();
 FILLCELL_X32 FILLER_310_3702 ();
 FILLCELL_X4 FILLER_310_3734 ();
 FILLCELL_X32 FILLER_311_1 ();
 FILLCELL_X32 FILLER_311_33 ();
 FILLCELL_X32 FILLER_311_65 ();
 FILLCELL_X32 FILLER_311_97 ();
 FILLCELL_X32 FILLER_311_129 ();
 FILLCELL_X32 FILLER_311_161 ();
 FILLCELL_X32 FILLER_311_193 ();
 FILLCELL_X32 FILLER_311_225 ();
 FILLCELL_X32 FILLER_311_257 ();
 FILLCELL_X32 FILLER_311_289 ();
 FILLCELL_X32 FILLER_311_321 ();
 FILLCELL_X32 FILLER_311_353 ();
 FILLCELL_X32 FILLER_311_385 ();
 FILLCELL_X32 FILLER_311_417 ();
 FILLCELL_X32 FILLER_311_449 ();
 FILLCELL_X32 FILLER_311_481 ();
 FILLCELL_X32 FILLER_311_513 ();
 FILLCELL_X32 FILLER_311_545 ();
 FILLCELL_X32 FILLER_311_577 ();
 FILLCELL_X32 FILLER_311_609 ();
 FILLCELL_X32 FILLER_311_641 ();
 FILLCELL_X32 FILLER_311_673 ();
 FILLCELL_X32 FILLER_311_705 ();
 FILLCELL_X32 FILLER_311_737 ();
 FILLCELL_X32 FILLER_311_769 ();
 FILLCELL_X32 FILLER_311_801 ();
 FILLCELL_X32 FILLER_311_833 ();
 FILLCELL_X32 FILLER_311_865 ();
 FILLCELL_X32 FILLER_311_897 ();
 FILLCELL_X32 FILLER_311_929 ();
 FILLCELL_X32 FILLER_311_961 ();
 FILLCELL_X32 FILLER_311_993 ();
 FILLCELL_X32 FILLER_311_1025 ();
 FILLCELL_X32 FILLER_311_1057 ();
 FILLCELL_X32 FILLER_311_1089 ();
 FILLCELL_X32 FILLER_311_1121 ();
 FILLCELL_X32 FILLER_311_1153 ();
 FILLCELL_X32 FILLER_311_1185 ();
 FILLCELL_X32 FILLER_311_1217 ();
 FILLCELL_X8 FILLER_311_1249 ();
 FILLCELL_X4 FILLER_311_1257 ();
 FILLCELL_X2 FILLER_311_1261 ();
 FILLCELL_X32 FILLER_311_1264 ();
 FILLCELL_X32 FILLER_311_1296 ();
 FILLCELL_X32 FILLER_311_1328 ();
 FILLCELL_X32 FILLER_311_1360 ();
 FILLCELL_X32 FILLER_311_1392 ();
 FILLCELL_X32 FILLER_311_1424 ();
 FILLCELL_X32 FILLER_311_1456 ();
 FILLCELL_X32 FILLER_311_1488 ();
 FILLCELL_X32 FILLER_311_1520 ();
 FILLCELL_X32 FILLER_311_1552 ();
 FILLCELL_X32 FILLER_311_1584 ();
 FILLCELL_X32 FILLER_311_1616 ();
 FILLCELL_X32 FILLER_311_1648 ();
 FILLCELL_X32 FILLER_311_1680 ();
 FILLCELL_X32 FILLER_311_1712 ();
 FILLCELL_X32 FILLER_311_1744 ();
 FILLCELL_X32 FILLER_311_1776 ();
 FILLCELL_X32 FILLER_311_1808 ();
 FILLCELL_X32 FILLER_311_1840 ();
 FILLCELL_X32 FILLER_311_1872 ();
 FILLCELL_X32 FILLER_311_1904 ();
 FILLCELL_X32 FILLER_311_1936 ();
 FILLCELL_X32 FILLER_311_1968 ();
 FILLCELL_X32 FILLER_311_2000 ();
 FILLCELL_X32 FILLER_311_2032 ();
 FILLCELL_X32 FILLER_311_2064 ();
 FILLCELL_X32 FILLER_311_2096 ();
 FILLCELL_X32 FILLER_311_2128 ();
 FILLCELL_X32 FILLER_311_2160 ();
 FILLCELL_X32 FILLER_311_2192 ();
 FILLCELL_X32 FILLER_311_2224 ();
 FILLCELL_X32 FILLER_311_2256 ();
 FILLCELL_X32 FILLER_311_2288 ();
 FILLCELL_X32 FILLER_311_2320 ();
 FILLCELL_X32 FILLER_311_2352 ();
 FILLCELL_X32 FILLER_311_2384 ();
 FILLCELL_X32 FILLER_311_2416 ();
 FILLCELL_X32 FILLER_311_2448 ();
 FILLCELL_X32 FILLER_311_2480 ();
 FILLCELL_X8 FILLER_311_2512 ();
 FILLCELL_X4 FILLER_311_2520 ();
 FILLCELL_X2 FILLER_311_2524 ();
 FILLCELL_X32 FILLER_311_2527 ();
 FILLCELL_X32 FILLER_311_2559 ();
 FILLCELL_X32 FILLER_311_2591 ();
 FILLCELL_X32 FILLER_311_2623 ();
 FILLCELL_X32 FILLER_311_2655 ();
 FILLCELL_X32 FILLER_311_2687 ();
 FILLCELL_X32 FILLER_311_2719 ();
 FILLCELL_X32 FILLER_311_2751 ();
 FILLCELL_X32 FILLER_311_2783 ();
 FILLCELL_X32 FILLER_311_2815 ();
 FILLCELL_X32 FILLER_311_2847 ();
 FILLCELL_X32 FILLER_311_2879 ();
 FILLCELL_X32 FILLER_311_2911 ();
 FILLCELL_X32 FILLER_311_2943 ();
 FILLCELL_X32 FILLER_311_2975 ();
 FILLCELL_X32 FILLER_311_3007 ();
 FILLCELL_X32 FILLER_311_3039 ();
 FILLCELL_X32 FILLER_311_3071 ();
 FILLCELL_X32 FILLER_311_3103 ();
 FILLCELL_X32 FILLER_311_3135 ();
 FILLCELL_X32 FILLER_311_3167 ();
 FILLCELL_X32 FILLER_311_3199 ();
 FILLCELL_X32 FILLER_311_3231 ();
 FILLCELL_X32 FILLER_311_3263 ();
 FILLCELL_X32 FILLER_311_3295 ();
 FILLCELL_X32 FILLER_311_3327 ();
 FILLCELL_X32 FILLER_311_3359 ();
 FILLCELL_X32 FILLER_311_3391 ();
 FILLCELL_X32 FILLER_311_3423 ();
 FILLCELL_X32 FILLER_311_3455 ();
 FILLCELL_X32 FILLER_311_3487 ();
 FILLCELL_X32 FILLER_311_3519 ();
 FILLCELL_X32 FILLER_311_3551 ();
 FILLCELL_X32 FILLER_311_3583 ();
 FILLCELL_X32 FILLER_311_3615 ();
 FILLCELL_X32 FILLER_311_3647 ();
 FILLCELL_X32 FILLER_311_3679 ();
 FILLCELL_X16 FILLER_311_3711 ();
 FILLCELL_X8 FILLER_311_3727 ();
 FILLCELL_X2 FILLER_311_3735 ();
 FILLCELL_X1 FILLER_311_3737 ();
 FILLCELL_X32 FILLER_312_1 ();
 FILLCELL_X32 FILLER_312_33 ();
 FILLCELL_X32 FILLER_312_65 ();
 FILLCELL_X32 FILLER_312_97 ();
 FILLCELL_X32 FILLER_312_129 ();
 FILLCELL_X32 FILLER_312_161 ();
 FILLCELL_X32 FILLER_312_193 ();
 FILLCELL_X32 FILLER_312_225 ();
 FILLCELL_X32 FILLER_312_257 ();
 FILLCELL_X32 FILLER_312_289 ();
 FILLCELL_X32 FILLER_312_321 ();
 FILLCELL_X32 FILLER_312_353 ();
 FILLCELL_X32 FILLER_312_385 ();
 FILLCELL_X32 FILLER_312_417 ();
 FILLCELL_X32 FILLER_312_449 ();
 FILLCELL_X32 FILLER_312_481 ();
 FILLCELL_X32 FILLER_312_513 ();
 FILLCELL_X32 FILLER_312_545 ();
 FILLCELL_X32 FILLER_312_577 ();
 FILLCELL_X16 FILLER_312_609 ();
 FILLCELL_X4 FILLER_312_625 ();
 FILLCELL_X2 FILLER_312_629 ();
 FILLCELL_X32 FILLER_312_632 ();
 FILLCELL_X32 FILLER_312_664 ();
 FILLCELL_X32 FILLER_312_696 ();
 FILLCELL_X32 FILLER_312_728 ();
 FILLCELL_X32 FILLER_312_760 ();
 FILLCELL_X32 FILLER_312_792 ();
 FILLCELL_X32 FILLER_312_824 ();
 FILLCELL_X32 FILLER_312_856 ();
 FILLCELL_X32 FILLER_312_888 ();
 FILLCELL_X32 FILLER_312_920 ();
 FILLCELL_X32 FILLER_312_952 ();
 FILLCELL_X32 FILLER_312_984 ();
 FILLCELL_X32 FILLER_312_1016 ();
 FILLCELL_X32 FILLER_312_1048 ();
 FILLCELL_X32 FILLER_312_1080 ();
 FILLCELL_X32 FILLER_312_1112 ();
 FILLCELL_X32 FILLER_312_1144 ();
 FILLCELL_X32 FILLER_312_1176 ();
 FILLCELL_X32 FILLER_312_1208 ();
 FILLCELL_X32 FILLER_312_1240 ();
 FILLCELL_X32 FILLER_312_1272 ();
 FILLCELL_X32 FILLER_312_1304 ();
 FILLCELL_X32 FILLER_312_1336 ();
 FILLCELL_X32 FILLER_312_1368 ();
 FILLCELL_X32 FILLER_312_1400 ();
 FILLCELL_X32 FILLER_312_1432 ();
 FILLCELL_X32 FILLER_312_1464 ();
 FILLCELL_X32 FILLER_312_1496 ();
 FILLCELL_X32 FILLER_312_1528 ();
 FILLCELL_X32 FILLER_312_1560 ();
 FILLCELL_X32 FILLER_312_1592 ();
 FILLCELL_X32 FILLER_312_1624 ();
 FILLCELL_X32 FILLER_312_1656 ();
 FILLCELL_X32 FILLER_312_1688 ();
 FILLCELL_X32 FILLER_312_1720 ();
 FILLCELL_X32 FILLER_312_1752 ();
 FILLCELL_X32 FILLER_312_1784 ();
 FILLCELL_X32 FILLER_312_1816 ();
 FILLCELL_X32 FILLER_312_1848 ();
 FILLCELL_X8 FILLER_312_1880 ();
 FILLCELL_X4 FILLER_312_1888 ();
 FILLCELL_X2 FILLER_312_1892 ();
 FILLCELL_X32 FILLER_312_1895 ();
 FILLCELL_X32 FILLER_312_1927 ();
 FILLCELL_X32 FILLER_312_1959 ();
 FILLCELL_X32 FILLER_312_1991 ();
 FILLCELL_X32 FILLER_312_2023 ();
 FILLCELL_X32 FILLER_312_2055 ();
 FILLCELL_X32 FILLER_312_2087 ();
 FILLCELL_X32 FILLER_312_2119 ();
 FILLCELL_X32 FILLER_312_2151 ();
 FILLCELL_X32 FILLER_312_2183 ();
 FILLCELL_X32 FILLER_312_2215 ();
 FILLCELL_X32 FILLER_312_2247 ();
 FILLCELL_X32 FILLER_312_2279 ();
 FILLCELL_X32 FILLER_312_2311 ();
 FILLCELL_X32 FILLER_312_2343 ();
 FILLCELL_X32 FILLER_312_2375 ();
 FILLCELL_X32 FILLER_312_2407 ();
 FILLCELL_X32 FILLER_312_2439 ();
 FILLCELL_X32 FILLER_312_2471 ();
 FILLCELL_X32 FILLER_312_2503 ();
 FILLCELL_X32 FILLER_312_2535 ();
 FILLCELL_X32 FILLER_312_2567 ();
 FILLCELL_X32 FILLER_312_2599 ();
 FILLCELL_X32 FILLER_312_2631 ();
 FILLCELL_X32 FILLER_312_2663 ();
 FILLCELL_X32 FILLER_312_2695 ();
 FILLCELL_X32 FILLER_312_2727 ();
 FILLCELL_X32 FILLER_312_2759 ();
 FILLCELL_X32 FILLER_312_2791 ();
 FILLCELL_X32 FILLER_312_2823 ();
 FILLCELL_X32 FILLER_312_2855 ();
 FILLCELL_X32 FILLER_312_2887 ();
 FILLCELL_X32 FILLER_312_2919 ();
 FILLCELL_X32 FILLER_312_2951 ();
 FILLCELL_X32 FILLER_312_2983 ();
 FILLCELL_X32 FILLER_312_3015 ();
 FILLCELL_X32 FILLER_312_3047 ();
 FILLCELL_X32 FILLER_312_3079 ();
 FILLCELL_X32 FILLER_312_3111 ();
 FILLCELL_X8 FILLER_312_3143 ();
 FILLCELL_X4 FILLER_312_3151 ();
 FILLCELL_X2 FILLER_312_3155 ();
 FILLCELL_X32 FILLER_312_3158 ();
 FILLCELL_X32 FILLER_312_3190 ();
 FILLCELL_X32 FILLER_312_3222 ();
 FILLCELL_X32 FILLER_312_3254 ();
 FILLCELL_X32 FILLER_312_3286 ();
 FILLCELL_X32 FILLER_312_3318 ();
 FILLCELL_X32 FILLER_312_3350 ();
 FILLCELL_X32 FILLER_312_3382 ();
 FILLCELL_X32 FILLER_312_3414 ();
 FILLCELL_X32 FILLER_312_3446 ();
 FILLCELL_X32 FILLER_312_3478 ();
 FILLCELL_X32 FILLER_312_3510 ();
 FILLCELL_X32 FILLER_312_3542 ();
 FILLCELL_X32 FILLER_312_3574 ();
 FILLCELL_X32 FILLER_312_3606 ();
 FILLCELL_X32 FILLER_312_3638 ();
 FILLCELL_X32 FILLER_312_3670 ();
 FILLCELL_X32 FILLER_312_3702 ();
 FILLCELL_X4 FILLER_312_3734 ();
 FILLCELL_X32 FILLER_313_1 ();
 FILLCELL_X32 FILLER_313_33 ();
 FILLCELL_X32 FILLER_313_65 ();
 FILLCELL_X32 FILLER_313_97 ();
 FILLCELL_X32 FILLER_313_129 ();
 FILLCELL_X32 FILLER_313_161 ();
 FILLCELL_X32 FILLER_313_193 ();
 FILLCELL_X32 FILLER_313_225 ();
 FILLCELL_X32 FILLER_313_257 ();
 FILLCELL_X32 FILLER_313_289 ();
 FILLCELL_X32 FILLER_313_321 ();
 FILLCELL_X32 FILLER_313_353 ();
 FILLCELL_X32 FILLER_313_385 ();
 FILLCELL_X32 FILLER_313_417 ();
 FILLCELL_X32 FILLER_313_449 ();
 FILLCELL_X32 FILLER_313_481 ();
 FILLCELL_X32 FILLER_313_513 ();
 FILLCELL_X32 FILLER_313_545 ();
 FILLCELL_X32 FILLER_313_577 ();
 FILLCELL_X32 FILLER_313_609 ();
 FILLCELL_X32 FILLER_313_641 ();
 FILLCELL_X32 FILLER_313_673 ();
 FILLCELL_X32 FILLER_313_705 ();
 FILLCELL_X32 FILLER_313_737 ();
 FILLCELL_X32 FILLER_313_769 ();
 FILLCELL_X32 FILLER_313_801 ();
 FILLCELL_X32 FILLER_313_833 ();
 FILLCELL_X32 FILLER_313_865 ();
 FILLCELL_X32 FILLER_313_897 ();
 FILLCELL_X32 FILLER_313_929 ();
 FILLCELL_X32 FILLER_313_961 ();
 FILLCELL_X32 FILLER_313_993 ();
 FILLCELL_X32 FILLER_313_1025 ();
 FILLCELL_X32 FILLER_313_1057 ();
 FILLCELL_X32 FILLER_313_1089 ();
 FILLCELL_X32 FILLER_313_1121 ();
 FILLCELL_X32 FILLER_313_1153 ();
 FILLCELL_X32 FILLER_313_1185 ();
 FILLCELL_X32 FILLER_313_1217 ();
 FILLCELL_X8 FILLER_313_1249 ();
 FILLCELL_X4 FILLER_313_1257 ();
 FILLCELL_X2 FILLER_313_1261 ();
 FILLCELL_X32 FILLER_313_1264 ();
 FILLCELL_X32 FILLER_313_1296 ();
 FILLCELL_X32 FILLER_313_1328 ();
 FILLCELL_X32 FILLER_313_1360 ();
 FILLCELL_X32 FILLER_313_1392 ();
 FILLCELL_X32 FILLER_313_1424 ();
 FILLCELL_X32 FILLER_313_1456 ();
 FILLCELL_X32 FILLER_313_1488 ();
 FILLCELL_X32 FILLER_313_1520 ();
 FILLCELL_X32 FILLER_313_1552 ();
 FILLCELL_X32 FILLER_313_1584 ();
 FILLCELL_X32 FILLER_313_1616 ();
 FILLCELL_X32 FILLER_313_1648 ();
 FILLCELL_X32 FILLER_313_1680 ();
 FILLCELL_X32 FILLER_313_1712 ();
 FILLCELL_X32 FILLER_313_1744 ();
 FILLCELL_X32 FILLER_313_1776 ();
 FILLCELL_X32 FILLER_313_1808 ();
 FILLCELL_X32 FILLER_313_1840 ();
 FILLCELL_X32 FILLER_313_1872 ();
 FILLCELL_X32 FILLER_313_1904 ();
 FILLCELL_X32 FILLER_313_1936 ();
 FILLCELL_X32 FILLER_313_1968 ();
 FILLCELL_X32 FILLER_313_2000 ();
 FILLCELL_X32 FILLER_313_2032 ();
 FILLCELL_X32 FILLER_313_2064 ();
 FILLCELL_X32 FILLER_313_2096 ();
 FILLCELL_X32 FILLER_313_2128 ();
 FILLCELL_X32 FILLER_313_2160 ();
 FILLCELL_X32 FILLER_313_2192 ();
 FILLCELL_X32 FILLER_313_2224 ();
 FILLCELL_X32 FILLER_313_2256 ();
 FILLCELL_X32 FILLER_313_2288 ();
 FILLCELL_X32 FILLER_313_2320 ();
 FILLCELL_X32 FILLER_313_2352 ();
 FILLCELL_X32 FILLER_313_2384 ();
 FILLCELL_X32 FILLER_313_2416 ();
 FILLCELL_X32 FILLER_313_2448 ();
 FILLCELL_X32 FILLER_313_2480 ();
 FILLCELL_X8 FILLER_313_2512 ();
 FILLCELL_X4 FILLER_313_2520 ();
 FILLCELL_X2 FILLER_313_2524 ();
 FILLCELL_X32 FILLER_313_2527 ();
 FILLCELL_X32 FILLER_313_2559 ();
 FILLCELL_X32 FILLER_313_2591 ();
 FILLCELL_X32 FILLER_313_2623 ();
 FILLCELL_X32 FILLER_313_2655 ();
 FILLCELL_X32 FILLER_313_2687 ();
 FILLCELL_X32 FILLER_313_2719 ();
 FILLCELL_X32 FILLER_313_2751 ();
 FILLCELL_X32 FILLER_313_2783 ();
 FILLCELL_X32 FILLER_313_2815 ();
 FILLCELL_X32 FILLER_313_2847 ();
 FILLCELL_X32 FILLER_313_2879 ();
 FILLCELL_X32 FILLER_313_2911 ();
 FILLCELL_X32 FILLER_313_2943 ();
 FILLCELL_X32 FILLER_313_2975 ();
 FILLCELL_X32 FILLER_313_3007 ();
 FILLCELL_X32 FILLER_313_3039 ();
 FILLCELL_X32 FILLER_313_3071 ();
 FILLCELL_X32 FILLER_313_3103 ();
 FILLCELL_X32 FILLER_313_3135 ();
 FILLCELL_X32 FILLER_313_3167 ();
 FILLCELL_X32 FILLER_313_3199 ();
 FILLCELL_X32 FILLER_313_3231 ();
 FILLCELL_X32 FILLER_313_3263 ();
 FILLCELL_X32 FILLER_313_3295 ();
 FILLCELL_X32 FILLER_313_3327 ();
 FILLCELL_X32 FILLER_313_3359 ();
 FILLCELL_X32 FILLER_313_3391 ();
 FILLCELL_X32 FILLER_313_3423 ();
 FILLCELL_X32 FILLER_313_3455 ();
 FILLCELL_X32 FILLER_313_3487 ();
 FILLCELL_X32 FILLER_313_3519 ();
 FILLCELL_X32 FILLER_313_3551 ();
 FILLCELL_X32 FILLER_313_3583 ();
 FILLCELL_X32 FILLER_313_3615 ();
 FILLCELL_X32 FILLER_313_3647 ();
 FILLCELL_X32 FILLER_313_3679 ();
 FILLCELL_X16 FILLER_313_3711 ();
 FILLCELL_X8 FILLER_313_3727 ();
 FILLCELL_X2 FILLER_313_3735 ();
 FILLCELL_X1 FILLER_313_3737 ();
 FILLCELL_X32 FILLER_314_1 ();
 FILLCELL_X32 FILLER_314_33 ();
 FILLCELL_X32 FILLER_314_65 ();
 FILLCELL_X32 FILLER_314_97 ();
 FILLCELL_X32 FILLER_314_129 ();
 FILLCELL_X32 FILLER_314_161 ();
 FILLCELL_X32 FILLER_314_193 ();
 FILLCELL_X32 FILLER_314_225 ();
 FILLCELL_X32 FILLER_314_257 ();
 FILLCELL_X32 FILLER_314_289 ();
 FILLCELL_X32 FILLER_314_321 ();
 FILLCELL_X32 FILLER_314_353 ();
 FILLCELL_X32 FILLER_314_385 ();
 FILLCELL_X32 FILLER_314_417 ();
 FILLCELL_X32 FILLER_314_449 ();
 FILLCELL_X32 FILLER_314_481 ();
 FILLCELL_X32 FILLER_314_513 ();
 FILLCELL_X32 FILLER_314_545 ();
 FILLCELL_X32 FILLER_314_577 ();
 FILLCELL_X16 FILLER_314_609 ();
 FILLCELL_X4 FILLER_314_625 ();
 FILLCELL_X2 FILLER_314_629 ();
 FILLCELL_X32 FILLER_314_632 ();
 FILLCELL_X32 FILLER_314_664 ();
 FILLCELL_X32 FILLER_314_696 ();
 FILLCELL_X32 FILLER_314_728 ();
 FILLCELL_X32 FILLER_314_760 ();
 FILLCELL_X32 FILLER_314_792 ();
 FILLCELL_X32 FILLER_314_824 ();
 FILLCELL_X32 FILLER_314_856 ();
 FILLCELL_X32 FILLER_314_888 ();
 FILLCELL_X32 FILLER_314_920 ();
 FILLCELL_X32 FILLER_314_952 ();
 FILLCELL_X32 FILLER_314_984 ();
 FILLCELL_X32 FILLER_314_1016 ();
 FILLCELL_X32 FILLER_314_1048 ();
 FILLCELL_X32 FILLER_314_1080 ();
 FILLCELL_X32 FILLER_314_1112 ();
 FILLCELL_X32 FILLER_314_1144 ();
 FILLCELL_X32 FILLER_314_1176 ();
 FILLCELL_X32 FILLER_314_1208 ();
 FILLCELL_X32 FILLER_314_1240 ();
 FILLCELL_X32 FILLER_314_1272 ();
 FILLCELL_X32 FILLER_314_1304 ();
 FILLCELL_X32 FILLER_314_1336 ();
 FILLCELL_X32 FILLER_314_1368 ();
 FILLCELL_X32 FILLER_314_1400 ();
 FILLCELL_X32 FILLER_314_1432 ();
 FILLCELL_X32 FILLER_314_1464 ();
 FILLCELL_X32 FILLER_314_1496 ();
 FILLCELL_X32 FILLER_314_1528 ();
 FILLCELL_X32 FILLER_314_1560 ();
 FILLCELL_X32 FILLER_314_1592 ();
 FILLCELL_X32 FILLER_314_1624 ();
 FILLCELL_X32 FILLER_314_1656 ();
 FILLCELL_X32 FILLER_314_1688 ();
 FILLCELL_X32 FILLER_314_1720 ();
 FILLCELL_X32 FILLER_314_1752 ();
 FILLCELL_X32 FILLER_314_1784 ();
 FILLCELL_X32 FILLER_314_1816 ();
 FILLCELL_X32 FILLER_314_1848 ();
 FILLCELL_X8 FILLER_314_1880 ();
 FILLCELL_X4 FILLER_314_1888 ();
 FILLCELL_X2 FILLER_314_1892 ();
 FILLCELL_X32 FILLER_314_1895 ();
 FILLCELL_X32 FILLER_314_1927 ();
 FILLCELL_X32 FILLER_314_1959 ();
 FILLCELL_X32 FILLER_314_1991 ();
 FILLCELL_X32 FILLER_314_2023 ();
 FILLCELL_X32 FILLER_314_2055 ();
 FILLCELL_X32 FILLER_314_2087 ();
 FILLCELL_X32 FILLER_314_2119 ();
 FILLCELL_X32 FILLER_314_2151 ();
 FILLCELL_X32 FILLER_314_2183 ();
 FILLCELL_X32 FILLER_314_2215 ();
 FILLCELL_X32 FILLER_314_2247 ();
 FILLCELL_X32 FILLER_314_2279 ();
 FILLCELL_X32 FILLER_314_2311 ();
 FILLCELL_X32 FILLER_314_2343 ();
 FILLCELL_X32 FILLER_314_2375 ();
 FILLCELL_X32 FILLER_314_2407 ();
 FILLCELL_X32 FILLER_314_2439 ();
 FILLCELL_X32 FILLER_314_2471 ();
 FILLCELL_X32 FILLER_314_2503 ();
 FILLCELL_X32 FILLER_314_2535 ();
 FILLCELL_X32 FILLER_314_2567 ();
 FILLCELL_X32 FILLER_314_2599 ();
 FILLCELL_X32 FILLER_314_2631 ();
 FILLCELL_X32 FILLER_314_2663 ();
 FILLCELL_X32 FILLER_314_2695 ();
 FILLCELL_X32 FILLER_314_2727 ();
 FILLCELL_X32 FILLER_314_2759 ();
 FILLCELL_X32 FILLER_314_2791 ();
 FILLCELL_X32 FILLER_314_2823 ();
 FILLCELL_X32 FILLER_314_2855 ();
 FILLCELL_X32 FILLER_314_2887 ();
 FILLCELL_X32 FILLER_314_2919 ();
 FILLCELL_X32 FILLER_314_2951 ();
 FILLCELL_X32 FILLER_314_2983 ();
 FILLCELL_X32 FILLER_314_3015 ();
 FILLCELL_X32 FILLER_314_3047 ();
 FILLCELL_X32 FILLER_314_3079 ();
 FILLCELL_X32 FILLER_314_3111 ();
 FILLCELL_X8 FILLER_314_3143 ();
 FILLCELL_X4 FILLER_314_3151 ();
 FILLCELL_X2 FILLER_314_3155 ();
 FILLCELL_X32 FILLER_314_3158 ();
 FILLCELL_X32 FILLER_314_3190 ();
 FILLCELL_X32 FILLER_314_3222 ();
 FILLCELL_X32 FILLER_314_3254 ();
 FILLCELL_X32 FILLER_314_3286 ();
 FILLCELL_X32 FILLER_314_3318 ();
 FILLCELL_X32 FILLER_314_3350 ();
 FILLCELL_X32 FILLER_314_3382 ();
 FILLCELL_X32 FILLER_314_3414 ();
 FILLCELL_X32 FILLER_314_3446 ();
 FILLCELL_X32 FILLER_314_3478 ();
 FILLCELL_X32 FILLER_314_3510 ();
 FILLCELL_X32 FILLER_314_3542 ();
 FILLCELL_X32 FILLER_314_3574 ();
 FILLCELL_X32 FILLER_314_3606 ();
 FILLCELL_X32 FILLER_314_3638 ();
 FILLCELL_X32 FILLER_314_3670 ();
 FILLCELL_X32 FILLER_314_3702 ();
 FILLCELL_X4 FILLER_314_3734 ();
 FILLCELL_X32 FILLER_315_1 ();
 FILLCELL_X32 FILLER_315_33 ();
 FILLCELL_X32 FILLER_315_65 ();
 FILLCELL_X32 FILLER_315_97 ();
 FILLCELL_X32 FILLER_315_129 ();
 FILLCELL_X32 FILLER_315_161 ();
 FILLCELL_X32 FILLER_315_193 ();
 FILLCELL_X32 FILLER_315_225 ();
 FILLCELL_X32 FILLER_315_257 ();
 FILLCELL_X32 FILLER_315_289 ();
 FILLCELL_X32 FILLER_315_321 ();
 FILLCELL_X32 FILLER_315_353 ();
 FILLCELL_X32 FILLER_315_385 ();
 FILLCELL_X32 FILLER_315_417 ();
 FILLCELL_X32 FILLER_315_449 ();
 FILLCELL_X32 FILLER_315_481 ();
 FILLCELL_X32 FILLER_315_513 ();
 FILLCELL_X32 FILLER_315_545 ();
 FILLCELL_X32 FILLER_315_577 ();
 FILLCELL_X32 FILLER_315_609 ();
 FILLCELL_X32 FILLER_315_641 ();
 FILLCELL_X32 FILLER_315_673 ();
 FILLCELL_X32 FILLER_315_705 ();
 FILLCELL_X32 FILLER_315_737 ();
 FILLCELL_X32 FILLER_315_769 ();
 FILLCELL_X32 FILLER_315_801 ();
 FILLCELL_X32 FILLER_315_833 ();
 FILLCELL_X32 FILLER_315_865 ();
 FILLCELL_X32 FILLER_315_897 ();
 FILLCELL_X32 FILLER_315_929 ();
 FILLCELL_X32 FILLER_315_961 ();
 FILLCELL_X32 FILLER_315_993 ();
 FILLCELL_X32 FILLER_315_1025 ();
 FILLCELL_X32 FILLER_315_1057 ();
 FILLCELL_X32 FILLER_315_1089 ();
 FILLCELL_X32 FILLER_315_1121 ();
 FILLCELL_X32 FILLER_315_1153 ();
 FILLCELL_X32 FILLER_315_1185 ();
 FILLCELL_X32 FILLER_315_1217 ();
 FILLCELL_X8 FILLER_315_1249 ();
 FILLCELL_X4 FILLER_315_1257 ();
 FILLCELL_X2 FILLER_315_1261 ();
 FILLCELL_X32 FILLER_315_1264 ();
 FILLCELL_X32 FILLER_315_1296 ();
 FILLCELL_X32 FILLER_315_1328 ();
 FILLCELL_X32 FILLER_315_1360 ();
 FILLCELL_X32 FILLER_315_1392 ();
 FILLCELL_X32 FILLER_315_1424 ();
 FILLCELL_X32 FILLER_315_1456 ();
 FILLCELL_X32 FILLER_315_1488 ();
 FILLCELL_X32 FILLER_315_1520 ();
 FILLCELL_X32 FILLER_315_1552 ();
 FILLCELL_X32 FILLER_315_1584 ();
 FILLCELL_X32 FILLER_315_1616 ();
 FILLCELL_X32 FILLER_315_1648 ();
 FILLCELL_X32 FILLER_315_1680 ();
 FILLCELL_X32 FILLER_315_1712 ();
 FILLCELL_X32 FILLER_315_1744 ();
 FILLCELL_X32 FILLER_315_1776 ();
 FILLCELL_X32 FILLER_315_1808 ();
 FILLCELL_X32 FILLER_315_1840 ();
 FILLCELL_X32 FILLER_315_1872 ();
 FILLCELL_X32 FILLER_315_1904 ();
 FILLCELL_X32 FILLER_315_1936 ();
 FILLCELL_X32 FILLER_315_1968 ();
 FILLCELL_X32 FILLER_315_2000 ();
 FILLCELL_X32 FILLER_315_2032 ();
 FILLCELL_X32 FILLER_315_2064 ();
 FILLCELL_X32 FILLER_315_2096 ();
 FILLCELL_X32 FILLER_315_2128 ();
 FILLCELL_X32 FILLER_315_2160 ();
 FILLCELL_X32 FILLER_315_2192 ();
 FILLCELL_X32 FILLER_315_2224 ();
 FILLCELL_X32 FILLER_315_2256 ();
 FILLCELL_X32 FILLER_315_2288 ();
 FILLCELL_X32 FILLER_315_2320 ();
 FILLCELL_X32 FILLER_315_2352 ();
 FILLCELL_X32 FILLER_315_2384 ();
 FILLCELL_X32 FILLER_315_2416 ();
 FILLCELL_X32 FILLER_315_2448 ();
 FILLCELL_X32 FILLER_315_2480 ();
 FILLCELL_X8 FILLER_315_2512 ();
 FILLCELL_X4 FILLER_315_2520 ();
 FILLCELL_X2 FILLER_315_2524 ();
 FILLCELL_X32 FILLER_315_2527 ();
 FILLCELL_X32 FILLER_315_2559 ();
 FILLCELL_X32 FILLER_315_2591 ();
 FILLCELL_X32 FILLER_315_2623 ();
 FILLCELL_X32 FILLER_315_2655 ();
 FILLCELL_X32 FILLER_315_2687 ();
 FILLCELL_X32 FILLER_315_2719 ();
 FILLCELL_X32 FILLER_315_2751 ();
 FILLCELL_X32 FILLER_315_2783 ();
 FILLCELL_X32 FILLER_315_2815 ();
 FILLCELL_X32 FILLER_315_2847 ();
 FILLCELL_X32 FILLER_315_2879 ();
 FILLCELL_X32 FILLER_315_2911 ();
 FILLCELL_X32 FILLER_315_2943 ();
 FILLCELL_X32 FILLER_315_2975 ();
 FILLCELL_X32 FILLER_315_3007 ();
 FILLCELL_X32 FILLER_315_3039 ();
 FILLCELL_X32 FILLER_315_3071 ();
 FILLCELL_X32 FILLER_315_3103 ();
 FILLCELL_X32 FILLER_315_3135 ();
 FILLCELL_X32 FILLER_315_3167 ();
 FILLCELL_X32 FILLER_315_3199 ();
 FILLCELL_X32 FILLER_315_3231 ();
 FILLCELL_X32 FILLER_315_3263 ();
 FILLCELL_X32 FILLER_315_3295 ();
 FILLCELL_X32 FILLER_315_3327 ();
 FILLCELL_X32 FILLER_315_3359 ();
 FILLCELL_X32 FILLER_315_3391 ();
 FILLCELL_X32 FILLER_315_3423 ();
 FILLCELL_X32 FILLER_315_3455 ();
 FILLCELL_X32 FILLER_315_3487 ();
 FILLCELL_X32 FILLER_315_3519 ();
 FILLCELL_X32 FILLER_315_3551 ();
 FILLCELL_X32 FILLER_315_3583 ();
 FILLCELL_X32 FILLER_315_3615 ();
 FILLCELL_X32 FILLER_315_3647 ();
 FILLCELL_X32 FILLER_315_3679 ();
 FILLCELL_X16 FILLER_315_3711 ();
 FILLCELL_X8 FILLER_315_3727 ();
 FILLCELL_X2 FILLER_315_3735 ();
 FILLCELL_X1 FILLER_315_3737 ();
 FILLCELL_X32 FILLER_316_1 ();
 FILLCELL_X32 FILLER_316_33 ();
 FILLCELL_X32 FILLER_316_65 ();
 FILLCELL_X32 FILLER_316_97 ();
 FILLCELL_X32 FILLER_316_129 ();
 FILLCELL_X32 FILLER_316_161 ();
 FILLCELL_X32 FILLER_316_193 ();
 FILLCELL_X32 FILLER_316_225 ();
 FILLCELL_X32 FILLER_316_257 ();
 FILLCELL_X32 FILLER_316_289 ();
 FILLCELL_X32 FILLER_316_321 ();
 FILLCELL_X32 FILLER_316_353 ();
 FILLCELL_X32 FILLER_316_385 ();
 FILLCELL_X32 FILLER_316_417 ();
 FILLCELL_X32 FILLER_316_449 ();
 FILLCELL_X32 FILLER_316_481 ();
 FILLCELL_X32 FILLER_316_513 ();
 FILLCELL_X32 FILLER_316_545 ();
 FILLCELL_X32 FILLER_316_577 ();
 FILLCELL_X16 FILLER_316_609 ();
 FILLCELL_X4 FILLER_316_625 ();
 FILLCELL_X2 FILLER_316_629 ();
 FILLCELL_X32 FILLER_316_632 ();
 FILLCELL_X32 FILLER_316_664 ();
 FILLCELL_X32 FILLER_316_696 ();
 FILLCELL_X32 FILLER_316_728 ();
 FILLCELL_X32 FILLER_316_760 ();
 FILLCELL_X32 FILLER_316_792 ();
 FILLCELL_X32 FILLER_316_824 ();
 FILLCELL_X32 FILLER_316_856 ();
 FILLCELL_X32 FILLER_316_888 ();
 FILLCELL_X32 FILLER_316_920 ();
 FILLCELL_X32 FILLER_316_952 ();
 FILLCELL_X32 FILLER_316_984 ();
 FILLCELL_X32 FILLER_316_1016 ();
 FILLCELL_X32 FILLER_316_1048 ();
 FILLCELL_X32 FILLER_316_1080 ();
 FILLCELL_X32 FILLER_316_1112 ();
 FILLCELL_X32 FILLER_316_1144 ();
 FILLCELL_X32 FILLER_316_1176 ();
 FILLCELL_X32 FILLER_316_1208 ();
 FILLCELL_X32 FILLER_316_1240 ();
 FILLCELL_X32 FILLER_316_1272 ();
 FILLCELL_X32 FILLER_316_1304 ();
 FILLCELL_X32 FILLER_316_1336 ();
 FILLCELL_X32 FILLER_316_1368 ();
 FILLCELL_X32 FILLER_316_1400 ();
 FILLCELL_X32 FILLER_316_1432 ();
 FILLCELL_X32 FILLER_316_1464 ();
 FILLCELL_X32 FILLER_316_1496 ();
 FILLCELL_X32 FILLER_316_1528 ();
 FILLCELL_X32 FILLER_316_1560 ();
 FILLCELL_X32 FILLER_316_1592 ();
 FILLCELL_X32 FILLER_316_1624 ();
 FILLCELL_X32 FILLER_316_1656 ();
 FILLCELL_X32 FILLER_316_1688 ();
 FILLCELL_X32 FILLER_316_1720 ();
 FILLCELL_X32 FILLER_316_1752 ();
 FILLCELL_X32 FILLER_316_1784 ();
 FILLCELL_X32 FILLER_316_1816 ();
 FILLCELL_X32 FILLER_316_1848 ();
 FILLCELL_X8 FILLER_316_1880 ();
 FILLCELL_X4 FILLER_316_1888 ();
 FILLCELL_X2 FILLER_316_1892 ();
 FILLCELL_X32 FILLER_316_1895 ();
 FILLCELL_X32 FILLER_316_1927 ();
 FILLCELL_X32 FILLER_316_1959 ();
 FILLCELL_X32 FILLER_316_1991 ();
 FILLCELL_X32 FILLER_316_2023 ();
 FILLCELL_X32 FILLER_316_2055 ();
 FILLCELL_X32 FILLER_316_2087 ();
 FILLCELL_X32 FILLER_316_2119 ();
 FILLCELL_X32 FILLER_316_2151 ();
 FILLCELL_X32 FILLER_316_2183 ();
 FILLCELL_X32 FILLER_316_2215 ();
 FILLCELL_X32 FILLER_316_2247 ();
 FILLCELL_X32 FILLER_316_2279 ();
 FILLCELL_X32 FILLER_316_2311 ();
 FILLCELL_X32 FILLER_316_2343 ();
 FILLCELL_X32 FILLER_316_2375 ();
 FILLCELL_X32 FILLER_316_2407 ();
 FILLCELL_X32 FILLER_316_2439 ();
 FILLCELL_X32 FILLER_316_2471 ();
 FILLCELL_X32 FILLER_316_2503 ();
 FILLCELL_X32 FILLER_316_2535 ();
 FILLCELL_X32 FILLER_316_2567 ();
 FILLCELL_X32 FILLER_316_2599 ();
 FILLCELL_X32 FILLER_316_2631 ();
 FILLCELL_X32 FILLER_316_2663 ();
 FILLCELL_X32 FILLER_316_2695 ();
 FILLCELL_X32 FILLER_316_2727 ();
 FILLCELL_X32 FILLER_316_2759 ();
 FILLCELL_X32 FILLER_316_2791 ();
 FILLCELL_X32 FILLER_316_2823 ();
 FILLCELL_X32 FILLER_316_2855 ();
 FILLCELL_X32 FILLER_316_2887 ();
 FILLCELL_X32 FILLER_316_2919 ();
 FILLCELL_X32 FILLER_316_2951 ();
 FILLCELL_X32 FILLER_316_2983 ();
 FILLCELL_X32 FILLER_316_3015 ();
 FILLCELL_X32 FILLER_316_3047 ();
 FILLCELL_X32 FILLER_316_3079 ();
 FILLCELL_X32 FILLER_316_3111 ();
 FILLCELL_X8 FILLER_316_3143 ();
 FILLCELL_X4 FILLER_316_3151 ();
 FILLCELL_X2 FILLER_316_3155 ();
 FILLCELL_X32 FILLER_316_3158 ();
 FILLCELL_X32 FILLER_316_3190 ();
 FILLCELL_X32 FILLER_316_3222 ();
 FILLCELL_X32 FILLER_316_3254 ();
 FILLCELL_X32 FILLER_316_3286 ();
 FILLCELL_X32 FILLER_316_3318 ();
 FILLCELL_X32 FILLER_316_3350 ();
 FILLCELL_X32 FILLER_316_3382 ();
 FILLCELL_X32 FILLER_316_3414 ();
 FILLCELL_X32 FILLER_316_3446 ();
 FILLCELL_X32 FILLER_316_3478 ();
 FILLCELL_X32 FILLER_316_3510 ();
 FILLCELL_X32 FILLER_316_3542 ();
 FILLCELL_X32 FILLER_316_3574 ();
 FILLCELL_X32 FILLER_316_3606 ();
 FILLCELL_X32 FILLER_316_3638 ();
 FILLCELL_X32 FILLER_316_3670 ();
 FILLCELL_X32 FILLER_316_3702 ();
 FILLCELL_X4 FILLER_316_3734 ();
 FILLCELL_X32 FILLER_317_1 ();
 FILLCELL_X32 FILLER_317_33 ();
 FILLCELL_X32 FILLER_317_65 ();
 FILLCELL_X32 FILLER_317_97 ();
 FILLCELL_X32 FILLER_317_129 ();
 FILLCELL_X32 FILLER_317_161 ();
 FILLCELL_X32 FILLER_317_193 ();
 FILLCELL_X32 FILLER_317_225 ();
 FILLCELL_X32 FILLER_317_257 ();
 FILLCELL_X32 FILLER_317_289 ();
 FILLCELL_X32 FILLER_317_321 ();
 FILLCELL_X32 FILLER_317_353 ();
 FILLCELL_X32 FILLER_317_385 ();
 FILLCELL_X32 FILLER_317_417 ();
 FILLCELL_X32 FILLER_317_449 ();
 FILLCELL_X32 FILLER_317_481 ();
 FILLCELL_X32 FILLER_317_513 ();
 FILLCELL_X32 FILLER_317_545 ();
 FILLCELL_X32 FILLER_317_577 ();
 FILLCELL_X32 FILLER_317_609 ();
 FILLCELL_X32 FILLER_317_641 ();
 FILLCELL_X32 FILLER_317_673 ();
 FILLCELL_X32 FILLER_317_705 ();
 FILLCELL_X32 FILLER_317_737 ();
 FILLCELL_X32 FILLER_317_769 ();
 FILLCELL_X32 FILLER_317_801 ();
 FILLCELL_X32 FILLER_317_833 ();
 FILLCELL_X32 FILLER_317_865 ();
 FILLCELL_X32 FILLER_317_897 ();
 FILLCELL_X32 FILLER_317_929 ();
 FILLCELL_X32 FILLER_317_961 ();
 FILLCELL_X32 FILLER_317_993 ();
 FILLCELL_X32 FILLER_317_1025 ();
 FILLCELL_X32 FILLER_317_1057 ();
 FILLCELL_X32 FILLER_317_1089 ();
 FILLCELL_X32 FILLER_317_1121 ();
 FILLCELL_X32 FILLER_317_1153 ();
 FILLCELL_X32 FILLER_317_1185 ();
 FILLCELL_X32 FILLER_317_1217 ();
 FILLCELL_X8 FILLER_317_1249 ();
 FILLCELL_X4 FILLER_317_1257 ();
 FILLCELL_X2 FILLER_317_1261 ();
 FILLCELL_X32 FILLER_317_1264 ();
 FILLCELL_X32 FILLER_317_1296 ();
 FILLCELL_X32 FILLER_317_1328 ();
 FILLCELL_X32 FILLER_317_1360 ();
 FILLCELL_X32 FILLER_317_1392 ();
 FILLCELL_X32 FILLER_317_1424 ();
 FILLCELL_X32 FILLER_317_1456 ();
 FILLCELL_X32 FILLER_317_1488 ();
 FILLCELL_X32 FILLER_317_1520 ();
 FILLCELL_X32 FILLER_317_1552 ();
 FILLCELL_X32 FILLER_317_1584 ();
 FILLCELL_X32 FILLER_317_1616 ();
 FILLCELL_X32 FILLER_317_1648 ();
 FILLCELL_X32 FILLER_317_1680 ();
 FILLCELL_X32 FILLER_317_1712 ();
 FILLCELL_X32 FILLER_317_1744 ();
 FILLCELL_X32 FILLER_317_1776 ();
 FILLCELL_X32 FILLER_317_1808 ();
 FILLCELL_X32 FILLER_317_1840 ();
 FILLCELL_X32 FILLER_317_1872 ();
 FILLCELL_X32 FILLER_317_1904 ();
 FILLCELL_X32 FILLER_317_1936 ();
 FILLCELL_X32 FILLER_317_1968 ();
 FILLCELL_X32 FILLER_317_2000 ();
 FILLCELL_X32 FILLER_317_2032 ();
 FILLCELL_X32 FILLER_317_2064 ();
 FILLCELL_X32 FILLER_317_2096 ();
 FILLCELL_X32 FILLER_317_2128 ();
 FILLCELL_X32 FILLER_317_2160 ();
 FILLCELL_X32 FILLER_317_2192 ();
 FILLCELL_X32 FILLER_317_2224 ();
 FILLCELL_X32 FILLER_317_2256 ();
 FILLCELL_X32 FILLER_317_2288 ();
 FILLCELL_X32 FILLER_317_2320 ();
 FILLCELL_X32 FILLER_317_2352 ();
 FILLCELL_X32 FILLER_317_2384 ();
 FILLCELL_X32 FILLER_317_2416 ();
 FILLCELL_X32 FILLER_317_2448 ();
 FILLCELL_X32 FILLER_317_2480 ();
 FILLCELL_X8 FILLER_317_2512 ();
 FILLCELL_X4 FILLER_317_2520 ();
 FILLCELL_X2 FILLER_317_2524 ();
 FILLCELL_X32 FILLER_317_2527 ();
 FILLCELL_X32 FILLER_317_2559 ();
 FILLCELL_X32 FILLER_317_2591 ();
 FILLCELL_X32 FILLER_317_2623 ();
 FILLCELL_X32 FILLER_317_2655 ();
 FILLCELL_X32 FILLER_317_2687 ();
 FILLCELL_X32 FILLER_317_2719 ();
 FILLCELL_X32 FILLER_317_2751 ();
 FILLCELL_X32 FILLER_317_2783 ();
 FILLCELL_X32 FILLER_317_2815 ();
 FILLCELL_X32 FILLER_317_2847 ();
 FILLCELL_X32 FILLER_317_2879 ();
 FILLCELL_X32 FILLER_317_2911 ();
 FILLCELL_X32 FILLER_317_2943 ();
 FILLCELL_X32 FILLER_317_2975 ();
 FILLCELL_X32 FILLER_317_3007 ();
 FILLCELL_X32 FILLER_317_3039 ();
 FILLCELL_X32 FILLER_317_3071 ();
 FILLCELL_X32 FILLER_317_3103 ();
 FILLCELL_X32 FILLER_317_3135 ();
 FILLCELL_X32 FILLER_317_3167 ();
 FILLCELL_X32 FILLER_317_3199 ();
 FILLCELL_X32 FILLER_317_3231 ();
 FILLCELL_X32 FILLER_317_3263 ();
 FILLCELL_X32 FILLER_317_3295 ();
 FILLCELL_X32 FILLER_317_3327 ();
 FILLCELL_X32 FILLER_317_3359 ();
 FILLCELL_X32 FILLER_317_3391 ();
 FILLCELL_X32 FILLER_317_3423 ();
 FILLCELL_X32 FILLER_317_3455 ();
 FILLCELL_X32 FILLER_317_3487 ();
 FILLCELL_X32 FILLER_317_3519 ();
 FILLCELL_X32 FILLER_317_3551 ();
 FILLCELL_X32 FILLER_317_3583 ();
 FILLCELL_X32 FILLER_317_3615 ();
 FILLCELL_X32 FILLER_317_3647 ();
 FILLCELL_X32 FILLER_317_3679 ();
 FILLCELL_X16 FILLER_317_3711 ();
 FILLCELL_X8 FILLER_317_3727 ();
 FILLCELL_X2 FILLER_317_3735 ();
 FILLCELL_X1 FILLER_317_3737 ();
 FILLCELL_X32 FILLER_318_1 ();
 FILLCELL_X32 FILLER_318_33 ();
 FILLCELL_X32 FILLER_318_65 ();
 FILLCELL_X32 FILLER_318_97 ();
 FILLCELL_X32 FILLER_318_129 ();
 FILLCELL_X32 FILLER_318_161 ();
 FILLCELL_X32 FILLER_318_193 ();
 FILLCELL_X32 FILLER_318_225 ();
 FILLCELL_X32 FILLER_318_257 ();
 FILLCELL_X32 FILLER_318_289 ();
 FILLCELL_X32 FILLER_318_321 ();
 FILLCELL_X32 FILLER_318_353 ();
 FILLCELL_X32 FILLER_318_385 ();
 FILLCELL_X32 FILLER_318_417 ();
 FILLCELL_X32 FILLER_318_449 ();
 FILLCELL_X32 FILLER_318_481 ();
 FILLCELL_X32 FILLER_318_513 ();
 FILLCELL_X32 FILLER_318_545 ();
 FILLCELL_X32 FILLER_318_577 ();
 FILLCELL_X16 FILLER_318_609 ();
 FILLCELL_X4 FILLER_318_625 ();
 FILLCELL_X2 FILLER_318_629 ();
 FILLCELL_X32 FILLER_318_632 ();
 FILLCELL_X32 FILLER_318_664 ();
 FILLCELL_X32 FILLER_318_696 ();
 FILLCELL_X32 FILLER_318_728 ();
 FILLCELL_X32 FILLER_318_760 ();
 FILLCELL_X32 FILLER_318_792 ();
 FILLCELL_X32 FILLER_318_824 ();
 FILLCELL_X32 FILLER_318_856 ();
 FILLCELL_X32 FILLER_318_888 ();
 FILLCELL_X32 FILLER_318_920 ();
 FILLCELL_X32 FILLER_318_952 ();
 FILLCELL_X32 FILLER_318_984 ();
 FILLCELL_X32 FILLER_318_1016 ();
 FILLCELL_X32 FILLER_318_1048 ();
 FILLCELL_X32 FILLER_318_1080 ();
 FILLCELL_X32 FILLER_318_1112 ();
 FILLCELL_X32 FILLER_318_1144 ();
 FILLCELL_X32 FILLER_318_1176 ();
 FILLCELL_X32 FILLER_318_1208 ();
 FILLCELL_X32 FILLER_318_1240 ();
 FILLCELL_X32 FILLER_318_1272 ();
 FILLCELL_X32 FILLER_318_1304 ();
 FILLCELL_X32 FILLER_318_1336 ();
 FILLCELL_X32 FILLER_318_1368 ();
 FILLCELL_X32 FILLER_318_1400 ();
 FILLCELL_X32 FILLER_318_1432 ();
 FILLCELL_X32 FILLER_318_1464 ();
 FILLCELL_X32 FILLER_318_1496 ();
 FILLCELL_X32 FILLER_318_1528 ();
 FILLCELL_X32 FILLER_318_1560 ();
 FILLCELL_X32 FILLER_318_1592 ();
 FILLCELL_X32 FILLER_318_1624 ();
 FILLCELL_X32 FILLER_318_1656 ();
 FILLCELL_X32 FILLER_318_1688 ();
 FILLCELL_X32 FILLER_318_1720 ();
 FILLCELL_X32 FILLER_318_1752 ();
 FILLCELL_X32 FILLER_318_1784 ();
 FILLCELL_X32 FILLER_318_1816 ();
 FILLCELL_X32 FILLER_318_1848 ();
 FILLCELL_X8 FILLER_318_1880 ();
 FILLCELL_X4 FILLER_318_1888 ();
 FILLCELL_X2 FILLER_318_1892 ();
 FILLCELL_X32 FILLER_318_1895 ();
 FILLCELL_X32 FILLER_318_1927 ();
 FILLCELL_X32 FILLER_318_1959 ();
 FILLCELL_X32 FILLER_318_1991 ();
 FILLCELL_X32 FILLER_318_2023 ();
 FILLCELL_X32 FILLER_318_2055 ();
 FILLCELL_X32 FILLER_318_2087 ();
 FILLCELL_X32 FILLER_318_2119 ();
 FILLCELL_X32 FILLER_318_2151 ();
 FILLCELL_X32 FILLER_318_2183 ();
 FILLCELL_X32 FILLER_318_2215 ();
 FILLCELL_X32 FILLER_318_2247 ();
 FILLCELL_X32 FILLER_318_2279 ();
 FILLCELL_X32 FILLER_318_2311 ();
 FILLCELL_X32 FILLER_318_2343 ();
 FILLCELL_X32 FILLER_318_2375 ();
 FILLCELL_X32 FILLER_318_2407 ();
 FILLCELL_X32 FILLER_318_2439 ();
 FILLCELL_X32 FILLER_318_2471 ();
 FILLCELL_X32 FILLER_318_2503 ();
 FILLCELL_X32 FILLER_318_2535 ();
 FILLCELL_X32 FILLER_318_2567 ();
 FILLCELL_X32 FILLER_318_2599 ();
 FILLCELL_X32 FILLER_318_2631 ();
 FILLCELL_X32 FILLER_318_2663 ();
 FILLCELL_X32 FILLER_318_2695 ();
 FILLCELL_X32 FILLER_318_2727 ();
 FILLCELL_X32 FILLER_318_2759 ();
 FILLCELL_X32 FILLER_318_2791 ();
 FILLCELL_X32 FILLER_318_2823 ();
 FILLCELL_X32 FILLER_318_2855 ();
 FILLCELL_X32 FILLER_318_2887 ();
 FILLCELL_X32 FILLER_318_2919 ();
 FILLCELL_X32 FILLER_318_2951 ();
 FILLCELL_X32 FILLER_318_2983 ();
 FILLCELL_X32 FILLER_318_3015 ();
 FILLCELL_X32 FILLER_318_3047 ();
 FILLCELL_X32 FILLER_318_3079 ();
 FILLCELL_X32 FILLER_318_3111 ();
 FILLCELL_X8 FILLER_318_3143 ();
 FILLCELL_X4 FILLER_318_3151 ();
 FILLCELL_X2 FILLER_318_3155 ();
 FILLCELL_X32 FILLER_318_3158 ();
 FILLCELL_X32 FILLER_318_3190 ();
 FILLCELL_X32 FILLER_318_3222 ();
 FILLCELL_X32 FILLER_318_3254 ();
 FILLCELL_X32 FILLER_318_3286 ();
 FILLCELL_X32 FILLER_318_3318 ();
 FILLCELL_X32 FILLER_318_3350 ();
 FILLCELL_X32 FILLER_318_3382 ();
 FILLCELL_X32 FILLER_318_3414 ();
 FILLCELL_X32 FILLER_318_3446 ();
 FILLCELL_X32 FILLER_318_3478 ();
 FILLCELL_X32 FILLER_318_3510 ();
 FILLCELL_X32 FILLER_318_3542 ();
 FILLCELL_X32 FILLER_318_3574 ();
 FILLCELL_X32 FILLER_318_3606 ();
 FILLCELL_X32 FILLER_318_3638 ();
 FILLCELL_X32 FILLER_318_3670 ();
 FILLCELL_X32 FILLER_318_3702 ();
 FILLCELL_X4 FILLER_318_3734 ();
 FILLCELL_X32 FILLER_319_1 ();
 FILLCELL_X32 FILLER_319_33 ();
 FILLCELL_X32 FILLER_319_65 ();
 FILLCELL_X32 FILLER_319_97 ();
 FILLCELL_X32 FILLER_319_129 ();
 FILLCELL_X32 FILLER_319_161 ();
 FILLCELL_X32 FILLER_319_193 ();
 FILLCELL_X32 FILLER_319_225 ();
 FILLCELL_X32 FILLER_319_257 ();
 FILLCELL_X32 FILLER_319_289 ();
 FILLCELL_X32 FILLER_319_321 ();
 FILLCELL_X32 FILLER_319_353 ();
 FILLCELL_X32 FILLER_319_385 ();
 FILLCELL_X32 FILLER_319_417 ();
 FILLCELL_X32 FILLER_319_449 ();
 FILLCELL_X32 FILLER_319_481 ();
 FILLCELL_X32 FILLER_319_513 ();
 FILLCELL_X32 FILLER_319_545 ();
 FILLCELL_X32 FILLER_319_577 ();
 FILLCELL_X32 FILLER_319_609 ();
 FILLCELL_X32 FILLER_319_641 ();
 FILLCELL_X32 FILLER_319_673 ();
 FILLCELL_X32 FILLER_319_705 ();
 FILLCELL_X32 FILLER_319_737 ();
 FILLCELL_X32 FILLER_319_769 ();
 FILLCELL_X32 FILLER_319_801 ();
 FILLCELL_X32 FILLER_319_833 ();
 FILLCELL_X32 FILLER_319_865 ();
 FILLCELL_X32 FILLER_319_897 ();
 FILLCELL_X32 FILLER_319_929 ();
 FILLCELL_X32 FILLER_319_961 ();
 FILLCELL_X32 FILLER_319_993 ();
 FILLCELL_X32 FILLER_319_1025 ();
 FILLCELL_X32 FILLER_319_1057 ();
 FILLCELL_X32 FILLER_319_1089 ();
 FILLCELL_X32 FILLER_319_1121 ();
 FILLCELL_X32 FILLER_319_1153 ();
 FILLCELL_X32 FILLER_319_1185 ();
 FILLCELL_X32 FILLER_319_1217 ();
 FILLCELL_X8 FILLER_319_1249 ();
 FILLCELL_X4 FILLER_319_1257 ();
 FILLCELL_X2 FILLER_319_1261 ();
 FILLCELL_X32 FILLER_319_1264 ();
 FILLCELL_X32 FILLER_319_1296 ();
 FILLCELL_X32 FILLER_319_1328 ();
 FILLCELL_X32 FILLER_319_1360 ();
 FILLCELL_X32 FILLER_319_1392 ();
 FILLCELL_X32 FILLER_319_1424 ();
 FILLCELL_X32 FILLER_319_1456 ();
 FILLCELL_X32 FILLER_319_1488 ();
 FILLCELL_X32 FILLER_319_1520 ();
 FILLCELL_X32 FILLER_319_1552 ();
 FILLCELL_X32 FILLER_319_1584 ();
 FILLCELL_X32 FILLER_319_1616 ();
 FILLCELL_X32 FILLER_319_1648 ();
 FILLCELL_X32 FILLER_319_1680 ();
 FILLCELL_X32 FILLER_319_1712 ();
 FILLCELL_X32 FILLER_319_1744 ();
 FILLCELL_X32 FILLER_319_1776 ();
 FILLCELL_X32 FILLER_319_1808 ();
 FILLCELL_X32 FILLER_319_1840 ();
 FILLCELL_X32 FILLER_319_1872 ();
 FILLCELL_X32 FILLER_319_1904 ();
 FILLCELL_X32 FILLER_319_1936 ();
 FILLCELL_X32 FILLER_319_1968 ();
 FILLCELL_X32 FILLER_319_2000 ();
 FILLCELL_X32 FILLER_319_2032 ();
 FILLCELL_X32 FILLER_319_2064 ();
 FILLCELL_X32 FILLER_319_2096 ();
 FILLCELL_X32 FILLER_319_2128 ();
 FILLCELL_X32 FILLER_319_2160 ();
 FILLCELL_X32 FILLER_319_2192 ();
 FILLCELL_X32 FILLER_319_2224 ();
 FILLCELL_X32 FILLER_319_2256 ();
 FILLCELL_X32 FILLER_319_2288 ();
 FILLCELL_X32 FILLER_319_2320 ();
 FILLCELL_X32 FILLER_319_2352 ();
 FILLCELL_X32 FILLER_319_2384 ();
 FILLCELL_X32 FILLER_319_2416 ();
 FILLCELL_X32 FILLER_319_2448 ();
 FILLCELL_X32 FILLER_319_2480 ();
 FILLCELL_X8 FILLER_319_2512 ();
 FILLCELL_X4 FILLER_319_2520 ();
 FILLCELL_X2 FILLER_319_2524 ();
 FILLCELL_X32 FILLER_319_2527 ();
 FILLCELL_X32 FILLER_319_2559 ();
 FILLCELL_X32 FILLER_319_2591 ();
 FILLCELL_X32 FILLER_319_2623 ();
 FILLCELL_X32 FILLER_319_2655 ();
 FILLCELL_X32 FILLER_319_2687 ();
 FILLCELL_X32 FILLER_319_2719 ();
 FILLCELL_X32 FILLER_319_2751 ();
 FILLCELL_X32 FILLER_319_2783 ();
 FILLCELL_X32 FILLER_319_2815 ();
 FILLCELL_X32 FILLER_319_2847 ();
 FILLCELL_X32 FILLER_319_2879 ();
 FILLCELL_X32 FILLER_319_2911 ();
 FILLCELL_X32 FILLER_319_2943 ();
 FILLCELL_X32 FILLER_319_2975 ();
 FILLCELL_X32 FILLER_319_3007 ();
 FILLCELL_X32 FILLER_319_3039 ();
 FILLCELL_X32 FILLER_319_3071 ();
 FILLCELL_X32 FILLER_319_3103 ();
 FILLCELL_X32 FILLER_319_3135 ();
 FILLCELL_X32 FILLER_319_3167 ();
 FILLCELL_X32 FILLER_319_3199 ();
 FILLCELL_X32 FILLER_319_3231 ();
 FILLCELL_X32 FILLER_319_3263 ();
 FILLCELL_X32 FILLER_319_3295 ();
 FILLCELL_X32 FILLER_319_3327 ();
 FILLCELL_X32 FILLER_319_3359 ();
 FILLCELL_X32 FILLER_319_3391 ();
 FILLCELL_X32 FILLER_319_3423 ();
 FILLCELL_X32 FILLER_319_3455 ();
 FILLCELL_X32 FILLER_319_3487 ();
 FILLCELL_X32 FILLER_319_3519 ();
 FILLCELL_X32 FILLER_319_3551 ();
 FILLCELL_X32 FILLER_319_3583 ();
 FILLCELL_X32 FILLER_319_3615 ();
 FILLCELL_X32 FILLER_319_3647 ();
 FILLCELL_X32 FILLER_319_3679 ();
 FILLCELL_X16 FILLER_319_3711 ();
 FILLCELL_X8 FILLER_319_3727 ();
 FILLCELL_X2 FILLER_319_3735 ();
 FILLCELL_X1 FILLER_319_3737 ();
 FILLCELL_X32 FILLER_320_1 ();
 FILLCELL_X32 FILLER_320_33 ();
 FILLCELL_X32 FILLER_320_65 ();
 FILLCELL_X32 FILLER_320_97 ();
 FILLCELL_X32 FILLER_320_129 ();
 FILLCELL_X32 FILLER_320_161 ();
 FILLCELL_X32 FILLER_320_193 ();
 FILLCELL_X32 FILLER_320_225 ();
 FILLCELL_X32 FILLER_320_257 ();
 FILLCELL_X32 FILLER_320_289 ();
 FILLCELL_X32 FILLER_320_321 ();
 FILLCELL_X32 FILLER_320_353 ();
 FILLCELL_X32 FILLER_320_385 ();
 FILLCELL_X32 FILLER_320_417 ();
 FILLCELL_X32 FILLER_320_449 ();
 FILLCELL_X32 FILLER_320_481 ();
 FILLCELL_X32 FILLER_320_513 ();
 FILLCELL_X32 FILLER_320_545 ();
 FILLCELL_X32 FILLER_320_577 ();
 FILLCELL_X16 FILLER_320_609 ();
 FILLCELL_X4 FILLER_320_625 ();
 FILLCELL_X2 FILLER_320_629 ();
 FILLCELL_X32 FILLER_320_632 ();
 FILLCELL_X32 FILLER_320_664 ();
 FILLCELL_X32 FILLER_320_696 ();
 FILLCELL_X32 FILLER_320_728 ();
 FILLCELL_X32 FILLER_320_760 ();
 FILLCELL_X32 FILLER_320_792 ();
 FILLCELL_X32 FILLER_320_824 ();
 FILLCELL_X32 FILLER_320_856 ();
 FILLCELL_X32 FILLER_320_888 ();
 FILLCELL_X32 FILLER_320_920 ();
 FILLCELL_X32 FILLER_320_952 ();
 FILLCELL_X32 FILLER_320_984 ();
 FILLCELL_X32 FILLER_320_1016 ();
 FILLCELL_X32 FILLER_320_1048 ();
 FILLCELL_X32 FILLER_320_1080 ();
 FILLCELL_X32 FILLER_320_1112 ();
 FILLCELL_X32 FILLER_320_1144 ();
 FILLCELL_X32 FILLER_320_1176 ();
 FILLCELL_X32 FILLER_320_1208 ();
 FILLCELL_X32 FILLER_320_1240 ();
 FILLCELL_X32 FILLER_320_1272 ();
 FILLCELL_X32 FILLER_320_1304 ();
 FILLCELL_X32 FILLER_320_1336 ();
 FILLCELL_X32 FILLER_320_1368 ();
 FILLCELL_X32 FILLER_320_1400 ();
 FILLCELL_X32 FILLER_320_1432 ();
 FILLCELL_X32 FILLER_320_1464 ();
 FILLCELL_X32 FILLER_320_1496 ();
 FILLCELL_X32 FILLER_320_1528 ();
 FILLCELL_X32 FILLER_320_1560 ();
 FILLCELL_X32 FILLER_320_1592 ();
 FILLCELL_X32 FILLER_320_1624 ();
 FILLCELL_X32 FILLER_320_1656 ();
 FILLCELL_X32 FILLER_320_1688 ();
 FILLCELL_X32 FILLER_320_1720 ();
 FILLCELL_X32 FILLER_320_1752 ();
 FILLCELL_X32 FILLER_320_1784 ();
 FILLCELL_X32 FILLER_320_1816 ();
 FILLCELL_X32 FILLER_320_1848 ();
 FILLCELL_X8 FILLER_320_1880 ();
 FILLCELL_X4 FILLER_320_1888 ();
 FILLCELL_X2 FILLER_320_1892 ();
 FILLCELL_X32 FILLER_320_1895 ();
 FILLCELL_X32 FILLER_320_1927 ();
 FILLCELL_X32 FILLER_320_1959 ();
 FILLCELL_X32 FILLER_320_1991 ();
 FILLCELL_X32 FILLER_320_2023 ();
 FILLCELL_X32 FILLER_320_2055 ();
 FILLCELL_X32 FILLER_320_2087 ();
 FILLCELL_X32 FILLER_320_2119 ();
 FILLCELL_X32 FILLER_320_2151 ();
 FILLCELL_X32 FILLER_320_2183 ();
 FILLCELL_X32 FILLER_320_2215 ();
 FILLCELL_X32 FILLER_320_2247 ();
 FILLCELL_X32 FILLER_320_2279 ();
 FILLCELL_X32 FILLER_320_2311 ();
 FILLCELL_X32 FILLER_320_2343 ();
 FILLCELL_X32 FILLER_320_2375 ();
 FILLCELL_X32 FILLER_320_2407 ();
 FILLCELL_X32 FILLER_320_2439 ();
 FILLCELL_X32 FILLER_320_2471 ();
 FILLCELL_X32 FILLER_320_2503 ();
 FILLCELL_X32 FILLER_320_2535 ();
 FILLCELL_X32 FILLER_320_2567 ();
 FILLCELL_X32 FILLER_320_2599 ();
 FILLCELL_X32 FILLER_320_2631 ();
 FILLCELL_X32 FILLER_320_2663 ();
 FILLCELL_X32 FILLER_320_2695 ();
 FILLCELL_X32 FILLER_320_2727 ();
 FILLCELL_X32 FILLER_320_2759 ();
 FILLCELL_X32 FILLER_320_2791 ();
 FILLCELL_X32 FILLER_320_2823 ();
 FILLCELL_X32 FILLER_320_2855 ();
 FILLCELL_X32 FILLER_320_2887 ();
 FILLCELL_X32 FILLER_320_2919 ();
 FILLCELL_X32 FILLER_320_2951 ();
 FILLCELL_X32 FILLER_320_2983 ();
 FILLCELL_X32 FILLER_320_3015 ();
 FILLCELL_X32 FILLER_320_3047 ();
 FILLCELL_X32 FILLER_320_3079 ();
 FILLCELL_X32 FILLER_320_3111 ();
 FILLCELL_X8 FILLER_320_3143 ();
 FILLCELL_X4 FILLER_320_3151 ();
 FILLCELL_X2 FILLER_320_3155 ();
 FILLCELL_X32 FILLER_320_3158 ();
 FILLCELL_X32 FILLER_320_3190 ();
 FILLCELL_X32 FILLER_320_3222 ();
 FILLCELL_X32 FILLER_320_3254 ();
 FILLCELL_X32 FILLER_320_3286 ();
 FILLCELL_X32 FILLER_320_3318 ();
 FILLCELL_X32 FILLER_320_3350 ();
 FILLCELL_X32 FILLER_320_3382 ();
 FILLCELL_X32 FILLER_320_3414 ();
 FILLCELL_X32 FILLER_320_3446 ();
 FILLCELL_X32 FILLER_320_3478 ();
 FILLCELL_X32 FILLER_320_3510 ();
 FILLCELL_X32 FILLER_320_3542 ();
 FILLCELL_X32 FILLER_320_3574 ();
 FILLCELL_X32 FILLER_320_3606 ();
 FILLCELL_X32 FILLER_320_3638 ();
 FILLCELL_X32 FILLER_320_3670 ();
 FILLCELL_X32 FILLER_320_3702 ();
 FILLCELL_X4 FILLER_320_3734 ();
 FILLCELL_X32 FILLER_321_1 ();
 FILLCELL_X32 FILLER_321_33 ();
 FILLCELL_X32 FILLER_321_65 ();
 FILLCELL_X32 FILLER_321_97 ();
 FILLCELL_X32 FILLER_321_129 ();
 FILLCELL_X32 FILLER_321_161 ();
 FILLCELL_X32 FILLER_321_193 ();
 FILLCELL_X32 FILLER_321_225 ();
 FILLCELL_X32 FILLER_321_257 ();
 FILLCELL_X32 FILLER_321_289 ();
 FILLCELL_X32 FILLER_321_321 ();
 FILLCELL_X32 FILLER_321_353 ();
 FILLCELL_X32 FILLER_321_385 ();
 FILLCELL_X32 FILLER_321_417 ();
 FILLCELL_X32 FILLER_321_449 ();
 FILLCELL_X32 FILLER_321_481 ();
 FILLCELL_X32 FILLER_321_513 ();
 FILLCELL_X32 FILLER_321_545 ();
 FILLCELL_X32 FILLER_321_577 ();
 FILLCELL_X32 FILLER_321_609 ();
 FILLCELL_X32 FILLER_321_641 ();
 FILLCELL_X32 FILLER_321_673 ();
 FILLCELL_X32 FILLER_321_705 ();
 FILLCELL_X32 FILLER_321_737 ();
 FILLCELL_X32 FILLER_321_769 ();
 FILLCELL_X32 FILLER_321_801 ();
 FILLCELL_X32 FILLER_321_833 ();
 FILLCELL_X32 FILLER_321_865 ();
 FILLCELL_X32 FILLER_321_897 ();
 FILLCELL_X32 FILLER_321_929 ();
 FILLCELL_X32 FILLER_321_961 ();
 FILLCELL_X32 FILLER_321_993 ();
 FILLCELL_X32 FILLER_321_1025 ();
 FILLCELL_X32 FILLER_321_1057 ();
 FILLCELL_X32 FILLER_321_1089 ();
 FILLCELL_X32 FILLER_321_1121 ();
 FILLCELL_X32 FILLER_321_1153 ();
 FILLCELL_X32 FILLER_321_1185 ();
 FILLCELL_X32 FILLER_321_1217 ();
 FILLCELL_X8 FILLER_321_1249 ();
 FILLCELL_X4 FILLER_321_1257 ();
 FILLCELL_X2 FILLER_321_1261 ();
 FILLCELL_X32 FILLER_321_1264 ();
 FILLCELL_X32 FILLER_321_1296 ();
 FILLCELL_X32 FILLER_321_1328 ();
 FILLCELL_X32 FILLER_321_1360 ();
 FILLCELL_X32 FILLER_321_1392 ();
 FILLCELL_X32 FILLER_321_1424 ();
 FILLCELL_X32 FILLER_321_1456 ();
 FILLCELL_X32 FILLER_321_1488 ();
 FILLCELL_X32 FILLER_321_1520 ();
 FILLCELL_X32 FILLER_321_1552 ();
 FILLCELL_X32 FILLER_321_1584 ();
 FILLCELL_X32 FILLER_321_1616 ();
 FILLCELL_X32 FILLER_321_1648 ();
 FILLCELL_X32 FILLER_321_1680 ();
 FILLCELL_X32 FILLER_321_1712 ();
 FILLCELL_X32 FILLER_321_1744 ();
 FILLCELL_X32 FILLER_321_1776 ();
 FILLCELL_X32 FILLER_321_1808 ();
 FILLCELL_X32 FILLER_321_1840 ();
 FILLCELL_X32 FILLER_321_1872 ();
 FILLCELL_X32 FILLER_321_1904 ();
 FILLCELL_X32 FILLER_321_1936 ();
 FILLCELL_X32 FILLER_321_1968 ();
 FILLCELL_X32 FILLER_321_2000 ();
 FILLCELL_X32 FILLER_321_2032 ();
 FILLCELL_X32 FILLER_321_2064 ();
 FILLCELL_X32 FILLER_321_2096 ();
 FILLCELL_X32 FILLER_321_2128 ();
 FILLCELL_X32 FILLER_321_2160 ();
 FILLCELL_X32 FILLER_321_2192 ();
 FILLCELL_X32 FILLER_321_2224 ();
 FILLCELL_X32 FILLER_321_2256 ();
 FILLCELL_X32 FILLER_321_2288 ();
 FILLCELL_X32 FILLER_321_2320 ();
 FILLCELL_X32 FILLER_321_2352 ();
 FILLCELL_X32 FILLER_321_2384 ();
 FILLCELL_X32 FILLER_321_2416 ();
 FILLCELL_X32 FILLER_321_2448 ();
 FILLCELL_X32 FILLER_321_2480 ();
 FILLCELL_X8 FILLER_321_2512 ();
 FILLCELL_X4 FILLER_321_2520 ();
 FILLCELL_X2 FILLER_321_2524 ();
 FILLCELL_X32 FILLER_321_2527 ();
 FILLCELL_X32 FILLER_321_2559 ();
 FILLCELL_X32 FILLER_321_2591 ();
 FILLCELL_X32 FILLER_321_2623 ();
 FILLCELL_X32 FILLER_321_2655 ();
 FILLCELL_X32 FILLER_321_2687 ();
 FILLCELL_X32 FILLER_321_2719 ();
 FILLCELL_X32 FILLER_321_2751 ();
 FILLCELL_X32 FILLER_321_2783 ();
 FILLCELL_X32 FILLER_321_2815 ();
 FILLCELL_X32 FILLER_321_2847 ();
 FILLCELL_X32 FILLER_321_2879 ();
 FILLCELL_X32 FILLER_321_2911 ();
 FILLCELL_X32 FILLER_321_2943 ();
 FILLCELL_X32 FILLER_321_2975 ();
 FILLCELL_X32 FILLER_321_3007 ();
 FILLCELL_X32 FILLER_321_3039 ();
 FILLCELL_X32 FILLER_321_3071 ();
 FILLCELL_X32 FILLER_321_3103 ();
 FILLCELL_X32 FILLER_321_3135 ();
 FILLCELL_X32 FILLER_321_3167 ();
 FILLCELL_X32 FILLER_321_3199 ();
 FILLCELL_X32 FILLER_321_3231 ();
 FILLCELL_X32 FILLER_321_3263 ();
 FILLCELL_X32 FILLER_321_3295 ();
 FILLCELL_X32 FILLER_321_3327 ();
 FILLCELL_X32 FILLER_321_3359 ();
 FILLCELL_X32 FILLER_321_3391 ();
 FILLCELL_X32 FILLER_321_3423 ();
 FILLCELL_X32 FILLER_321_3455 ();
 FILLCELL_X32 FILLER_321_3487 ();
 FILLCELL_X32 FILLER_321_3519 ();
 FILLCELL_X32 FILLER_321_3551 ();
 FILLCELL_X32 FILLER_321_3583 ();
 FILLCELL_X32 FILLER_321_3615 ();
 FILLCELL_X32 FILLER_321_3647 ();
 FILLCELL_X32 FILLER_321_3679 ();
 FILLCELL_X16 FILLER_321_3711 ();
 FILLCELL_X8 FILLER_321_3727 ();
 FILLCELL_X2 FILLER_321_3735 ();
 FILLCELL_X1 FILLER_321_3737 ();
 FILLCELL_X32 FILLER_322_1 ();
 FILLCELL_X32 FILLER_322_33 ();
 FILLCELL_X32 FILLER_322_65 ();
 FILLCELL_X32 FILLER_322_97 ();
 FILLCELL_X32 FILLER_322_129 ();
 FILLCELL_X32 FILLER_322_161 ();
 FILLCELL_X32 FILLER_322_193 ();
 FILLCELL_X32 FILLER_322_225 ();
 FILLCELL_X32 FILLER_322_257 ();
 FILLCELL_X32 FILLER_322_289 ();
 FILLCELL_X32 FILLER_322_321 ();
 FILLCELL_X32 FILLER_322_353 ();
 FILLCELL_X32 FILLER_322_385 ();
 FILLCELL_X32 FILLER_322_417 ();
 FILLCELL_X32 FILLER_322_449 ();
 FILLCELL_X32 FILLER_322_481 ();
 FILLCELL_X32 FILLER_322_513 ();
 FILLCELL_X32 FILLER_322_545 ();
 FILLCELL_X32 FILLER_322_577 ();
 FILLCELL_X16 FILLER_322_609 ();
 FILLCELL_X4 FILLER_322_625 ();
 FILLCELL_X2 FILLER_322_629 ();
 FILLCELL_X32 FILLER_322_632 ();
 FILLCELL_X32 FILLER_322_664 ();
 FILLCELL_X32 FILLER_322_696 ();
 FILLCELL_X32 FILLER_322_728 ();
 FILLCELL_X32 FILLER_322_760 ();
 FILLCELL_X32 FILLER_322_792 ();
 FILLCELL_X32 FILLER_322_824 ();
 FILLCELL_X32 FILLER_322_856 ();
 FILLCELL_X32 FILLER_322_888 ();
 FILLCELL_X32 FILLER_322_920 ();
 FILLCELL_X32 FILLER_322_952 ();
 FILLCELL_X32 FILLER_322_984 ();
 FILLCELL_X32 FILLER_322_1016 ();
 FILLCELL_X32 FILLER_322_1048 ();
 FILLCELL_X32 FILLER_322_1080 ();
 FILLCELL_X32 FILLER_322_1112 ();
 FILLCELL_X32 FILLER_322_1144 ();
 FILLCELL_X32 FILLER_322_1176 ();
 FILLCELL_X32 FILLER_322_1208 ();
 FILLCELL_X32 FILLER_322_1240 ();
 FILLCELL_X32 FILLER_322_1272 ();
 FILLCELL_X32 FILLER_322_1304 ();
 FILLCELL_X32 FILLER_322_1336 ();
 FILLCELL_X32 FILLER_322_1368 ();
 FILLCELL_X32 FILLER_322_1400 ();
 FILLCELL_X32 FILLER_322_1432 ();
 FILLCELL_X32 FILLER_322_1464 ();
 FILLCELL_X32 FILLER_322_1496 ();
 FILLCELL_X32 FILLER_322_1528 ();
 FILLCELL_X32 FILLER_322_1560 ();
 FILLCELL_X32 FILLER_322_1592 ();
 FILLCELL_X32 FILLER_322_1624 ();
 FILLCELL_X32 FILLER_322_1656 ();
 FILLCELL_X32 FILLER_322_1688 ();
 FILLCELL_X32 FILLER_322_1720 ();
 FILLCELL_X32 FILLER_322_1752 ();
 FILLCELL_X32 FILLER_322_1784 ();
 FILLCELL_X32 FILLER_322_1816 ();
 FILLCELL_X32 FILLER_322_1848 ();
 FILLCELL_X8 FILLER_322_1880 ();
 FILLCELL_X4 FILLER_322_1888 ();
 FILLCELL_X2 FILLER_322_1892 ();
 FILLCELL_X32 FILLER_322_1895 ();
 FILLCELL_X32 FILLER_322_1927 ();
 FILLCELL_X32 FILLER_322_1959 ();
 FILLCELL_X32 FILLER_322_1991 ();
 FILLCELL_X32 FILLER_322_2023 ();
 FILLCELL_X32 FILLER_322_2055 ();
 FILLCELL_X32 FILLER_322_2087 ();
 FILLCELL_X32 FILLER_322_2119 ();
 FILLCELL_X32 FILLER_322_2151 ();
 FILLCELL_X32 FILLER_322_2183 ();
 FILLCELL_X32 FILLER_322_2215 ();
 FILLCELL_X32 FILLER_322_2247 ();
 FILLCELL_X32 FILLER_322_2279 ();
 FILLCELL_X32 FILLER_322_2311 ();
 FILLCELL_X32 FILLER_322_2343 ();
 FILLCELL_X32 FILLER_322_2375 ();
 FILLCELL_X32 FILLER_322_2407 ();
 FILLCELL_X32 FILLER_322_2439 ();
 FILLCELL_X32 FILLER_322_2471 ();
 FILLCELL_X32 FILLER_322_2503 ();
 FILLCELL_X32 FILLER_322_2535 ();
 FILLCELL_X32 FILLER_322_2567 ();
 FILLCELL_X32 FILLER_322_2599 ();
 FILLCELL_X32 FILLER_322_2631 ();
 FILLCELL_X32 FILLER_322_2663 ();
 FILLCELL_X32 FILLER_322_2695 ();
 FILLCELL_X32 FILLER_322_2727 ();
 FILLCELL_X32 FILLER_322_2759 ();
 FILLCELL_X32 FILLER_322_2791 ();
 FILLCELL_X32 FILLER_322_2823 ();
 FILLCELL_X32 FILLER_322_2855 ();
 FILLCELL_X32 FILLER_322_2887 ();
 FILLCELL_X32 FILLER_322_2919 ();
 FILLCELL_X32 FILLER_322_2951 ();
 FILLCELL_X32 FILLER_322_2983 ();
 FILLCELL_X32 FILLER_322_3015 ();
 FILLCELL_X32 FILLER_322_3047 ();
 FILLCELL_X32 FILLER_322_3079 ();
 FILLCELL_X32 FILLER_322_3111 ();
 FILLCELL_X8 FILLER_322_3143 ();
 FILLCELL_X4 FILLER_322_3151 ();
 FILLCELL_X2 FILLER_322_3155 ();
 FILLCELL_X32 FILLER_322_3158 ();
 FILLCELL_X32 FILLER_322_3190 ();
 FILLCELL_X32 FILLER_322_3222 ();
 FILLCELL_X32 FILLER_322_3254 ();
 FILLCELL_X32 FILLER_322_3286 ();
 FILLCELL_X32 FILLER_322_3318 ();
 FILLCELL_X32 FILLER_322_3350 ();
 FILLCELL_X32 FILLER_322_3382 ();
 FILLCELL_X32 FILLER_322_3414 ();
 FILLCELL_X32 FILLER_322_3446 ();
 FILLCELL_X32 FILLER_322_3478 ();
 FILLCELL_X32 FILLER_322_3510 ();
 FILLCELL_X32 FILLER_322_3542 ();
 FILLCELL_X32 FILLER_322_3574 ();
 FILLCELL_X32 FILLER_322_3606 ();
 FILLCELL_X32 FILLER_322_3638 ();
 FILLCELL_X32 FILLER_322_3670 ();
 FILLCELL_X32 FILLER_322_3702 ();
 FILLCELL_X4 FILLER_322_3734 ();
 FILLCELL_X32 FILLER_323_1 ();
 FILLCELL_X32 FILLER_323_33 ();
 FILLCELL_X32 FILLER_323_65 ();
 FILLCELL_X32 FILLER_323_97 ();
 FILLCELL_X32 FILLER_323_129 ();
 FILLCELL_X32 FILLER_323_161 ();
 FILLCELL_X32 FILLER_323_193 ();
 FILLCELL_X32 FILLER_323_225 ();
 FILLCELL_X32 FILLER_323_257 ();
 FILLCELL_X32 FILLER_323_289 ();
 FILLCELL_X32 FILLER_323_321 ();
 FILLCELL_X32 FILLER_323_353 ();
 FILLCELL_X32 FILLER_323_385 ();
 FILLCELL_X32 FILLER_323_417 ();
 FILLCELL_X32 FILLER_323_449 ();
 FILLCELL_X32 FILLER_323_481 ();
 FILLCELL_X32 FILLER_323_513 ();
 FILLCELL_X32 FILLER_323_545 ();
 FILLCELL_X32 FILLER_323_577 ();
 FILLCELL_X32 FILLER_323_609 ();
 FILLCELL_X32 FILLER_323_641 ();
 FILLCELL_X32 FILLER_323_673 ();
 FILLCELL_X32 FILLER_323_705 ();
 FILLCELL_X32 FILLER_323_737 ();
 FILLCELL_X32 FILLER_323_769 ();
 FILLCELL_X32 FILLER_323_801 ();
 FILLCELL_X32 FILLER_323_833 ();
 FILLCELL_X32 FILLER_323_865 ();
 FILLCELL_X32 FILLER_323_897 ();
 FILLCELL_X32 FILLER_323_929 ();
 FILLCELL_X32 FILLER_323_961 ();
 FILLCELL_X32 FILLER_323_993 ();
 FILLCELL_X32 FILLER_323_1025 ();
 FILLCELL_X32 FILLER_323_1057 ();
 FILLCELL_X32 FILLER_323_1089 ();
 FILLCELL_X32 FILLER_323_1121 ();
 FILLCELL_X32 FILLER_323_1153 ();
 FILLCELL_X32 FILLER_323_1185 ();
 FILLCELL_X32 FILLER_323_1217 ();
 FILLCELL_X8 FILLER_323_1249 ();
 FILLCELL_X4 FILLER_323_1257 ();
 FILLCELL_X2 FILLER_323_1261 ();
 FILLCELL_X32 FILLER_323_1264 ();
 FILLCELL_X32 FILLER_323_1296 ();
 FILLCELL_X32 FILLER_323_1328 ();
 FILLCELL_X32 FILLER_323_1360 ();
 FILLCELL_X32 FILLER_323_1392 ();
 FILLCELL_X32 FILLER_323_1424 ();
 FILLCELL_X32 FILLER_323_1456 ();
 FILLCELL_X32 FILLER_323_1488 ();
 FILLCELL_X32 FILLER_323_1520 ();
 FILLCELL_X32 FILLER_323_1552 ();
 FILLCELL_X32 FILLER_323_1584 ();
 FILLCELL_X32 FILLER_323_1616 ();
 FILLCELL_X32 FILLER_323_1648 ();
 FILLCELL_X32 FILLER_323_1680 ();
 FILLCELL_X32 FILLER_323_1712 ();
 FILLCELL_X32 FILLER_323_1744 ();
 FILLCELL_X32 FILLER_323_1776 ();
 FILLCELL_X32 FILLER_323_1808 ();
 FILLCELL_X32 FILLER_323_1840 ();
 FILLCELL_X32 FILLER_323_1872 ();
 FILLCELL_X32 FILLER_323_1904 ();
 FILLCELL_X32 FILLER_323_1936 ();
 FILLCELL_X32 FILLER_323_1968 ();
 FILLCELL_X32 FILLER_323_2000 ();
 FILLCELL_X32 FILLER_323_2032 ();
 FILLCELL_X32 FILLER_323_2064 ();
 FILLCELL_X32 FILLER_323_2096 ();
 FILLCELL_X32 FILLER_323_2128 ();
 FILLCELL_X32 FILLER_323_2160 ();
 FILLCELL_X32 FILLER_323_2192 ();
 FILLCELL_X32 FILLER_323_2224 ();
 FILLCELL_X32 FILLER_323_2256 ();
 FILLCELL_X32 FILLER_323_2288 ();
 FILLCELL_X32 FILLER_323_2320 ();
 FILLCELL_X32 FILLER_323_2352 ();
 FILLCELL_X32 FILLER_323_2384 ();
 FILLCELL_X32 FILLER_323_2416 ();
 FILLCELL_X32 FILLER_323_2448 ();
 FILLCELL_X32 FILLER_323_2480 ();
 FILLCELL_X8 FILLER_323_2512 ();
 FILLCELL_X4 FILLER_323_2520 ();
 FILLCELL_X2 FILLER_323_2524 ();
 FILLCELL_X32 FILLER_323_2527 ();
 FILLCELL_X32 FILLER_323_2559 ();
 FILLCELL_X32 FILLER_323_2591 ();
 FILLCELL_X32 FILLER_323_2623 ();
 FILLCELL_X32 FILLER_323_2655 ();
 FILLCELL_X32 FILLER_323_2687 ();
 FILLCELL_X32 FILLER_323_2719 ();
 FILLCELL_X32 FILLER_323_2751 ();
 FILLCELL_X32 FILLER_323_2783 ();
 FILLCELL_X32 FILLER_323_2815 ();
 FILLCELL_X32 FILLER_323_2847 ();
 FILLCELL_X32 FILLER_323_2879 ();
 FILLCELL_X32 FILLER_323_2911 ();
 FILLCELL_X32 FILLER_323_2943 ();
 FILLCELL_X32 FILLER_323_2975 ();
 FILLCELL_X32 FILLER_323_3007 ();
 FILLCELL_X32 FILLER_323_3039 ();
 FILLCELL_X32 FILLER_323_3071 ();
 FILLCELL_X32 FILLER_323_3103 ();
 FILLCELL_X32 FILLER_323_3135 ();
 FILLCELL_X32 FILLER_323_3167 ();
 FILLCELL_X32 FILLER_323_3199 ();
 FILLCELL_X32 FILLER_323_3231 ();
 FILLCELL_X32 FILLER_323_3263 ();
 FILLCELL_X32 FILLER_323_3295 ();
 FILLCELL_X32 FILLER_323_3327 ();
 FILLCELL_X32 FILLER_323_3359 ();
 FILLCELL_X32 FILLER_323_3391 ();
 FILLCELL_X32 FILLER_323_3423 ();
 FILLCELL_X32 FILLER_323_3455 ();
 FILLCELL_X32 FILLER_323_3487 ();
 FILLCELL_X32 FILLER_323_3519 ();
 FILLCELL_X32 FILLER_323_3551 ();
 FILLCELL_X32 FILLER_323_3583 ();
 FILLCELL_X32 FILLER_323_3615 ();
 FILLCELL_X32 FILLER_323_3647 ();
 FILLCELL_X32 FILLER_323_3679 ();
 FILLCELL_X16 FILLER_323_3711 ();
 FILLCELL_X8 FILLER_323_3727 ();
 FILLCELL_X2 FILLER_323_3735 ();
 FILLCELL_X1 FILLER_323_3737 ();
 FILLCELL_X32 FILLER_324_1 ();
 FILLCELL_X32 FILLER_324_33 ();
 FILLCELL_X32 FILLER_324_65 ();
 FILLCELL_X32 FILLER_324_97 ();
 FILLCELL_X32 FILLER_324_129 ();
 FILLCELL_X32 FILLER_324_161 ();
 FILLCELL_X32 FILLER_324_193 ();
 FILLCELL_X32 FILLER_324_225 ();
 FILLCELL_X32 FILLER_324_257 ();
 FILLCELL_X32 FILLER_324_289 ();
 FILLCELL_X32 FILLER_324_321 ();
 FILLCELL_X32 FILLER_324_353 ();
 FILLCELL_X32 FILLER_324_385 ();
 FILLCELL_X32 FILLER_324_417 ();
 FILLCELL_X32 FILLER_324_449 ();
 FILLCELL_X32 FILLER_324_481 ();
 FILLCELL_X32 FILLER_324_513 ();
 FILLCELL_X32 FILLER_324_545 ();
 FILLCELL_X32 FILLER_324_577 ();
 FILLCELL_X16 FILLER_324_609 ();
 FILLCELL_X4 FILLER_324_625 ();
 FILLCELL_X2 FILLER_324_629 ();
 FILLCELL_X32 FILLER_324_632 ();
 FILLCELL_X32 FILLER_324_664 ();
 FILLCELL_X32 FILLER_324_696 ();
 FILLCELL_X32 FILLER_324_728 ();
 FILLCELL_X32 FILLER_324_760 ();
 FILLCELL_X32 FILLER_324_792 ();
 FILLCELL_X32 FILLER_324_824 ();
 FILLCELL_X32 FILLER_324_856 ();
 FILLCELL_X32 FILLER_324_888 ();
 FILLCELL_X32 FILLER_324_920 ();
 FILLCELL_X32 FILLER_324_952 ();
 FILLCELL_X32 FILLER_324_984 ();
 FILLCELL_X32 FILLER_324_1016 ();
 FILLCELL_X32 FILLER_324_1048 ();
 FILLCELL_X32 FILLER_324_1080 ();
 FILLCELL_X32 FILLER_324_1112 ();
 FILLCELL_X32 FILLER_324_1144 ();
 FILLCELL_X32 FILLER_324_1176 ();
 FILLCELL_X32 FILLER_324_1208 ();
 FILLCELL_X32 FILLER_324_1240 ();
 FILLCELL_X32 FILLER_324_1272 ();
 FILLCELL_X32 FILLER_324_1304 ();
 FILLCELL_X32 FILLER_324_1336 ();
 FILLCELL_X32 FILLER_324_1368 ();
 FILLCELL_X32 FILLER_324_1400 ();
 FILLCELL_X32 FILLER_324_1432 ();
 FILLCELL_X32 FILLER_324_1464 ();
 FILLCELL_X32 FILLER_324_1496 ();
 FILLCELL_X32 FILLER_324_1528 ();
 FILLCELL_X32 FILLER_324_1560 ();
 FILLCELL_X32 FILLER_324_1592 ();
 FILLCELL_X32 FILLER_324_1624 ();
 FILLCELL_X32 FILLER_324_1656 ();
 FILLCELL_X32 FILLER_324_1688 ();
 FILLCELL_X32 FILLER_324_1720 ();
 FILLCELL_X32 FILLER_324_1752 ();
 FILLCELL_X32 FILLER_324_1784 ();
 FILLCELL_X32 FILLER_324_1816 ();
 FILLCELL_X32 FILLER_324_1848 ();
 FILLCELL_X8 FILLER_324_1880 ();
 FILLCELL_X4 FILLER_324_1888 ();
 FILLCELL_X2 FILLER_324_1892 ();
 FILLCELL_X32 FILLER_324_1895 ();
 FILLCELL_X32 FILLER_324_1927 ();
 FILLCELL_X32 FILLER_324_1959 ();
 FILLCELL_X32 FILLER_324_1991 ();
 FILLCELL_X32 FILLER_324_2023 ();
 FILLCELL_X32 FILLER_324_2055 ();
 FILLCELL_X32 FILLER_324_2087 ();
 FILLCELL_X32 FILLER_324_2119 ();
 FILLCELL_X32 FILLER_324_2151 ();
 FILLCELL_X32 FILLER_324_2183 ();
 FILLCELL_X32 FILLER_324_2215 ();
 FILLCELL_X32 FILLER_324_2247 ();
 FILLCELL_X32 FILLER_324_2279 ();
 FILLCELL_X32 FILLER_324_2311 ();
 FILLCELL_X32 FILLER_324_2343 ();
 FILLCELL_X32 FILLER_324_2375 ();
 FILLCELL_X32 FILLER_324_2407 ();
 FILLCELL_X32 FILLER_324_2439 ();
 FILLCELL_X32 FILLER_324_2471 ();
 FILLCELL_X32 FILLER_324_2503 ();
 FILLCELL_X32 FILLER_324_2535 ();
 FILLCELL_X32 FILLER_324_2567 ();
 FILLCELL_X32 FILLER_324_2599 ();
 FILLCELL_X32 FILLER_324_2631 ();
 FILLCELL_X32 FILLER_324_2663 ();
 FILLCELL_X32 FILLER_324_2695 ();
 FILLCELL_X32 FILLER_324_2727 ();
 FILLCELL_X32 FILLER_324_2759 ();
 FILLCELL_X32 FILLER_324_2791 ();
 FILLCELL_X32 FILLER_324_2823 ();
 FILLCELL_X32 FILLER_324_2855 ();
 FILLCELL_X32 FILLER_324_2887 ();
 FILLCELL_X32 FILLER_324_2919 ();
 FILLCELL_X32 FILLER_324_2951 ();
 FILLCELL_X32 FILLER_324_2983 ();
 FILLCELL_X32 FILLER_324_3015 ();
 FILLCELL_X32 FILLER_324_3047 ();
 FILLCELL_X32 FILLER_324_3079 ();
 FILLCELL_X32 FILLER_324_3111 ();
 FILLCELL_X8 FILLER_324_3143 ();
 FILLCELL_X4 FILLER_324_3151 ();
 FILLCELL_X2 FILLER_324_3155 ();
 FILLCELL_X32 FILLER_324_3158 ();
 FILLCELL_X32 FILLER_324_3190 ();
 FILLCELL_X32 FILLER_324_3222 ();
 FILLCELL_X32 FILLER_324_3254 ();
 FILLCELL_X32 FILLER_324_3286 ();
 FILLCELL_X32 FILLER_324_3318 ();
 FILLCELL_X32 FILLER_324_3350 ();
 FILLCELL_X32 FILLER_324_3382 ();
 FILLCELL_X32 FILLER_324_3414 ();
 FILLCELL_X32 FILLER_324_3446 ();
 FILLCELL_X32 FILLER_324_3478 ();
 FILLCELL_X32 FILLER_324_3510 ();
 FILLCELL_X32 FILLER_324_3542 ();
 FILLCELL_X32 FILLER_324_3574 ();
 FILLCELL_X32 FILLER_324_3606 ();
 FILLCELL_X32 FILLER_324_3638 ();
 FILLCELL_X32 FILLER_324_3670 ();
 FILLCELL_X32 FILLER_324_3702 ();
 FILLCELL_X4 FILLER_324_3734 ();
 FILLCELL_X32 FILLER_325_1 ();
 FILLCELL_X32 FILLER_325_33 ();
 FILLCELL_X32 FILLER_325_65 ();
 FILLCELL_X32 FILLER_325_97 ();
 FILLCELL_X32 FILLER_325_129 ();
 FILLCELL_X32 FILLER_325_161 ();
 FILLCELL_X32 FILLER_325_193 ();
 FILLCELL_X32 FILLER_325_225 ();
 FILLCELL_X32 FILLER_325_257 ();
 FILLCELL_X32 FILLER_325_289 ();
 FILLCELL_X32 FILLER_325_321 ();
 FILLCELL_X32 FILLER_325_353 ();
 FILLCELL_X32 FILLER_325_385 ();
 FILLCELL_X32 FILLER_325_417 ();
 FILLCELL_X32 FILLER_325_449 ();
 FILLCELL_X32 FILLER_325_481 ();
 FILLCELL_X32 FILLER_325_513 ();
 FILLCELL_X32 FILLER_325_545 ();
 FILLCELL_X32 FILLER_325_577 ();
 FILLCELL_X32 FILLER_325_609 ();
 FILLCELL_X32 FILLER_325_641 ();
 FILLCELL_X32 FILLER_325_673 ();
 FILLCELL_X32 FILLER_325_705 ();
 FILLCELL_X32 FILLER_325_737 ();
 FILLCELL_X32 FILLER_325_769 ();
 FILLCELL_X32 FILLER_325_801 ();
 FILLCELL_X32 FILLER_325_833 ();
 FILLCELL_X32 FILLER_325_865 ();
 FILLCELL_X32 FILLER_325_897 ();
 FILLCELL_X32 FILLER_325_929 ();
 FILLCELL_X32 FILLER_325_961 ();
 FILLCELL_X32 FILLER_325_993 ();
 FILLCELL_X32 FILLER_325_1025 ();
 FILLCELL_X32 FILLER_325_1057 ();
 FILLCELL_X32 FILLER_325_1089 ();
 FILLCELL_X32 FILLER_325_1121 ();
 FILLCELL_X32 FILLER_325_1153 ();
 FILLCELL_X32 FILLER_325_1185 ();
 FILLCELL_X32 FILLER_325_1217 ();
 FILLCELL_X8 FILLER_325_1249 ();
 FILLCELL_X4 FILLER_325_1257 ();
 FILLCELL_X2 FILLER_325_1261 ();
 FILLCELL_X32 FILLER_325_1264 ();
 FILLCELL_X32 FILLER_325_1296 ();
 FILLCELL_X32 FILLER_325_1328 ();
 FILLCELL_X32 FILLER_325_1360 ();
 FILLCELL_X32 FILLER_325_1392 ();
 FILLCELL_X32 FILLER_325_1424 ();
 FILLCELL_X32 FILLER_325_1456 ();
 FILLCELL_X32 FILLER_325_1488 ();
 FILLCELL_X32 FILLER_325_1520 ();
 FILLCELL_X32 FILLER_325_1552 ();
 FILLCELL_X32 FILLER_325_1584 ();
 FILLCELL_X32 FILLER_325_1616 ();
 FILLCELL_X32 FILLER_325_1648 ();
 FILLCELL_X32 FILLER_325_1680 ();
 FILLCELL_X32 FILLER_325_1712 ();
 FILLCELL_X32 FILLER_325_1744 ();
 FILLCELL_X32 FILLER_325_1776 ();
 FILLCELL_X32 FILLER_325_1808 ();
 FILLCELL_X32 FILLER_325_1840 ();
 FILLCELL_X32 FILLER_325_1872 ();
 FILLCELL_X32 FILLER_325_1904 ();
 FILLCELL_X32 FILLER_325_1936 ();
 FILLCELL_X32 FILLER_325_1968 ();
 FILLCELL_X32 FILLER_325_2000 ();
 FILLCELL_X32 FILLER_325_2032 ();
 FILLCELL_X32 FILLER_325_2064 ();
 FILLCELL_X32 FILLER_325_2096 ();
 FILLCELL_X32 FILLER_325_2128 ();
 FILLCELL_X32 FILLER_325_2160 ();
 FILLCELL_X32 FILLER_325_2192 ();
 FILLCELL_X32 FILLER_325_2224 ();
 FILLCELL_X32 FILLER_325_2256 ();
 FILLCELL_X32 FILLER_325_2288 ();
 FILLCELL_X32 FILLER_325_2320 ();
 FILLCELL_X32 FILLER_325_2352 ();
 FILLCELL_X32 FILLER_325_2384 ();
 FILLCELL_X32 FILLER_325_2416 ();
 FILLCELL_X32 FILLER_325_2448 ();
 FILLCELL_X32 FILLER_325_2480 ();
 FILLCELL_X8 FILLER_325_2512 ();
 FILLCELL_X4 FILLER_325_2520 ();
 FILLCELL_X2 FILLER_325_2524 ();
 FILLCELL_X32 FILLER_325_2527 ();
 FILLCELL_X32 FILLER_325_2559 ();
 FILLCELL_X32 FILLER_325_2591 ();
 FILLCELL_X32 FILLER_325_2623 ();
 FILLCELL_X32 FILLER_325_2655 ();
 FILLCELL_X32 FILLER_325_2687 ();
 FILLCELL_X32 FILLER_325_2719 ();
 FILLCELL_X32 FILLER_325_2751 ();
 FILLCELL_X32 FILLER_325_2783 ();
 FILLCELL_X32 FILLER_325_2815 ();
 FILLCELL_X32 FILLER_325_2847 ();
 FILLCELL_X32 FILLER_325_2879 ();
 FILLCELL_X32 FILLER_325_2911 ();
 FILLCELL_X32 FILLER_325_2943 ();
 FILLCELL_X32 FILLER_325_2975 ();
 FILLCELL_X32 FILLER_325_3007 ();
 FILLCELL_X32 FILLER_325_3039 ();
 FILLCELL_X32 FILLER_325_3071 ();
 FILLCELL_X32 FILLER_325_3103 ();
 FILLCELL_X32 FILLER_325_3135 ();
 FILLCELL_X32 FILLER_325_3167 ();
 FILLCELL_X32 FILLER_325_3199 ();
 FILLCELL_X32 FILLER_325_3231 ();
 FILLCELL_X32 FILLER_325_3263 ();
 FILLCELL_X32 FILLER_325_3295 ();
 FILLCELL_X32 FILLER_325_3327 ();
 FILLCELL_X32 FILLER_325_3359 ();
 FILLCELL_X32 FILLER_325_3391 ();
 FILLCELL_X32 FILLER_325_3423 ();
 FILLCELL_X32 FILLER_325_3455 ();
 FILLCELL_X32 FILLER_325_3487 ();
 FILLCELL_X32 FILLER_325_3519 ();
 FILLCELL_X32 FILLER_325_3551 ();
 FILLCELL_X32 FILLER_325_3583 ();
 FILLCELL_X32 FILLER_325_3615 ();
 FILLCELL_X32 FILLER_325_3647 ();
 FILLCELL_X32 FILLER_325_3679 ();
 FILLCELL_X16 FILLER_325_3711 ();
 FILLCELL_X8 FILLER_325_3727 ();
 FILLCELL_X2 FILLER_325_3735 ();
 FILLCELL_X1 FILLER_325_3737 ();
 FILLCELL_X32 FILLER_326_1 ();
 FILLCELL_X32 FILLER_326_33 ();
 FILLCELL_X32 FILLER_326_65 ();
 FILLCELL_X32 FILLER_326_97 ();
 FILLCELL_X32 FILLER_326_129 ();
 FILLCELL_X32 FILLER_326_161 ();
 FILLCELL_X32 FILLER_326_193 ();
 FILLCELL_X32 FILLER_326_225 ();
 FILLCELL_X32 FILLER_326_257 ();
 FILLCELL_X32 FILLER_326_289 ();
 FILLCELL_X32 FILLER_326_321 ();
 FILLCELL_X32 FILLER_326_353 ();
 FILLCELL_X32 FILLER_326_385 ();
 FILLCELL_X32 FILLER_326_417 ();
 FILLCELL_X32 FILLER_326_449 ();
 FILLCELL_X32 FILLER_326_481 ();
 FILLCELL_X32 FILLER_326_513 ();
 FILLCELL_X32 FILLER_326_545 ();
 FILLCELL_X32 FILLER_326_577 ();
 FILLCELL_X16 FILLER_326_609 ();
 FILLCELL_X4 FILLER_326_625 ();
 FILLCELL_X2 FILLER_326_629 ();
 FILLCELL_X32 FILLER_326_632 ();
 FILLCELL_X32 FILLER_326_664 ();
 FILLCELL_X32 FILLER_326_696 ();
 FILLCELL_X32 FILLER_326_728 ();
 FILLCELL_X32 FILLER_326_760 ();
 FILLCELL_X32 FILLER_326_792 ();
 FILLCELL_X32 FILLER_326_824 ();
 FILLCELL_X32 FILLER_326_856 ();
 FILLCELL_X32 FILLER_326_888 ();
 FILLCELL_X32 FILLER_326_920 ();
 FILLCELL_X32 FILLER_326_952 ();
 FILLCELL_X32 FILLER_326_984 ();
 FILLCELL_X32 FILLER_326_1016 ();
 FILLCELL_X32 FILLER_326_1048 ();
 FILLCELL_X32 FILLER_326_1080 ();
 FILLCELL_X32 FILLER_326_1112 ();
 FILLCELL_X32 FILLER_326_1144 ();
 FILLCELL_X32 FILLER_326_1176 ();
 FILLCELL_X32 FILLER_326_1208 ();
 FILLCELL_X32 FILLER_326_1240 ();
 FILLCELL_X32 FILLER_326_1272 ();
 FILLCELL_X32 FILLER_326_1304 ();
 FILLCELL_X32 FILLER_326_1336 ();
 FILLCELL_X32 FILLER_326_1368 ();
 FILLCELL_X32 FILLER_326_1400 ();
 FILLCELL_X32 FILLER_326_1432 ();
 FILLCELL_X32 FILLER_326_1464 ();
 FILLCELL_X32 FILLER_326_1496 ();
 FILLCELL_X32 FILLER_326_1528 ();
 FILLCELL_X32 FILLER_326_1560 ();
 FILLCELL_X32 FILLER_326_1592 ();
 FILLCELL_X32 FILLER_326_1624 ();
 FILLCELL_X32 FILLER_326_1656 ();
 FILLCELL_X32 FILLER_326_1688 ();
 FILLCELL_X32 FILLER_326_1720 ();
 FILLCELL_X32 FILLER_326_1752 ();
 FILLCELL_X32 FILLER_326_1784 ();
 FILLCELL_X32 FILLER_326_1816 ();
 FILLCELL_X32 FILLER_326_1848 ();
 FILLCELL_X8 FILLER_326_1880 ();
 FILLCELL_X4 FILLER_326_1888 ();
 FILLCELL_X2 FILLER_326_1892 ();
 FILLCELL_X32 FILLER_326_1895 ();
 FILLCELL_X32 FILLER_326_1927 ();
 FILLCELL_X32 FILLER_326_1959 ();
 FILLCELL_X32 FILLER_326_1991 ();
 FILLCELL_X32 FILLER_326_2023 ();
 FILLCELL_X32 FILLER_326_2055 ();
 FILLCELL_X32 FILLER_326_2087 ();
 FILLCELL_X32 FILLER_326_2119 ();
 FILLCELL_X32 FILLER_326_2151 ();
 FILLCELL_X32 FILLER_326_2183 ();
 FILLCELL_X32 FILLER_326_2215 ();
 FILLCELL_X32 FILLER_326_2247 ();
 FILLCELL_X32 FILLER_326_2279 ();
 FILLCELL_X32 FILLER_326_2311 ();
 FILLCELL_X32 FILLER_326_2343 ();
 FILLCELL_X32 FILLER_326_2375 ();
 FILLCELL_X32 FILLER_326_2407 ();
 FILLCELL_X32 FILLER_326_2439 ();
 FILLCELL_X32 FILLER_326_2471 ();
 FILLCELL_X32 FILLER_326_2503 ();
 FILLCELL_X32 FILLER_326_2535 ();
 FILLCELL_X32 FILLER_326_2567 ();
 FILLCELL_X32 FILLER_326_2599 ();
 FILLCELL_X32 FILLER_326_2631 ();
 FILLCELL_X32 FILLER_326_2663 ();
 FILLCELL_X32 FILLER_326_2695 ();
 FILLCELL_X32 FILLER_326_2727 ();
 FILLCELL_X32 FILLER_326_2759 ();
 FILLCELL_X32 FILLER_326_2791 ();
 FILLCELL_X32 FILLER_326_2823 ();
 FILLCELL_X32 FILLER_326_2855 ();
 FILLCELL_X32 FILLER_326_2887 ();
 FILLCELL_X32 FILLER_326_2919 ();
 FILLCELL_X32 FILLER_326_2951 ();
 FILLCELL_X32 FILLER_326_2983 ();
 FILLCELL_X32 FILLER_326_3015 ();
 FILLCELL_X32 FILLER_326_3047 ();
 FILLCELL_X32 FILLER_326_3079 ();
 FILLCELL_X32 FILLER_326_3111 ();
 FILLCELL_X8 FILLER_326_3143 ();
 FILLCELL_X4 FILLER_326_3151 ();
 FILLCELL_X2 FILLER_326_3155 ();
 FILLCELL_X32 FILLER_326_3158 ();
 FILLCELL_X32 FILLER_326_3190 ();
 FILLCELL_X32 FILLER_326_3222 ();
 FILLCELL_X32 FILLER_326_3254 ();
 FILLCELL_X32 FILLER_326_3286 ();
 FILLCELL_X32 FILLER_326_3318 ();
 FILLCELL_X32 FILLER_326_3350 ();
 FILLCELL_X32 FILLER_326_3382 ();
 FILLCELL_X32 FILLER_326_3414 ();
 FILLCELL_X32 FILLER_326_3446 ();
 FILLCELL_X32 FILLER_326_3478 ();
 FILLCELL_X32 FILLER_326_3510 ();
 FILLCELL_X32 FILLER_326_3542 ();
 FILLCELL_X32 FILLER_326_3574 ();
 FILLCELL_X32 FILLER_326_3606 ();
 FILLCELL_X32 FILLER_326_3638 ();
 FILLCELL_X32 FILLER_326_3670 ();
 FILLCELL_X32 FILLER_326_3702 ();
 FILLCELL_X4 FILLER_326_3734 ();
 FILLCELL_X32 FILLER_327_1 ();
 FILLCELL_X32 FILLER_327_33 ();
 FILLCELL_X32 FILLER_327_65 ();
 FILLCELL_X32 FILLER_327_97 ();
 FILLCELL_X32 FILLER_327_129 ();
 FILLCELL_X32 FILLER_327_161 ();
 FILLCELL_X32 FILLER_327_193 ();
 FILLCELL_X32 FILLER_327_225 ();
 FILLCELL_X32 FILLER_327_257 ();
 FILLCELL_X32 FILLER_327_289 ();
 FILLCELL_X32 FILLER_327_321 ();
 FILLCELL_X32 FILLER_327_353 ();
 FILLCELL_X32 FILLER_327_385 ();
 FILLCELL_X32 FILLER_327_417 ();
 FILLCELL_X32 FILLER_327_449 ();
 FILLCELL_X32 FILLER_327_481 ();
 FILLCELL_X32 FILLER_327_513 ();
 FILLCELL_X32 FILLER_327_545 ();
 FILLCELL_X32 FILLER_327_577 ();
 FILLCELL_X32 FILLER_327_609 ();
 FILLCELL_X32 FILLER_327_641 ();
 FILLCELL_X32 FILLER_327_673 ();
 FILLCELL_X32 FILLER_327_705 ();
 FILLCELL_X32 FILLER_327_737 ();
 FILLCELL_X32 FILLER_327_769 ();
 FILLCELL_X32 FILLER_327_801 ();
 FILLCELL_X32 FILLER_327_833 ();
 FILLCELL_X32 FILLER_327_865 ();
 FILLCELL_X32 FILLER_327_897 ();
 FILLCELL_X32 FILLER_327_929 ();
 FILLCELL_X32 FILLER_327_961 ();
 FILLCELL_X32 FILLER_327_993 ();
 FILLCELL_X32 FILLER_327_1025 ();
 FILLCELL_X32 FILLER_327_1057 ();
 FILLCELL_X32 FILLER_327_1089 ();
 FILLCELL_X32 FILLER_327_1121 ();
 FILLCELL_X32 FILLER_327_1153 ();
 FILLCELL_X32 FILLER_327_1185 ();
 FILLCELL_X32 FILLER_327_1217 ();
 FILLCELL_X8 FILLER_327_1249 ();
 FILLCELL_X4 FILLER_327_1257 ();
 FILLCELL_X2 FILLER_327_1261 ();
 FILLCELL_X32 FILLER_327_1264 ();
 FILLCELL_X32 FILLER_327_1296 ();
 FILLCELL_X32 FILLER_327_1328 ();
 FILLCELL_X32 FILLER_327_1360 ();
 FILLCELL_X32 FILLER_327_1392 ();
 FILLCELL_X32 FILLER_327_1424 ();
 FILLCELL_X32 FILLER_327_1456 ();
 FILLCELL_X32 FILLER_327_1488 ();
 FILLCELL_X32 FILLER_327_1520 ();
 FILLCELL_X32 FILLER_327_1552 ();
 FILLCELL_X32 FILLER_327_1584 ();
 FILLCELL_X32 FILLER_327_1616 ();
 FILLCELL_X32 FILLER_327_1648 ();
 FILLCELL_X32 FILLER_327_1680 ();
 FILLCELL_X32 FILLER_327_1712 ();
 FILLCELL_X32 FILLER_327_1744 ();
 FILLCELL_X32 FILLER_327_1776 ();
 FILLCELL_X32 FILLER_327_1808 ();
 FILLCELL_X32 FILLER_327_1840 ();
 FILLCELL_X32 FILLER_327_1872 ();
 FILLCELL_X32 FILLER_327_1904 ();
 FILLCELL_X32 FILLER_327_1936 ();
 FILLCELL_X32 FILLER_327_1968 ();
 FILLCELL_X32 FILLER_327_2000 ();
 FILLCELL_X32 FILLER_327_2032 ();
 FILLCELL_X32 FILLER_327_2064 ();
 FILLCELL_X32 FILLER_327_2096 ();
 FILLCELL_X32 FILLER_327_2128 ();
 FILLCELL_X32 FILLER_327_2160 ();
 FILLCELL_X32 FILLER_327_2192 ();
 FILLCELL_X32 FILLER_327_2224 ();
 FILLCELL_X32 FILLER_327_2256 ();
 FILLCELL_X32 FILLER_327_2288 ();
 FILLCELL_X32 FILLER_327_2320 ();
 FILLCELL_X32 FILLER_327_2352 ();
 FILLCELL_X32 FILLER_327_2384 ();
 FILLCELL_X32 FILLER_327_2416 ();
 FILLCELL_X32 FILLER_327_2448 ();
 FILLCELL_X32 FILLER_327_2480 ();
 FILLCELL_X8 FILLER_327_2512 ();
 FILLCELL_X4 FILLER_327_2520 ();
 FILLCELL_X2 FILLER_327_2524 ();
 FILLCELL_X32 FILLER_327_2527 ();
 FILLCELL_X32 FILLER_327_2559 ();
 FILLCELL_X32 FILLER_327_2591 ();
 FILLCELL_X32 FILLER_327_2623 ();
 FILLCELL_X32 FILLER_327_2655 ();
 FILLCELL_X32 FILLER_327_2687 ();
 FILLCELL_X32 FILLER_327_2719 ();
 FILLCELL_X32 FILLER_327_2751 ();
 FILLCELL_X32 FILLER_327_2783 ();
 FILLCELL_X32 FILLER_327_2815 ();
 FILLCELL_X32 FILLER_327_2847 ();
 FILLCELL_X32 FILLER_327_2879 ();
 FILLCELL_X32 FILLER_327_2911 ();
 FILLCELL_X32 FILLER_327_2943 ();
 FILLCELL_X32 FILLER_327_2975 ();
 FILLCELL_X32 FILLER_327_3007 ();
 FILLCELL_X32 FILLER_327_3039 ();
 FILLCELL_X32 FILLER_327_3071 ();
 FILLCELL_X32 FILLER_327_3103 ();
 FILLCELL_X32 FILLER_327_3135 ();
 FILLCELL_X32 FILLER_327_3167 ();
 FILLCELL_X32 FILLER_327_3199 ();
 FILLCELL_X32 FILLER_327_3231 ();
 FILLCELL_X32 FILLER_327_3263 ();
 FILLCELL_X32 FILLER_327_3295 ();
 FILLCELL_X32 FILLER_327_3327 ();
 FILLCELL_X32 FILLER_327_3359 ();
 FILLCELL_X32 FILLER_327_3391 ();
 FILLCELL_X32 FILLER_327_3423 ();
 FILLCELL_X32 FILLER_327_3455 ();
 FILLCELL_X32 FILLER_327_3487 ();
 FILLCELL_X32 FILLER_327_3519 ();
 FILLCELL_X32 FILLER_327_3551 ();
 FILLCELL_X32 FILLER_327_3583 ();
 FILLCELL_X32 FILLER_327_3615 ();
 FILLCELL_X32 FILLER_327_3647 ();
 FILLCELL_X32 FILLER_327_3679 ();
 FILLCELL_X16 FILLER_327_3711 ();
 FILLCELL_X8 FILLER_327_3727 ();
 FILLCELL_X2 FILLER_327_3735 ();
 FILLCELL_X1 FILLER_327_3737 ();
 FILLCELL_X32 FILLER_328_1 ();
 FILLCELL_X32 FILLER_328_33 ();
 FILLCELL_X32 FILLER_328_65 ();
 FILLCELL_X32 FILLER_328_97 ();
 FILLCELL_X32 FILLER_328_129 ();
 FILLCELL_X32 FILLER_328_161 ();
 FILLCELL_X32 FILLER_328_193 ();
 FILLCELL_X32 FILLER_328_225 ();
 FILLCELL_X32 FILLER_328_257 ();
 FILLCELL_X32 FILLER_328_289 ();
 FILLCELL_X32 FILLER_328_321 ();
 FILLCELL_X32 FILLER_328_353 ();
 FILLCELL_X32 FILLER_328_385 ();
 FILLCELL_X32 FILLER_328_417 ();
 FILLCELL_X32 FILLER_328_449 ();
 FILLCELL_X32 FILLER_328_481 ();
 FILLCELL_X32 FILLER_328_513 ();
 FILLCELL_X32 FILLER_328_545 ();
 FILLCELL_X32 FILLER_328_577 ();
 FILLCELL_X16 FILLER_328_609 ();
 FILLCELL_X4 FILLER_328_625 ();
 FILLCELL_X2 FILLER_328_629 ();
 FILLCELL_X32 FILLER_328_632 ();
 FILLCELL_X32 FILLER_328_664 ();
 FILLCELL_X32 FILLER_328_696 ();
 FILLCELL_X32 FILLER_328_728 ();
 FILLCELL_X32 FILLER_328_760 ();
 FILLCELL_X32 FILLER_328_792 ();
 FILLCELL_X32 FILLER_328_824 ();
 FILLCELL_X32 FILLER_328_856 ();
 FILLCELL_X32 FILLER_328_888 ();
 FILLCELL_X32 FILLER_328_920 ();
 FILLCELL_X32 FILLER_328_952 ();
 FILLCELL_X32 FILLER_328_984 ();
 FILLCELL_X32 FILLER_328_1016 ();
 FILLCELL_X32 FILLER_328_1048 ();
 FILLCELL_X32 FILLER_328_1080 ();
 FILLCELL_X32 FILLER_328_1112 ();
 FILLCELL_X32 FILLER_328_1144 ();
 FILLCELL_X32 FILLER_328_1176 ();
 FILLCELL_X32 FILLER_328_1208 ();
 FILLCELL_X32 FILLER_328_1240 ();
 FILLCELL_X32 FILLER_328_1272 ();
 FILLCELL_X32 FILLER_328_1304 ();
 FILLCELL_X32 FILLER_328_1336 ();
 FILLCELL_X32 FILLER_328_1368 ();
 FILLCELL_X32 FILLER_328_1400 ();
 FILLCELL_X32 FILLER_328_1432 ();
 FILLCELL_X32 FILLER_328_1464 ();
 FILLCELL_X32 FILLER_328_1496 ();
 FILLCELL_X32 FILLER_328_1528 ();
 FILLCELL_X32 FILLER_328_1560 ();
 FILLCELL_X32 FILLER_328_1592 ();
 FILLCELL_X32 FILLER_328_1624 ();
 FILLCELL_X32 FILLER_328_1656 ();
 FILLCELL_X32 FILLER_328_1688 ();
 FILLCELL_X32 FILLER_328_1720 ();
 FILLCELL_X32 FILLER_328_1752 ();
 FILLCELL_X32 FILLER_328_1784 ();
 FILLCELL_X32 FILLER_328_1816 ();
 FILLCELL_X32 FILLER_328_1848 ();
 FILLCELL_X8 FILLER_328_1880 ();
 FILLCELL_X4 FILLER_328_1888 ();
 FILLCELL_X2 FILLER_328_1892 ();
 FILLCELL_X32 FILLER_328_1895 ();
 FILLCELL_X32 FILLER_328_1927 ();
 FILLCELL_X32 FILLER_328_1959 ();
 FILLCELL_X32 FILLER_328_1991 ();
 FILLCELL_X32 FILLER_328_2023 ();
 FILLCELL_X32 FILLER_328_2055 ();
 FILLCELL_X32 FILLER_328_2087 ();
 FILLCELL_X32 FILLER_328_2119 ();
 FILLCELL_X32 FILLER_328_2151 ();
 FILLCELL_X32 FILLER_328_2183 ();
 FILLCELL_X32 FILLER_328_2215 ();
 FILLCELL_X32 FILLER_328_2247 ();
 FILLCELL_X32 FILLER_328_2279 ();
 FILLCELL_X32 FILLER_328_2311 ();
 FILLCELL_X32 FILLER_328_2343 ();
 FILLCELL_X32 FILLER_328_2375 ();
 FILLCELL_X32 FILLER_328_2407 ();
 FILLCELL_X32 FILLER_328_2439 ();
 FILLCELL_X32 FILLER_328_2471 ();
 FILLCELL_X32 FILLER_328_2503 ();
 FILLCELL_X32 FILLER_328_2535 ();
 FILLCELL_X32 FILLER_328_2567 ();
 FILLCELL_X32 FILLER_328_2599 ();
 FILLCELL_X32 FILLER_328_2631 ();
 FILLCELL_X32 FILLER_328_2663 ();
 FILLCELL_X32 FILLER_328_2695 ();
 FILLCELL_X32 FILLER_328_2727 ();
 FILLCELL_X32 FILLER_328_2759 ();
 FILLCELL_X32 FILLER_328_2791 ();
 FILLCELL_X32 FILLER_328_2823 ();
 FILLCELL_X32 FILLER_328_2855 ();
 FILLCELL_X32 FILLER_328_2887 ();
 FILLCELL_X32 FILLER_328_2919 ();
 FILLCELL_X32 FILLER_328_2951 ();
 FILLCELL_X32 FILLER_328_2983 ();
 FILLCELL_X32 FILLER_328_3015 ();
 FILLCELL_X32 FILLER_328_3047 ();
 FILLCELL_X32 FILLER_328_3079 ();
 FILLCELL_X32 FILLER_328_3111 ();
 FILLCELL_X8 FILLER_328_3143 ();
 FILLCELL_X4 FILLER_328_3151 ();
 FILLCELL_X2 FILLER_328_3155 ();
 FILLCELL_X32 FILLER_328_3158 ();
 FILLCELL_X32 FILLER_328_3190 ();
 FILLCELL_X32 FILLER_328_3222 ();
 FILLCELL_X32 FILLER_328_3254 ();
 FILLCELL_X32 FILLER_328_3286 ();
 FILLCELL_X32 FILLER_328_3318 ();
 FILLCELL_X32 FILLER_328_3350 ();
 FILLCELL_X32 FILLER_328_3382 ();
 FILLCELL_X32 FILLER_328_3414 ();
 FILLCELL_X32 FILLER_328_3446 ();
 FILLCELL_X32 FILLER_328_3478 ();
 FILLCELL_X32 FILLER_328_3510 ();
 FILLCELL_X32 FILLER_328_3542 ();
 FILLCELL_X32 FILLER_328_3574 ();
 FILLCELL_X32 FILLER_328_3606 ();
 FILLCELL_X32 FILLER_328_3638 ();
 FILLCELL_X32 FILLER_328_3670 ();
 FILLCELL_X32 FILLER_328_3702 ();
 FILLCELL_X4 FILLER_328_3734 ();
 FILLCELL_X32 FILLER_329_1 ();
 FILLCELL_X32 FILLER_329_33 ();
 FILLCELL_X32 FILLER_329_65 ();
 FILLCELL_X32 FILLER_329_97 ();
 FILLCELL_X32 FILLER_329_129 ();
 FILLCELL_X32 FILLER_329_161 ();
 FILLCELL_X32 FILLER_329_193 ();
 FILLCELL_X32 FILLER_329_225 ();
 FILLCELL_X32 FILLER_329_257 ();
 FILLCELL_X32 FILLER_329_289 ();
 FILLCELL_X32 FILLER_329_321 ();
 FILLCELL_X32 FILLER_329_353 ();
 FILLCELL_X32 FILLER_329_385 ();
 FILLCELL_X32 FILLER_329_417 ();
 FILLCELL_X32 FILLER_329_449 ();
 FILLCELL_X32 FILLER_329_481 ();
 FILLCELL_X32 FILLER_329_513 ();
 FILLCELL_X32 FILLER_329_545 ();
 FILLCELL_X32 FILLER_329_577 ();
 FILLCELL_X32 FILLER_329_609 ();
 FILLCELL_X32 FILLER_329_641 ();
 FILLCELL_X32 FILLER_329_673 ();
 FILLCELL_X32 FILLER_329_705 ();
 FILLCELL_X32 FILLER_329_737 ();
 FILLCELL_X32 FILLER_329_769 ();
 FILLCELL_X32 FILLER_329_801 ();
 FILLCELL_X32 FILLER_329_833 ();
 FILLCELL_X32 FILLER_329_865 ();
 FILLCELL_X32 FILLER_329_897 ();
 FILLCELL_X32 FILLER_329_929 ();
 FILLCELL_X32 FILLER_329_961 ();
 FILLCELL_X32 FILLER_329_993 ();
 FILLCELL_X32 FILLER_329_1025 ();
 FILLCELL_X32 FILLER_329_1057 ();
 FILLCELL_X32 FILLER_329_1089 ();
 FILLCELL_X32 FILLER_329_1121 ();
 FILLCELL_X32 FILLER_329_1153 ();
 FILLCELL_X32 FILLER_329_1185 ();
 FILLCELL_X32 FILLER_329_1217 ();
 FILLCELL_X8 FILLER_329_1249 ();
 FILLCELL_X4 FILLER_329_1257 ();
 FILLCELL_X2 FILLER_329_1261 ();
 FILLCELL_X32 FILLER_329_1264 ();
 FILLCELL_X32 FILLER_329_1296 ();
 FILLCELL_X32 FILLER_329_1328 ();
 FILLCELL_X32 FILLER_329_1360 ();
 FILLCELL_X32 FILLER_329_1392 ();
 FILLCELL_X32 FILLER_329_1424 ();
 FILLCELL_X32 FILLER_329_1456 ();
 FILLCELL_X32 FILLER_329_1488 ();
 FILLCELL_X32 FILLER_329_1520 ();
 FILLCELL_X32 FILLER_329_1552 ();
 FILLCELL_X32 FILLER_329_1584 ();
 FILLCELL_X32 FILLER_329_1616 ();
 FILLCELL_X32 FILLER_329_1648 ();
 FILLCELL_X32 FILLER_329_1680 ();
 FILLCELL_X32 FILLER_329_1712 ();
 FILLCELL_X32 FILLER_329_1744 ();
 FILLCELL_X32 FILLER_329_1776 ();
 FILLCELL_X32 FILLER_329_1808 ();
 FILLCELL_X32 FILLER_329_1840 ();
 FILLCELL_X32 FILLER_329_1872 ();
 FILLCELL_X32 FILLER_329_1904 ();
 FILLCELL_X32 FILLER_329_1936 ();
 FILLCELL_X32 FILLER_329_1968 ();
 FILLCELL_X32 FILLER_329_2000 ();
 FILLCELL_X32 FILLER_329_2032 ();
 FILLCELL_X32 FILLER_329_2064 ();
 FILLCELL_X32 FILLER_329_2096 ();
 FILLCELL_X32 FILLER_329_2128 ();
 FILLCELL_X32 FILLER_329_2160 ();
 FILLCELL_X32 FILLER_329_2192 ();
 FILLCELL_X32 FILLER_329_2224 ();
 FILLCELL_X32 FILLER_329_2256 ();
 FILLCELL_X32 FILLER_329_2288 ();
 FILLCELL_X32 FILLER_329_2320 ();
 FILLCELL_X32 FILLER_329_2352 ();
 FILLCELL_X32 FILLER_329_2384 ();
 FILLCELL_X32 FILLER_329_2416 ();
 FILLCELL_X32 FILLER_329_2448 ();
 FILLCELL_X32 FILLER_329_2480 ();
 FILLCELL_X8 FILLER_329_2512 ();
 FILLCELL_X4 FILLER_329_2520 ();
 FILLCELL_X2 FILLER_329_2524 ();
 FILLCELL_X32 FILLER_329_2527 ();
 FILLCELL_X32 FILLER_329_2559 ();
 FILLCELL_X32 FILLER_329_2591 ();
 FILLCELL_X32 FILLER_329_2623 ();
 FILLCELL_X32 FILLER_329_2655 ();
 FILLCELL_X32 FILLER_329_2687 ();
 FILLCELL_X32 FILLER_329_2719 ();
 FILLCELL_X32 FILLER_329_2751 ();
 FILLCELL_X32 FILLER_329_2783 ();
 FILLCELL_X32 FILLER_329_2815 ();
 FILLCELL_X32 FILLER_329_2847 ();
 FILLCELL_X32 FILLER_329_2879 ();
 FILLCELL_X32 FILLER_329_2911 ();
 FILLCELL_X32 FILLER_329_2943 ();
 FILLCELL_X32 FILLER_329_2975 ();
 FILLCELL_X32 FILLER_329_3007 ();
 FILLCELL_X32 FILLER_329_3039 ();
 FILLCELL_X32 FILLER_329_3071 ();
 FILLCELL_X32 FILLER_329_3103 ();
 FILLCELL_X32 FILLER_329_3135 ();
 FILLCELL_X32 FILLER_329_3167 ();
 FILLCELL_X32 FILLER_329_3199 ();
 FILLCELL_X32 FILLER_329_3231 ();
 FILLCELL_X32 FILLER_329_3263 ();
 FILLCELL_X32 FILLER_329_3295 ();
 FILLCELL_X32 FILLER_329_3327 ();
 FILLCELL_X32 FILLER_329_3359 ();
 FILLCELL_X32 FILLER_329_3391 ();
 FILLCELL_X32 FILLER_329_3423 ();
 FILLCELL_X32 FILLER_329_3455 ();
 FILLCELL_X32 FILLER_329_3487 ();
 FILLCELL_X32 FILLER_329_3519 ();
 FILLCELL_X32 FILLER_329_3551 ();
 FILLCELL_X32 FILLER_329_3583 ();
 FILLCELL_X32 FILLER_329_3615 ();
 FILLCELL_X32 FILLER_329_3647 ();
 FILLCELL_X32 FILLER_329_3679 ();
 FILLCELL_X16 FILLER_329_3711 ();
 FILLCELL_X8 FILLER_329_3727 ();
 FILLCELL_X2 FILLER_329_3735 ();
 FILLCELL_X1 FILLER_329_3737 ();
 FILLCELL_X32 FILLER_330_1 ();
 FILLCELL_X32 FILLER_330_33 ();
 FILLCELL_X32 FILLER_330_65 ();
 FILLCELL_X32 FILLER_330_97 ();
 FILLCELL_X32 FILLER_330_129 ();
 FILLCELL_X32 FILLER_330_161 ();
 FILLCELL_X32 FILLER_330_193 ();
 FILLCELL_X32 FILLER_330_225 ();
 FILLCELL_X32 FILLER_330_257 ();
 FILLCELL_X32 FILLER_330_289 ();
 FILLCELL_X32 FILLER_330_321 ();
 FILLCELL_X32 FILLER_330_353 ();
 FILLCELL_X32 FILLER_330_385 ();
 FILLCELL_X32 FILLER_330_417 ();
 FILLCELL_X32 FILLER_330_449 ();
 FILLCELL_X32 FILLER_330_481 ();
 FILLCELL_X32 FILLER_330_513 ();
 FILLCELL_X32 FILLER_330_545 ();
 FILLCELL_X32 FILLER_330_577 ();
 FILLCELL_X16 FILLER_330_609 ();
 FILLCELL_X4 FILLER_330_625 ();
 FILLCELL_X2 FILLER_330_629 ();
 FILLCELL_X32 FILLER_330_632 ();
 FILLCELL_X32 FILLER_330_664 ();
 FILLCELL_X32 FILLER_330_696 ();
 FILLCELL_X32 FILLER_330_728 ();
 FILLCELL_X32 FILLER_330_760 ();
 FILLCELL_X32 FILLER_330_792 ();
 FILLCELL_X32 FILLER_330_824 ();
 FILLCELL_X32 FILLER_330_856 ();
 FILLCELL_X32 FILLER_330_888 ();
 FILLCELL_X32 FILLER_330_920 ();
 FILLCELL_X32 FILLER_330_952 ();
 FILLCELL_X32 FILLER_330_984 ();
 FILLCELL_X32 FILLER_330_1016 ();
 FILLCELL_X32 FILLER_330_1048 ();
 FILLCELL_X32 FILLER_330_1080 ();
 FILLCELL_X32 FILLER_330_1112 ();
 FILLCELL_X32 FILLER_330_1144 ();
 FILLCELL_X32 FILLER_330_1176 ();
 FILLCELL_X32 FILLER_330_1208 ();
 FILLCELL_X32 FILLER_330_1240 ();
 FILLCELL_X32 FILLER_330_1272 ();
 FILLCELL_X32 FILLER_330_1304 ();
 FILLCELL_X32 FILLER_330_1336 ();
 FILLCELL_X32 FILLER_330_1368 ();
 FILLCELL_X32 FILLER_330_1400 ();
 FILLCELL_X32 FILLER_330_1432 ();
 FILLCELL_X32 FILLER_330_1464 ();
 FILLCELL_X32 FILLER_330_1496 ();
 FILLCELL_X32 FILLER_330_1528 ();
 FILLCELL_X32 FILLER_330_1560 ();
 FILLCELL_X32 FILLER_330_1592 ();
 FILLCELL_X32 FILLER_330_1624 ();
 FILLCELL_X32 FILLER_330_1656 ();
 FILLCELL_X32 FILLER_330_1688 ();
 FILLCELL_X32 FILLER_330_1720 ();
 FILLCELL_X32 FILLER_330_1752 ();
 FILLCELL_X32 FILLER_330_1784 ();
 FILLCELL_X32 FILLER_330_1816 ();
 FILLCELL_X32 FILLER_330_1848 ();
 FILLCELL_X8 FILLER_330_1880 ();
 FILLCELL_X4 FILLER_330_1888 ();
 FILLCELL_X2 FILLER_330_1892 ();
 FILLCELL_X32 FILLER_330_1895 ();
 FILLCELL_X32 FILLER_330_1927 ();
 FILLCELL_X32 FILLER_330_1959 ();
 FILLCELL_X32 FILLER_330_1991 ();
 FILLCELL_X32 FILLER_330_2023 ();
 FILLCELL_X32 FILLER_330_2055 ();
 FILLCELL_X32 FILLER_330_2087 ();
 FILLCELL_X32 FILLER_330_2119 ();
 FILLCELL_X32 FILLER_330_2151 ();
 FILLCELL_X32 FILLER_330_2183 ();
 FILLCELL_X32 FILLER_330_2215 ();
 FILLCELL_X32 FILLER_330_2247 ();
 FILLCELL_X32 FILLER_330_2279 ();
 FILLCELL_X32 FILLER_330_2311 ();
 FILLCELL_X32 FILLER_330_2343 ();
 FILLCELL_X32 FILLER_330_2375 ();
 FILLCELL_X32 FILLER_330_2407 ();
 FILLCELL_X32 FILLER_330_2439 ();
 FILLCELL_X32 FILLER_330_2471 ();
 FILLCELL_X32 FILLER_330_2503 ();
 FILLCELL_X32 FILLER_330_2535 ();
 FILLCELL_X32 FILLER_330_2567 ();
 FILLCELL_X32 FILLER_330_2599 ();
 FILLCELL_X32 FILLER_330_2631 ();
 FILLCELL_X32 FILLER_330_2663 ();
 FILLCELL_X32 FILLER_330_2695 ();
 FILLCELL_X32 FILLER_330_2727 ();
 FILLCELL_X32 FILLER_330_2759 ();
 FILLCELL_X32 FILLER_330_2791 ();
 FILLCELL_X32 FILLER_330_2823 ();
 FILLCELL_X32 FILLER_330_2855 ();
 FILLCELL_X32 FILLER_330_2887 ();
 FILLCELL_X32 FILLER_330_2919 ();
 FILLCELL_X32 FILLER_330_2951 ();
 FILLCELL_X32 FILLER_330_2983 ();
 FILLCELL_X32 FILLER_330_3015 ();
 FILLCELL_X32 FILLER_330_3047 ();
 FILLCELL_X32 FILLER_330_3079 ();
 FILLCELL_X32 FILLER_330_3111 ();
 FILLCELL_X8 FILLER_330_3143 ();
 FILLCELL_X4 FILLER_330_3151 ();
 FILLCELL_X2 FILLER_330_3155 ();
 FILLCELL_X32 FILLER_330_3158 ();
 FILLCELL_X32 FILLER_330_3190 ();
 FILLCELL_X32 FILLER_330_3222 ();
 FILLCELL_X32 FILLER_330_3254 ();
 FILLCELL_X32 FILLER_330_3286 ();
 FILLCELL_X32 FILLER_330_3318 ();
 FILLCELL_X32 FILLER_330_3350 ();
 FILLCELL_X32 FILLER_330_3382 ();
 FILLCELL_X32 FILLER_330_3414 ();
 FILLCELL_X32 FILLER_330_3446 ();
 FILLCELL_X32 FILLER_330_3478 ();
 FILLCELL_X32 FILLER_330_3510 ();
 FILLCELL_X32 FILLER_330_3542 ();
 FILLCELL_X32 FILLER_330_3574 ();
 FILLCELL_X32 FILLER_330_3606 ();
 FILLCELL_X32 FILLER_330_3638 ();
 FILLCELL_X32 FILLER_330_3670 ();
 FILLCELL_X32 FILLER_330_3702 ();
 FILLCELL_X4 FILLER_330_3734 ();
 FILLCELL_X32 FILLER_331_1 ();
 FILLCELL_X32 FILLER_331_33 ();
 FILLCELL_X32 FILLER_331_65 ();
 FILLCELL_X32 FILLER_331_97 ();
 FILLCELL_X32 FILLER_331_129 ();
 FILLCELL_X32 FILLER_331_161 ();
 FILLCELL_X32 FILLER_331_193 ();
 FILLCELL_X32 FILLER_331_225 ();
 FILLCELL_X32 FILLER_331_257 ();
 FILLCELL_X32 FILLER_331_289 ();
 FILLCELL_X32 FILLER_331_321 ();
 FILLCELL_X32 FILLER_331_353 ();
 FILLCELL_X32 FILLER_331_385 ();
 FILLCELL_X32 FILLER_331_417 ();
 FILLCELL_X32 FILLER_331_449 ();
 FILLCELL_X32 FILLER_331_481 ();
 FILLCELL_X32 FILLER_331_513 ();
 FILLCELL_X32 FILLER_331_545 ();
 FILLCELL_X32 FILLER_331_577 ();
 FILLCELL_X32 FILLER_331_609 ();
 FILLCELL_X32 FILLER_331_641 ();
 FILLCELL_X32 FILLER_331_673 ();
 FILLCELL_X32 FILLER_331_705 ();
 FILLCELL_X32 FILLER_331_737 ();
 FILLCELL_X32 FILLER_331_769 ();
 FILLCELL_X32 FILLER_331_801 ();
 FILLCELL_X32 FILLER_331_833 ();
 FILLCELL_X32 FILLER_331_865 ();
 FILLCELL_X32 FILLER_331_897 ();
 FILLCELL_X32 FILLER_331_929 ();
 FILLCELL_X32 FILLER_331_961 ();
 FILLCELL_X32 FILLER_331_993 ();
 FILLCELL_X32 FILLER_331_1025 ();
 FILLCELL_X32 FILLER_331_1057 ();
 FILLCELL_X32 FILLER_331_1089 ();
 FILLCELL_X32 FILLER_331_1121 ();
 FILLCELL_X32 FILLER_331_1153 ();
 FILLCELL_X32 FILLER_331_1185 ();
 FILLCELL_X32 FILLER_331_1217 ();
 FILLCELL_X8 FILLER_331_1249 ();
 FILLCELL_X4 FILLER_331_1257 ();
 FILLCELL_X2 FILLER_331_1261 ();
 FILLCELL_X32 FILLER_331_1264 ();
 FILLCELL_X32 FILLER_331_1296 ();
 FILLCELL_X32 FILLER_331_1328 ();
 FILLCELL_X32 FILLER_331_1360 ();
 FILLCELL_X32 FILLER_331_1392 ();
 FILLCELL_X32 FILLER_331_1424 ();
 FILLCELL_X32 FILLER_331_1456 ();
 FILLCELL_X32 FILLER_331_1488 ();
 FILLCELL_X32 FILLER_331_1520 ();
 FILLCELL_X32 FILLER_331_1552 ();
 FILLCELL_X32 FILLER_331_1584 ();
 FILLCELL_X32 FILLER_331_1616 ();
 FILLCELL_X32 FILLER_331_1648 ();
 FILLCELL_X32 FILLER_331_1680 ();
 FILLCELL_X32 FILLER_331_1712 ();
 FILLCELL_X32 FILLER_331_1744 ();
 FILLCELL_X32 FILLER_331_1776 ();
 FILLCELL_X32 FILLER_331_1808 ();
 FILLCELL_X32 FILLER_331_1840 ();
 FILLCELL_X32 FILLER_331_1872 ();
 FILLCELL_X32 FILLER_331_1904 ();
 FILLCELL_X32 FILLER_331_1936 ();
 FILLCELL_X32 FILLER_331_1968 ();
 FILLCELL_X32 FILLER_331_2000 ();
 FILLCELL_X32 FILLER_331_2032 ();
 FILLCELL_X32 FILLER_331_2064 ();
 FILLCELL_X32 FILLER_331_2096 ();
 FILLCELL_X32 FILLER_331_2128 ();
 FILLCELL_X32 FILLER_331_2160 ();
 FILLCELL_X32 FILLER_331_2192 ();
 FILLCELL_X32 FILLER_331_2224 ();
 FILLCELL_X32 FILLER_331_2256 ();
 FILLCELL_X32 FILLER_331_2288 ();
 FILLCELL_X32 FILLER_331_2320 ();
 FILLCELL_X32 FILLER_331_2352 ();
 FILLCELL_X32 FILLER_331_2384 ();
 FILLCELL_X32 FILLER_331_2416 ();
 FILLCELL_X32 FILLER_331_2448 ();
 FILLCELL_X32 FILLER_331_2480 ();
 FILLCELL_X8 FILLER_331_2512 ();
 FILLCELL_X4 FILLER_331_2520 ();
 FILLCELL_X2 FILLER_331_2524 ();
 FILLCELL_X32 FILLER_331_2527 ();
 FILLCELL_X32 FILLER_331_2559 ();
 FILLCELL_X32 FILLER_331_2591 ();
 FILLCELL_X32 FILLER_331_2623 ();
 FILLCELL_X32 FILLER_331_2655 ();
 FILLCELL_X32 FILLER_331_2687 ();
 FILLCELL_X32 FILLER_331_2719 ();
 FILLCELL_X32 FILLER_331_2751 ();
 FILLCELL_X32 FILLER_331_2783 ();
 FILLCELL_X32 FILLER_331_2815 ();
 FILLCELL_X32 FILLER_331_2847 ();
 FILLCELL_X32 FILLER_331_2879 ();
 FILLCELL_X32 FILLER_331_2911 ();
 FILLCELL_X32 FILLER_331_2943 ();
 FILLCELL_X32 FILLER_331_2975 ();
 FILLCELL_X32 FILLER_331_3007 ();
 FILLCELL_X32 FILLER_331_3039 ();
 FILLCELL_X32 FILLER_331_3071 ();
 FILLCELL_X32 FILLER_331_3103 ();
 FILLCELL_X32 FILLER_331_3135 ();
 FILLCELL_X32 FILLER_331_3167 ();
 FILLCELL_X32 FILLER_331_3199 ();
 FILLCELL_X32 FILLER_331_3231 ();
 FILLCELL_X32 FILLER_331_3263 ();
 FILLCELL_X32 FILLER_331_3295 ();
 FILLCELL_X32 FILLER_331_3327 ();
 FILLCELL_X32 FILLER_331_3359 ();
 FILLCELL_X32 FILLER_331_3391 ();
 FILLCELL_X32 FILLER_331_3423 ();
 FILLCELL_X32 FILLER_331_3455 ();
 FILLCELL_X32 FILLER_331_3487 ();
 FILLCELL_X32 FILLER_331_3519 ();
 FILLCELL_X32 FILLER_331_3551 ();
 FILLCELL_X32 FILLER_331_3583 ();
 FILLCELL_X32 FILLER_331_3615 ();
 FILLCELL_X32 FILLER_331_3647 ();
 FILLCELL_X32 FILLER_331_3679 ();
 FILLCELL_X16 FILLER_331_3711 ();
 FILLCELL_X8 FILLER_331_3727 ();
 FILLCELL_X2 FILLER_331_3735 ();
 FILLCELL_X1 FILLER_331_3737 ();
 FILLCELL_X32 FILLER_332_1 ();
 FILLCELL_X32 FILLER_332_33 ();
 FILLCELL_X32 FILLER_332_65 ();
 FILLCELL_X32 FILLER_332_97 ();
 FILLCELL_X32 FILLER_332_129 ();
 FILLCELL_X32 FILLER_332_161 ();
 FILLCELL_X32 FILLER_332_193 ();
 FILLCELL_X32 FILLER_332_225 ();
 FILLCELL_X32 FILLER_332_257 ();
 FILLCELL_X32 FILLER_332_289 ();
 FILLCELL_X32 FILLER_332_321 ();
 FILLCELL_X32 FILLER_332_353 ();
 FILLCELL_X32 FILLER_332_385 ();
 FILLCELL_X32 FILLER_332_417 ();
 FILLCELL_X32 FILLER_332_449 ();
 FILLCELL_X32 FILLER_332_481 ();
 FILLCELL_X32 FILLER_332_513 ();
 FILLCELL_X32 FILLER_332_545 ();
 FILLCELL_X32 FILLER_332_577 ();
 FILLCELL_X16 FILLER_332_609 ();
 FILLCELL_X4 FILLER_332_625 ();
 FILLCELL_X2 FILLER_332_629 ();
 FILLCELL_X32 FILLER_332_632 ();
 FILLCELL_X32 FILLER_332_664 ();
 FILLCELL_X32 FILLER_332_696 ();
 FILLCELL_X32 FILLER_332_728 ();
 FILLCELL_X32 FILLER_332_760 ();
 FILLCELL_X32 FILLER_332_792 ();
 FILLCELL_X32 FILLER_332_824 ();
 FILLCELL_X32 FILLER_332_856 ();
 FILLCELL_X32 FILLER_332_888 ();
 FILLCELL_X32 FILLER_332_920 ();
 FILLCELL_X32 FILLER_332_952 ();
 FILLCELL_X32 FILLER_332_984 ();
 FILLCELL_X32 FILLER_332_1016 ();
 FILLCELL_X32 FILLER_332_1048 ();
 FILLCELL_X32 FILLER_332_1080 ();
 FILLCELL_X32 FILLER_332_1112 ();
 FILLCELL_X32 FILLER_332_1144 ();
 FILLCELL_X32 FILLER_332_1176 ();
 FILLCELL_X32 FILLER_332_1208 ();
 FILLCELL_X32 FILLER_332_1240 ();
 FILLCELL_X32 FILLER_332_1272 ();
 FILLCELL_X32 FILLER_332_1304 ();
 FILLCELL_X32 FILLER_332_1336 ();
 FILLCELL_X32 FILLER_332_1368 ();
 FILLCELL_X32 FILLER_332_1400 ();
 FILLCELL_X32 FILLER_332_1432 ();
 FILLCELL_X32 FILLER_332_1464 ();
 FILLCELL_X32 FILLER_332_1496 ();
 FILLCELL_X32 FILLER_332_1528 ();
 FILLCELL_X32 FILLER_332_1560 ();
 FILLCELL_X32 FILLER_332_1592 ();
 FILLCELL_X32 FILLER_332_1624 ();
 FILLCELL_X32 FILLER_332_1656 ();
 FILLCELL_X32 FILLER_332_1688 ();
 FILLCELL_X32 FILLER_332_1720 ();
 FILLCELL_X32 FILLER_332_1752 ();
 FILLCELL_X32 FILLER_332_1784 ();
 FILLCELL_X32 FILLER_332_1816 ();
 FILLCELL_X32 FILLER_332_1848 ();
 FILLCELL_X8 FILLER_332_1880 ();
 FILLCELL_X4 FILLER_332_1888 ();
 FILLCELL_X2 FILLER_332_1892 ();
 FILLCELL_X32 FILLER_332_1895 ();
 FILLCELL_X32 FILLER_332_1927 ();
 FILLCELL_X32 FILLER_332_1959 ();
 FILLCELL_X32 FILLER_332_1991 ();
 FILLCELL_X32 FILLER_332_2023 ();
 FILLCELL_X32 FILLER_332_2055 ();
 FILLCELL_X32 FILLER_332_2087 ();
 FILLCELL_X32 FILLER_332_2119 ();
 FILLCELL_X32 FILLER_332_2151 ();
 FILLCELL_X32 FILLER_332_2183 ();
 FILLCELL_X32 FILLER_332_2215 ();
 FILLCELL_X32 FILLER_332_2247 ();
 FILLCELL_X32 FILLER_332_2279 ();
 FILLCELL_X32 FILLER_332_2311 ();
 FILLCELL_X32 FILLER_332_2343 ();
 FILLCELL_X32 FILLER_332_2375 ();
 FILLCELL_X32 FILLER_332_2407 ();
 FILLCELL_X32 FILLER_332_2439 ();
 FILLCELL_X32 FILLER_332_2471 ();
 FILLCELL_X32 FILLER_332_2503 ();
 FILLCELL_X32 FILLER_332_2535 ();
 FILLCELL_X32 FILLER_332_2567 ();
 FILLCELL_X32 FILLER_332_2599 ();
 FILLCELL_X32 FILLER_332_2631 ();
 FILLCELL_X32 FILLER_332_2663 ();
 FILLCELL_X32 FILLER_332_2695 ();
 FILLCELL_X32 FILLER_332_2727 ();
 FILLCELL_X32 FILLER_332_2759 ();
 FILLCELL_X32 FILLER_332_2791 ();
 FILLCELL_X32 FILLER_332_2823 ();
 FILLCELL_X32 FILLER_332_2855 ();
 FILLCELL_X32 FILLER_332_2887 ();
 FILLCELL_X32 FILLER_332_2919 ();
 FILLCELL_X32 FILLER_332_2951 ();
 FILLCELL_X32 FILLER_332_2983 ();
 FILLCELL_X32 FILLER_332_3015 ();
 FILLCELL_X32 FILLER_332_3047 ();
 FILLCELL_X32 FILLER_332_3079 ();
 FILLCELL_X32 FILLER_332_3111 ();
 FILLCELL_X8 FILLER_332_3143 ();
 FILLCELL_X4 FILLER_332_3151 ();
 FILLCELL_X2 FILLER_332_3155 ();
 FILLCELL_X32 FILLER_332_3158 ();
 FILLCELL_X32 FILLER_332_3190 ();
 FILLCELL_X32 FILLER_332_3222 ();
 FILLCELL_X32 FILLER_332_3254 ();
 FILLCELL_X32 FILLER_332_3286 ();
 FILLCELL_X32 FILLER_332_3318 ();
 FILLCELL_X32 FILLER_332_3350 ();
 FILLCELL_X32 FILLER_332_3382 ();
 FILLCELL_X32 FILLER_332_3414 ();
 FILLCELL_X32 FILLER_332_3446 ();
 FILLCELL_X32 FILLER_332_3478 ();
 FILLCELL_X32 FILLER_332_3510 ();
 FILLCELL_X32 FILLER_332_3542 ();
 FILLCELL_X32 FILLER_332_3574 ();
 FILLCELL_X32 FILLER_332_3606 ();
 FILLCELL_X32 FILLER_332_3638 ();
 FILLCELL_X32 FILLER_332_3670 ();
 FILLCELL_X32 FILLER_332_3702 ();
 FILLCELL_X4 FILLER_332_3734 ();
 FILLCELL_X32 FILLER_333_1 ();
 FILLCELL_X32 FILLER_333_33 ();
 FILLCELL_X32 FILLER_333_65 ();
 FILLCELL_X32 FILLER_333_97 ();
 FILLCELL_X32 FILLER_333_129 ();
 FILLCELL_X32 FILLER_333_161 ();
 FILLCELL_X32 FILLER_333_193 ();
 FILLCELL_X32 FILLER_333_225 ();
 FILLCELL_X32 FILLER_333_257 ();
 FILLCELL_X32 FILLER_333_289 ();
 FILLCELL_X32 FILLER_333_321 ();
 FILLCELL_X32 FILLER_333_353 ();
 FILLCELL_X32 FILLER_333_385 ();
 FILLCELL_X32 FILLER_333_417 ();
 FILLCELL_X32 FILLER_333_449 ();
 FILLCELL_X32 FILLER_333_481 ();
 FILLCELL_X32 FILLER_333_513 ();
 FILLCELL_X32 FILLER_333_545 ();
 FILLCELL_X32 FILLER_333_577 ();
 FILLCELL_X32 FILLER_333_609 ();
 FILLCELL_X32 FILLER_333_641 ();
 FILLCELL_X32 FILLER_333_673 ();
 FILLCELL_X32 FILLER_333_705 ();
 FILLCELL_X32 FILLER_333_737 ();
 FILLCELL_X32 FILLER_333_769 ();
 FILLCELL_X32 FILLER_333_801 ();
 FILLCELL_X32 FILLER_333_833 ();
 FILLCELL_X32 FILLER_333_865 ();
 FILLCELL_X32 FILLER_333_897 ();
 FILLCELL_X32 FILLER_333_929 ();
 FILLCELL_X32 FILLER_333_961 ();
 FILLCELL_X32 FILLER_333_993 ();
 FILLCELL_X32 FILLER_333_1025 ();
 FILLCELL_X32 FILLER_333_1057 ();
 FILLCELL_X32 FILLER_333_1089 ();
 FILLCELL_X32 FILLER_333_1121 ();
 FILLCELL_X32 FILLER_333_1153 ();
 FILLCELL_X32 FILLER_333_1185 ();
 FILLCELL_X32 FILLER_333_1217 ();
 FILLCELL_X8 FILLER_333_1249 ();
 FILLCELL_X4 FILLER_333_1257 ();
 FILLCELL_X2 FILLER_333_1261 ();
 FILLCELL_X32 FILLER_333_1264 ();
 FILLCELL_X32 FILLER_333_1296 ();
 FILLCELL_X32 FILLER_333_1328 ();
 FILLCELL_X32 FILLER_333_1360 ();
 FILLCELL_X32 FILLER_333_1392 ();
 FILLCELL_X32 FILLER_333_1424 ();
 FILLCELL_X32 FILLER_333_1456 ();
 FILLCELL_X32 FILLER_333_1488 ();
 FILLCELL_X32 FILLER_333_1520 ();
 FILLCELL_X32 FILLER_333_1552 ();
 FILLCELL_X32 FILLER_333_1584 ();
 FILLCELL_X32 FILLER_333_1616 ();
 FILLCELL_X32 FILLER_333_1648 ();
 FILLCELL_X32 FILLER_333_1680 ();
 FILLCELL_X32 FILLER_333_1712 ();
 FILLCELL_X32 FILLER_333_1744 ();
 FILLCELL_X32 FILLER_333_1776 ();
 FILLCELL_X32 FILLER_333_1808 ();
 FILLCELL_X32 FILLER_333_1840 ();
 FILLCELL_X32 FILLER_333_1872 ();
 FILLCELL_X32 FILLER_333_1904 ();
 FILLCELL_X32 FILLER_333_1936 ();
 FILLCELL_X32 FILLER_333_1968 ();
 FILLCELL_X32 FILLER_333_2000 ();
 FILLCELL_X32 FILLER_333_2032 ();
 FILLCELL_X32 FILLER_333_2064 ();
 FILLCELL_X32 FILLER_333_2096 ();
 FILLCELL_X32 FILLER_333_2128 ();
 FILLCELL_X32 FILLER_333_2160 ();
 FILLCELL_X32 FILLER_333_2192 ();
 FILLCELL_X32 FILLER_333_2224 ();
 FILLCELL_X32 FILLER_333_2256 ();
 FILLCELL_X32 FILLER_333_2288 ();
 FILLCELL_X32 FILLER_333_2320 ();
 FILLCELL_X32 FILLER_333_2352 ();
 FILLCELL_X32 FILLER_333_2384 ();
 FILLCELL_X32 FILLER_333_2416 ();
 FILLCELL_X32 FILLER_333_2448 ();
 FILLCELL_X32 FILLER_333_2480 ();
 FILLCELL_X8 FILLER_333_2512 ();
 FILLCELL_X4 FILLER_333_2520 ();
 FILLCELL_X2 FILLER_333_2524 ();
 FILLCELL_X32 FILLER_333_2527 ();
 FILLCELL_X32 FILLER_333_2559 ();
 FILLCELL_X32 FILLER_333_2591 ();
 FILLCELL_X32 FILLER_333_2623 ();
 FILLCELL_X32 FILLER_333_2655 ();
 FILLCELL_X32 FILLER_333_2687 ();
 FILLCELL_X32 FILLER_333_2719 ();
 FILLCELL_X32 FILLER_333_2751 ();
 FILLCELL_X32 FILLER_333_2783 ();
 FILLCELL_X32 FILLER_333_2815 ();
 FILLCELL_X32 FILLER_333_2847 ();
 FILLCELL_X32 FILLER_333_2879 ();
 FILLCELL_X32 FILLER_333_2911 ();
 FILLCELL_X32 FILLER_333_2943 ();
 FILLCELL_X32 FILLER_333_2975 ();
 FILLCELL_X32 FILLER_333_3007 ();
 FILLCELL_X32 FILLER_333_3039 ();
 FILLCELL_X32 FILLER_333_3071 ();
 FILLCELL_X32 FILLER_333_3103 ();
 FILLCELL_X32 FILLER_333_3135 ();
 FILLCELL_X32 FILLER_333_3167 ();
 FILLCELL_X32 FILLER_333_3199 ();
 FILLCELL_X32 FILLER_333_3231 ();
 FILLCELL_X32 FILLER_333_3263 ();
 FILLCELL_X32 FILLER_333_3295 ();
 FILLCELL_X32 FILLER_333_3327 ();
 FILLCELL_X32 FILLER_333_3359 ();
 FILLCELL_X32 FILLER_333_3391 ();
 FILLCELL_X32 FILLER_333_3423 ();
 FILLCELL_X32 FILLER_333_3455 ();
 FILLCELL_X32 FILLER_333_3487 ();
 FILLCELL_X32 FILLER_333_3519 ();
 FILLCELL_X32 FILLER_333_3551 ();
 FILLCELL_X32 FILLER_333_3583 ();
 FILLCELL_X32 FILLER_333_3615 ();
 FILLCELL_X32 FILLER_333_3647 ();
 FILLCELL_X32 FILLER_333_3679 ();
 FILLCELL_X16 FILLER_333_3711 ();
 FILLCELL_X8 FILLER_333_3727 ();
 FILLCELL_X2 FILLER_333_3735 ();
 FILLCELL_X1 FILLER_333_3737 ();
 FILLCELL_X32 FILLER_334_1 ();
 FILLCELL_X32 FILLER_334_33 ();
 FILLCELL_X32 FILLER_334_65 ();
 FILLCELL_X32 FILLER_334_97 ();
 FILLCELL_X32 FILLER_334_129 ();
 FILLCELL_X32 FILLER_334_161 ();
 FILLCELL_X32 FILLER_334_193 ();
 FILLCELL_X32 FILLER_334_225 ();
 FILLCELL_X32 FILLER_334_257 ();
 FILLCELL_X32 FILLER_334_289 ();
 FILLCELL_X32 FILLER_334_321 ();
 FILLCELL_X32 FILLER_334_353 ();
 FILLCELL_X32 FILLER_334_385 ();
 FILLCELL_X32 FILLER_334_417 ();
 FILLCELL_X32 FILLER_334_449 ();
 FILLCELL_X32 FILLER_334_481 ();
 FILLCELL_X32 FILLER_334_513 ();
 FILLCELL_X32 FILLER_334_545 ();
 FILLCELL_X32 FILLER_334_577 ();
 FILLCELL_X16 FILLER_334_609 ();
 FILLCELL_X4 FILLER_334_625 ();
 FILLCELL_X2 FILLER_334_629 ();
 FILLCELL_X32 FILLER_334_632 ();
 FILLCELL_X32 FILLER_334_664 ();
 FILLCELL_X32 FILLER_334_696 ();
 FILLCELL_X32 FILLER_334_728 ();
 FILLCELL_X32 FILLER_334_760 ();
 FILLCELL_X32 FILLER_334_792 ();
 FILLCELL_X32 FILLER_334_824 ();
 FILLCELL_X32 FILLER_334_856 ();
 FILLCELL_X32 FILLER_334_888 ();
 FILLCELL_X32 FILLER_334_920 ();
 FILLCELL_X32 FILLER_334_952 ();
 FILLCELL_X32 FILLER_334_984 ();
 FILLCELL_X32 FILLER_334_1016 ();
 FILLCELL_X32 FILLER_334_1048 ();
 FILLCELL_X32 FILLER_334_1080 ();
 FILLCELL_X32 FILLER_334_1112 ();
 FILLCELL_X32 FILLER_334_1144 ();
 FILLCELL_X32 FILLER_334_1176 ();
 FILLCELL_X32 FILLER_334_1208 ();
 FILLCELL_X32 FILLER_334_1240 ();
 FILLCELL_X32 FILLER_334_1272 ();
 FILLCELL_X32 FILLER_334_1304 ();
 FILLCELL_X32 FILLER_334_1336 ();
 FILLCELL_X32 FILLER_334_1368 ();
 FILLCELL_X32 FILLER_334_1400 ();
 FILLCELL_X32 FILLER_334_1432 ();
 FILLCELL_X32 FILLER_334_1464 ();
 FILLCELL_X32 FILLER_334_1496 ();
 FILLCELL_X32 FILLER_334_1528 ();
 FILLCELL_X32 FILLER_334_1560 ();
 FILLCELL_X32 FILLER_334_1592 ();
 FILLCELL_X32 FILLER_334_1624 ();
 FILLCELL_X32 FILLER_334_1656 ();
 FILLCELL_X32 FILLER_334_1688 ();
 FILLCELL_X32 FILLER_334_1720 ();
 FILLCELL_X32 FILLER_334_1752 ();
 FILLCELL_X32 FILLER_334_1784 ();
 FILLCELL_X32 FILLER_334_1816 ();
 FILLCELL_X32 FILLER_334_1848 ();
 FILLCELL_X8 FILLER_334_1880 ();
 FILLCELL_X4 FILLER_334_1888 ();
 FILLCELL_X2 FILLER_334_1892 ();
 FILLCELL_X32 FILLER_334_1895 ();
 FILLCELL_X32 FILLER_334_1927 ();
 FILLCELL_X32 FILLER_334_1959 ();
 FILLCELL_X32 FILLER_334_1991 ();
 FILLCELL_X32 FILLER_334_2023 ();
 FILLCELL_X32 FILLER_334_2055 ();
 FILLCELL_X32 FILLER_334_2087 ();
 FILLCELL_X32 FILLER_334_2119 ();
 FILLCELL_X32 FILLER_334_2151 ();
 FILLCELL_X32 FILLER_334_2183 ();
 FILLCELL_X32 FILLER_334_2215 ();
 FILLCELL_X32 FILLER_334_2247 ();
 FILLCELL_X32 FILLER_334_2279 ();
 FILLCELL_X32 FILLER_334_2311 ();
 FILLCELL_X32 FILLER_334_2343 ();
 FILLCELL_X32 FILLER_334_2375 ();
 FILLCELL_X32 FILLER_334_2407 ();
 FILLCELL_X32 FILLER_334_2439 ();
 FILLCELL_X32 FILLER_334_2471 ();
 FILLCELL_X32 FILLER_334_2503 ();
 FILLCELL_X32 FILLER_334_2535 ();
 FILLCELL_X32 FILLER_334_2567 ();
 FILLCELL_X32 FILLER_334_2599 ();
 FILLCELL_X32 FILLER_334_2631 ();
 FILLCELL_X32 FILLER_334_2663 ();
 FILLCELL_X32 FILLER_334_2695 ();
 FILLCELL_X32 FILLER_334_2727 ();
 FILLCELL_X32 FILLER_334_2759 ();
 FILLCELL_X32 FILLER_334_2791 ();
 FILLCELL_X32 FILLER_334_2823 ();
 FILLCELL_X32 FILLER_334_2855 ();
 FILLCELL_X32 FILLER_334_2887 ();
 FILLCELL_X32 FILLER_334_2919 ();
 FILLCELL_X32 FILLER_334_2951 ();
 FILLCELL_X32 FILLER_334_2983 ();
 FILLCELL_X32 FILLER_334_3015 ();
 FILLCELL_X32 FILLER_334_3047 ();
 FILLCELL_X32 FILLER_334_3079 ();
 FILLCELL_X32 FILLER_334_3111 ();
 FILLCELL_X8 FILLER_334_3143 ();
 FILLCELL_X4 FILLER_334_3151 ();
 FILLCELL_X2 FILLER_334_3155 ();
 FILLCELL_X32 FILLER_334_3158 ();
 FILLCELL_X32 FILLER_334_3190 ();
 FILLCELL_X32 FILLER_334_3222 ();
 FILLCELL_X32 FILLER_334_3254 ();
 FILLCELL_X32 FILLER_334_3286 ();
 FILLCELL_X32 FILLER_334_3318 ();
 FILLCELL_X32 FILLER_334_3350 ();
 FILLCELL_X32 FILLER_334_3382 ();
 FILLCELL_X32 FILLER_334_3414 ();
 FILLCELL_X32 FILLER_334_3446 ();
 FILLCELL_X32 FILLER_334_3478 ();
 FILLCELL_X32 FILLER_334_3510 ();
 FILLCELL_X32 FILLER_334_3542 ();
 FILLCELL_X32 FILLER_334_3574 ();
 FILLCELL_X32 FILLER_334_3606 ();
 FILLCELL_X32 FILLER_334_3638 ();
 FILLCELL_X32 FILLER_334_3670 ();
 FILLCELL_X32 FILLER_334_3702 ();
 FILLCELL_X4 FILLER_334_3734 ();
 FILLCELL_X32 FILLER_335_1 ();
 FILLCELL_X32 FILLER_335_33 ();
 FILLCELL_X32 FILLER_335_65 ();
 FILLCELL_X32 FILLER_335_97 ();
 FILLCELL_X32 FILLER_335_129 ();
 FILLCELL_X32 FILLER_335_161 ();
 FILLCELL_X32 FILLER_335_193 ();
 FILLCELL_X32 FILLER_335_225 ();
 FILLCELL_X32 FILLER_335_257 ();
 FILLCELL_X32 FILLER_335_289 ();
 FILLCELL_X32 FILLER_335_321 ();
 FILLCELL_X32 FILLER_335_353 ();
 FILLCELL_X32 FILLER_335_385 ();
 FILLCELL_X32 FILLER_335_417 ();
 FILLCELL_X32 FILLER_335_449 ();
 FILLCELL_X32 FILLER_335_481 ();
 FILLCELL_X32 FILLER_335_513 ();
 FILLCELL_X32 FILLER_335_545 ();
 FILLCELL_X32 FILLER_335_577 ();
 FILLCELL_X32 FILLER_335_609 ();
 FILLCELL_X32 FILLER_335_641 ();
 FILLCELL_X32 FILLER_335_673 ();
 FILLCELL_X32 FILLER_335_705 ();
 FILLCELL_X32 FILLER_335_737 ();
 FILLCELL_X32 FILLER_335_769 ();
 FILLCELL_X32 FILLER_335_801 ();
 FILLCELL_X32 FILLER_335_833 ();
 FILLCELL_X32 FILLER_335_865 ();
 FILLCELL_X32 FILLER_335_897 ();
 FILLCELL_X32 FILLER_335_929 ();
 FILLCELL_X32 FILLER_335_961 ();
 FILLCELL_X32 FILLER_335_993 ();
 FILLCELL_X32 FILLER_335_1025 ();
 FILLCELL_X32 FILLER_335_1057 ();
 FILLCELL_X32 FILLER_335_1089 ();
 FILLCELL_X32 FILLER_335_1121 ();
 FILLCELL_X32 FILLER_335_1153 ();
 FILLCELL_X32 FILLER_335_1185 ();
 FILLCELL_X32 FILLER_335_1217 ();
 FILLCELL_X8 FILLER_335_1249 ();
 FILLCELL_X4 FILLER_335_1257 ();
 FILLCELL_X2 FILLER_335_1261 ();
 FILLCELL_X32 FILLER_335_1264 ();
 FILLCELL_X32 FILLER_335_1296 ();
 FILLCELL_X32 FILLER_335_1328 ();
 FILLCELL_X32 FILLER_335_1360 ();
 FILLCELL_X32 FILLER_335_1392 ();
 FILLCELL_X32 FILLER_335_1424 ();
 FILLCELL_X32 FILLER_335_1456 ();
 FILLCELL_X32 FILLER_335_1488 ();
 FILLCELL_X32 FILLER_335_1520 ();
 FILLCELL_X32 FILLER_335_1552 ();
 FILLCELL_X32 FILLER_335_1584 ();
 FILLCELL_X32 FILLER_335_1616 ();
 FILLCELL_X32 FILLER_335_1648 ();
 FILLCELL_X32 FILLER_335_1680 ();
 FILLCELL_X32 FILLER_335_1712 ();
 FILLCELL_X32 FILLER_335_1744 ();
 FILLCELL_X32 FILLER_335_1776 ();
 FILLCELL_X32 FILLER_335_1808 ();
 FILLCELL_X32 FILLER_335_1840 ();
 FILLCELL_X32 FILLER_335_1872 ();
 FILLCELL_X32 FILLER_335_1904 ();
 FILLCELL_X32 FILLER_335_1936 ();
 FILLCELL_X32 FILLER_335_1968 ();
 FILLCELL_X32 FILLER_335_2000 ();
 FILLCELL_X32 FILLER_335_2032 ();
 FILLCELL_X32 FILLER_335_2064 ();
 FILLCELL_X32 FILLER_335_2096 ();
 FILLCELL_X32 FILLER_335_2128 ();
 FILLCELL_X32 FILLER_335_2160 ();
 FILLCELL_X32 FILLER_335_2192 ();
 FILLCELL_X32 FILLER_335_2224 ();
 FILLCELL_X32 FILLER_335_2256 ();
 FILLCELL_X32 FILLER_335_2288 ();
 FILLCELL_X32 FILLER_335_2320 ();
 FILLCELL_X32 FILLER_335_2352 ();
 FILLCELL_X32 FILLER_335_2384 ();
 FILLCELL_X32 FILLER_335_2416 ();
 FILLCELL_X32 FILLER_335_2448 ();
 FILLCELL_X32 FILLER_335_2480 ();
 FILLCELL_X8 FILLER_335_2512 ();
 FILLCELL_X4 FILLER_335_2520 ();
 FILLCELL_X2 FILLER_335_2524 ();
 FILLCELL_X32 FILLER_335_2527 ();
 FILLCELL_X32 FILLER_335_2559 ();
 FILLCELL_X32 FILLER_335_2591 ();
 FILLCELL_X32 FILLER_335_2623 ();
 FILLCELL_X32 FILLER_335_2655 ();
 FILLCELL_X32 FILLER_335_2687 ();
 FILLCELL_X32 FILLER_335_2719 ();
 FILLCELL_X32 FILLER_335_2751 ();
 FILLCELL_X32 FILLER_335_2783 ();
 FILLCELL_X32 FILLER_335_2815 ();
 FILLCELL_X32 FILLER_335_2847 ();
 FILLCELL_X32 FILLER_335_2879 ();
 FILLCELL_X32 FILLER_335_2911 ();
 FILLCELL_X32 FILLER_335_2943 ();
 FILLCELL_X32 FILLER_335_2975 ();
 FILLCELL_X32 FILLER_335_3007 ();
 FILLCELL_X32 FILLER_335_3039 ();
 FILLCELL_X32 FILLER_335_3071 ();
 FILLCELL_X32 FILLER_335_3103 ();
 FILLCELL_X32 FILLER_335_3135 ();
 FILLCELL_X32 FILLER_335_3167 ();
 FILLCELL_X32 FILLER_335_3199 ();
 FILLCELL_X32 FILLER_335_3231 ();
 FILLCELL_X32 FILLER_335_3263 ();
 FILLCELL_X32 FILLER_335_3295 ();
 FILLCELL_X32 FILLER_335_3327 ();
 FILLCELL_X32 FILLER_335_3359 ();
 FILLCELL_X32 FILLER_335_3391 ();
 FILLCELL_X32 FILLER_335_3423 ();
 FILLCELL_X32 FILLER_335_3455 ();
 FILLCELL_X32 FILLER_335_3487 ();
 FILLCELL_X32 FILLER_335_3519 ();
 FILLCELL_X32 FILLER_335_3551 ();
 FILLCELL_X32 FILLER_335_3583 ();
 FILLCELL_X32 FILLER_335_3615 ();
 FILLCELL_X32 FILLER_335_3647 ();
 FILLCELL_X32 FILLER_335_3679 ();
 FILLCELL_X16 FILLER_335_3711 ();
 FILLCELL_X8 FILLER_335_3727 ();
 FILLCELL_X2 FILLER_335_3735 ();
 FILLCELL_X1 FILLER_335_3737 ();
 FILLCELL_X32 FILLER_336_1 ();
 FILLCELL_X32 FILLER_336_33 ();
 FILLCELL_X32 FILLER_336_65 ();
 FILLCELL_X32 FILLER_336_97 ();
 FILLCELL_X32 FILLER_336_129 ();
 FILLCELL_X32 FILLER_336_161 ();
 FILLCELL_X32 FILLER_336_193 ();
 FILLCELL_X32 FILLER_336_225 ();
 FILLCELL_X32 FILLER_336_257 ();
 FILLCELL_X32 FILLER_336_289 ();
 FILLCELL_X32 FILLER_336_321 ();
 FILLCELL_X32 FILLER_336_353 ();
 FILLCELL_X32 FILLER_336_385 ();
 FILLCELL_X32 FILLER_336_417 ();
 FILLCELL_X32 FILLER_336_449 ();
 FILLCELL_X32 FILLER_336_481 ();
 FILLCELL_X32 FILLER_336_513 ();
 FILLCELL_X32 FILLER_336_545 ();
 FILLCELL_X32 FILLER_336_577 ();
 FILLCELL_X16 FILLER_336_609 ();
 FILLCELL_X4 FILLER_336_625 ();
 FILLCELL_X2 FILLER_336_629 ();
 FILLCELL_X32 FILLER_336_632 ();
 FILLCELL_X32 FILLER_336_664 ();
 FILLCELL_X32 FILLER_336_696 ();
 FILLCELL_X32 FILLER_336_728 ();
 FILLCELL_X32 FILLER_336_760 ();
 FILLCELL_X32 FILLER_336_792 ();
 FILLCELL_X32 FILLER_336_824 ();
 FILLCELL_X32 FILLER_336_856 ();
 FILLCELL_X32 FILLER_336_888 ();
 FILLCELL_X32 FILLER_336_920 ();
 FILLCELL_X32 FILLER_336_952 ();
 FILLCELL_X32 FILLER_336_984 ();
 FILLCELL_X32 FILLER_336_1016 ();
 FILLCELL_X32 FILLER_336_1048 ();
 FILLCELL_X32 FILLER_336_1080 ();
 FILLCELL_X32 FILLER_336_1112 ();
 FILLCELL_X32 FILLER_336_1144 ();
 FILLCELL_X32 FILLER_336_1176 ();
 FILLCELL_X32 FILLER_336_1208 ();
 FILLCELL_X32 FILLER_336_1240 ();
 FILLCELL_X32 FILLER_336_1272 ();
 FILLCELL_X32 FILLER_336_1304 ();
 FILLCELL_X32 FILLER_336_1336 ();
 FILLCELL_X32 FILLER_336_1368 ();
 FILLCELL_X32 FILLER_336_1400 ();
 FILLCELL_X32 FILLER_336_1432 ();
 FILLCELL_X32 FILLER_336_1464 ();
 FILLCELL_X32 FILLER_336_1496 ();
 FILLCELL_X32 FILLER_336_1528 ();
 FILLCELL_X32 FILLER_336_1560 ();
 FILLCELL_X32 FILLER_336_1592 ();
 FILLCELL_X32 FILLER_336_1624 ();
 FILLCELL_X32 FILLER_336_1656 ();
 FILLCELL_X32 FILLER_336_1688 ();
 FILLCELL_X32 FILLER_336_1720 ();
 FILLCELL_X32 FILLER_336_1752 ();
 FILLCELL_X32 FILLER_336_1784 ();
 FILLCELL_X32 FILLER_336_1816 ();
 FILLCELL_X32 FILLER_336_1848 ();
 FILLCELL_X8 FILLER_336_1880 ();
 FILLCELL_X4 FILLER_336_1888 ();
 FILLCELL_X2 FILLER_336_1892 ();
 FILLCELL_X32 FILLER_336_1895 ();
 FILLCELL_X32 FILLER_336_1927 ();
 FILLCELL_X32 FILLER_336_1959 ();
 FILLCELL_X32 FILLER_336_1991 ();
 FILLCELL_X32 FILLER_336_2023 ();
 FILLCELL_X32 FILLER_336_2055 ();
 FILLCELL_X32 FILLER_336_2087 ();
 FILLCELL_X32 FILLER_336_2119 ();
 FILLCELL_X32 FILLER_336_2151 ();
 FILLCELL_X32 FILLER_336_2183 ();
 FILLCELL_X32 FILLER_336_2215 ();
 FILLCELL_X32 FILLER_336_2247 ();
 FILLCELL_X32 FILLER_336_2279 ();
 FILLCELL_X32 FILLER_336_2311 ();
 FILLCELL_X32 FILLER_336_2343 ();
 FILLCELL_X32 FILLER_336_2375 ();
 FILLCELL_X32 FILLER_336_2407 ();
 FILLCELL_X32 FILLER_336_2439 ();
 FILLCELL_X32 FILLER_336_2471 ();
 FILLCELL_X32 FILLER_336_2503 ();
 FILLCELL_X32 FILLER_336_2535 ();
 FILLCELL_X32 FILLER_336_2567 ();
 FILLCELL_X32 FILLER_336_2599 ();
 FILLCELL_X32 FILLER_336_2631 ();
 FILLCELL_X32 FILLER_336_2663 ();
 FILLCELL_X32 FILLER_336_2695 ();
 FILLCELL_X32 FILLER_336_2727 ();
 FILLCELL_X32 FILLER_336_2759 ();
 FILLCELL_X32 FILLER_336_2791 ();
 FILLCELL_X32 FILLER_336_2823 ();
 FILLCELL_X32 FILLER_336_2855 ();
 FILLCELL_X32 FILLER_336_2887 ();
 FILLCELL_X32 FILLER_336_2919 ();
 FILLCELL_X32 FILLER_336_2951 ();
 FILLCELL_X32 FILLER_336_2983 ();
 FILLCELL_X32 FILLER_336_3015 ();
 FILLCELL_X32 FILLER_336_3047 ();
 FILLCELL_X32 FILLER_336_3079 ();
 FILLCELL_X32 FILLER_336_3111 ();
 FILLCELL_X8 FILLER_336_3143 ();
 FILLCELL_X4 FILLER_336_3151 ();
 FILLCELL_X2 FILLER_336_3155 ();
 FILLCELL_X32 FILLER_336_3158 ();
 FILLCELL_X32 FILLER_336_3190 ();
 FILLCELL_X32 FILLER_336_3222 ();
 FILLCELL_X32 FILLER_336_3254 ();
 FILLCELL_X32 FILLER_336_3286 ();
 FILLCELL_X32 FILLER_336_3318 ();
 FILLCELL_X32 FILLER_336_3350 ();
 FILLCELL_X32 FILLER_336_3382 ();
 FILLCELL_X32 FILLER_336_3414 ();
 FILLCELL_X32 FILLER_336_3446 ();
 FILLCELL_X32 FILLER_336_3478 ();
 FILLCELL_X32 FILLER_336_3510 ();
 FILLCELL_X32 FILLER_336_3542 ();
 FILLCELL_X32 FILLER_336_3574 ();
 FILLCELL_X32 FILLER_336_3606 ();
 FILLCELL_X32 FILLER_336_3638 ();
 FILLCELL_X32 FILLER_336_3670 ();
 FILLCELL_X32 FILLER_336_3702 ();
 FILLCELL_X4 FILLER_336_3734 ();
 FILLCELL_X32 FILLER_337_1 ();
 FILLCELL_X32 FILLER_337_33 ();
 FILLCELL_X32 FILLER_337_65 ();
 FILLCELL_X32 FILLER_337_97 ();
 FILLCELL_X32 FILLER_337_129 ();
 FILLCELL_X32 FILLER_337_161 ();
 FILLCELL_X32 FILLER_337_193 ();
 FILLCELL_X32 FILLER_337_225 ();
 FILLCELL_X32 FILLER_337_257 ();
 FILLCELL_X32 FILLER_337_289 ();
 FILLCELL_X32 FILLER_337_321 ();
 FILLCELL_X32 FILLER_337_353 ();
 FILLCELL_X32 FILLER_337_385 ();
 FILLCELL_X32 FILLER_337_417 ();
 FILLCELL_X32 FILLER_337_449 ();
 FILLCELL_X32 FILLER_337_481 ();
 FILLCELL_X32 FILLER_337_513 ();
 FILLCELL_X32 FILLER_337_545 ();
 FILLCELL_X32 FILLER_337_577 ();
 FILLCELL_X32 FILLER_337_609 ();
 FILLCELL_X32 FILLER_337_641 ();
 FILLCELL_X32 FILLER_337_673 ();
 FILLCELL_X32 FILLER_337_705 ();
 FILLCELL_X32 FILLER_337_737 ();
 FILLCELL_X32 FILLER_337_769 ();
 FILLCELL_X32 FILLER_337_801 ();
 FILLCELL_X32 FILLER_337_833 ();
 FILLCELL_X32 FILLER_337_865 ();
 FILLCELL_X32 FILLER_337_897 ();
 FILLCELL_X32 FILLER_337_929 ();
 FILLCELL_X32 FILLER_337_961 ();
 FILLCELL_X32 FILLER_337_993 ();
 FILLCELL_X32 FILLER_337_1025 ();
 FILLCELL_X32 FILLER_337_1057 ();
 FILLCELL_X32 FILLER_337_1089 ();
 FILLCELL_X32 FILLER_337_1121 ();
 FILLCELL_X32 FILLER_337_1153 ();
 FILLCELL_X32 FILLER_337_1185 ();
 FILLCELL_X32 FILLER_337_1217 ();
 FILLCELL_X8 FILLER_337_1249 ();
 FILLCELL_X4 FILLER_337_1257 ();
 FILLCELL_X2 FILLER_337_1261 ();
 FILLCELL_X32 FILLER_337_1264 ();
 FILLCELL_X32 FILLER_337_1296 ();
 FILLCELL_X32 FILLER_337_1328 ();
 FILLCELL_X32 FILLER_337_1360 ();
 FILLCELL_X32 FILLER_337_1392 ();
 FILLCELL_X32 FILLER_337_1424 ();
 FILLCELL_X32 FILLER_337_1456 ();
 FILLCELL_X32 FILLER_337_1488 ();
 FILLCELL_X32 FILLER_337_1520 ();
 FILLCELL_X32 FILLER_337_1552 ();
 FILLCELL_X32 FILLER_337_1584 ();
 FILLCELL_X32 FILLER_337_1616 ();
 FILLCELL_X32 FILLER_337_1648 ();
 FILLCELL_X32 FILLER_337_1680 ();
 FILLCELL_X32 FILLER_337_1712 ();
 FILLCELL_X32 FILLER_337_1744 ();
 FILLCELL_X32 FILLER_337_1776 ();
 FILLCELL_X32 FILLER_337_1808 ();
 FILLCELL_X32 FILLER_337_1840 ();
 FILLCELL_X32 FILLER_337_1872 ();
 FILLCELL_X32 FILLER_337_1904 ();
 FILLCELL_X32 FILLER_337_1936 ();
 FILLCELL_X32 FILLER_337_1968 ();
 FILLCELL_X32 FILLER_337_2000 ();
 FILLCELL_X32 FILLER_337_2032 ();
 FILLCELL_X32 FILLER_337_2064 ();
 FILLCELL_X32 FILLER_337_2096 ();
 FILLCELL_X32 FILLER_337_2128 ();
 FILLCELL_X32 FILLER_337_2160 ();
 FILLCELL_X32 FILLER_337_2192 ();
 FILLCELL_X32 FILLER_337_2224 ();
 FILLCELL_X32 FILLER_337_2256 ();
 FILLCELL_X32 FILLER_337_2288 ();
 FILLCELL_X32 FILLER_337_2320 ();
 FILLCELL_X32 FILLER_337_2352 ();
 FILLCELL_X32 FILLER_337_2384 ();
 FILLCELL_X32 FILLER_337_2416 ();
 FILLCELL_X32 FILLER_337_2448 ();
 FILLCELL_X32 FILLER_337_2480 ();
 FILLCELL_X8 FILLER_337_2512 ();
 FILLCELL_X4 FILLER_337_2520 ();
 FILLCELL_X2 FILLER_337_2524 ();
 FILLCELL_X32 FILLER_337_2527 ();
 FILLCELL_X32 FILLER_337_2559 ();
 FILLCELL_X32 FILLER_337_2591 ();
 FILLCELL_X32 FILLER_337_2623 ();
 FILLCELL_X32 FILLER_337_2655 ();
 FILLCELL_X32 FILLER_337_2687 ();
 FILLCELL_X32 FILLER_337_2719 ();
 FILLCELL_X32 FILLER_337_2751 ();
 FILLCELL_X32 FILLER_337_2783 ();
 FILLCELL_X32 FILLER_337_2815 ();
 FILLCELL_X32 FILLER_337_2847 ();
 FILLCELL_X32 FILLER_337_2879 ();
 FILLCELL_X32 FILLER_337_2911 ();
 FILLCELL_X32 FILLER_337_2943 ();
 FILLCELL_X32 FILLER_337_2975 ();
 FILLCELL_X32 FILLER_337_3007 ();
 FILLCELL_X32 FILLER_337_3039 ();
 FILLCELL_X32 FILLER_337_3071 ();
 FILLCELL_X32 FILLER_337_3103 ();
 FILLCELL_X32 FILLER_337_3135 ();
 FILLCELL_X32 FILLER_337_3167 ();
 FILLCELL_X32 FILLER_337_3199 ();
 FILLCELL_X32 FILLER_337_3231 ();
 FILLCELL_X32 FILLER_337_3263 ();
 FILLCELL_X32 FILLER_337_3295 ();
 FILLCELL_X32 FILLER_337_3327 ();
 FILLCELL_X32 FILLER_337_3359 ();
 FILLCELL_X32 FILLER_337_3391 ();
 FILLCELL_X32 FILLER_337_3423 ();
 FILLCELL_X32 FILLER_337_3455 ();
 FILLCELL_X32 FILLER_337_3487 ();
 FILLCELL_X32 FILLER_337_3519 ();
 FILLCELL_X32 FILLER_337_3551 ();
 FILLCELL_X32 FILLER_337_3583 ();
 FILLCELL_X32 FILLER_337_3615 ();
 FILLCELL_X32 FILLER_337_3647 ();
 FILLCELL_X32 FILLER_337_3679 ();
 FILLCELL_X16 FILLER_337_3711 ();
 FILLCELL_X8 FILLER_337_3727 ();
 FILLCELL_X2 FILLER_337_3735 ();
 FILLCELL_X1 FILLER_337_3737 ();
 FILLCELL_X32 FILLER_338_1 ();
 FILLCELL_X32 FILLER_338_33 ();
 FILLCELL_X32 FILLER_338_65 ();
 FILLCELL_X32 FILLER_338_97 ();
 FILLCELL_X32 FILLER_338_129 ();
 FILLCELL_X32 FILLER_338_161 ();
 FILLCELL_X32 FILLER_338_193 ();
 FILLCELL_X32 FILLER_338_225 ();
 FILLCELL_X32 FILLER_338_257 ();
 FILLCELL_X32 FILLER_338_289 ();
 FILLCELL_X32 FILLER_338_321 ();
 FILLCELL_X32 FILLER_338_353 ();
 FILLCELL_X32 FILLER_338_385 ();
 FILLCELL_X32 FILLER_338_417 ();
 FILLCELL_X32 FILLER_338_449 ();
 FILLCELL_X32 FILLER_338_481 ();
 FILLCELL_X32 FILLER_338_513 ();
 FILLCELL_X32 FILLER_338_545 ();
 FILLCELL_X32 FILLER_338_577 ();
 FILLCELL_X16 FILLER_338_609 ();
 FILLCELL_X4 FILLER_338_625 ();
 FILLCELL_X2 FILLER_338_629 ();
 FILLCELL_X32 FILLER_338_632 ();
 FILLCELL_X32 FILLER_338_664 ();
 FILLCELL_X32 FILLER_338_696 ();
 FILLCELL_X32 FILLER_338_728 ();
 FILLCELL_X32 FILLER_338_760 ();
 FILLCELL_X32 FILLER_338_792 ();
 FILLCELL_X32 FILLER_338_824 ();
 FILLCELL_X32 FILLER_338_856 ();
 FILLCELL_X32 FILLER_338_888 ();
 FILLCELL_X32 FILLER_338_920 ();
 FILLCELL_X32 FILLER_338_952 ();
 FILLCELL_X32 FILLER_338_984 ();
 FILLCELL_X32 FILLER_338_1016 ();
 FILLCELL_X32 FILLER_338_1048 ();
 FILLCELL_X32 FILLER_338_1080 ();
 FILLCELL_X32 FILLER_338_1112 ();
 FILLCELL_X32 FILLER_338_1144 ();
 FILLCELL_X32 FILLER_338_1176 ();
 FILLCELL_X32 FILLER_338_1208 ();
 FILLCELL_X32 FILLER_338_1240 ();
 FILLCELL_X32 FILLER_338_1272 ();
 FILLCELL_X32 FILLER_338_1304 ();
 FILLCELL_X32 FILLER_338_1336 ();
 FILLCELL_X32 FILLER_338_1368 ();
 FILLCELL_X32 FILLER_338_1400 ();
 FILLCELL_X32 FILLER_338_1432 ();
 FILLCELL_X32 FILLER_338_1464 ();
 FILLCELL_X32 FILLER_338_1496 ();
 FILLCELL_X32 FILLER_338_1528 ();
 FILLCELL_X32 FILLER_338_1560 ();
 FILLCELL_X32 FILLER_338_1592 ();
 FILLCELL_X32 FILLER_338_1624 ();
 FILLCELL_X32 FILLER_338_1656 ();
 FILLCELL_X32 FILLER_338_1688 ();
 FILLCELL_X32 FILLER_338_1720 ();
 FILLCELL_X32 FILLER_338_1752 ();
 FILLCELL_X32 FILLER_338_1784 ();
 FILLCELL_X32 FILLER_338_1816 ();
 FILLCELL_X32 FILLER_338_1848 ();
 FILLCELL_X8 FILLER_338_1880 ();
 FILLCELL_X4 FILLER_338_1888 ();
 FILLCELL_X2 FILLER_338_1892 ();
 FILLCELL_X32 FILLER_338_1895 ();
 FILLCELL_X32 FILLER_338_1927 ();
 FILLCELL_X32 FILLER_338_1959 ();
 FILLCELL_X32 FILLER_338_1991 ();
 FILLCELL_X32 FILLER_338_2023 ();
 FILLCELL_X32 FILLER_338_2055 ();
 FILLCELL_X32 FILLER_338_2087 ();
 FILLCELL_X32 FILLER_338_2119 ();
 FILLCELL_X32 FILLER_338_2151 ();
 FILLCELL_X32 FILLER_338_2183 ();
 FILLCELL_X32 FILLER_338_2215 ();
 FILLCELL_X32 FILLER_338_2247 ();
 FILLCELL_X32 FILLER_338_2279 ();
 FILLCELL_X32 FILLER_338_2311 ();
 FILLCELL_X32 FILLER_338_2343 ();
 FILLCELL_X32 FILLER_338_2375 ();
 FILLCELL_X32 FILLER_338_2407 ();
 FILLCELL_X32 FILLER_338_2439 ();
 FILLCELL_X32 FILLER_338_2471 ();
 FILLCELL_X32 FILLER_338_2503 ();
 FILLCELL_X32 FILLER_338_2535 ();
 FILLCELL_X32 FILLER_338_2567 ();
 FILLCELL_X32 FILLER_338_2599 ();
 FILLCELL_X32 FILLER_338_2631 ();
 FILLCELL_X32 FILLER_338_2663 ();
 FILLCELL_X32 FILLER_338_2695 ();
 FILLCELL_X32 FILLER_338_2727 ();
 FILLCELL_X32 FILLER_338_2759 ();
 FILLCELL_X32 FILLER_338_2791 ();
 FILLCELL_X32 FILLER_338_2823 ();
 FILLCELL_X32 FILLER_338_2855 ();
 FILLCELL_X32 FILLER_338_2887 ();
 FILLCELL_X32 FILLER_338_2919 ();
 FILLCELL_X32 FILLER_338_2951 ();
 FILLCELL_X32 FILLER_338_2983 ();
 FILLCELL_X32 FILLER_338_3015 ();
 FILLCELL_X32 FILLER_338_3047 ();
 FILLCELL_X32 FILLER_338_3079 ();
 FILLCELL_X32 FILLER_338_3111 ();
 FILLCELL_X8 FILLER_338_3143 ();
 FILLCELL_X4 FILLER_338_3151 ();
 FILLCELL_X2 FILLER_338_3155 ();
 FILLCELL_X32 FILLER_338_3158 ();
 FILLCELL_X32 FILLER_338_3190 ();
 FILLCELL_X32 FILLER_338_3222 ();
 FILLCELL_X32 FILLER_338_3254 ();
 FILLCELL_X32 FILLER_338_3286 ();
 FILLCELL_X32 FILLER_338_3318 ();
 FILLCELL_X32 FILLER_338_3350 ();
 FILLCELL_X32 FILLER_338_3382 ();
 FILLCELL_X32 FILLER_338_3414 ();
 FILLCELL_X32 FILLER_338_3446 ();
 FILLCELL_X32 FILLER_338_3478 ();
 FILLCELL_X32 FILLER_338_3510 ();
 FILLCELL_X32 FILLER_338_3542 ();
 FILLCELL_X32 FILLER_338_3574 ();
 FILLCELL_X32 FILLER_338_3606 ();
 FILLCELL_X32 FILLER_338_3638 ();
 FILLCELL_X32 FILLER_338_3670 ();
 FILLCELL_X32 FILLER_338_3702 ();
 FILLCELL_X4 FILLER_338_3734 ();
 FILLCELL_X32 FILLER_339_1 ();
 FILLCELL_X32 FILLER_339_33 ();
 FILLCELL_X32 FILLER_339_65 ();
 FILLCELL_X32 FILLER_339_97 ();
 FILLCELL_X32 FILLER_339_129 ();
 FILLCELL_X32 FILLER_339_161 ();
 FILLCELL_X32 FILLER_339_193 ();
 FILLCELL_X32 FILLER_339_225 ();
 FILLCELL_X32 FILLER_339_257 ();
 FILLCELL_X32 FILLER_339_289 ();
 FILLCELL_X32 FILLER_339_321 ();
 FILLCELL_X32 FILLER_339_353 ();
 FILLCELL_X32 FILLER_339_385 ();
 FILLCELL_X32 FILLER_339_417 ();
 FILLCELL_X32 FILLER_339_449 ();
 FILLCELL_X32 FILLER_339_481 ();
 FILLCELL_X32 FILLER_339_513 ();
 FILLCELL_X32 FILLER_339_545 ();
 FILLCELL_X32 FILLER_339_577 ();
 FILLCELL_X32 FILLER_339_609 ();
 FILLCELL_X32 FILLER_339_641 ();
 FILLCELL_X32 FILLER_339_673 ();
 FILLCELL_X32 FILLER_339_705 ();
 FILLCELL_X32 FILLER_339_737 ();
 FILLCELL_X32 FILLER_339_769 ();
 FILLCELL_X32 FILLER_339_801 ();
 FILLCELL_X32 FILLER_339_833 ();
 FILLCELL_X32 FILLER_339_865 ();
 FILLCELL_X32 FILLER_339_897 ();
 FILLCELL_X32 FILLER_339_929 ();
 FILLCELL_X32 FILLER_339_961 ();
 FILLCELL_X32 FILLER_339_993 ();
 FILLCELL_X32 FILLER_339_1025 ();
 FILLCELL_X32 FILLER_339_1057 ();
 FILLCELL_X32 FILLER_339_1089 ();
 FILLCELL_X32 FILLER_339_1121 ();
 FILLCELL_X32 FILLER_339_1153 ();
 FILLCELL_X32 FILLER_339_1185 ();
 FILLCELL_X32 FILLER_339_1217 ();
 FILLCELL_X8 FILLER_339_1249 ();
 FILLCELL_X4 FILLER_339_1257 ();
 FILLCELL_X2 FILLER_339_1261 ();
 FILLCELL_X32 FILLER_339_1264 ();
 FILLCELL_X32 FILLER_339_1296 ();
 FILLCELL_X32 FILLER_339_1328 ();
 FILLCELL_X32 FILLER_339_1360 ();
 FILLCELL_X32 FILLER_339_1392 ();
 FILLCELL_X32 FILLER_339_1424 ();
 FILLCELL_X32 FILLER_339_1456 ();
 FILLCELL_X32 FILLER_339_1488 ();
 FILLCELL_X32 FILLER_339_1520 ();
 FILLCELL_X32 FILLER_339_1552 ();
 FILLCELL_X32 FILLER_339_1584 ();
 FILLCELL_X32 FILLER_339_1616 ();
 FILLCELL_X32 FILLER_339_1648 ();
 FILLCELL_X32 FILLER_339_1680 ();
 FILLCELL_X32 FILLER_339_1712 ();
 FILLCELL_X32 FILLER_339_1744 ();
 FILLCELL_X32 FILLER_339_1776 ();
 FILLCELL_X32 FILLER_339_1808 ();
 FILLCELL_X32 FILLER_339_1840 ();
 FILLCELL_X32 FILLER_339_1872 ();
 FILLCELL_X32 FILLER_339_1904 ();
 FILLCELL_X32 FILLER_339_1936 ();
 FILLCELL_X32 FILLER_339_1968 ();
 FILLCELL_X32 FILLER_339_2000 ();
 FILLCELL_X32 FILLER_339_2032 ();
 FILLCELL_X32 FILLER_339_2064 ();
 FILLCELL_X32 FILLER_339_2096 ();
 FILLCELL_X32 FILLER_339_2128 ();
 FILLCELL_X32 FILLER_339_2160 ();
 FILLCELL_X32 FILLER_339_2192 ();
 FILLCELL_X32 FILLER_339_2224 ();
 FILLCELL_X32 FILLER_339_2256 ();
 FILLCELL_X32 FILLER_339_2288 ();
 FILLCELL_X32 FILLER_339_2320 ();
 FILLCELL_X32 FILLER_339_2352 ();
 FILLCELL_X32 FILLER_339_2384 ();
 FILLCELL_X32 FILLER_339_2416 ();
 FILLCELL_X32 FILLER_339_2448 ();
 FILLCELL_X32 FILLER_339_2480 ();
 FILLCELL_X8 FILLER_339_2512 ();
 FILLCELL_X4 FILLER_339_2520 ();
 FILLCELL_X2 FILLER_339_2524 ();
 FILLCELL_X32 FILLER_339_2527 ();
 FILLCELL_X32 FILLER_339_2559 ();
 FILLCELL_X32 FILLER_339_2591 ();
 FILLCELL_X32 FILLER_339_2623 ();
 FILLCELL_X32 FILLER_339_2655 ();
 FILLCELL_X32 FILLER_339_2687 ();
 FILLCELL_X32 FILLER_339_2719 ();
 FILLCELL_X32 FILLER_339_2751 ();
 FILLCELL_X32 FILLER_339_2783 ();
 FILLCELL_X32 FILLER_339_2815 ();
 FILLCELL_X32 FILLER_339_2847 ();
 FILLCELL_X32 FILLER_339_2879 ();
 FILLCELL_X32 FILLER_339_2911 ();
 FILLCELL_X32 FILLER_339_2943 ();
 FILLCELL_X32 FILLER_339_2975 ();
 FILLCELL_X32 FILLER_339_3007 ();
 FILLCELL_X32 FILLER_339_3039 ();
 FILLCELL_X32 FILLER_339_3071 ();
 FILLCELL_X32 FILLER_339_3103 ();
 FILLCELL_X32 FILLER_339_3135 ();
 FILLCELL_X32 FILLER_339_3167 ();
 FILLCELL_X32 FILLER_339_3199 ();
 FILLCELL_X32 FILLER_339_3231 ();
 FILLCELL_X32 FILLER_339_3263 ();
 FILLCELL_X32 FILLER_339_3295 ();
 FILLCELL_X32 FILLER_339_3327 ();
 FILLCELL_X32 FILLER_339_3359 ();
 FILLCELL_X32 FILLER_339_3391 ();
 FILLCELL_X32 FILLER_339_3423 ();
 FILLCELL_X32 FILLER_339_3455 ();
 FILLCELL_X32 FILLER_339_3487 ();
 FILLCELL_X32 FILLER_339_3519 ();
 FILLCELL_X32 FILLER_339_3551 ();
 FILLCELL_X32 FILLER_339_3583 ();
 FILLCELL_X32 FILLER_339_3615 ();
 FILLCELL_X32 FILLER_339_3647 ();
 FILLCELL_X32 FILLER_339_3679 ();
 FILLCELL_X16 FILLER_339_3711 ();
 FILLCELL_X8 FILLER_339_3727 ();
 FILLCELL_X2 FILLER_339_3735 ();
 FILLCELL_X1 FILLER_339_3737 ();
 FILLCELL_X32 FILLER_340_1 ();
 FILLCELL_X32 FILLER_340_33 ();
 FILLCELL_X32 FILLER_340_65 ();
 FILLCELL_X32 FILLER_340_97 ();
 FILLCELL_X32 FILLER_340_129 ();
 FILLCELL_X32 FILLER_340_161 ();
 FILLCELL_X32 FILLER_340_193 ();
 FILLCELL_X32 FILLER_340_225 ();
 FILLCELL_X32 FILLER_340_257 ();
 FILLCELL_X32 FILLER_340_289 ();
 FILLCELL_X32 FILLER_340_321 ();
 FILLCELL_X32 FILLER_340_353 ();
 FILLCELL_X32 FILLER_340_385 ();
 FILLCELL_X32 FILLER_340_417 ();
 FILLCELL_X32 FILLER_340_449 ();
 FILLCELL_X32 FILLER_340_481 ();
 FILLCELL_X32 FILLER_340_513 ();
 FILLCELL_X32 FILLER_340_545 ();
 FILLCELL_X32 FILLER_340_577 ();
 FILLCELL_X16 FILLER_340_609 ();
 FILLCELL_X4 FILLER_340_625 ();
 FILLCELL_X2 FILLER_340_629 ();
 FILLCELL_X32 FILLER_340_632 ();
 FILLCELL_X32 FILLER_340_664 ();
 FILLCELL_X32 FILLER_340_696 ();
 FILLCELL_X32 FILLER_340_728 ();
 FILLCELL_X32 FILLER_340_760 ();
 FILLCELL_X32 FILLER_340_792 ();
 FILLCELL_X32 FILLER_340_824 ();
 FILLCELL_X32 FILLER_340_856 ();
 FILLCELL_X32 FILLER_340_888 ();
 FILLCELL_X32 FILLER_340_920 ();
 FILLCELL_X32 FILLER_340_952 ();
 FILLCELL_X32 FILLER_340_984 ();
 FILLCELL_X32 FILLER_340_1016 ();
 FILLCELL_X32 FILLER_340_1048 ();
 FILLCELL_X32 FILLER_340_1080 ();
 FILLCELL_X32 FILLER_340_1112 ();
 FILLCELL_X32 FILLER_340_1144 ();
 FILLCELL_X32 FILLER_340_1176 ();
 FILLCELL_X32 FILLER_340_1208 ();
 FILLCELL_X32 FILLER_340_1240 ();
 FILLCELL_X32 FILLER_340_1272 ();
 FILLCELL_X32 FILLER_340_1304 ();
 FILLCELL_X32 FILLER_340_1336 ();
 FILLCELL_X32 FILLER_340_1368 ();
 FILLCELL_X32 FILLER_340_1400 ();
 FILLCELL_X32 FILLER_340_1432 ();
 FILLCELL_X32 FILLER_340_1464 ();
 FILLCELL_X32 FILLER_340_1496 ();
 FILLCELL_X32 FILLER_340_1528 ();
 FILLCELL_X32 FILLER_340_1560 ();
 FILLCELL_X32 FILLER_340_1592 ();
 FILLCELL_X32 FILLER_340_1624 ();
 FILLCELL_X32 FILLER_340_1656 ();
 FILLCELL_X32 FILLER_340_1688 ();
 FILLCELL_X32 FILLER_340_1720 ();
 FILLCELL_X32 FILLER_340_1752 ();
 FILLCELL_X32 FILLER_340_1784 ();
 FILLCELL_X32 FILLER_340_1816 ();
 FILLCELL_X32 FILLER_340_1848 ();
 FILLCELL_X8 FILLER_340_1880 ();
 FILLCELL_X4 FILLER_340_1888 ();
 FILLCELL_X2 FILLER_340_1892 ();
 FILLCELL_X32 FILLER_340_1895 ();
 FILLCELL_X32 FILLER_340_1927 ();
 FILLCELL_X32 FILLER_340_1959 ();
 FILLCELL_X32 FILLER_340_1991 ();
 FILLCELL_X32 FILLER_340_2023 ();
 FILLCELL_X32 FILLER_340_2055 ();
 FILLCELL_X32 FILLER_340_2087 ();
 FILLCELL_X32 FILLER_340_2119 ();
 FILLCELL_X32 FILLER_340_2151 ();
 FILLCELL_X32 FILLER_340_2183 ();
 FILLCELL_X32 FILLER_340_2215 ();
 FILLCELL_X32 FILLER_340_2247 ();
 FILLCELL_X32 FILLER_340_2279 ();
 FILLCELL_X32 FILLER_340_2311 ();
 FILLCELL_X32 FILLER_340_2343 ();
 FILLCELL_X32 FILLER_340_2375 ();
 FILLCELL_X32 FILLER_340_2407 ();
 FILLCELL_X32 FILLER_340_2439 ();
 FILLCELL_X32 FILLER_340_2471 ();
 FILLCELL_X32 FILLER_340_2503 ();
 FILLCELL_X32 FILLER_340_2535 ();
 FILLCELL_X32 FILLER_340_2567 ();
 FILLCELL_X32 FILLER_340_2599 ();
 FILLCELL_X32 FILLER_340_2631 ();
 FILLCELL_X32 FILLER_340_2663 ();
 FILLCELL_X32 FILLER_340_2695 ();
 FILLCELL_X32 FILLER_340_2727 ();
 FILLCELL_X32 FILLER_340_2759 ();
 FILLCELL_X32 FILLER_340_2791 ();
 FILLCELL_X32 FILLER_340_2823 ();
 FILLCELL_X32 FILLER_340_2855 ();
 FILLCELL_X32 FILLER_340_2887 ();
 FILLCELL_X32 FILLER_340_2919 ();
 FILLCELL_X32 FILLER_340_2951 ();
 FILLCELL_X32 FILLER_340_2983 ();
 FILLCELL_X32 FILLER_340_3015 ();
 FILLCELL_X32 FILLER_340_3047 ();
 FILLCELL_X32 FILLER_340_3079 ();
 FILLCELL_X32 FILLER_340_3111 ();
 FILLCELL_X8 FILLER_340_3143 ();
 FILLCELL_X4 FILLER_340_3151 ();
 FILLCELL_X2 FILLER_340_3155 ();
 FILLCELL_X32 FILLER_340_3158 ();
 FILLCELL_X32 FILLER_340_3190 ();
 FILLCELL_X32 FILLER_340_3222 ();
 FILLCELL_X32 FILLER_340_3254 ();
 FILLCELL_X32 FILLER_340_3286 ();
 FILLCELL_X32 FILLER_340_3318 ();
 FILLCELL_X32 FILLER_340_3350 ();
 FILLCELL_X32 FILLER_340_3382 ();
 FILLCELL_X32 FILLER_340_3414 ();
 FILLCELL_X32 FILLER_340_3446 ();
 FILLCELL_X32 FILLER_340_3478 ();
 FILLCELL_X32 FILLER_340_3510 ();
 FILLCELL_X32 FILLER_340_3542 ();
 FILLCELL_X32 FILLER_340_3574 ();
 FILLCELL_X32 FILLER_340_3606 ();
 FILLCELL_X32 FILLER_340_3638 ();
 FILLCELL_X32 FILLER_340_3670 ();
 FILLCELL_X32 FILLER_340_3702 ();
 FILLCELL_X4 FILLER_340_3734 ();
 FILLCELL_X32 FILLER_341_1 ();
 FILLCELL_X32 FILLER_341_33 ();
 FILLCELL_X32 FILLER_341_65 ();
 FILLCELL_X32 FILLER_341_97 ();
 FILLCELL_X32 FILLER_341_129 ();
 FILLCELL_X32 FILLER_341_161 ();
 FILLCELL_X32 FILLER_341_193 ();
 FILLCELL_X32 FILLER_341_225 ();
 FILLCELL_X32 FILLER_341_257 ();
 FILLCELL_X32 FILLER_341_289 ();
 FILLCELL_X32 FILLER_341_321 ();
 FILLCELL_X32 FILLER_341_353 ();
 FILLCELL_X32 FILLER_341_385 ();
 FILLCELL_X32 FILLER_341_417 ();
 FILLCELL_X32 FILLER_341_449 ();
 FILLCELL_X32 FILLER_341_481 ();
 FILLCELL_X32 FILLER_341_513 ();
 FILLCELL_X32 FILLER_341_545 ();
 FILLCELL_X32 FILLER_341_577 ();
 FILLCELL_X32 FILLER_341_609 ();
 FILLCELL_X32 FILLER_341_641 ();
 FILLCELL_X32 FILLER_341_673 ();
 FILLCELL_X32 FILLER_341_705 ();
 FILLCELL_X32 FILLER_341_737 ();
 FILLCELL_X32 FILLER_341_769 ();
 FILLCELL_X32 FILLER_341_801 ();
 FILLCELL_X32 FILLER_341_833 ();
 FILLCELL_X32 FILLER_341_865 ();
 FILLCELL_X32 FILLER_341_897 ();
 FILLCELL_X32 FILLER_341_929 ();
 FILLCELL_X32 FILLER_341_961 ();
 FILLCELL_X32 FILLER_341_993 ();
 FILLCELL_X32 FILLER_341_1025 ();
 FILLCELL_X32 FILLER_341_1057 ();
 FILLCELL_X32 FILLER_341_1089 ();
 FILLCELL_X32 FILLER_341_1121 ();
 FILLCELL_X32 FILLER_341_1153 ();
 FILLCELL_X32 FILLER_341_1185 ();
 FILLCELL_X32 FILLER_341_1217 ();
 FILLCELL_X8 FILLER_341_1249 ();
 FILLCELL_X4 FILLER_341_1257 ();
 FILLCELL_X2 FILLER_341_1261 ();
 FILLCELL_X32 FILLER_341_1264 ();
 FILLCELL_X32 FILLER_341_1296 ();
 FILLCELL_X32 FILLER_341_1328 ();
 FILLCELL_X32 FILLER_341_1360 ();
 FILLCELL_X32 FILLER_341_1392 ();
 FILLCELL_X32 FILLER_341_1424 ();
 FILLCELL_X32 FILLER_341_1456 ();
 FILLCELL_X32 FILLER_341_1488 ();
 FILLCELL_X32 FILLER_341_1520 ();
 FILLCELL_X32 FILLER_341_1552 ();
 FILLCELL_X32 FILLER_341_1584 ();
 FILLCELL_X32 FILLER_341_1616 ();
 FILLCELL_X32 FILLER_341_1648 ();
 FILLCELL_X32 FILLER_341_1680 ();
 FILLCELL_X32 FILLER_341_1712 ();
 FILLCELL_X32 FILLER_341_1744 ();
 FILLCELL_X32 FILLER_341_1776 ();
 FILLCELL_X32 FILLER_341_1808 ();
 FILLCELL_X32 FILLER_341_1840 ();
 FILLCELL_X32 FILLER_341_1872 ();
 FILLCELL_X32 FILLER_341_1904 ();
 FILLCELL_X32 FILLER_341_1936 ();
 FILLCELL_X32 FILLER_341_1968 ();
 FILLCELL_X32 FILLER_341_2000 ();
 FILLCELL_X32 FILLER_341_2032 ();
 FILLCELL_X32 FILLER_341_2064 ();
 FILLCELL_X32 FILLER_341_2096 ();
 FILLCELL_X32 FILLER_341_2128 ();
 FILLCELL_X32 FILLER_341_2160 ();
 FILLCELL_X32 FILLER_341_2192 ();
 FILLCELL_X32 FILLER_341_2224 ();
 FILLCELL_X32 FILLER_341_2256 ();
 FILLCELL_X32 FILLER_341_2288 ();
 FILLCELL_X32 FILLER_341_2320 ();
 FILLCELL_X32 FILLER_341_2352 ();
 FILLCELL_X32 FILLER_341_2384 ();
 FILLCELL_X32 FILLER_341_2416 ();
 FILLCELL_X32 FILLER_341_2448 ();
 FILLCELL_X32 FILLER_341_2480 ();
 FILLCELL_X8 FILLER_341_2512 ();
 FILLCELL_X4 FILLER_341_2520 ();
 FILLCELL_X2 FILLER_341_2524 ();
 FILLCELL_X32 FILLER_341_2527 ();
 FILLCELL_X32 FILLER_341_2559 ();
 FILLCELL_X32 FILLER_341_2591 ();
 FILLCELL_X32 FILLER_341_2623 ();
 FILLCELL_X32 FILLER_341_2655 ();
 FILLCELL_X32 FILLER_341_2687 ();
 FILLCELL_X32 FILLER_341_2719 ();
 FILLCELL_X32 FILLER_341_2751 ();
 FILLCELL_X32 FILLER_341_2783 ();
 FILLCELL_X32 FILLER_341_2815 ();
 FILLCELL_X32 FILLER_341_2847 ();
 FILLCELL_X32 FILLER_341_2879 ();
 FILLCELL_X32 FILLER_341_2911 ();
 FILLCELL_X32 FILLER_341_2943 ();
 FILLCELL_X32 FILLER_341_2975 ();
 FILLCELL_X32 FILLER_341_3007 ();
 FILLCELL_X32 FILLER_341_3039 ();
 FILLCELL_X32 FILLER_341_3071 ();
 FILLCELL_X32 FILLER_341_3103 ();
 FILLCELL_X32 FILLER_341_3135 ();
 FILLCELL_X32 FILLER_341_3167 ();
 FILLCELL_X32 FILLER_341_3199 ();
 FILLCELL_X32 FILLER_341_3231 ();
 FILLCELL_X32 FILLER_341_3263 ();
 FILLCELL_X32 FILLER_341_3295 ();
 FILLCELL_X32 FILLER_341_3327 ();
 FILLCELL_X32 FILLER_341_3359 ();
 FILLCELL_X32 FILLER_341_3391 ();
 FILLCELL_X32 FILLER_341_3423 ();
 FILLCELL_X32 FILLER_341_3455 ();
 FILLCELL_X32 FILLER_341_3487 ();
 FILLCELL_X32 FILLER_341_3519 ();
 FILLCELL_X32 FILLER_341_3551 ();
 FILLCELL_X32 FILLER_341_3583 ();
 FILLCELL_X32 FILLER_341_3615 ();
 FILLCELL_X32 FILLER_341_3647 ();
 FILLCELL_X32 FILLER_341_3679 ();
 FILLCELL_X16 FILLER_341_3711 ();
 FILLCELL_X8 FILLER_341_3727 ();
 FILLCELL_X2 FILLER_341_3735 ();
 FILLCELL_X1 FILLER_341_3737 ();
 FILLCELL_X32 FILLER_342_1 ();
 FILLCELL_X32 FILLER_342_33 ();
 FILLCELL_X32 FILLER_342_65 ();
 FILLCELL_X32 FILLER_342_97 ();
 FILLCELL_X32 FILLER_342_129 ();
 FILLCELL_X32 FILLER_342_161 ();
 FILLCELL_X32 FILLER_342_193 ();
 FILLCELL_X32 FILLER_342_225 ();
 FILLCELL_X32 FILLER_342_257 ();
 FILLCELL_X32 FILLER_342_289 ();
 FILLCELL_X32 FILLER_342_321 ();
 FILLCELL_X32 FILLER_342_353 ();
 FILLCELL_X32 FILLER_342_385 ();
 FILLCELL_X32 FILLER_342_417 ();
 FILLCELL_X32 FILLER_342_449 ();
 FILLCELL_X32 FILLER_342_481 ();
 FILLCELL_X32 FILLER_342_513 ();
 FILLCELL_X32 FILLER_342_545 ();
 FILLCELL_X32 FILLER_342_577 ();
 FILLCELL_X16 FILLER_342_609 ();
 FILLCELL_X4 FILLER_342_625 ();
 FILLCELL_X2 FILLER_342_629 ();
 FILLCELL_X32 FILLER_342_632 ();
 FILLCELL_X32 FILLER_342_664 ();
 FILLCELL_X32 FILLER_342_696 ();
 FILLCELL_X32 FILLER_342_728 ();
 FILLCELL_X32 FILLER_342_760 ();
 FILLCELL_X32 FILLER_342_792 ();
 FILLCELL_X32 FILLER_342_824 ();
 FILLCELL_X32 FILLER_342_856 ();
 FILLCELL_X32 FILLER_342_888 ();
 FILLCELL_X32 FILLER_342_920 ();
 FILLCELL_X32 FILLER_342_952 ();
 FILLCELL_X32 FILLER_342_984 ();
 FILLCELL_X32 FILLER_342_1016 ();
 FILLCELL_X32 FILLER_342_1048 ();
 FILLCELL_X32 FILLER_342_1080 ();
 FILLCELL_X32 FILLER_342_1112 ();
 FILLCELL_X32 FILLER_342_1144 ();
 FILLCELL_X32 FILLER_342_1176 ();
 FILLCELL_X32 FILLER_342_1208 ();
 FILLCELL_X32 FILLER_342_1240 ();
 FILLCELL_X32 FILLER_342_1272 ();
 FILLCELL_X32 FILLER_342_1304 ();
 FILLCELL_X32 FILLER_342_1336 ();
 FILLCELL_X32 FILLER_342_1368 ();
 FILLCELL_X32 FILLER_342_1400 ();
 FILLCELL_X32 FILLER_342_1432 ();
 FILLCELL_X32 FILLER_342_1464 ();
 FILLCELL_X32 FILLER_342_1496 ();
 FILLCELL_X32 FILLER_342_1528 ();
 FILLCELL_X32 FILLER_342_1560 ();
 FILLCELL_X32 FILLER_342_1592 ();
 FILLCELL_X32 FILLER_342_1624 ();
 FILLCELL_X32 FILLER_342_1656 ();
 FILLCELL_X32 FILLER_342_1688 ();
 FILLCELL_X32 FILLER_342_1720 ();
 FILLCELL_X32 FILLER_342_1752 ();
 FILLCELL_X32 FILLER_342_1784 ();
 FILLCELL_X32 FILLER_342_1816 ();
 FILLCELL_X32 FILLER_342_1848 ();
 FILLCELL_X8 FILLER_342_1880 ();
 FILLCELL_X4 FILLER_342_1888 ();
 FILLCELL_X2 FILLER_342_1892 ();
 FILLCELL_X32 FILLER_342_1895 ();
 FILLCELL_X32 FILLER_342_1927 ();
 FILLCELL_X32 FILLER_342_1959 ();
 FILLCELL_X32 FILLER_342_1991 ();
 FILLCELL_X32 FILLER_342_2023 ();
 FILLCELL_X32 FILLER_342_2055 ();
 FILLCELL_X32 FILLER_342_2087 ();
 FILLCELL_X32 FILLER_342_2119 ();
 FILLCELL_X32 FILLER_342_2151 ();
 FILLCELL_X32 FILLER_342_2183 ();
 FILLCELL_X32 FILLER_342_2215 ();
 FILLCELL_X32 FILLER_342_2247 ();
 FILLCELL_X32 FILLER_342_2279 ();
 FILLCELL_X32 FILLER_342_2311 ();
 FILLCELL_X32 FILLER_342_2343 ();
 FILLCELL_X32 FILLER_342_2375 ();
 FILLCELL_X32 FILLER_342_2407 ();
 FILLCELL_X32 FILLER_342_2439 ();
 FILLCELL_X32 FILLER_342_2471 ();
 FILLCELL_X32 FILLER_342_2503 ();
 FILLCELL_X32 FILLER_342_2535 ();
 FILLCELL_X32 FILLER_342_2567 ();
 FILLCELL_X32 FILLER_342_2599 ();
 FILLCELL_X32 FILLER_342_2631 ();
 FILLCELL_X32 FILLER_342_2663 ();
 FILLCELL_X32 FILLER_342_2695 ();
 FILLCELL_X32 FILLER_342_2727 ();
 FILLCELL_X32 FILLER_342_2759 ();
 FILLCELL_X32 FILLER_342_2791 ();
 FILLCELL_X32 FILLER_342_2823 ();
 FILLCELL_X32 FILLER_342_2855 ();
 FILLCELL_X32 FILLER_342_2887 ();
 FILLCELL_X32 FILLER_342_2919 ();
 FILLCELL_X32 FILLER_342_2951 ();
 FILLCELL_X32 FILLER_342_2983 ();
 FILLCELL_X32 FILLER_342_3015 ();
 FILLCELL_X32 FILLER_342_3047 ();
 FILLCELL_X32 FILLER_342_3079 ();
 FILLCELL_X32 FILLER_342_3111 ();
 FILLCELL_X8 FILLER_342_3143 ();
 FILLCELL_X4 FILLER_342_3151 ();
 FILLCELL_X2 FILLER_342_3155 ();
 FILLCELL_X32 FILLER_342_3158 ();
 FILLCELL_X32 FILLER_342_3190 ();
 FILLCELL_X32 FILLER_342_3222 ();
 FILLCELL_X32 FILLER_342_3254 ();
 FILLCELL_X32 FILLER_342_3286 ();
 FILLCELL_X32 FILLER_342_3318 ();
 FILLCELL_X32 FILLER_342_3350 ();
 FILLCELL_X32 FILLER_342_3382 ();
 FILLCELL_X32 FILLER_342_3414 ();
 FILLCELL_X32 FILLER_342_3446 ();
 FILLCELL_X32 FILLER_342_3478 ();
 FILLCELL_X32 FILLER_342_3510 ();
 FILLCELL_X32 FILLER_342_3542 ();
 FILLCELL_X32 FILLER_342_3574 ();
 FILLCELL_X32 FILLER_342_3606 ();
 FILLCELL_X32 FILLER_342_3638 ();
 FILLCELL_X32 FILLER_342_3670 ();
 FILLCELL_X32 FILLER_342_3702 ();
 FILLCELL_X4 FILLER_342_3734 ();
 FILLCELL_X32 FILLER_343_1 ();
 FILLCELL_X32 FILLER_343_33 ();
 FILLCELL_X32 FILLER_343_65 ();
 FILLCELL_X32 FILLER_343_97 ();
 FILLCELL_X32 FILLER_343_129 ();
 FILLCELL_X32 FILLER_343_161 ();
 FILLCELL_X32 FILLER_343_193 ();
 FILLCELL_X32 FILLER_343_225 ();
 FILLCELL_X32 FILLER_343_257 ();
 FILLCELL_X32 FILLER_343_289 ();
 FILLCELL_X32 FILLER_343_321 ();
 FILLCELL_X32 FILLER_343_353 ();
 FILLCELL_X32 FILLER_343_385 ();
 FILLCELL_X32 FILLER_343_417 ();
 FILLCELL_X32 FILLER_343_449 ();
 FILLCELL_X32 FILLER_343_481 ();
 FILLCELL_X32 FILLER_343_513 ();
 FILLCELL_X32 FILLER_343_545 ();
 FILLCELL_X32 FILLER_343_577 ();
 FILLCELL_X32 FILLER_343_609 ();
 FILLCELL_X32 FILLER_343_641 ();
 FILLCELL_X32 FILLER_343_673 ();
 FILLCELL_X32 FILLER_343_705 ();
 FILLCELL_X32 FILLER_343_737 ();
 FILLCELL_X32 FILLER_343_769 ();
 FILLCELL_X32 FILLER_343_801 ();
 FILLCELL_X32 FILLER_343_833 ();
 FILLCELL_X32 FILLER_343_865 ();
 FILLCELL_X32 FILLER_343_897 ();
 FILLCELL_X32 FILLER_343_929 ();
 FILLCELL_X32 FILLER_343_961 ();
 FILLCELL_X32 FILLER_343_993 ();
 FILLCELL_X32 FILLER_343_1025 ();
 FILLCELL_X32 FILLER_343_1057 ();
 FILLCELL_X32 FILLER_343_1089 ();
 FILLCELL_X32 FILLER_343_1121 ();
 FILLCELL_X32 FILLER_343_1153 ();
 FILLCELL_X32 FILLER_343_1185 ();
 FILLCELL_X32 FILLER_343_1217 ();
 FILLCELL_X8 FILLER_343_1249 ();
 FILLCELL_X4 FILLER_343_1257 ();
 FILLCELL_X2 FILLER_343_1261 ();
 FILLCELL_X32 FILLER_343_1264 ();
 FILLCELL_X32 FILLER_343_1296 ();
 FILLCELL_X32 FILLER_343_1328 ();
 FILLCELL_X32 FILLER_343_1360 ();
 FILLCELL_X32 FILLER_343_1392 ();
 FILLCELL_X32 FILLER_343_1424 ();
 FILLCELL_X32 FILLER_343_1456 ();
 FILLCELL_X32 FILLER_343_1488 ();
 FILLCELL_X32 FILLER_343_1520 ();
 FILLCELL_X32 FILLER_343_1552 ();
 FILLCELL_X32 FILLER_343_1584 ();
 FILLCELL_X32 FILLER_343_1616 ();
 FILLCELL_X32 FILLER_343_1648 ();
 FILLCELL_X32 FILLER_343_1680 ();
 FILLCELL_X32 FILLER_343_1712 ();
 FILLCELL_X32 FILLER_343_1744 ();
 FILLCELL_X32 FILLER_343_1776 ();
 FILLCELL_X32 FILLER_343_1808 ();
 FILLCELL_X32 FILLER_343_1840 ();
 FILLCELL_X32 FILLER_343_1872 ();
 FILLCELL_X32 FILLER_343_1904 ();
 FILLCELL_X32 FILLER_343_1936 ();
 FILLCELL_X32 FILLER_343_1968 ();
 FILLCELL_X32 FILLER_343_2000 ();
 FILLCELL_X32 FILLER_343_2032 ();
 FILLCELL_X32 FILLER_343_2064 ();
 FILLCELL_X32 FILLER_343_2096 ();
 FILLCELL_X32 FILLER_343_2128 ();
 FILLCELL_X32 FILLER_343_2160 ();
 FILLCELL_X32 FILLER_343_2192 ();
 FILLCELL_X32 FILLER_343_2224 ();
 FILLCELL_X32 FILLER_343_2256 ();
 FILLCELL_X32 FILLER_343_2288 ();
 FILLCELL_X32 FILLER_343_2320 ();
 FILLCELL_X32 FILLER_343_2352 ();
 FILLCELL_X32 FILLER_343_2384 ();
 FILLCELL_X32 FILLER_343_2416 ();
 FILLCELL_X32 FILLER_343_2448 ();
 FILLCELL_X32 FILLER_343_2480 ();
 FILLCELL_X8 FILLER_343_2512 ();
 FILLCELL_X4 FILLER_343_2520 ();
 FILLCELL_X2 FILLER_343_2524 ();
 FILLCELL_X32 FILLER_343_2527 ();
 FILLCELL_X32 FILLER_343_2559 ();
 FILLCELL_X32 FILLER_343_2591 ();
 FILLCELL_X32 FILLER_343_2623 ();
 FILLCELL_X32 FILLER_343_2655 ();
 FILLCELL_X32 FILLER_343_2687 ();
 FILLCELL_X32 FILLER_343_2719 ();
 FILLCELL_X32 FILLER_343_2751 ();
 FILLCELL_X32 FILLER_343_2783 ();
 FILLCELL_X32 FILLER_343_2815 ();
 FILLCELL_X32 FILLER_343_2847 ();
 FILLCELL_X32 FILLER_343_2879 ();
 FILLCELL_X32 FILLER_343_2911 ();
 FILLCELL_X32 FILLER_343_2943 ();
 FILLCELL_X32 FILLER_343_2975 ();
 FILLCELL_X32 FILLER_343_3007 ();
 FILLCELL_X32 FILLER_343_3039 ();
 FILLCELL_X32 FILLER_343_3071 ();
 FILLCELL_X32 FILLER_343_3103 ();
 FILLCELL_X32 FILLER_343_3135 ();
 FILLCELL_X32 FILLER_343_3167 ();
 FILLCELL_X32 FILLER_343_3199 ();
 FILLCELL_X32 FILLER_343_3231 ();
 FILLCELL_X32 FILLER_343_3263 ();
 FILLCELL_X32 FILLER_343_3295 ();
 FILLCELL_X32 FILLER_343_3327 ();
 FILLCELL_X32 FILLER_343_3359 ();
 FILLCELL_X32 FILLER_343_3391 ();
 FILLCELL_X32 FILLER_343_3423 ();
 FILLCELL_X32 FILLER_343_3455 ();
 FILLCELL_X32 FILLER_343_3487 ();
 FILLCELL_X32 FILLER_343_3519 ();
 FILLCELL_X32 FILLER_343_3551 ();
 FILLCELL_X32 FILLER_343_3583 ();
 FILLCELL_X32 FILLER_343_3615 ();
 FILLCELL_X32 FILLER_343_3647 ();
 FILLCELL_X32 FILLER_343_3679 ();
 FILLCELL_X16 FILLER_343_3711 ();
 FILLCELL_X8 FILLER_343_3727 ();
 FILLCELL_X2 FILLER_343_3735 ();
 FILLCELL_X1 FILLER_343_3737 ();
 FILLCELL_X32 FILLER_344_1 ();
 FILLCELL_X32 FILLER_344_33 ();
 FILLCELL_X32 FILLER_344_65 ();
 FILLCELL_X32 FILLER_344_97 ();
 FILLCELL_X32 FILLER_344_129 ();
 FILLCELL_X32 FILLER_344_161 ();
 FILLCELL_X32 FILLER_344_193 ();
 FILLCELL_X32 FILLER_344_225 ();
 FILLCELL_X32 FILLER_344_257 ();
 FILLCELL_X32 FILLER_344_289 ();
 FILLCELL_X32 FILLER_344_321 ();
 FILLCELL_X32 FILLER_344_353 ();
 FILLCELL_X32 FILLER_344_385 ();
 FILLCELL_X32 FILLER_344_417 ();
 FILLCELL_X32 FILLER_344_449 ();
 FILLCELL_X32 FILLER_344_481 ();
 FILLCELL_X32 FILLER_344_513 ();
 FILLCELL_X32 FILLER_344_545 ();
 FILLCELL_X32 FILLER_344_577 ();
 FILLCELL_X16 FILLER_344_609 ();
 FILLCELL_X4 FILLER_344_625 ();
 FILLCELL_X2 FILLER_344_629 ();
 FILLCELL_X32 FILLER_344_632 ();
 FILLCELL_X32 FILLER_344_664 ();
 FILLCELL_X32 FILLER_344_696 ();
 FILLCELL_X32 FILLER_344_728 ();
 FILLCELL_X32 FILLER_344_760 ();
 FILLCELL_X32 FILLER_344_792 ();
 FILLCELL_X32 FILLER_344_824 ();
 FILLCELL_X32 FILLER_344_856 ();
 FILLCELL_X32 FILLER_344_888 ();
 FILLCELL_X32 FILLER_344_920 ();
 FILLCELL_X32 FILLER_344_952 ();
 FILLCELL_X32 FILLER_344_984 ();
 FILLCELL_X32 FILLER_344_1016 ();
 FILLCELL_X32 FILLER_344_1048 ();
 FILLCELL_X32 FILLER_344_1080 ();
 FILLCELL_X32 FILLER_344_1112 ();
 FILLCELL_X32 FILLER_344_1144 ();
 FILLCELL_X32 FILLER_344_1176 ();
 FILLCELL_X32 FILLER_344_1208 ();
 FILLCELL_X32 FILLER_344_1240 ();
 FILLCELL_X32 FILLER_344_1272 ();
 FILLCELL_X32 FILLER_344_1304 ();
 FILLCELL_X32 FILLER_344_1336 ();
 FILLCELL_X32 FILLER_344_1368 ();
 FILLCELL_X32 FILLER_344_1400 ();
 FILLCELL_X32 FILLER_344_1432 ();
 FILLCELL_X32 FILLER_344_1464 ();
 FILLCELL_X32 FILLER_344_1496 ();
 FILLCELL_X32 FILLER_344_1528 ();
 FILLCELL_X32 FILLER_344_1560 ();
 FILLCELL_X32 FILLER_344_1592 ();
 FILLCELL_X32 FILLER_344_1624 ();
 FILLCELL_X32 FILLER_344_1656 ();
 FILLCELL_X32 FILLER_344_1688 ();
 FILLCELL_X32 FILLER_344_1720 ();
 FILLCELL_X32 FILLER_344_1752 ();
 FILLCELL_X32 FILLER_344_1784 ();
 FILLCELL_X32 FILLER_344_1816 ();
 FILLCELL_X32 FILLER_344_1848 ();
 FILLCELL_X8 FILLER_344_1880 ();
 FILLCELL_X4 FILLER_344_1888 ();
 FILLCELL_X2 FILLER_344_1892 ();
 FILLCELL_X32 FILLER_344_1895 ();
 FILLCELL_X32 FILLER_344_1927 ();
 FILLCELL_X32 FILLER_344_1959 ();
 FILLCELL_X32 FILLER_344_1991 ();
 FILLCELL_X32 FILLER_344_2023 ();
 FILLCELL_X32 FILLER_344_2055 ();
 FILLCELL_X32 FILLER_344_2087 ();
 FILLCELL_X32 FILLER_344_2119 ();
 FILLCELL_X32 FILLER_344_2151 ();
 FILLCELL_X32 FILLER_344_2183 ();
 FILLCELL_X32 FILLER_344_2215 ();
 FILLCELL_X32 FILLER_344_2247 ();
 FILLCELL_X32 FILLER_344_2279 ();
 FILLCELL_X32 FILLER_344_2311 ();
 FILLCELL_X32 FILLER_344_2343 ();
 FILLCELL_X32 FILLER_344_2375 ();
 FILLCELL_X32 FILLER_344_2407 ();
 FILLCELL_X32 FILLER_344_2439 ();
 FILLCELL_X32 FILLER_344_2471 ();
 FILLCELL_X32 FILLER_344_2503 ();
 FILLCELL_X32 FILLER_344_2535 ();
 FILLCELL_X32 FILLER_344_2567 ();
 FILLCELL_X32 FILLER_344_2599 ();
 FILLCELL_X32 FILLER_344_2631 ();
 FILLCELL_X32 FILLER_344_2663 ();
 FILLCELL_X32 FILLER_344_2695 ();
 FILLCELL_X32 FILLER_344_2727 ();
 FILLCELL_X32 FILLER_344_2759 ();
 FILLCELL_X32 FILLER_344_2791 ();
 FILLCELL_X32 FILLER_344_2823 ();
 FILLCELL_X32 FILLER_344_2855 ();
 FILLCELL_X32 FILLER_344_2887 ();
 FILLCELL_X32 FILLER_344_2919 ();
 FILLCELL_X32 FILLER_344_2951 ();
 FILLCELL_X32 FILLER_344_2983 ();
 FILLCELL_X32 FILLER_344_3015 ();
 FILLCELL_X32 FILLER_344_3047 ();
 FILLCELL_X32 FILLER_344_3079 ();
 FILLCELL_X32 FILLER_344_3111 ();
 FILLCELL_X8 FILLER_344_3143 ();
 FILLCELL_X4 FILLER_344_3151 ();
 FILLCELL_X2 FILLER_344_3155 ();
 FILLCELL_X32 FILLER_344_3158 ();
 FILLCELL_X32 FILLER_344_3190 ();
 FILLCELL_X32 FILLER_344_3222 ();
 FILLCELL_X32 FILLER_344_3254 ();
 FILLCELL_X32 FILLER_344_3286 ();
 FILLCELL_X32 FILLER_344_3318 ();
 FILLCELL_X32 FILLER_344_3350 ();
 FILLCELL_X32 FILLER_344_3382 ();
 FILLCELL_X32 FILLER_344_3414 ();
 FILLCELL_X32 FILLER_344_3446 ();
 FILLCELL_X32 FILLER_344_3478 ();
 FILLCELL_X32 FILLER_344_3510 ();
 FILLCELL_X32 FILLER_344_3542 ();
 FILLCELL_X32 FILLER_344_3574 ();
 FILLCELL_X32 FILLER_344_3606 ();
 FILLCELL_X32 FILLER_344_3638 ();
 FILLCELL_X32 FILLER_344_3670 ();
 FILLCELL_X32 FILLER_344_3702 ();
 FILLCELL_X4 FILLER_344_3734 ();
 FILLCELL_X32 FILLER_345_1 ();
 FILLCELL_X32 FILLER_345_33 ();
 FILLCELL_X32 FILLER_345_65 ();
 FILLCELL_X32 FILLER_345_97 ();
 FILLCELL_X32 FILLER_345_129 ();
 FILLCELL_X32 FILLER_345_161 ();
 FILLCELL_X32 FILLER_345_193 ();
 FILLCELL_X32 FILLER_345_225 ();
 FILLCELL_X32 FILLER_345_257 ();
 FILLCELL_X32 FILLER_345_289 ();
 FILLCELL_X32 FILLER_345_321 ();
 FILLCELL_X32 FILLER_345_353 ();
 FILLCELL_X32 FILLER_345_385 ();
 FILLCELL_X32 FILLER_345_417 ();
 FILLCELL_X32 FILLER_345_449 ();
 FILLCELL_X32 FILLER_345_481 ();
 FILLCELL_X32 FILLER_345_513 ();
 FILLCELL_X32 FILLER_345_545 ();
 FILLCELL_X32 FILLER_345_577 ();
 FILLCELL_X32 FILLER_345_609 ();
 FILLCELL_X32 FILLER_345_641 ();
 FILLCELL_X32 FILLER_345_673 ();
 FILLCELL_X32 FILLER_345_705 ();
 FILLCELL_X32 FILLER_345_737 ();
 FILLCELL_X32 FILLER_345_769 ();
 FILLCELL_X32 FILLER_345_801 ();
 FILLCELL_X32 FILLER_345_833 ();
 FILLCELL_X32 FILLER_345_865 ();
 FILLCELL_X32 FILLER_345_897 ();
 FILLCELL_X32 FILLER_345_929 ();
 FILLCELL_X32 FILLER_345_961 ();
 FILLCELL_X32 FILLER_345_993 ();
 FILLCELL_X32 FILLER_345_1025 ();
 FILLCELL_X32 FILLER_345_1057 ();
 FILLCELL_X32 FILLER_345_1089 ();
 FILLCELL_X32 FILLER_345_1121 ();
 FILLCELL_X32 FILLER_345_1153 ();
 FILLCELL_X32 FILLER_345_1185 ();
 FILLCELL_X32 FILLER_345_1217 ();
 FILLCELL_X8 FILLER_345_1249 ();
 FILLCELL_X4 FILLER_345_1257 ();
 FILLCELL_X2 FILLER_345_1261 ();
 FILLCELL_X32 FILLER_345_1264 ();
 FILLCELL_X32 FILLER_345_1296 ();
 FILLCELL_X32 FILLER_345_1328 ();
 FILLCELL_X32 FILLER_345_1360 ();
 FILLCELL_X32 FILLER_345_1392 ();
 FILLCELL_X32 FILLER_345_1424 ();
 FILLCELL_X32 FILLER_345_1456 ();
 FILLCELL_X32 FILLER_345_1488 ();
 FILLCELL_X32 FILLER_345_1520 ();
 FILLCELL_X32 FILLER_345_1552 ();
 FILLCELL_X32 FILLER_345_1584 ();
 FILLCELL_X32 FILLER_345_1616 ();
 FILLCELL_X32 FILLER_345_1648 ();
 FILLCELL_X32 FILLER_345_1680 ();
 FILLCELL_X32 FILLER_345_1712 ();
 FILLCELL_X32 FILLER_345_1744 ();
 FILLCELL_X32 FILLER_345_1776 ();
 FILLCELL_X32 FILLER_345_1808 ();
 FILLCELL_X32 FILLER_345_1840 ();
 FILLCELL_X32 FILLER_345_1872 ();
 FILLCELL_X32 FILLER_345_1904 ();
 FILLCELL_X32 FILLER_345_1936 ();
 FILLCELL_X32 FILLER_345_1968 ();
 FILLCELL_X32 FILLER_345_2000 ();
 FILLCELL_X32 FILLER_345_2032 ();
 FILLCELL_X32 FILLER_345_2064 ();
 FILLCELL_X32 FILLER_345_2096 ();
 FILLCELL_X32 FILLER_345_2128 ();
 FILLCELL_X32 FILLER_345_2160 ();
 FILLCELL_X32 FILLER_345_2192 ();
 FILLCELL_X32 FILLER_345_2224 ();
 FILLCELL_X32 FILLER_345_2256 ();
 FILLCELL_X32 FILLER_345_2288 ();
 FILLCELL_X32 FILLER_345_2320 ();
 FILLCELL_X32 FILLER_345_2352 ();
 FILLCELL_X32 FILLER_345_2384 ();
 FILLCELL_X32 FILLER_345_2416 ();
 FILLCELL_X32 FILLER_345_2448 ();
 FILLCELL_X32 FILLER_345_2480 ();
 FILLCELL_X8 FILLER_345_2512 ();
 FILLCELL_X4 FILLER_345_2520 ();
 FILLCELL_X2 FILLER_345_2524 ();
 FILLCELL_X32 FILLER_345_2527 ();
 FILLCELL_X32 FILLER_345_2559 ();
 FILLCELL_X32 FILLER_345_2591 ();
 FILLCELL_X32 FILLER_345_2623 ();
 FILLCELL_X32 FILLER_345_2655 ();
 FILLCELL_X32 FILLER_345_2687 ();
 FILLCELL_X32 FILLER_345_2719 ();
 FILLCELL_X32 FILLER_345_2751 ();
 FILLCELL_X32 FILLER_345_2783 ();
 FILLCELL_X32 FILLER_345_2815 ();
 FILLCELL_X32 FILLER_345_2847 ();
 FILLCELL_X32 FILLER_345_2879 ();
 FILLCELL_X32 FILLER_345_2911 ();
 FILLCELL_X32 FILLER_345_2943 ();
 FILLCELL_X32 FILLER_345_2975 ();
 FILLCELL_X32 FILLER_345_3007 ();
 FILLCELL_X32 FILLER_345_3039 ();
 FILLCELL_X32 FILLER_345_3071 ();
 FILLCELL_X32 FILLER_345_3103 ();
 FILLCELL_X32 FILLER_345_3135 ();
 FILLCELL_X32 FILLER_345_3167 ();
 FILLCELL_X32 FILLER_345_3199 ();
 FILLCELL_X32 FILLER_345_3231 ();
 FILLCELL_X32 FILLER_345_3263 ();
 FILLCELL_X32 FILLER_345_3295 ();
 FILLCELL_X32 FILLER_345_3327 ();
 FILLCELL_X32 FILLER_345_3359 ();
 FILLCELL_X32 FILLER_345_3391 ();
 FILLCELL_X32 FILLER_345_3423 ();
 FILLCELL_X32 FILLER_345_3455 ();
 FILLCELL_X32 FILLER_345_3487 ();
 FILLCELL_X32 FILLER_345_3519 ();
 FILLCELL_X32 FILLER_345_3551 ();
 FILLCELL_X32 FILLER_345_3583 ();
 FILLCELL_X32 FILLER_345_3615 ();
 FILLCELL_X32 FILLER_345_3647 ();
 FILLCELL_X32 FILLER_345_3679 ();
 FILLCELL_X16 FILLER_345_3711 ();
 FILLCELL_X8 FILLER_345_3727 ();
 FILLCELL_X2 FILLER_345_3735 ();
 FILLCELL_X1 FILLER_345_3737 ();
 FILLCELL_X32 FILLER_346_1 ();
 FILLCELL_X32 FILLER_346_33 ();
 FILLCELL_X32 FILLER_346_65 ();
 FILLCELL_X32 FILLER_346_97 ();
 FILLCELL_X32 FILLER_346_129 ();
 FILLCELL_X32 FILLER_346_161 ();
 FILLCELL_X32 FILLER_346_193 ();
 FILLCELL_X32 FILLER_346_225 ();
 FILLCELL_X32 FILLER_346_257 ();
 FILLCELL_X32 FILLER_346_289 ();
 FILLCELL_X32 FILLER_346_321 ();
 FILLCELL_X32 FILLER_346_353 ();
 FILLCELL_X32 FILLER_346_385 ();
 FILLCELL_X32 FILLER_346_417 ();
 FILLCELL_X32 FILLER_346_449 ();
 FILLCELL_X32 FILLER_346_481 ();
 FILLCELL_X32 FILLER_346_513 ();
 FILLCELL_X32 FILLER_346_545 ();
 FILLCELL_X32 FILLER_346_577 ();
 FILLCELL_X16 FILLER_346_609 ();
 FILLCELL_X4 FILLER_346_625 ();
 FILLCELL_X2 FILLER_346_629 ();
 FILLCELL_X32 FILLER_346_632 ();
 FILLCELL_X32 FILLER_346_664 ();
 FILLCELL_X32 FILLER_346_696 ();
 FILLCELL_X32 FILLER_346_728 ();
 FILLCELL_X32 FILLER_346_760 ();
 FILLCELL_X32 FILLER_346_792 ();
 FILLCELL_X32 FILLER_346_824 ();
 FILLCELL_X32 FILLER_346_856 ();
 FILLCELL_X32 FILLER_346_888 ();
 FILLCELL_X32 FILLER_346_920 ();
 FILLCELL_X32 FILLER_346_952 ();
 FILLCELL_X32 FILLER_346_984 ();
 FILLCELL_X32 FILLER_346_1016 ();
 FILLCELL_X32 FILLER_346_1048 ();
 FILLCELL_X32 FILLER_346_1080 ();
 FILLCELL_X32 FILLER_346_1112 ();
 FILLCELL_X32 FILLER_346_1144 ();
 FILLCELL_X32 FILLER_346_1176 ();
 FILLCELL_X32 FILLER_346_1208 ();
 FILLCELL_X32 FILLER_346_1240 ();
 FILLCELL_X32 FILLER_346_1272 ();
 FILLCELL_X32 FILLER_346_1304 ();
 FILLCELL_X32 FILLER_346_1336 ();
 FILLCELL_X32 FILLER_346_1368 ();
 FILLCELL_X32 FILLER_346_1400 ();
 FILLCELL_X32 FILLER_346_1432 ();
 FILLCELL_X32 FILLER_346_1464 ();
 FILLCELL_X32 FILLER_346_1496 ();
 FILLCELL_X32 FILLER_346_1528 ();
 FILLCELL_X32 FILLER_346_1560 ();
 FILLCELL_X32 FILLER_346_1592 ();
 FILLCELL_X32 FILLER_346_1624 ();
 FILLCELL_X32 FILLER_346_1656 ();
 FILLCELL_X32 FILLER_346_1688 ();
 FILLCELL_X32 FILLER_346_1720 ();
 FILLCELL_X32 FILLER_346_1752 ();
 FILLCELL_X32 FILLER_346_1784 ();
 FILLCELL_X32 FILLER_346_1816 ();
 FILLCELL_X32 FILLER_346_1848 ();
 FILLCELL_X8 FILLER_346_1880 ();
 FILLCELL_X4 FILLER_346_1888 ();
 FILLCELL_X2 FILLER_346_1892 ();
 FILLCELL_X32 FILLER_346_1895 ();
 FILLCELL_X32 FILLER_346_1927 ();
 FILLCELL_X32 FILLER_346_1959 ();
 FILLCELL_X32 FILLER_346_1991 ();
 FILLCELL_X32 FILLER_346_2023 ();
 FILLCELL_X32 FILLER_346_2055 ();
 FILLCELL_X32 FILLER_346_2087 ();
 FILLCELL_X32 FILLER_346_2119 ();
 FILLCELL_X32 FILLER_346_2151 ();
 FILLCELL_X32 FILLER_346_2183 ();
 FILLCELL_X32 FILLER_346_2215 ();
 FILLCELL_X32 FILLER_346_2247 ();
 FILLCELL_X32 FILLER_346_2279 ();
 FILLCELL_X32 FILLER_346_2311 ();
 FILLCELL_X32 FILLER_346_2343 ();
 FILLCELL_X32 FILLER_346_2375 ();
 FILLCELL_X32 FILLER_346_2407 ();
 FILLCELL_X32 FILLER_346_2439 ();
 FILLCELL_X32 FILLER_346_2471 ();
 FILLCELL_X32 FILLER_346_2503 ();
 FILLCELL_X32 FILLER_346_2535 ();
 FILLCELL_X32 FILLER_346_2567 ();
 FILLCELL_X32 FILLER_346_2599 ();
 FILLCELL_X32 FILLER_346_2631 ();
 FILLCELL_X32 FILLER_346_2663 ();
 FILLCELL_X32 FILLER_346_2695 ();
 FILLCELL_X32 FILLER_346_2727 ();
 FILLCELL_X32 FILLER_346_2759 ();
 FILLCELL_X32 FILLER_346_2791 ();
 FILLCELL_X32 FILLER_346_2823 ();
 FILLCELL_X32 FILLER_346_2855 ();
 FILLCELL_X32 FILLER_346_2887 ();
 FILLCELL_X32 FILLER_346_2919 ();
 FILLCELL_X32 FILLER_346_2951 ();
 FILLCELL_X32 FILLER_346_2983 ();
 FILLCELL_X32 FILLER_346_3015 ();
 FILLCELL_X32 FILLER_346_3047 ();
 FILLCELL_X32 FILLER_346_3079 ();
 FILLCELL_X32 FILLER_346_3111 ();
 FILLCELL_X8 FILLER_346_3143 ();
 FILLCELL_X4 FILLER_346_3151 ();
 FILLCELL_X2 FILLER_346_3155 ();
 FILLCELL_X32 FILLER_346_3158 ();
 FILLCELL_X32 FILLER_346_3190 ();
 FILLCELL_X32 FILLER_346_3222 ();
 FILLCELL_X32 FILLER_346_3254 ();
 FILLCELL_X32 FILLER_346_3286 ();
 FILLCELL_X32 FILLER_346_3318 ();
 FILLCELL_X32 FILLER_346_3350 ();
 FILLCELL_X32 FILLER_346_3382 ();
 FILLCELL_X32 FILLER_346_3414 ();
 FILLCELL_X32 FILLER_346_3446 ();
 FILLCELL_X32 FILLER_346_3478 ();
 FILLCELL_X32 FILLER_346_3510 ();
 FILLCELL_X32 FILLER_346_3542 ();
 FILLCELL_X32 FILLER_346_3574 ();
 FILLCELL_X32 FILLER_346_3606 ();
 FILLCELL_X32 FILLER_346_3638 ();
 FILLCELL_X32 FILLER_346_3670 ();
 FILLCELL_X32 FILLER_346_3702 ();
 FILLCELL_X4 FILLER_346_3734 ();
 FILLCELL_X32 FILLER_347_1 ();
 FILLCELL_X32 FILLER_347_33 ();
 FILLCELL_X32 FILLER_347_65 ();
 FILLCELL_X32 FILLER_347_97 ();
 FILLCELL_X32 FILLER_347_129 ();
 FILLCELL_X32 FILLER_347_161 ();
 FILLCELL_X32 FILLER_347_193 ();
 FILLCELL_X32 FILLER_347_225 ();
 FILLCELL_X32 FILLER_347_257 ();
 FILLCELL_X32 FILLER_347_289 ();
 FILLCELL_X32 FILLER_347_321 ();
 FILLCELL_X32 FILLER_347_353 ();
 FILLCELL_X32 FILLER_347_385 ();
 FILLCELL_X32 FILLER_347_417 ();
 FILLCELL_X32 FILLER_347_449 ();
 FILLCELL_X32 FILLER_347_481 ();
 FILLCELL_X32 FILLER_347_513 ();
 FILLCELL_X32 FILLER_347_545 ();
 FILLCELL_X32 FILLER_347_577 ();
 FILLCELL_X32 FILLER_347_609 ();
 FILLCELL_X32 FILLER_347_641 ();
 FILLCELL_X32 FILLER_347_673 ();
 FILLCELL_X32 FILLER_347_705 ();
 FILLCELL_X32 FILLER_347_737 ();
 FILLCELL_X32 FILLER_347_769 ();
 FILLCELL_X32 FILLER_347_801 ();
 FILLCELL_X32 FILLER_347_833 ();
 FILLCELL_X32 FILLER_347_865 ();
 FILLCELL_X32 FILLER_347_897 ();
 FILLCELL_X32 FILLER_347_929 ();
 FILLCELL_X32 FILLER_347_961 ();
 FILLCELL_X32 FILLER_347_993 ();
 FILLCELL_X32 FILLER_347_1025 ();
 FILLCELL_X32 FILLER_347_1057 ();
 FILLCELL_X32 FILLER_347_1089 ();
 FILLCELL_X32 FILLER_347_1121 ();
 FILLCELL_X32 FILLER_347_1153 ();
 FILLCELL_X32 FILLER_347_1185 ();
 FILLCELL_X32 FILLER_347_1217 ();
 FILLCELL_X8 FILLER_347_1249 ();
 FILLCELL_X4 FILLER_347_1257 ();
 FILLCELL_X2 FILLER_347_1261 ();
 FILLCELL_X32 FILLER_347_1264 ();
 FILLCELL_X32 FILLER_347_1296 ();
 FILLCELL_X32 FILLER_347_1328 ();
 FILLCELL_X32 FILLER_347_1360 ();
 FILLCELL_X32 FILLER_347_1392 ();
 FILLCELL_X32 FILLER_347_1424 ();
 FILLCELL_X32 FILLER_347_1456 ();
 FILLCELL_X32 FILLER_347_1488 ();
 FILLCELL_X32 FILLER_347_1520 ();
 FILLCELL_X32 FILLER_347_1552 ();
 FILLCELL_X32 FILLER_347_1584 ();
 FILLCELL_X32 FILLER_347_1616 ();
 FILLCELL_X32 FILLER_347_1648 ();
 FILLCELL_X32 FILLER_347_1680 ();
 FILLCELL_X32 FILLER_347_1712 ();
 FILLCELL_X32 FILLER_347_1744 ();
 FILLCELL_X32 FILLER_347_1776 ();
 FILLCELL_X32 FILLER_347_1808 ();
 FILLCELL_X32 FILLER_347_1840 ();
 FILLCELL_X32 FILLER_347_1872 ();
 FILLCELL_X32 FILLER_347_1904 ();
 FILLCELL_X32 FILLER_347_1936 ();
 FILLCELL_X32 FILLER_347_1968 ();
 FILLCELL_X32 FILLER_347_2000 ();
 FILLCELL_X32 FILLER_347_2032 ();
 FILLCELL_X32 FILLER_347_2064 ();
 FILLCELL_X32 FILLER_347_2096 ();
 FILLCELL_X32 FILLER_347_2128 ();
 FILLCELL_X32 FILLER_347_2160 ();
 FILLCELL_X32 FILLER_347_2192 ();
 FILLCELL_X32 FILLER_347_2224 ();
 FILLCELL_X32 FILLER_347_2256 ();
 FILLCELL_X32 FILLER_347_2288 ();
 FILLCELL_X32 FILLER_347_2320 ();
 FILLCELL_X32 FILLER_347_2352 ();
 FILLCELL_X32 FILLER_347_2384 ();
 FILLCELL_X32 FILLER_347_2416 ();
 FILLCELL_X32 FILLER_347_2448 ();
 FILLCELL_X32 FILLER_347_2480 ();
 FILLCELL_X8 FILLER_347_2512 ();
 FILLCELL_X4 FILLER_347_2520 ();
 FILLCELL_X2 FILLER_347_2524 ();
 FILLCELL_X32 FILLER_347_2527 ();
 FILLCELL_X32 FILLER_347_2559 ();
 FILLCELL_X32 FILLER_347_2591 ();
 FILLCELL_X32 FILLER_347_2623 ();
 FILLCELL_X32 FILLER_347_2655 ();
 FILLCELL_X32 FILLER_347_2687 ();
 FILLCELL_X32 FILLER_347_2719 ();
 FILLCELL_X32 FILLER_347_2751 ();
 FILLCELL_X32 FILLER_347_2783 ();
 FILLCELL_X32 FILLER_347_2815 ();
 FILLCELL_X32 FILLER_347_2847 ();
 FILLCELL_X32 FILLER_347_2879 ();
 FILLCELL_X32 FILLER_347_2911 ();
 FILLCELL_X32 FILLER_347_2943 ();
 FILLCELL_X32 FILLER_347_2975 ();
 FILLCELL_X32 FILLER_347_3007 ();
 FILLCELL_X32 FILLER_347_3039 ();
 FILLCELL_X32 FILLER_347_3071 ();
 FILLCELL_X32 FILLER_347_3103 ();
 FILLCELL_X32 FILLER_347_3135 ();
 FILLCELL_X32 FILLER_347_3167 ();
 FILLCELL_X32 FILLER_347_3199 ();
 FILLCELL_X32 FILLER_347_3231 ();
 FILLCELL_X32 FILLER_347_3263 ();
 FILLCELL_X32 FILLER_347_3295 ();
 FILLCELL_X32 FILLER_347_3327 ();
 FILLCELL_X32 FILLER_347_3359 ();
 FILLCELL_X32 FILLER_347_3391 ();
 FILLCELL_X32 FILLER_347_3423 ();
 FILLCELL_X32 FILLER_347_3455 ();
 FILLCELL_X32 FILLER_347_3487 ();
 FILLCELL_X32 FILLER_347_3519 ();
 FILLCELL_X32 FILLER_347_3551 ();
 FILLCELL_X32 FILLER_347_3583 ();
 FILLCELL_X32 FILLER_347_3615 ();
 FILLCELL_X32 FILLER_347_3647 ();
 FILLCELL_X32 FILLER_347_3679 ();
 FILLCELL_X16 FILLER_347_3711 ();
 FILLCELL_X8 FILLER_347_3727 ();
 FILLCELL_X2 FILLER_347_3735 ();
 FILLCELL_X1 FILLER_347_3737 ();
 FILLCELL_X32 FILLER_348_1 ();
 FILLCELL_X32 FILLER_348_33 ();
 FILLCELL_X32 FILLER_348_65 ();
 FILLCELL_X32 FILLER_348_97 ();
 FILLCELL_X32 FILLER_348_129 ();
 FILLCELL_X32 FILLER_348_161 ();
 FILLCELL_X32 FILLER_348_193 ();
 FILLCELL_X32 FILLER_348_225 ();
 FILLCELL_X32 FILLER_348_257 ();
 FILLCELL_X32 FILLER_348_289 ();
 FILLCELL_X32 FILLER_348_321 ();
 FILLCELL_X32 FILLER_348_353 ();
 FILLCELL_X32 FILLER_348_385 ();
 FILLCELL_X32 FILLER_348_417 ();
 FILLCELL_X32 FILLER_348_449 ();
 FILLCELL_X32 FILLER_348_481 ();
 FILLCELL_X32 FILLER_348_513 ();
 FILLCELL_X32 FILLER_348_545 ();
 FILLCELL_X32 FILLER_348_577 ();
 FILLCELL_X16 FILLER_348_609 ();
 FILLCELL_X4 FILLER_348_625 ();
 FILLCELL_X2 FILLER_348_629 ();
 FILLCELL_X32 FILLER_348_632 ();
 FILLCELL_X32 FILLER_348_664 ();
 FILLCELL_X32 FILLER_348_696 ();
 FILLCELL_X32 FILLER_348_728 ();
 FILLCELL_X32 FILLER_348_760 ();
 FILLCELL_X32 FILLER_348_792 ();
 FILLCELL_X32 FILLER_348_824 ();
 FILLCELL_X32 FILLER_348_856 ();
 FILLCELL_X32 FILLER_348_888 ();
 FILLCELL_X32 FILLER_348_920 ();
 FILLCELL_X32 FILLER_348_952 ();
 FILLCELL_X32 FILLER_348_984 ();
 FILLCELL_X32 FILLER_348_1016 ();
 FILLCELL_X32 FILLER_348_1048 ();
 FILLCELL_X32 FILLER_348_1080 ();
 FILLCELL_X32 FILLER_348_1112 ();
 FILLCELL_X32 FILLER_348_1144 ();
 FILLCELL_X32 FILLER_348_1176 ();
 FILLCELL_X32 FILLER_348_1208 ();
 FILLCELL_X32 FILLER_348_1240 ();
 FILLCELL_X32 FILLER_348_1272 ();
 FILLCELL_X32 FILLER_348_1304 ();
 FILLCELL_X32 FILLER_348_1336 ();
 FILLCELL_X32 FILLER_348_1368 ();
 FILLCELL_X32 FILLER_348_1400 ();
 FILLCELL_X32 FILLER_348_1432 ();
 FILLCELL_X32 FILLER_348_1464 ();
 FILLCELL_X32 FILLER_348_1496 ();
 FILLCELL_X32 FILLER_348_1528 ();
 FILLCELL_X32 FILLER_348_1560 ();
 FILLCELL_X32 FILLER_348_1592 ();
 FILLCELL_X32 FILLER_348_1624 ();
 FILLCELL_X32 FILLER_348_1656 ();
 FILLCELL_X32 FILLER_348_1688 ();
 FILLCELL_X32 FILLER_348_1720 ();
 FILLCELL_X32 FILLER_348_1752 ();
 FILLCELL_X32 FILLER_348_1784 ();
 FILLCELL_X32 FILLER_348_1816 ();
 FILLCELL_X32 FILLER_348_1848 ();
 FILLCELL_X8 FILLER_348_1880 ();
 FILLCELL_X4 FILLER_348_1888 ();
 FILLCELL_X2 FILLER_348_1892 ();
 FILLCELL_X32 FILLER_348_1895 ();
 FILLCELL_X32 FILLER_348_1927 ();
 FILLCELL_X32 FILLER_348_1959 ();
 FILLCELL_X32 FILLER_348_1991 ();
 FILLCELL_X32 FILLER_348_2023 ();
 FILLCELL_X32 FILLER_348_2055 ();
 FILLCELL_X32 FILLER_348_2087 ();
 FILLCELL_X32 FILLER_348_2119 ();
 FILLCELL_X32 FILLER_348_2151 ();
 FILLCELL_X32 FILLER_348_2183 ();
 FILLCELL_X32 FILLER_348_2215 ();
 FILLCELL_X32 FILLER_348_2247 ();
 FILLCELL_X32 FILLER_348_2279 ();
 FILLCELL_X32 FILLER_348_2311 ();
 FILLCELL_X32 FILLER_348_2343 ();
 FILLCELL_X32 FILLER_348_2375 ();
 FILLCELL_X32 FILLER_348_2407 ();
 FILLCELL_X32 FILLER_348_2439 ();
 FILLCELL_X32 FILLER_348_2471 ();
 FILLCELL_X32 FILLER_348_2503 ();
 FILLCELL_X32 FILLER_348_2535 ();
 FILLCELL_X32 FILLER_348_2567 ();
 FILLCELL_X32 FILLER_348_2599 ();
 FILLCELL_X32 FILLER_348_2631 ();
 FILLCELL_X32 FILLER_348_2663 ();
 FILLCELL_X32 FILLER_348_2695 ();
 FILLCELL_X32 FILLER_348_2727 ();
 FILLCELL_X32 FILLER_348_2759 ();
 FILLCELL_X32 FILLER_348_2791 ();
 FILLCELL_X32 FILLER_348_2823 ();
 FILLCELL_X32 FILLER_348_2855 ();
 FILLCELL_X32 FILLER_348_2887 ();
 FILLCELL_X32 FILLER_348_2919 ();
 FILLCELL_X32 FILLER_348_2951 ();
 FILLCELL_X32 FILLER_348_2983 ();
 FILLCELL_X32 FILLER_348_3015 ();
 FILLCELL_X32 FILLER_348_3047 ();
 FILLCELL_X32 FILLER_348_3079 ();
 FILLCELL_X32 FILLER_348_3111 ();
 FILLCELL_X8 FILLER_348_3143 ();
 FILLCELL_X4 FILLER_348_3151 ();
 FILLCELL_X2 FILLER_348_3155 ();
 FILLCELL_X32 FILLER_348_3158 ();
 FILLCELL_X32 FILLER_348_3190 ();
 FILLCELL_X32 FILLER_348_3222 ();
 FILLCELL_X32 FILLER_348_3254 ();
 FILLCELL_X32 FILLER_348_3286 ();
 FILLCELL_X32 FILLER_348_3318 ();
 FILLCELL_X32 FILLER_348_3350 ();
 FILLCELL_X32 FILLER_348_3382 ();
 FILLCELL_X32 FILLER_348_3414 ();
 FILLCELL_X32 FILLER_348_3446 ();
 FILLCELL_X32 FILLER_348_3478 ();
 FILLCELL_X32 FILLER_348_3510 ();
 FILLCELL_X32 FILLER_348_3542 ();
 FILLCELL_X32 FILLER_348_3574 ();
 FILLCELL_X32 FILLER_348_3606 ();
 FILLCELL_X32 FILLER_348_3638 ();
 FILLCELL_X32 FILLER_348_3670 ();
 FILLCELL_X32 FILLER_348_3702 ();
 FILLCELL_X4 FILLER_348_3734 ();
 FILLCELL_X32 FILLER_349_1 ();
 FILLCELL_X32 FILLER_349_33 ();
 FILLCELL_X32 FILLER_349_65 ();
 FILLCELL_X32 FILLER_349_97 ();
 FILLCELL_X32 FILLER_349_129 ();
 FILLCELL_X32 FILLER_349_161 ();
 FILLCELL_X32 FILLER_349_193 ();
 FILLCELL_X32 FILLER_349_225 ();
 FILLCELL_X32 FILLER_349_257 ();
 FILLCELL_X32 FILLER_349_289 ();
 FILLCELL_X32 FILLER_349_321 ();
 FILLCELL_X32 FILLER_349_353 ();
 FILLCELL_X32 FILLER_349_385 ();
 FILLCELL_X32 FILLER_349_417 ();
 FILLCELL_X32 FILLER_349_449 ();
 FILLCELL_X32 FILLER_349_481 ();
 FILLCELL_X32 FILLER_349_513 ();
 FILLCELL_X32 FILLER_349_545 ();
 FILLCELL_X32 FILLER_349_577 ();
 FILLCELL_X32 FILLER_349_609 ();
 FILLCELL_X32 FILLER_349_641 ();
 FILLCELL_X32 FILLER_349_673 ();
 FILLCELL_X32 FILLER_349_705 ();
 FILLCELL_X32 FILLER_349_737 ();
 FILLCELL_X32 FILLER_349_769 ();
 FILLCELL_X32 FILLER_349_801 ();
 FILLCELL_X32 FILLER_349_833 ();
 FILLCELL_X32 FILLER_349_865 ();
 FILLCELL_X32 FILLER_349_897 ();
 FILLCELL_X32 FILLER_349_929 ();
 FILLCELL_X32 FILLER_349_961 ();
 FILLCELL_X32 FILLER_349_993 ();
 FILLCELL_X32 FILLER_349_1025 ();
 FILLCELL_X32 FILLER_349_1057 ();
 FILLCELL_X32 FILLER_349_1089 ();
 FILLCELL_X32 FILLER_349_1121 ();
 FILLCELL_X32 FILLER_349_1153 ();
 FILLCELL_X32 FILLER_349_1185 ();
 FILLCELL_X32 FILLER_349_1217 ();
 FILLCELL_X8 FILLER_349_1249 ();
 FILLCELL_X4 FILLER_349_1257 ();
 FILLCELL_X2 FILLER_349_1261 ();
 FILLCELL_X32 FILLER_349_1264 ();
 FILLCELL_X32 FILLER_349_1296 ();
 FILLCELL_X32 FILLER_349_1328 ();
 FILLCELL_X32 FILLER_349_1360 ();
 FILLCELL_X32 FILLER_349_1392 ();
 FILLCELL_X32 FILLER_349_1424 ();
 FILLCELL_X32 FILLER_349_1456 ();
 FILLCELL_X32 FILLER_349_1488 ();
 FILLCELL_X32 FILLER_349_1520 ();
 FILLCELL_X32 FILLER_349_1552 ();
 FILLCELL_X32 FILLER_349_1584 ();
 FILLCELL_X32 FILLER_349_1616 ();
 FILLCELL_X32 FILLER_349_1648 ();
 FILLCELL_X32 FILLER_349_1680 ();
 FILLCELL_X32 FILLER_349_1712 ();
 FILLCELL_X32 FILLER_349_1744 ();
 FILLCELL_X32 FILLER_349_1776 ();
 FILLCELL_X32 FILLER_349_1808 ();
 FILLCELL_X32 FILLER_349_1840 ();
 FILLCELL_X32 FILLER_349_1872 ();
 FILLCELL_X32 FILLER_349_1904 ();
 FILLCELL_X32 FILLER_349_1936 ();
 FILLCELL_X32 FILLER_349_1968 ();
 FILLCELL_X32 FILLER_349_2000 ();
 FILLCELL_X32 FILLER_349_2032 ();
 FILLCELL_X32 FILLER_349_2064 ();
 FILLCELL_X32 FILLER_349_2096 ();
 FILLCELL_X32 FILLER_349_2128 ();
 FILLCELL_X32 FILLER_349_2160 ();
 FILLCELL_X32 FILLER_349_2192 ();
 FILLCELL_X32 FILLER_349_2224 ();
 FILLCELL_X32 FILLER_349_2256 ();
 FILLCELL_X32 FILLER_349_2288 ();
 FILLCELL_X32 FILLER_349_2320 ();
 FILLCELL_X32 FILLER_349_2352 ();
 FILLCELL_X32 FILLER_349_2384 ();
 FILLCELL_X32 FILLER_349_2416 ();
 FILLCELL_X32 FILLER_349_2448 ();
 FILLCELL_X32 FILLER_349_2480 ();
 FILLCELL_X8 FILLER_349_2512 ();
 FILLCELL_X4 FILLER_349_2520 ();
 FILLCELL_X2 FILLER_349_2524 ();
 FILLCELL_X32 FILLER_349_2527 ();
 FILLCELL_X32 FILLER_349_2559 ();
 FILLCELL_X32 FILLER_349_2591 ();
 FILLCELL_X32 FILLER_349_2623 ();
 FILLCELL_X32 FILLER_349_2655 ();
 FILLCELL_X32 FILLER_349_2687 ();
 FILLCELL_X32 FILLER_349_2719 ();
 FILLCELL_X32 FILLER_349_2751 ();
 FILLCELL_X32 FILLER_349_2783 ();
 FILLCELL_X32 FILLER_349_2815 ();
 FILLCELL_X32 FILLER_349_2847 ();
 FILLCELL_X32 FILLER_349_2879 ();
 FILLCELL_X32 FILLER_349_2911 ();
 FILLCELL_X32 FILLER_349_2943 ();
 FILLCELL_X32 FILLER_349_2975 ();
 FILLCELL_X32 FILLER_349_3007 ();
 FILLCELL_X32 FILLER_349_3039 ();
 FILLCELL_X32 FILLER_349_3071 ();
 FILLCELL_X32 FILLER_349_3103 ();
 FILLCELL_X32 FILLER_349_3135 ();
 FILLCELL_X32 FILLER_349_3167 ();
 FILLCELL_X32 FILLER_349_3199 ();
 FILLCELL_X32 FILLER_349_3231 ();
 FILLCELL_X32 FILLER_349_3263 ();
 FILLCELL_X32 FILLER_349_3295 ();
 FILLCELL_X32 FILLER_349_3327 ();
 FILLCELL_X32 FILLER_349_3359 ();
 FILLCELL_X32 FILLER_349_3391 ();
 FILLCELL_X32 FILLER_349_3423 ();
 FILLCELL_X32 FILLER_349_3455 ();
 FILLCELL_X32 FILLER_349_3487 ();
 FILLCELL_X32 FILLER_349_3519 ();
 FILLCELL_X32 FILLER_349_3551 ();
 FILLCELL_X32 FILLER_349_3583 ();
 FILLCELL_X32 FILLER_349_3615 ();
 FILLCELL_X32 FILLER_349_3647 ();
 FILLCELL_X32 FILLER_349_3679 ();
 FILLCELL_X16 FILLER_349_3711 ();
 FILLCELL_X8 FILLER_349_3727 ();
 FILLCELL_X2 FILLER_349_3735 ();
 FILLCELL_X1 FILLER_349_3737 ();
 FILLCELL_X32 FILLER_350_1 ();
 FILLCELL_X32 FILLER_350_33 ();
 FILLCELL_X32 FILLER_350_65 ();
 FILLCELL_X32 FILLER_350_97 ();
 FILLCELL_X32 FILLER_350_129 ();
 FILLCELL_X32 FILLER_350_161 ();
 FILLCELL_X32 FILLER_350_193 ();
 FILLCELL_X32 FILLER_350_225 ();
 FILLCELL_X32 FILLER_350_257 ();
 FILLCELL_X32 FILLER_350_289 ();
 FILLCELL_X32 FILLER_350_321 ();
 FILLCELL_X32 FILLER_350_353 ();
 FILLCELL_X32 FILLER_350_385 ();
 FILLCELL_X32 FILLER_350_417 ();
 FILLCELL_X32 FILLER_350_449 ();
 FILLCELL_X32 FILLER_350_481 ();
 FILLCELL_X32 FILLER_350_513 ();
 FILLCELL_X32 FILLER_350_545 ();
 FILLCELL_X32 FILLER_350_577 ();
 FILLCELL_X16 FILLER_350_609 ();
 FILLCELL_X4 FILLER_350_625 ();
 FILLCELL_X2 FILLER_350_629 ();
 FILLCELL_X32 FILLER_350_632 ();
 FILLCELL_X32 FILLER_350_664 ();
 FILLCELL_X32 FILLER_350_696 ();
 FILLCELL_X32 FILLER_350_728 ();
 FILLCELL_X32 FILLER_350_760 ();
 FILLCELL_X32 FILLER_350_792 ();
 FILLCELL_X32 FILLER_350_824 ();
 FILLCELL_X32 FILLER_350_856 ();
 FILLCELL_X32 FILLER_350_888 ();
 FILLCELL_X32 FILLER_350_920 ();
 FILLCELL_X32 FILLER_350_952 ();
 FILLCELL_X32 FILLER_350_984 ();
 FILLCELL_X32 FILLER_350_1016 ();
 FILLCELL_X32 FILLER_350_1048 ();
 FILLCELL_X32 FILLER_350_1080 ();
 FILLCELL_X32 FILLER_350_1112 ();
 FILLCELL_X32 FILLER_350_1144 ();
 FILLCELL_X32 FILLER_350_1176 ();
 FILLCELL_X32 FILLER_350_1208 ();
 FILLCELL_X32 FILLER_350_1240 ();
 FILLCELL_X32 FILLER_350_1272 ();
 FILLCELL_X32 FILLER_350_1304 ();
 FILLCELL_X32 FILLER_350_1336 ();
 FILLCELL_X32 FILLER_350_1368 ();
 FILLCELL_X32 FILLER_350_1400 ();
 FILLCELL_X32 FILLER_350_1432 ();
 FILLCELL_X32 FILLER_350_1464 ();
 FILLCELL_X32 FILLER_350_1496 ();
 FILLCELL_X32 FILLER_350_1528 ();
 FILLCELL_X32 FILLER_350_1560 ();
 FILLCELL_X32 FILLER_350_1592 ();
 FILLCELL_X32 FILLER_350_1624 ();
 FILLCELL_X32 FILLER_350_1656 ();
 FILLCELL_X32 FILLER_350_1688 ();
 FILLCELL_X32 FILLER_350_1720 ();
 FILLCELL_X32 FILLER_350_1752 ();
 FILLCELL_X32 FILLER_350_1784 ();
 FILLCELL_X32 FILLER_350_1816 ();
 FILLCELL_X32 FILLER_350_1848 ();
 FILLCELL_X8 FILLER_350_1880 ();
 FILLCELL_X4 FILLER_350_1888 ();
 FILLCELL_X2 FILLER_350_1892 ();
 FILLCELL_X32 FILLER_350_1895 ();
 FILLCELL_X32 FILLER_350_1927 ();
 FILLCELL_X32 FILLER_350_1959 ();
 FILLCELL_X32 FILLER_350_1991 ();
 FILLCELL_X32 FILLER_350_2023 ();
 FILLCELL_X32 FILLER_350_2055 ();
 FILLCELL_X32 FILLER_350_2087 ();
 FILLCELL_X32 FILLER_350_2119 ();
 FILLCELL_X32 FILLER_350_2151 ();
 FILLCELL_X32 FILLER_350_2183 ();
 FILLCELL_X32 FILLER_350_2215 ();
 FILLCELL_X32 FILLER_350_2247 ();
 FILLCELL_X32 FILLER_350_2279 ();
 FILLCELL_X32 FILLER_350_2311 ();
 FILLCELL_X32 FILLER_350_2343 ();
 FILLCELL_X32 FILLER_350_2375 ();
 FILLCELL_X32 FILLER_350_2407 ();
 FILLCELL_X32 FILLER_350_2439 ();
 FILLCELL_X32 FILLER_350_2471 ();
 FILLCELL_X32 FILLER_350_2503 ();
 FILLCELL_X32 FILLER_350_2535 ();
 FILLCELL_X32 FILLER_350_2567 ();
 FILLCELL_X32 FILLER_350_2599 ();
 FILLCELL_X32 FILLER_350_2631 ();
 FILLCELL_X32 FILLER_350_2663 ();
 FILLCELL_X32 FILLER_350_2695 ();
 FILLCELL_X32 FILLER_350_2727 ();
 FILLCELL_X32 FILLER_350_2759 ();
 FILLCELL_X32 FILLER_350_2791 ();
 FILLCELL_X32 FILLER_350_2823 ();
 FILLCELL_X32 FILLER_350_2855 ();
 FILLCELL_X32 FILLER_350_2887 ();
 FILLCELL_X32 FILLER_350_2919 ();
 FILLCELL_X32 FILLER_350_2951 ();
 FILLCELL_X32 FILLER_350_2983 ();
 FILLCELL_X32 FILLER_350_3015 ();
 FILLCELL_X32 FILLER_350_3047 ();
 FILLCELL_X32 FILLER_350_3079 ();
 FILLCELL_X32 FILLER_350_3111 ();
 FILLCELL_X8 FILLER_350_3143 ();
 FILLCELL_X4 FILLER_350_3151 ();
 FILLCELL_X2 FILLER_350_3155 ();
 FILLCELL_X32 FILLER_350_3158 ();
 FILLCELL_X32 FILLER_350_3190 ();
 FILLCELL_X32 FILLER_350_3222 ();
 FILLCELL_X32 FILLER_350_3254 ();
 FILLCELL_X32 FILLER_350_3286 ();
 FILLCELL_X32 FILLER_350_3318 ();
 FILLCELL_X32 FILLER_350_3350 ();
 FILLCELL_X32 FILLER_350_3382 ();
 FILLCELL_X32 FILLER_350_3414 ();
 FILLCELL_X32 FILLER_350_3446 ();
 FILLCELL_X32 FILLER_350_3478 ();
 FILLCELL_X32 FILLER_350_3510 ();
 FILLCELL_X32 FILLER_350_3542 ();
 FILLCELL_X32 FILLER_350_3574 ();
 FILLCELL_X32 FILLER_350_3606 ();
 FILLCELL_X32 FILLER_350_3638 ();
 FILLCELL_X32 FILLER_350_3670 ();
 FILLCELL_X32 FILLER_350_3702 ();
 FILLCELL_X4 FILLER_350_3734 ();
 FILLCELL_X32 FILLER_351_1 ();
 FILLCELL_X32 FILLER_351_33 ();
 FILLCELL_X32 FILLER_351_65 ();
 FILLCELL_X32 FILLER_351_97 ();
 FILLCELL_X32 FILLER_351_129 ();
 FILLCELL_X32 FILLER_351_161 ();
 FILLCELL_X32 FILLER_351_193 ();
 FILLCELL_X32 FILLER_351_225 ();
 FILLCELL_X32 FILLER_351_257 ();
 FILLCELL_X32 FILLER_351_289 ();
 FILLCELL_X32 FILLER_351_321 ();
 FILLCELL_X32 FILLER_351_353 ();
 FILLCELL_X32 FILLER_351_385 ();
 FILLCELL_X32 FILLER_351_417 ();
 FILLCELL_X32 FILLER_351_449 ();
 FILLCELL_X32 FILLER_351_481 ();
 FILLCELL_X32 FILLER_351_513 ();
 FILLCELL_X32 FILLER_351_545 ();
 FILLCELL_X32 FILLER_351_577 ();
 FILLCELL_X32 FILLER_351_609 ();
 FILLCELL_X32 FILLER_351_641 ();
 FILLCELL_X32 FILLER_351_673 ();
 FILLCELL_X32 FILLER_351_705 ();
 FILLCELL_X32 FILLER_351_737 ();
 FILLCELL_X32 FILLER_351_769 ();
 FILLCELL_X32 FILLER_351_801 ();
 FILLCELL_X32 FILLER_351_833 ();
 FILLCELL_X32 FILLER_351_865 ();
 FILLCELL_X32 FILLER_351_897 ();
 FILLCELL_X32 FILLER_351_929 ();
 FILLCELL_X32 FILLER_351_961 ();
 FILLCELL_X32 FILLER_351_993 ();
 FILLCELL_X32 FILLER_351_1025 ();
 FILLCELL_X32 FILLER_351_1057 ();
 FILLCELL_X32 FILLER_351_1089 ();
 FILLCELL_X32 FILLER_351_1121 ();
 FILLCELL_X32 FILLER_351_1153 ();
 FILLCELL_X32 FILLER_351_1185 ();
 FILLCELL_X32 FILLER_351_1217 ();
 FILLCELL_X8 FILLER_351_1249 ();
 FILLCELL_X4 FILLER_351_1257 ();
 FILLCELL_X2 FILLER_351_1261 ();
 FILLCELL_X32 FILLER_351_1264 ();
 FILLCELL_X32 FILLER_351_1296 ();
 FILLCELL_X32 FILLER_351_1328 ();
 FILLCELL_X32 FILLER_351_1360 ();
 FILLCELL_X32 FILLER_351_1392 ();
 FILLCELL_X32 FILLER_351_1424 ();
 FILLCELL_X32 FILLER_351_1456 ();
 FILLCELL_X32 FILLER_351_1488 ();
 FILLCELL_X32 FILLER_351_1520 ();
 FILLCELL_X32 FILLER_351_1552 ();
 FILLCELL_X32 FILLER_351_1584 ();
 FILLCELL_X32 FILLER_351_1616 ();
 FILLCELL_X32 FILLER_351_1648 ();
 FILLCELL_X32 FILLER_351_1680 ();
 FILLCELL_X32 FILLER_351_1712 ();
 FILLCELL_X32 FILLER_351_1744 ();
 FILLCELL_X32 FILLER_351_1776 ();
 FILLCELL_X32 FILLER_351_1808 ();
 FILLCELL_X32 FILLER_351_1840 ();
 FILLCELL_X32 FILLER_351_1872 ();
 FILLCELL_X32 FILLER_351_1904 ();
 FILLCELL_X32 FILLER_351_1936 ();
 FILLCELL_X32 FILLER_351_1968 ();
 FILLCELL_X32 FILLER_351_2000 ();
 FILLCELL_X32 FILLER_351_2032 ();
 FILLCELL_X32 FILLER_351_2064 ();
 FILLCELL_X32 FILLER_351_2096 ();
 FILLCELL_X32 FILLER_351_2128 ();
 FILLCELL_X32 FILLER_351_2160 ();
 FILLCELL_X32 FILLER_351_2192 ();
 FILLCELL_X32 FILLER_351_2224 ();
 FILLCELL_X32 FILLER_351_2256 ();
 FILLCELL_X32 FILLER_351_2288 ();
 FILLCELL_X32 FILLER_351_2320 ();
 FILLCELL_X32 FILLER_351_2352 ();
 FILLCELL_X32 FILLER_351_2384 ();
 FILLCELL_X32 FILLER_351_2416 ();
 FILLCELL_X32 FILLER_351_2448 ();
 FILLCELL_X32 FILLER_351_2480 ();
 FILLCELL_X8 FILLER_351_2512 ();
 FILLCELL_X4 FILLER_351_2520 ();
 FILLCELL_X2 FILLER_351_2524 ();
 FILLCELL_X32 FILLER_351_2527 ();
 FILLCELL_X32 FILLER_351_2559 ();
 FILLCELL_X32 FILLER_351_2591 ();
 FILLCELL_X32 FILLER_351_2623 ();
 FILLCELL_X32 FILLER_351_2655 ();
 FILLCELL_X32 FILLER_351_2687 ();
 FILLCELL_X32 FILLER_351_2719 ();
 FILLCELL_X32 FILLER_351_2751 ();
 FILLCELL_X32 FILLER_351_2783 ();
 FILLCELL_X32 FILLER_351_2815 ();
 FILLCELL_X32 FILLER_351_2847 ();
 FILLCELL_X32 FILLER_351_2879 ();
 FILLCELL_X32 FILLER_351_2911 ();
 FILLCELL_X32 FILLER_351_2943 ();
 FILLCELL_X32 FILLER_351_2975 ();
 FILLCELL_X32 FILLER_351_3007 ();
 FILLCELL_X32 FILLER_351_3039 ();
 FILLCELL_X32 FILLER_351_3071 ();
 FILLCELL_X32 FILLER_351_3103 ();
 FILLCELL_X32 FILLER_351_3135 ();
 FILLCELL_X32 FILLER_351_3167 ();
 FILLCELL_X32 FILLER_351_3199 ();
 FILLCELL_X32 FILLER_351_3231 ();
 FILLCELL_X32 FILLER_351_3263 ();
 FILLCELL_X32 FILLER_351_3295 ();
 FILLCELL_X32 FILLER_351_3327 ();
 FILLCELL_X32 FILLER_351_3359 ();
 FILLCELL_X32 FILLER_351_3391 ();
 FILLCELL_X32 FILLER_351_3423 ();
 FILLCELL_X32 FILLER_351_3455 ();
 FILLCELL_X32 FILLER_351_3487 ();
 FILLCELL_X32 FILLER_351_3519 ();
 FILLCELL_X32 FILLER_351_3551 ();
 FILLCELL_X32 FILLER_351_3583 ();
 FILLCELL_X32 FILLER_351_3615 ();
 FILLCELL_X32 FILLER_351_3647 ();
 FILLCELL_X32 FILLER_351_3679 ();
 FILLCELL_X16 FILLER_351_3711 ();
 FILLCELL_X8 FILLER_351_3727 ();
 FILLCELL_X2 FILLER_351_3735 ();
 FILLCELL_X1 FILLER_351_3737 ();
 FILLCELL_X32 FILLER_352_1 ();
 FILLCELL_X32 FILLER_352_33 ();
 FILLCELL_X32 FILLER_352_65 ();
 FILLCELL_X32 FILLER_352_97 ();
 FILLCELL_X32 FILLER_352_129 ();
 FILLCELL_X32 FILLER_352_161 ();
 FILLCELL_X32 FILLER_352_193 ();
 FILLCELL_X32 FILLER_352_225 ();
 FILLCELL_X32 FILLER_352_257 ();
 FILLCELL_X32 FILLER_352_289 ();
 FILLCELL_X32 FILLER_352_321 ();
 FILLCELL_X32 FILLER_352_353 ();
 FILLCELL_X32 FILLER_352_385 ();
 FILLCELL_X32 FILLER_352_417 ();
 FILLCELL_X32 FILLER_352_449 ();
 FILLCELL_X32 FILLER_352_481 ();
 FILLCELL_X32 FILLER_352_513 ();
 FILLCELL_X32 FILLER_352_545 ();
 FILLCELL_X32 FILLER_352_577 ();
 FILLCELL_X16 FILLER_352_609 ();
 FILLCELL_X4 FILLER_352_625 ();
 FILLCELL_X2 FILLER_352_629 ();
 FILLCELL_X32 FILLER_352_632 ();
 FILLCELL_X32 FILLER_352_664 ();
 FILLCELL_X32 FILLER_352_696 ();
 FILLCELL_X32 FILLER_352_728 ();
 FILLCELL_X32 FILLER_352_760 ();
 FILLCELL_X32 FILLER_352_792 ();
 FILLCELL_X32 FILLER_352_824 ();
 FILLCELL_X32 FILLER_352_856 ();
 FILLCELL_X32 FILLER_352_888 ();
 FILLCELL_X32 FILLER_352_920 ();
 FILLCELL_X32 FILLER_352_952 ();
 FILLCELL_X32 FILLER_352_984 ();
 FILLCELL_X32 FILLER_352_1016 ();
 FILLCELL_X32 FILLER_352_1048 ();
 FILLCELL_X32 FILLER_352_1080 ();
 FILLCELL_X32 FILLER_352_1112 ();
 FILLCELL_X32 FILLER_352_1144 ();
 FILLCELL_X32 FILLER_352_1176 ();
 FILLCELL_X32 FILLER_352_1208 ();
 FILLCELL_X32 FILLER_352_1240 ();
 FILLCELL_X32 FILLER_352_1272 ();
 FILLCELL_X32 FILLER_352_1304 ();
 FILLCELL_X32 FILLER_352_1336 ();
 FILLCELL_X32 FILLER_352_1368 ();
 FILLCELL_X32 FILLER_352_1400 ();
 FILLCELL_X32 FILLER_352_1432 ();
 FILLCELL_X32 FILLER_352_1464 ();
 FILLCELL_X32 FILLER_352_1496 ();
 FILLCELL_X32 FILLER_352_1528 ();
 FILLCELL_X32 FILLER_352_1560 ();
 FILLCELL_X32 FILLER_352_1592 ();
 FILLCELL_X32 FILLER_352_1624 ();
 FILLCELL_X32 FILLER_352_1656 ();
 FILLCELL_X32 FILLER_352_1688 ();
 FILLCELL_X32 FILLER_352_1720 ();
 FILLCELL_X32 FILLER_352_1752 ();
 FILLCELL_X32 FILLER_352_1784 ();
 FILLCELL_X32 FILLER_352_1816 ();
 FILLCELL_X32 FILLER_352_1848 ();
 FILLCELL_X8 FILLER_352_1880 ();
 FILLCELL_X4 FILLER_352_1888 ();
 FILLCELL_X2 FILLER_352_1892 ();
 FILLCELL_X32 FILLER_352_1895 ();
 FILLCELL_X32 FILLER_352_1927 ();
 FILLCELL_X32 FILLER_352_1959 ();
 FILLCELL_X32 FILLER_352_1991 ();
 FILLCELL_X32 FILLER_352_2023 ();
 FILLCELL_X32 FILLER_352_2055 ();
 FILLCELL_X32 FILLER_352_2087 ();
 FILLCELL_X32 FILLER_352_2119 ();
 FILLCELL_X32 FILLER_352_2151 ();
 FILLCELL_X32 FILLER_352_2183 ();
 FILLCELL_X32 FILLER_352_2215 ();
 FILLCELL_X32 FILLER_352_2247 ();
 FILLCELL_X32 FILLER_352_2279 ();
 FILLCELL_X32 FILLER_352_2311 ();
 FILLCELL_X32 FILLER_352_2343 ();
 FILLCELL_X32 FILLER_352_2375 ();
 FILLCELL_X32 FILLER_352_2407 ();
 FILLCELL_X32 FILLER_352_2439 ();
 FILLCELL_X32 FILLER_352_2471 ();
 FILLCELL_X32 FILLER_352_2503 ();
 FILLCELL_X32 FILLER_352_2535 ();
 FILLCELL_X32 FILLER_352_2567 ();
 FILLCELL_X32 FILLER_352_2599 ();
 FILLCELL_X32 FILLER_352_2631 ();
 FILLCELL_X32 FILLER_352_2663 ();
 FILLCELL_X32 FILLER_352_2695 ();
 FILLCELL_X32 FILLER_352_2727 ();
 FILLCELL_X32 FILLER_352_2759 ();
 FILLCELL_X32 FILLER_352_2791 ();
 FILLCELL_X32 FILLER_352_2823 ();
 FILLCELL_X32 FILLER_352_2855 ();
 FILLCELL_X32 FILLER_352_2887 ();
 FILLCELL_X32 FILLER_352_2919 ();
 FILLCELL_X32 FILLER_352_2951 ();
 FILLCELL_X32 FILLER_352_2983 ();
 FILLCELL_X32 FILLER_352_3015 ();
 FILLCELL_X32 FILLER_352_3047 ();
 FILLCELL_X32 FILLER_352_3079 ();
 FILLCELL_X32 FILLER_352_3111 ();
 FILLCELL_X8 FILLER_352_3143 ();
 FILLCELL_X4 FILLER_352_3151 ();
 FILLCELL_X2 FILLER_352_3155 ();
 FILLCELL_X32 FILLER_352_3158 ();
 FILLCELL_X32 FILLER_352_3190 ();
 FILLCELL_X32 FILLER_352_3222 ();
 FILLCELL_X32 FILLER_352_3254 ();
 FILLCELL_X32 FILLER_352_3286 ();
 FILLCELL_X32 FILLER_352_3318 ();
 FILLCELL_X32 FILLER_352_3350 ();
 FILLCELL_X32 FILLER_352_3382 ();
 FILLCELL_X32 FILLER_352_3414 ();
 FILLCELL_X32 FILLER_352_3446 ();
 FILLCELL_X32 FILLER_352_3478 ();
 FILLCELL_X32 FILLER_352_3510 ();
 FILLCELL_X32 FILLER_352_3542 ();
 FILLCELL_X32 FILLER_352_3574 ();
 FILLCELL_X32 FILLER_352_3606 ();
 FILLCELL_X32 FILLER_352_3638 ();
 FILLCELL_X32 FILLER_352_3670 ();
 FILLCELL_X32 FILLER_352_3702 ();
 FILLCELL_X4 FILLER_352_3734 ();
 FILLCELL_X32 FILLER_353_1 ();
 FILLCELL_X32 FILLER_353_33 ();
 FILLCELL_X32 FILLER_353_65 ();
 FILLCELL_X32 FILLER_353_97 ();
 FILLCELL_X32 FILLER_353_129 ();
 FILLCELL_X32 FILLER_353_161 ();
 FILLCELL_X32 FILLER_353_193 ();
 FILLCELL_X32 FILLER_353_225 ();
 FILLCELL_X32 FILLER_353_257 ();
 FILLCELL_X32 FILLER_353_289 ();
 FILLCELL_X32 FILLER_353_321 ();
 FILLCELL_X32 FILLER_353_353 ();
 FILLCELL_X32 FILLER_353_385 ();
 FILLCELL_X32 FILLER_353_417 ();
 FILLCELL_X32 FILLER_353_449 ();
 FILLCELL_X32 FILLER_353_481 ();
 FILLCELL_X32 FILLER_353_513 ();
 FILLCELL_X32 FILLER_353_545 ();
 FILLCELL_X32 FILLER_353_577 ();
 FILLCELL_X32 FILLER_353_609 ();
 FILLCELL_X32 FILLER_353_641 ();
 FILLCELL_X32 FILLER_353_673 ();
 FILLCELL_X32 FILLER_353_705 ();
 FILLCELL_X32 FILLER_353_737 ();
 FILLCELL_X32 FILLER_353_769 ();
 FILLCELL_X32 FILLER_353_801 ();
 FILLCELL_X32 FILLER_353_833 ();
 FILLCELL_X32 FILLER_353_865 ();
 FILLCELL_X32 FILLER_353_897 ();
 FILLCELL_X32 FILLER_353_929 ();
 FILLCELL_X32 FILLER_353_961 ();
 FILLCELL_X32 FILLER_353_993 ();
 FILLCELL_X32 FILLER_353_1025 ();
 FILLCELL_X32 FILLER_353_1057 ();
 FILLCELL_X32 FILLER_353_1089 ();
 FILLCELL_X32 FILLER_353_1121 ();
 FILLCELL_X32 FILLER_353_1153 ();
 FILLCELL_X32 FILLER_353_1185 ();
 FILLCELL_X32 FILLER_353_1217 ();
 FILLCELL_X8 FILLER_353_1249 ();
 FILLCELL_X4 FILLER_353_1257 ();
 FILLCELL_X2 FILLER_353_1261 ();
 FILLCELL_X32 FILLER_353_1264 ();
 FILLCELL_X32 FILLER_353_1296 ();
 FILLCELL_X32 FILLER_353_1328 ();
 FILLCELL_X32 FILLER_353_1360 ();
 FILLCELL_X32 FILLER_353_1392 ();
 FILLCELL_X32 FILLER_353_1424 ();
 FILLCELL_X32 FILLER_353_1456 ();
 FILLCELL_X32 FILLER_353_1488 ();
 FILLCELL_X32 FILLER_353_1520 ();
 FILLCELL_X32 FILLER_353_1552 ();
 FILLCELL_X32 FILLER_353_1584 ();
 FILLCELL_X32 FILLER_353_1616 ();
 FILLCELL_X32 FILLER_353_1648 ();
 FILLCELL_X32 FILLER_353_1680 ();
 FILLCELL_X32 FILLER_353_1712 ();
 FILLCELL_X32 FILLER_353_1744 ();
 FILLCELL_X32 FILLER_353_1776 ();
 FILLCELL_X32 FILLER_353_1808 ();
 FILLCELL_X32 FILLER_353_1840 ();
 FILLCELL_X32 FILLER_353_1872 ();
 FILLCELL_X32 FILLER_353_1904 ();
 FILLCELL_X32 FILLER_353_1936 ();
 FILLCELL_X32 FILLER_353_1968 ();
 FILLCELL_X32 FILLER_353_2000 ();
 FILLCELL_X32 FILLER_353_2032 ();
 FILLCELL_X32 FILLER_353_2064 ();
 FILLCELL_X32 FILLER_353_2096 ();
 FILLCELL_X32 FILLER_353_2128 ();
 FILLCELL_X32 FILLER_353_2160 ();
 FILLCELL_X32 FILLER_353_2192 ();
 FILLCELL_X32 FILLER_353_2224 ();
 FILLCELL_X32 FILLER_353_2256 ();
 FILLCELL_X32 FILLER_353_2288 ();
 FILLCELL_X32 FILLER_353_2320 ();
 FILLCELL_X32 FILLER_353_2352 ();
 FILLCELL_X32 FILLER_353_2384 ();
 FILLCELL_X32 FILLER_353_2416 ();
 FILLCELL_X32 FILLER_353_2448 ();
 FILLCELL_X32 FILLER_353_2480 ();
 FILLCELL_X8 FILLER_353_2512 ();
 FILLCELL_X4 FILLER_353_2520 ();
 FILLCELL_X2 FILLER_353_2524 ();
 FILLCELL_X32 FILLER_353_2527 ();
 FILLCELL_X32 FILLER_353_2559 ();
 FILLCELL_X32 FILLER_353_2591 ();
 FILLCELL_X32 FILLER_353_2623 ();
 FILLCELL_X32 FILLER_353_2655 ();
 FILLCELL_X32 FILLER_353_2687 ();
 FILLCELL_X32 FILLER_353_2719 ();
 FILLCELL_X32 FILLER_353_2751 ();
 FILLCELL_X32 FILLER_353_2783 ();
 FILLCELL_X32 FILLER_353_2815 ();
 FILLCELL_X32 FILLER_353_2847 ();
 FILLCELL_X32 FILLER_353_2879 ();
 FILLCELL_X32 FILLER_353_2911 ();
 FILLCELL_X32 FILLER_353_2943 ();
 FILLCELL_X32 FILLER_353_2975 ();
 FILLCELL_X32 FILLER_353_3007 ();
 FILLCELL_X32 FILLER_353_3039 ();
 FILLCELL_X32 FILLER_353_3071 ();
 FILLCELL_X32 FILLER_353_3103 ();
 FILLCELL_X32 FILLER_353_3135 ();
 FILLCELL_X32 FILLER_353_3167 ();
 FILLCELL_X32 FILLER_353_3199 ();
 FILLCELL_X32 FILLER_353_3231 ();
 FILLCELL_X32 FILLER_353_3263 ();
 FILLCELL_X32 FILLER_353_3295 ();
 FILLCELL_X32 FILLER_353_3327 ();
 FILLCELL_X32 FILLER_353_3359 ();
 FILLCELL_X32 FILLER_353_3391 ();
 FILLCELL_X32 FILLER_353_3423 ();
 FILLCELL_X32 FILLER_353_3455 ();
 FILLCELL_X32 FILLER_353_3487 ();
 FILLCELL_X32 FILLER_353_3519 ();
 FILLCELL_X32 FILLER_353_3551 ();
 FILLCELL_X32 FILLER_353_3583 ();
 FILLCELL_X32 FILLER_353_3615 ();
 FILLCELL_X32 FILLER_353_3647 ();
 FILLCELL_X32 FILLER_353_3679 ();
 FILLCELL_X16 FILLER_353_3711 ();
 FILLCELL_X8 FILLER_353_3727 ();
 FILLCELL_X2 FILLER_353_3735 ();
 FILLCELL_X1 FILLER_353_3737 ();
 FILLCELL_X32 FILLER_354_1 ();
 FILLCELL_X32 FILLER_354_33 ();
 FILLCELL_X32 FILLER_354_65 ();
 FILLCELL_X32 FILLER_354_97 ();
 FILLCELL_X32 FILLER_354_129 ();
 FILLCELL_X32 FILLER_354_161 ();
 FILLCELL_X32 FILLER_354_193 ();
 FILLCELL_X32 FILLER_354_225 ();
 FILLCELL_X32 FILLER_354_257 ();
 FILLCELL_X32 FILLER_354_289 ();
 FILLCELL_X32 FILLER_354_321 ();
 FILLCELL_X32 FILLER_354_353 ();
 FILLCELL_X32 FILLER_354_385 ();
 FILLCELL_X32 FILLER_354_417 ();
 FILLCELL_X32 FILLER_354_449 ();
 FILLCELL_X32 FILLER_354_481 ();
 FILLCELL_X32 FILLER_354_513 ();
 FILLCELL_X32 FILLER_354_545 ();
 FILLCELL_X32 FILLER_354_577 ();
 FILLCELL_X16 FILLER_354_609 ();
 FILLCELL_X4 FILLER_354_625 ();
 FILLCELL_X2 FILLER_354_629 ();
 FILLCELL_X32 FILLER_354_632 ();
 FILLCELL_X32 FILLER_354_664 ();
 FILLCELL_X32 FILLER_354_696 ();
 FILLCELL_X32 FILLER_354_728 ();
 FILLCELL_X32 FILLER_354_760 ();
 FILLCELL_X32 FILLER_354_792 ();
 FILLCELL_X32 FILLER_354_824 ();
 FILLCELL_X32 FILLER_354_856 ();
 FILLCELL_X32 FILLER_354_888 ();
 FILLCELL_X32 FILLER_354_920 ();
 FILLCELL_X32 FILLER_354_952 ();
 FILLCELL_X32 FILLER_354_984 ();
 FILLCELL_X32 FILLER_354_1016 ();
 FILLCELL_X32 FILLER_354_1048 ();
 FILLCELL_X32 FILLER_354_1080 ();
 FILLCELL_X32 FILLER_354_1112 ();
 FILLCELL_X32 FILLER_354_1144 ();
 FILLCELL_X32 FILLER_354_1176 ();
 FILLCELL_X32 FILLER_354_1208 ();
 FILLCELL_X32 FILLER_354_1240 ();
 FILLCELL_X32 FILLER_354_1272 ();
 FILLCELL_X32 FILLER_354_1304 ();
 FILLCELL_X32 FILLER_354_1336 ();
 FILLCELL_X32 FILLER_354_1368 ();
 FILLCELL_X32 FILLER_354_1400 ();
 FILLCELL_X32 FILLER_354_1432 ();
 FILLCELL_X32 FILLER_354_1464 ();
 FILLCELL_X32 FILLER_354_1496 ();
 FILLCELL_X32 FILLER_354_1528 ();
 FILLCELL_X32 FILLER_354_1560 ();
 FILLCELL_X32 FILLER_354_1592 ();
 FILLCELL_X32 FILLER_354_1624 ();
 FILLCELL_X32 FILLER_354_1656 ();
 FILLCELL_X32 FILLER_354_1688 ();
 FILLCELL_X32 FILLER_354_1720 ();
 FILLCELL_X32 FILLER_354_1752 ();
 FILLCELL_X32 FILLER_354_1784 ();
 FILLCELL_X32 FILLER_354_1816 ();
 FILLCELL_X32 FILLER_354_1848 ();
 FILLCELL_X8 FILLER_354_1880 ();
 FILLCELL_X4 FILLER_354_1888 ();
 FILLCELL_X2 FILLER_354_1892 ();
 FILLCELL_X32 FILLER_354_1895 ();
 FILLCELL_X32 FILLER_354_1927 ();
 FILLCELL_X32 FILLER_354_1959 ();
 FILLCELL_X32 FILLER_354_1991 ();
 FILLCELL_X32 FILLER_354_2023 ();
 FILLCELL_X32 FILLER_354_2055 ();
 FILLCELL_X32 FILLER_354_2087 ();
 FILLCELL_X32 FILLER_354_2119 ();
 FILLCELL_X32 FILLER_354_2151 ();
 FILLCELL_X32 FILLER_354_2183 ();
 FILLCELL_X32 FILLER_354_2215 ();
 FILLCELL_X32 FILLER_354_2247 ();
 FILLCELL_X32 FILLER_354_2279 ();
 FILLCELL_X32 FILLER_354_2311 ();
 FILLCELL_X32 FILLER_354_2343 ();
 FILLCELL_X32 FILLER_354_2375 ();
 FILLCELL_X32 FILLER_354_2407 ();
 FILLCELL_X32 FILLER_354_2439 ();
 FILLCELL_X32 FILLER_354_2471 ();
 FILLCELL_X32 FILLER_354_2503 ();
 FILLCELL_X32 FILLER_354_2535 ();
 FILLCELL_X32 FILLER_354_2567 ();
 FILLCELL_X32 FILLER_354_2599 ();
 FILLCELL_X32 FILLER_354_2631 ();
 FILLCELL_X32 FILLER_354_2663 ();
 FILLCELL_X32 FILLER_354_2695 ();
 FILLCELL_X32 FILLER_354_2727 ();
 FILLCELL_X32 FILLER_354_2759 ();
 FILLCELL_X32 FILLER_354_2791 ();
 FILLCELL_X32 FILLER_354_2823 ();
 FILLCELL_X32 FILLER_354_2855 ();
 FILLCELL_X32 FILLER_354_2887 ();
 FILLCELL_X32 FILLER_354_2919 ();
 FILLCELL_X32 FILLER_354_2951 ();
 FILLCELL_X32 FILLER_354_2983 ();
 FILLCELL_X32 FILLER_354_3015 ();
 FILLCELL_X32 FILLER_354_3047 ();
 FILLCELL_X32 FILLER_354_3079 ();
 FILLCELL_X32 FILLER_354_3111 ();
 FILLCELL_X8 FILLER_354_3143 ();
 FILLCELL_X4 FILLER_354_3151 ();
 FILLCELL_X2 FILLER_354_3155 ();
 FILLCELL_X32 FILLER_354_3158 ();
 FILLCELL_X32 FILLER_354_3190 ();
 FILLCELL_X32 FILLER_354_3222 ();
 FILLCELL_X32 FILLER_354_3254 ();
 FILLCELL_X32 FILLER_354_3286 ();
 FILLCELL_X32 FILLER_354_3318 ();
 FILLCELL_X32 FILLER_354_3350 ();
 FILLCELL_X32 FILLER_354_3382 ();
 FILLCELL_X32 FILLER_354_3414 ();
 FILLCELL_X32 FILLER_354_3446 ();
 FILLCELL_X32 FILLER_354_3478 ();
 FILLCELL_X32 FILLER_354_3510 ();
 FILLCELL_X32 FILLER_354_3542 ();
 FILLCELL_X32 FILLER_354_3574 ();
 FILLCELL_X32 FILLER_354_3606 ();
 FILLCELL_X32 FILLER_354_3638 ();
 FILLCELL_X32 FILLER_354_3670 ();
 FILLCELL_X32 FILLER_354_3702 ();
 FILLCELL_X4 FILLER_354_3734 ();
 FILLCELL_X32 FILLER_355_1 ();
 FILLCELL_X32 FILLER_355_33 ();
 FILLCELL_X32 FILLER_355_65 ();
 FILLCELL_X32 FILLER_355_97 ();
 FILLCELL_X32 FILLER_355_129 ();
 FILLCELL_X32 FILLER_355_161 ();
 FILLCELL_X32 FILLER_355_193 ();
 FILLCELL_X32 FILLER_355_225 ();
 FILLCELL_X32 FILLER_355_257 ();
 FILLCELL_X32 FILLER_355_289 ();
 FILLCELL_X32 FILLER_355_321 ();
 FILLCELL_X32 FILLER_355_353 ();
 FILLCELL_X32 FILLER_355_385 ();
 FILLCELL_X32 FILLER_355_417 ();
 FILLCELL_X32 FILLER_355_449 ();
 FILLCELL_X32 FILLER_355_481 ();
 FILLCELL_X32 FILLER_355_513 ();
 FILLCELL_X32 FILLER_355_545 ();
 FILLCELL_X32 FILLER_355_577 ();
 FILLCELL_X32 FILLER_355_609 ();
 FILLCELL_X32 FILLER_355_641 ();
 FILLCELL_X32 FILLER_355_673 ();
 FILLCELL_X32 FILLER_355_705 ();
 FILLCELL_X32 FILLER_355_737 ();
 FILLCELL_X32 FILLER_355_769 ();
 FILLCELL_X32 FILLER_355_801 ();
 FILLCELL_X32 FILLER_355_833 ();
 FILLCELL_X32 FILLER_355_865 ();
 FILLCELL_X32 FILLER_355_897 ();
 FILLCELL_X32 FILLER_355_929 ();
 FILLCELL_X32 FILLER_355_961 ();
 FILLCELL_X32 FILLER_355_993 ();
 FILLCELL_X32 FILLER_355_1025 ();
 FILLCELL_X32 FILLER_355_1057 ();
 FILLCELL_X32 FILLER_355_1089 ();
 FILLCELL_X32 FILLER_355_1121 ();
 FILLCELL_X32 FILLER_355_1153 ();
 FILLCELL_X32 FILLER_355_1185 ();
 FILLCELL_X32 FILLER_355_1217 ();
 FILLCELL_X8 FILLER_355_1249 ();
 FILLCELL_X4 FILLER_355_1257 ();
 FILLCELL_X2 FILLER_355_1261 ();
 FILLCELL_X32 FILLER_355_1264 ();
 FILLCELL_X32 FILLER_355_1296 ();
 FILLCELL_X32 FILLER_355_1328 ();
 FILLCELL_X32 FILLER_355_1360 ();
 FILLCELL_X32 FILLER_355_1392 ();
 FILLCELL_X32 FILLER_355_1424 ();
 FILLCELL_X32 FILLER_355_1456 ();
 FILLCELL_X32 FILLER_355_1488 ();
 FILLCELL_X32 FILLER_355_1520 ();
 FILLCELL_X32 FILLER_355_1552 ();
 FILLCELL_X32 FILLER_355_1584 ();
 FILLCELL_X32 FILLER_355_1616 ();
 FILLCELL_X32 FILLER_355_1648 ();
 FILLCELL_X32 FILLER_355_1680 ();
 FILLCELL_X32 FILLER_355_1712 ();
 FILLCELL_X32 FILLER_355_1744 ();
 FILLCELL_X32 FILLER_355_1776 ();
 FILLCELL_X32 FILLER_355_1808 ();
 FILLCELL_X32 FILLER_355_1840 ();
 FILLCELL_X32 FILLER_355_1872 ();
 FILLCELL_X32 FILLER_355_1904 ();
 FILLCELL_X32 FILLER_355_1936 ();
 FILLCELL_X32 FILLER_355_1968 ();
 FILLCELL_X32 FILLER_355_2000 ();
 FILLCELL_X32 FILLER_355_2032 ();
 FILLCELL_X32 FILLER_355_2064 ();
 FILLCELL_X32 FILLER_355_2096 ();
 FILLCELL_X32 FILLER_355_2128 ();
 FILLCELL_X32 FILLER_355_2160 ();
 FILLCELL_X32 FILLER_355_2192 ();
 FILLCELL_X32 FILLER_355_2224 ();
 FILLCELL_X32 FILLER_355_2256 ();
 FILLCELL_X32 FILLER_355_2288 ();
 FILLCELL_X32 FILLER_355_2320 ();
 FILLCELL_X32 FILLER_355_2352 ();
 FILLCELL_X32 FILLER_355_2384 ();
 FILLCELL_X32 FILLER_355_2416 ();
 FILLCELL_X32 FILLER_355_2448 ();
 FILLCELL_X32 FILLER_355_2480 ();
 FILLCELL_X8 FILLER_355_2512 ();
 FILLCELL_X4 FILLER_355_2520 ();
 FILLCELL_X2 FILLER_355_2524 ();
 FILLCELL_X32 FILLER_355_2527 ();
 FILLCELL_X32 FILLER_355_2559 ();
 FILLCELL_X32 FILLER_355_2591 ();
 FILLCELL_X32 FILLER_355_2623 ();
 FILLCELL_X32 FILLER_355_2655 ();
 FILLCELL_X32 FILLER_355_2687 ();
 FILLCELL_X32 FILLER_355_2719 ();
 FILLCELL_X32 FILLER_355_2751 ();
 FILLCELL_X32 FILLER_355_2783 ();
 FILLCELL_X32 FILLER_355_2815 ();
 FILLCELL_X32 FILLER_355_2847 ();
 FILLCELL_X32 FILLER_355_2879 ();
 FILLCELL_X32 FILLER_355_2911 ();
 FILLCELL_X32 FILLER_355_2943 ();
 FILLCELL_X32 FILLER_355_2975 ();
 FILLCELL_X32 FILLER_355_3007 ();
 FILLCELL_X32 FILLER_355_3039 ();
 FILLCELL_X32 FILLER_355_3071 ();
 FILLCELL_X32 FILLER_355_3103 ();
 FILLCELL_X32 FILLER_355_3135 ();
 FILLCELL_X32 FILLER_355_3167 ();
 FILLCELL_X32 FILLER_355_3199 ();
 FILLCELL_X32 FILLER_355_3231 ();
 FILLCELL_X32 FILLER_355_3263 ();
 FILLCELL_X32 FILLER_355_3295 ();
 FILLCELL_X32 FILLER_355_3327 ();
 FILLCELL_X32 FILLER_355_3359 ();
 FILLCELL_X32 FILLER_355_3391 ();
 FILLCELL_X32 FILLER_355_3423 ();
 FILLCELL_X32 FILLER_355_3455 ();
 FILLCELL_X32 FILLER_355_3487 ();
 FILLCELL_X32 FILLER_355_3519 ();
 FILLCELL_X32 FILLER_355_3551 ();
 FILLCELL_X32 FILLER_355_3583 ();
 FILLCELL_X32 FILLER_355_3615 ();
 FILLCELL_X32 FILLER_355_3647 ();
 FILLCELL_X32 FILLER_355_3679 ();
 FILLCELL_X16 FILLER_355_3711 ();
 FILLCELL_X8 FILLER_355_3727 ();
 FILLCELL_X2 FILLER_355_3735 ();
 FILLCELL_X1 FILLER_355_3737 ();
 FILLCELL_X32 FILLER_356_1 ();
 FILLCELL_X32 FILLER_356_33 ();
 FILLCELL_X32 FILLER_356_65 ();
 FILLCELL_X32 FILLER_356_97 ();
 FILLCELL_X32 FILLER_356_129 ();
 FILLCELL_X32 FILLER_356_161 ();
 FILLCELL_X32 FILLER_356_193 ();
 FILLCELL_X32 FILLER_356_225 ();
 FILLCELL_X32 FILLER_356_257 ();
 FILLCELL_X32 FILLER_356_289 ();
 FILLCELL_X32 FILLER_356_321 ();
 FILLCELL_X32 FILLER_356_353 ();
 FILLCELL_X32 FILLER_356_385 ();
 FILLCELL_X32 FILLER_356_417 ();
 FILLCELL_X32 FILLER_356_449 ();
 FILLCELL_X32 FILLER_356_481 ();
 FILLCELL_X32 FILLER_356_513 ();
 FILLCELL_X32 FILLER_356_545 ();
 FILLCELL_X32 FILLER_356_577 ();
 FILLCELL_X16 FILLER_356_609 ();
 FILLCELL_X4 FILLER_356_625 ();
 FILLCELL_X2 FILLER_356_629 ();
 FILLCELL_X32 FILLER_356_632 ();
 FILLCELL_X32 FILLER_356_664 ();
 FILLCELL_X32 FILLER_356_696 ();
 FILLCELL_X32 FILLER_356_728 ();
 FILLCELL_X32 FILLER_356_760 ();
 FILLCELL_X32 FILLER_356_792 ();
 FILLCELL_X32 FILLER_356_824 ();
 FILLCELL_X32 FILLER_356_856 ();
 FILLCELL_X32 FILLER_356_888 ();
 FILLCELL_X32 FILLER_356_920 ();
 FILLCELL_X32 FILLER_356_952 ();
 FILLCELL_X32 FILLER_356_984 ();
 FILLCELL_X32 FILLER_356_1016 ();
 FILLCELL_X32 FILLER_356_1048 ();
 FILLCELL_X32 FILLER_356_1080 ();
 FILLCELL_X32 FILLER_356_1112 ();
 FILLCELL_X32 FILLER_356_1144 ();
 FILLCELL_X32 FILLER_356_1176 ();
 FILLCELL_X32 FILLER_356_1208 ();
 FILLCELL_X32 FILLER_356_1240 ();
 FILLCELL_X32 FILLER_356_1272 ();
 FILLCELL_X32 FILLER_356_1304 ();
 FILLCELL_X32 FILLER_356_1336 ();
 FILLCELL_X32 FILLER_356_1368 ();
 FILLCELL_X32 FILLER_356_1400 ();
 FILLCELL_X32 FILLER_356_1432 ();
 FILLCELL_X32 FILLER_356_1464 ();
 FILLCELL_X32 FILLER_356_1496 ();
 FILLCELL_X32 FILLER_356_1528 ();
 FILLCELL_X32 FILLER_356_1560 ();
 FILLCELL_X32 FILLER_356_1592 ();
 FILLCELL_X32 FILLER_356_1624 ();
 FILLCELL_X32 FILLER_356_1656 ();
 FILLCELL_X32 FILLER_356_1688 ();
 FILLCELL_X32 FILLER_356_1720 ();
 FILLCELL_X32 FILLER_356_1752 ();
 FILLCELL_X32 FILLER_356_1784 ();
 FILLCELL_X32 FILLER_356_1816 ();
 FILLCELL_X32 FILLER_356_1848 ();
 FILLCELL_X8 FILLER_356_1880 ();
 FILLCELL_X4 FILLER_356_1888 ();
 FILLCELL_X2 FILLER_356_1892 ();
 FILLCELL_X32 FILLER_356_1895 ();
 FILLCELL_X32 FILLER_356_1927 ();
 FILLCELL_X32 FILLER_356_1959 ();
 FILLCELL_X32 FILLER_356_1991 ();
 FILLCELL_X32 FILLER_356_2023 ();
 FILLCELL_X32 FILLER_356_2055 ();
 FILLCELL_X32 FILLER_356_2087 ();
 FILLCELL_X32 FILLER_356_2119 ();
 FILLCELL_X32 FILLER_356_2151 ();
 FILLCELL_X32 FILLER_356_2183 ();
 FILLCELL_X32 FILLER_356_2215 ();
 FILLCELL_X32 FILLER_356_2247 ();
 FILLCELL_X32 FILLER_356_2279 ();
 FILLCELL_X32 FILLER_356_2311 ();
 FILLCELL_X32 FILLER_356_2343 ();
 FILLCELL_X32 FILLER_356_2375 ();
 FILLCELL_X32 FILLER_356_2407 ();
 FILLCELL_X32 FILLER_356_2439 ();
 FILLCELL_X32 FILLER_356_2471 ();
 FILLCELL_X32 FILLER_356_2503 ();
 FILLCELL_X32 FILLER_356_2535 ();
 FILLCELL_X32 FILLER_356_2567 ();
 FILLCELL_X32 FILLER_356_2599 ();
 FILLCELL_X32 FILLER_356_2631 ();
 FILLCELL_X32 FILLER_356_2663 ();
 FILLCELL_X32 FILLER_356_2695 ();
 FILLCELL_X32 FILLER_356_2727 ();
 FILLCELL_X32 FILLER_356_2759 ();
 FILLCELL_X32 FILLER_356_2791 ();
 FILLCELL_X32 FILLER_356_2823 ();
 FILLCELL_X32 FILLER_356_2855 ();
 FILLCELL_X32 FILLER_356_2887 ();
 FILLCELL_X32 FILLER_356_2919 ();
 FILLCELL_X32 FILLER_356_2951 ();
 FILLCELL_X32 FILLER_356_2983 ();
 FILLCELL_X32 FILLER_356_3015 ();
 FILLCELL_X32 FILLER_356_3047 ();
 FILLCELL_X32 FILLER_356_3079 ();
 FILLCELL_X32 FILLER_356_3111 ();
 FILLCELL_X8 FILLER_356_3143 ();
 FILLCELL_X4 FILLER_356_3151 ();
 FILLCELL_X2 FILLER_356_3155 ();
 FILLCELL_X32 FILLER_356_3158 ();
 FILLCELL_X32 FILLER_356_3190 ();
 FILLCELL_X32 FILLER_356_3222 ();
 FILLCELL_X32 FILLER_356_3254 ();
 FILLCELL_X32 FILLER_356_3286 ();
 FILLCELL_X32 FILLER_356_3318 ();
 FILLCELL_X32 FILLER_356_3350 ();
 FILLCELL_X32 FILLER_356_3382 ();
 FILLCELL_X32 FILLER_356_3414 ();
 FILLCELL_X32 FILLER_356_3446 ();
 FILLCELL_X32 FILLER_356_3478 ();
 FILLCELL_X32 FILLER_356_3510 ();
 FILLCELL_X32 FILLER_356_3542 ();
 FILLCELL_X32 FILLER_356_3574 ();
 FILLCELL_X32 FILLER_356_3606 ();
 FILLCELL_X32 FILLER_356_3638 ();
 FILLCELL_X32 FILLER_356_3670 ();
 FILLCELL_X32 FILLER_356_3702 ();
 FILLCELL_X4 FILLER_356_3734 ();
 FILLCELL_X32 FILLER_357_1 ();
 FILLCELL_X32 FILLER_357_33 ();
 FILLCELL_X32 FILLER_357_65 ();
 FILLCELL_X32 FILLER_357_97 ();
 FILLCELL_X32 FILLER_357_129 ();
 FILLCELL_X32 FILLER_357_161 ();
 FILLCELL_X32 FILLER_357_193 ();
 FILLCELL_X32 FILLER_357_225 ();
 FILLCELL_X32 FILLER_357_257 ();
 FILLCELL_X32 FILLER_357_289 ();
 FILLCELL_X32 FILLER_357_321 ();
 FILLCELL_X32 FILLER_357_353 ();
 FILLCELL_X32 FILLER_357_385 ();
 FILLCELL_X32 FILLER_357_417 ();
 FILLCELL_X32 FILLER_357_449 ();
 FILLCELL_X32 FILLER_357_481 ();
 FILLCELL_X32 FILLER_357_513 ();
 FILLCELL_X32 FILLER_357_545 ();
 FILLCELL_X32 FILLER_357_577 ();
 FILLCELL_X32 FILLER_357_609 ();
 FILLCELL_X32 FILLER_357_641 ();
 FILLCELL_X32 FILLER_357_673 ();
 FILLCELL_X32 FILLER_357_705 ();
 FILLCELL_X32 FILLER_357_737 ();
 FILLCELL_X32 FILLER_357_769 ();
 FILLCELL_X32 FILLER_357_801 ();
 FILLCELL_X32 FILLER_357_833 ();
 FILLCELL_X32 FILLER_357_865 ();
 FILLCELL_X32 FILLER_357_897 ();
 FILLCELL_X32 FILLER_357_929 ();
 FILLCELL_X32 FILLER_357_961 ();
 FILLCELL_X32 FILLER_357_993 ();
 FILLCELL_X32 FILLER_357_1025 ();
 FILLCELL_X32 FILLER_357_1057 ();
 FILLCELL_X32 FILLER_357_1089 ();
 FILLCELL_X32 FILLER_357_1121 ();
 FILLCELL_X32 FILLER_357_1153 ();
 FILLCELL_X32 FILLER_357_1185 ();
 FILLCELL_X32 FILLER_357_1217 ();
 FILLCELL_X8 FILLER_357_1249 ();
 FILLCELL_X4 FILLER_357_1257 ();
 FILLCELL_X2 FILLER_357_1261 ();
 FILLCELL_X32 FILLER_357_1264 ();
 FILLCELL_X32 FILLER_357_1296 ();
 FILLCELL_X32 FILLER_357_1328 ();
 FILLCELL_X32 FILLER_357_1360 ();
 FILLCELL_X32 FILLER_357_1392 ();
 FILLCELL_X32 FILLER_357_1424 ();
 FILLCELL_X32 FILLER_357_1456 ();
 FILLCELL_X32 FILLER_357_1488 ();
 FILLCELL_X32 FILLER_357_1520 ();
 FILLCELL_X32 FILLER_357_1552 ();
 FILLCELL_X32 FILLER_357_1584 ();
 FILLCELL_X32 FILLER_357_1616 ();
 FILLCELL_X32 FILLER_357_1648 ();
 FILLCELL_X32 FILLER_357_1680 ();
 FILLCELL_X32 FILLER_357_1712 ();
 FILLCELL_X32 FILLER_357_1744 ();
 FILLCELL_X32 FILLER_357_1776 ();
 FILLCELL_X32 FILLER_357_1808 ();
 FILLCELL_X32 FILLER_357_1840 ();
 FILLCELL_X32 FILLER_357_1872 ();
 FILLCELL_X32 FILLER_357_1904 ();
 FILLCELL_X32 FILLER_357_1936 ();
 FILLCELL_X32 FILLER_357_1968 ();
 FILLCELL_X32 FILLER_357_2000 ();
 FILLCELL_X32 FILLER_357_2032 ();
 FILLCELL_X32 FILLER_357_2064 ();
 FILLCELL_X32 FILLER_357_2096 ();
 FILLCELL_X32 FILLER_357_2128 ();
 FILLCELL_X32 FILLER_357_2160 ();
 FILLCELL_X32 FILLER_357_2192 ();
 FILLCELL_X32 FILLER_357_2224 ();
 FILLCELL_X32 FILLER_357_2256 ();
 FILLCELL_X32 FILLER_357_2288 ();
 FILLCELL_X32 FILLER_357_2320 ();
 FILLCELL_X32 FILLER_357_2352 ();
 FILLCELL_X32 FILLER_357_2384 ();
 FILLCELL_X32 FILLER_357_2416 ();
 FILLCELL_X32 FILLER_357_2448 ();
 FILLCELL_X32 FILLER_357_2480 ();
 FILLCELL_X8 FILLER_357_2512 ();
 FILLCELL_X4 FILLER_357_2520 ();
 FILLCELL_X2 FILLER_357_2524 ();
 FILLCELL_X32 FILLER_357_2527 ();
 FILLCELL_X32 FILLER_357_2559 ();
 FILLCELL_X32 FILLER_357_2591 ();
 FILLCELL_X32 FILLER_357_2623 ();
 FILLCELL_X32 FILLER_357_2655 ();
 FILLCELL_X32 FILLER_357_2687 ();
 FILLCELL_X32 FILLER_357_2719 ();
 FILLCELL_X32 FILLER_357_2751 ();
 FILLCELL_X32 FILLER_357_2783 ();
 FILLCELL_X32 FILLER_357_2815 ();
 FILLCELL_X32 FILLER_357_2847 ();
 FILLCELL_X32 FILLER_357_2879 ();
 FILLCELL_X32 FILLER_357_2911 ();
 FILLCELL_X32 FILLER_357_2943 ();
 FILLCELL_X32 FILLER_357_2975 ();
 FILLCELL_X32 FILLER_357_3007 ();
 FILLCELL_X32 FILLER_357_3039 ();
 FILLCELL_X32 FILLER_357_3071 ();
 FILLCELL_X32 FILLER_357_3103 ();
 FILLCELL_X32 FILLER_357_3135 ();
 FILLCELL_X32 FILLER_357_3167 ();
 FILLCELL_X32 FILLER_357_3199 ();
 FILLCELL_X32 FILLER_357_3231 ();
 FILLCELL_X32 FILLER_357_3263 ();
 FILLCELL_X32 FILLER_357_3295 ();
 FILLCELL_X32 FILLER_357_3327 ();
 FILLCELL_X32 FILLER_357_3359 ();
 FILLCELL_X32 FILLER_357_3391 ();
 FILLCELL_X32 FILLER_357_3423 ();
 FILLCELL_X32 FILLER_357_3455 ();
 FILLCELL_X32 FILLER_357_3487 ();
 FILLCELL_X32 FILLER_357_3519 ();
 FILLCELL_X32 FILLER_357_3551 ();
 FILLCELL_X32 FILLER_357_3583 ();
 FILLCELL_X32 FILLER_357_3615 ();
 FILLCELL_X32 FILLER_357_3647 ();
 FILLCELL_X32 FILLER_357_3679 ();
 FILLCELL_X16 FILLER_357_3711 ();
 FILLCELL_X8 FILLER_357_3727 ();
 FILLCELL_X2 FILLER_357_3735 ();
 FILLCELL_X1 FILLER_357_3737 ();
 FILLCELL_X32 FILLER_358_1 ();
 FILLCELL_X32 FILLER_358_33 ();
 FILLCELL_X32 FILLER_358_65 ();
 FILLCELL_X32 FILLER_358_97 ();
 FILLCELL_X32 FILLER_358_129 ();
 FILLCELL_X32 FILLER_358_161 ();
 FILLCELL_X32 FILLER_358_193 ();
 FILLCELL_X32 FILLER_358_225 ();
 FILLCELL_X32 FILLER_358_257 ();
 FILLCELL_X32 FILLER_358_289 ();
 FILLCELL_X32 FILLER_358_321 ();
 FILLCELL_X32 FILLER_358_353 ();
 FILLCELL_X32 FILLER_358_385 ();
 FILLCELL_X32 FILLER_358_417 ();
 FILLCELL_X32 FILLER_358_449 ();
 FILLCELL_X32 FILLER_358_481 ();
 FILLCELL_X32 FILLER_358_513 ();
 FILLCELL_X32 FILLER_358_545 ();
 FILLCELL_X32 FILLER_358_577 ();
 FILLCELL_X16 FILLER_358_609 ();
 FILLCELL_X4 FILLER_358_625 ();
 FILLCELL_X2 FILLER_358_629 ();
 FILLCELL_X32 FILLER_358_632 ();
 FILLCELL_X32 FILLER_358_664 ();
 FILLCELL_X32 FILLER_358_696 ();
 FILLCELL_X32 FILLER_358_728 ();
 FILLCELL_X32 FILLER_358_760 ();
 FILLCELL_X32 FILLER_358_792 ();
 FILLCELL_X32 FILLER_358_824 ();
 FILLCELL_X32 FILLER_358_856 ();
 FILLCELL_X32 FILLER_358_888 ();
 FILLCELL_X32 FILLER_358_920 ();
 FILLCELL_X32 FILLER_358_952 ();
 FILLCELL_X32 FILLER_358_984 ();
 FILLCELL_X32 FILLER_358_1016 ();
 FILLCELL_X32 FILLER_358_1048 ();
 FILLCELL_X32 FILLER_358_1080 ();
 FILLCELL_X32 FILLER_358_1112 ();
 FILLCELL_X32 FILLER_358_1144 ();
 FILLCELL_X32 FILLER_358_1176 ();
 FILLCELL_X32 FILLER_358_1208 ();
 FILLCELL_X32 FILLER_358_1240 ();
 FILLCELL_X32 FILLER_358_1272 ();
 FILLCELL_X32 FILLER_358_1304 ();
 FILLCELL_X32 FILLER_358_1336 ();
 FILLCELL_X32 FILLER_358_1368 ();
 FILLCELL_X32 FILLER_358_1400 ();
 FILLCELL_X32 FILLER_358_1432 ();
 FILLCELL_X32 FILLER_358_1464 ();
 FILLCELL_X32 FILLER_358_1496 ();
 FILLCELL_X32 FILLER_358_1528 ();
 FILLCELL_X32 FILLER_358_1560 ();
 FILLCELL_X32 FILLER_358_1592 ();
 FILLCELL_X32 FILLER_358_1624 ();
 FILLCELL_X32 FILLER_358_1656 ();
 FILLCELL_X32 FILLER_358_1688 ();
 FILLCELL_X32 FILLER_358_1720 ();
 FILLCELL_X32 FILLER_358_1752 ();
 FILLCELL_X32 FILLER_358_1784 ();
 FILLCELL_X32 FILLER_358_1816 ();
 FILLCELL_X32 FILLER_358_1848 ();
 FILLCELL_X8 FILLER_358_1880 ();
 FILLCELL_X4 FILLER_358_1888 ();
 FILLCELL_X2 FILLER_358_1892 ();
 FILLCELL_X32 FILLER_358_1895 ();
 FILLCELL_X32 FILLER_358_1927 ();
 FILLCELL_X32 FILLER_358_1959 ();
 FILLCELL_X32 FILLER_358_1991 ();
 FILLCELL_X32 FILLER_358_2023 ();
 FILLCELL_X32 FILLER_358_2055 ();
 FILLCELL_X32 FILLER_358_2087 ();
 FILLCELL_X32 FILLER_358_2119 ();
 FILLCELL_X32 FILLER_358_2151 ();
 FILLCELL_X32 FILLER_358_2183 ();
 FILLCELL_X32 FILLER_358_2215 ();
 FILLCELL_X32 FILLER_358_2247 ();
 FILLCELL_X32 FILLER_358_2279 ();
 FILLCELL_X32 FILLER_358_2311 ();
 FILLCELL_X32 FILLER_358_2343 ();
 FILLCELL_X32 FILLER_358_2375 ();
 FILLCELL_X32 FILLER_358_2407 ();
 FILLCELL_X32 FILLER_358_2439 ();
 FILLCELL_X32 FILLER_358_2471 ();
 FILLCELL_X32 FILLER_358_2503 ();
 FILLCELL_X32 FILLER_358_2535 ();
 FILLCELL_X32 FILLER_358_2567 ();
 FILLCELL_X32 FILLER_358_2599 ();
 FILLCELL_X32 FILLER_358_2631 ();
 FILLCELL_X32 FILLER_358_2663 ();
 FILLCELL_X32 FILLER_358_2695 ();
 FILLCELL_X32 FILLER_358_2727 ();
 FILLCELL_X32 FILLER_358_2759 ();
 FILLCELL_X32 FILLER_358_2791 ();
 FILLCELL_X32 FILLER_358_2823 ();
 FILLCELL_X32 FILLER_358_2855 ();
 FILLCELL_X32 FILLER_358_2887 ();
 FILLCELL_X32 FILLER_358_2919 ();
 FILLCELL_X32 FILLER_358_2951 ();
 FILLCELL_X32 FILLER_358_2983 ();
 FILLCELL_X32 FILLER_358_3015 ();
 FILLCELL_X32 FILLER_358_3047 ();
 FILLCELL_X32 FILLER_358_3079 ();
 FILLCELL_X32 FILLER_358_3111 ();
 FILLCELL_X8 FILLER_358_3143 ();
 FILLCELL_X4 FILLER_358_3151 ();
 FILLCELL_X2 FILLER_358_3155 ();
 FILLCELL_X32 FILLER_358_3158 ();
 FILLCELL_X32 FILLER_358_3190 ();
 FILLCELL_X32 FILLER_358_3222 ();
 FILLCELL_X32 FILLER_358_3254 ();
 FILLCELL_X32 FILLER_358_3286 ();
 FILLCELL_X32 FILLER_358_3318 ();
 FILLCELL_X32 FILLER_358_3350 ();
 FILLCELL_X32 FILLER_358_3382 ();
 FILLCELL_X32 FILLER_358_3414 ();
 FILLCELL_X32 FILLER_358_3446 ();
 FILLCELL_X32 FILLER_358_3478 ();
 FILLCELL_X32 FILLER_358_3510 ();
 FILLCELL_X32 FILLER_358_3542 ();
 FILLCELL_X32 FILLER_358_3574 ();
 FILLCELL_X32 FILLER_358_3606 ();
 FILLCELL_X32 FILLER_358_3638 ();
 FILLCELL_X32 FILLER_358_3670 ();
 FILLCELL_X32 FILLER_358_3702 ();
 FILLCELL_X4 FILLER_358_3734 ();
 FILLCELL_X32 FILLER_359_1 ();
 FILLCELL_X32 FILLER_359_33 ();
 FILLCELL_X32 FILLER_359_65 ();
 FILLCELL_X32 FILLER_359_97 ();
 FILLCELL_X32 FILLER_359_129 ();
 FILLCELL_X32 FILLER_359_161 ();
 FILLCELL_X32 FILLER_359_193 ();
 FILLCELL_X32 FILLER_359_225 ();
 FILLCELL_X32 FILLER_359_257 ();
 FILLCELL_X32 FILLER_359_289 ();
 FILLCELL_X32 FILLER_359_321 ();
 FILLCELL_X32 FILLER_359_353 ();
 FILLCELL_X32 FILLER_359_385 ();
 FILLCELL_X32 FILLER_359_417 ();
 FILLCELL_X32 FILLER_359_449 ();
 FILLCELL_X32 FILLER_359_481 ();
 FILLCELL_X32 FILLER_359_513 ();
 FILLCELL_X32 FILLER_359_545 ();
 FILLCELL_X32 FILLER_359_577 ();
 FILLCELL_X32 FILLER_359_609 ();
 FILLCELL_X32 FILLER_359_641 ();
 FILLCELL_X32 FILLER_359_673 ();
 FILLCELL_X32 FILLER_359_705 ();
 FILLCELL_X32 FILLER_359_737 ();
 FILLCELL_X32 FILLER_359_769 ();
 FILLCELL_X32 FILLER_359_801 ();
 FILLCELL_X32 FILLER_359_833 ();
 FILLCELL_X32 FILLER_359_865 ();
 FILLCELL_X32 FILLER_359_897 ();
 FILLCELL_X32 FILLER_359_929 ();
 FILLCELL_X32 FILLER_359_961 ();
 FILLCELL_X32 FILLER_359_993 ();
 FILLCELL_X32 FILLER_359_1025 ();
 FILLCELL_X32 FILLER_359_1057 ();
 FILLCELL_X32 FILLER_359_1089 ();
 FILLCELL_X32 FILLER_359_1121 ();
 FILLCELL_X32 FILLER_359_1153 ();
 FILLCELL_X32 FILLER_359_1185 ();
 FILLCELL_X32 FILLER_359_1217 ();
 FILLCELL_X8 FILLER_359_1249 ();
 FILLCELL_X4 FILLER_359_1257 ();
 FILLCELL_X2 FILLER_359_1261 ();
 FILLCELL_X32 FILLER_359_1264 ();
 FILLCELL_X32 FILLER_359_1296 ();
 FILLCELL_X32 FILLER_359_1328 ();
 FILLCELL_X32 FILLER_359_1360 ();
 FILLCELL_X32 FILLER_359_1392 ();
 FILLCELL_X32 FILLER_359_1424 ();
 FILLCELL_X32 FILLER_359_1456 ();
 FILLCELL_X32 FILLER_359_1488 ();
 FILLCELL_X32 FILLER_359_1520 ();
 FILLCELL_X32 FILLER_359_1552 ();
 FILLCELL_X32 FILLER_359_1584 ();
 FILLCELL_X32 FILLER_359_1616 ();
 FILLCELL_X32 FILLER_359_1648 ();
 FILLCELL_X32 FILLER_359_1680 ();
 FILLCELL_X32 FILLER_359_1712 ();
 FILLCELL_X32 FILLER_359_1744 ();
 FILLCELL_X32 FILLER_359_1776 ();
 FILLCELL_X32 FILLER_359_1808 ();
 FILLCELL_X32 FILLER_359_1840 ();
 FILLCELL_X32 FILLER_359_1872 ();
 FILLCELL_X32 FILLER_359_1904 ();
 FILLCELL_X32 FILLER_359_1936 ();
 FILLCELL_X32 FILLER_359_1968 ();
 FILLCELL_X32 FILLER_359_2000 ();
 FILLCELL_X32 FILLER_359_2032 ();
 FILLCELL_X32 FILLER_359_2064 ();
 FILLCELL_X32 FILLER_359_2096 ();
 FILLCELL_X32 FILLER_359_2128 ();
 FILLCELL_X32 FILLER_359_2160 ();
 FILLCELL_X32 FILLER_359_2192 ();
 FILLCELL_X32 FILLER_359_2224 ();
 FILLCELL_X32 FILLER_359_2256 ();
 FILLCELL_X32 FILLER_359_2288 ();
 FILLCELL_X32 FILLER_359_2320 ();
 FILLCELL_X32 FILLER_359_2352 ();
 FILLCELL_X32 FILLER_359_2384 ();
 FILLCELL_X32 FILLER_359_2416 ();
 FILLCELL_X32 FILLER_359_2448 ();
 FILLCELL_X32 FILLER_359_2480 ();
 FILLCELL_X8 FILLER_359_2512 ();
 FILLCELL_X4 FILLER_359_2520 ();
 FILLCELL_X2 FILLER_359_2524 ();
 FILLCELL_X32 FILLER_359_2527 ();
 FILLCELL_X32 FILLER_359_2559 ();
 FILLCELL_X32 FILLER_359_2591 ();
 FILLCELL_X32 FILLER_359_2623 ();
 FILLCELL_X32 FILLER_359_2655 ();
 FILLCELL_X32 FILLER_359_2687 ();
 FILLCELL_X32 FILLER_359_2719 ();
 FILLCELL_X32 FILLER_359_2751 ();
 FILLCELL_X32 FILLER_359_2783 ();
 FILLCELL_X32 FILLER_359_2815 ();
 FILLCELL_X32 FILLER_359_2847 ();
 FILLCELL_X32 FILLER_359_2879 ();
 FILLCELL_X32 FILLER_359_2911 ();
 FILLCELL_X32 FILLER_359_2943 ();
 FILLCELL_X32 FILLER_359_2975 ();
 FILLCELL_X32 FILLER_359_3007 ();
 FILLCELL_X32 FILLER_359_3039 ();
 FILLCELL_X32 FILLER_359_3071 ();
 FILLCELL_X32 FILLER_359_3103 ();
 FILLCELL_X32 FILLER_359_3135 ();
 FILLCELL_X32 FILLER_359_3167 ();
 FILLCELL_X32 FILLER_359_3199 ();
 FILLCELL_X32 FILLER_359_3231 ();
 FILLCELL_X32 FILLER_359_3263 ();
 FILLCELL_X32 FILLER_359_3295 ();
 FILLCELL_X32 FILLER_359_3327 ();
 FILLCELL_X32 FILLER_359_3359 ();
 FILLCELL_X32 FILLER_359_3391 ();
 FILLCELL_X32 FILLER_359_3423 ();
 FILLCELL_X32 FILLER_359_3455 ();
 FILLCELL_X32 FILLER_359_3487 ();
 FILLCELL_X32 FILLER_359_3519 ();
 FILLCELL_X32 FILLER_359_3551 ();
 FILLCELL_X32 FILLER_359_3583 ();
 FILLCELL_X32 FILLER_359_3615 ();
 FILLCELL_X32 FILLER_359_3647 ();
 FILLCELL_X32 FILLER_359_3679 ();
 FILLCELL_X16 FILLER_359_3711 ();
 FILLCELL_X8 FILLER_359_3727 ();
 FILLCELL_X2 FILLER_359_3735 ();
 FILLCELL_X1 FILLER_359_3737 ();
 FILLCELL_X32 FILLER_360_1 ();
 FILLCELL_X32 FILLER_360_33 ();
 FILLCELL_X32 FILLER_360_65 ();
 FILLCELL_X32 FILLER_360_97 ();
 FILLCELL_X32 FILLER_360_129 ();
 FILLCELL_X32 FILLER_360_161 ();
 FILLCELL_X32 FILLER_360_193 ();
 FILLCELL_X32 FILLER_360_225 ();
 FILLCELL_X32 FILLER_360_257 ();
 FILLCELL_X32 FILLER_360_289 ();
 FILLCELL_X32 FILLER_360_321 ();
 FILLCELL_X32 FILLER_360_353 ();
 FILLCELL_X32 FILLER_360_385 ();
 FILLCELL_X32 FILLER_360_417 ();
 FILLCELL_X32 FILLER_360_449 ();
 FILLCELL_X32 FILLER_360_481 ();
 FILLCELL_X32 FILLER_360_513 ();
 FILLCELL_X32 FILLER_360_545 ();
 FILLCELL_X32 FILLER_360_577 ();
 FILLCELL_X16 FILLER_360_609 ();
 FILLCELL_X4 FILLER_360_625 ();
 FILLCELL_X2 FILLER_360_629 ();
 FILLCELL_X32 FILLER_360_632 ();
 FILLCELL_X32 FILLER_360_664 ();
 FILLCELL_X32 FILLER_360_696 ();
 FILLCELL_X32 FILLER_360_728 ();
 FILLCELL_X32 FILLER_360_760 ();
 FILLCELL_X32 FILLER_360_792 ();
 FILLCELL_X32 FILLER_360_824 ();
 FILLCELL_X32 FILLER_360_856 ();
 FILLCELL_X32 FILLER_360_888 ();
 FILLCELL_X32 FILLER_360_920 ();
 FILLCELL_X32 FILLER_360_952 ();
 FILLCELL_X32 FILLER_360_984 ();
 FILLCELL_X32 FILLER_360_1016 ();
 FILLCELL_X32 FILLER_360_1048 ();
 FILLCELL_X32 FILLER_360_1080 ();
 FILLCELL_X32 FILLER_360_1112 ();
 FILLCELL_X32 FILLER_360_1144 ();
 FILLCELL_X32 FILLER_360_1176 ();
 FILLCELL_X32 FILLER_360_1208 ();
 FILLCELL_X32 FILLER_360_1240 ();
 FILLCELL_X32 FILLER_360_1272 ();
 FILLCELL_X32 FILLER_360_1304 ();
 FILLCELL_X32 FILLER_360_1336 ();
 FILLCELL_X32 FILLER_360_1368 ();
 FILLCELL_X32 FILLER_360_1400 ();
 FILLCELL_X32 FILLER_360_1432 ();
 FILLCELL_X32 FILLER_360_1464 ();
 FILLCELL_X32 FILLER_360_1496 ();
 FILLCELL_X32 FILLER_360_1528 ();
 FILLCELL_X32 FILLER_360_1560 ();
 FILLCELL_X32 FILLER_360_1592 ();
 FILLCELL_X32 FILLER_360_1624 ();
 FILLCELL_X32 FILLER_360_1656 ();
 FILLCELL_X32 FILLER_360_1688 ();
 FILLCELL_X32 FILLER_360_1720 ();
 FILLCELL_X32 FILLER_360_1752 ();
 FILLCELL_X32 FILLER_360_1784 ();
 FILLCELL_X32 FILLER_360_1816 ();
 FILLCELL_X32 FILLER_360_1848 ();
 FILLCELL_X8 FILLER_360_1880 ();
 FILLCELL_X4 FILLER_360_1888 ();
 FILLCELL_X2 FILLER_360_1892 ();
 FILLCELL_X32 FILLER_360_1895 ();
 FILLCELL_X32 FILLER_360_1927 ();
 FILLCELL_X32 FILLER_360_1959 ();
 FILLCELL_X32 FILLER_360_1991 ();
 FILLCELL_X32 FILLER_360_2023 ();
 FILLCELL_X32 FILLER_360_2055 ();
 FILLCELL_X32 FILLER_360_2087 ();
 FILLCELL_X32 FILLER_360_2119 ();
 FILLCELL_X32 FILLER_360_2151 ();
 FILLCELL_X32 FILLER_360_2183 ();
 FILLCELL_X32 FILLER_360_2215 ();
 FILLCELL_X32 FILLER_360_2247 ();
 FILLCELL_X32 FILLER_360_2279 ();
 FILLCELL_X32 FILLER_360_2311 ();
 FILLCELL_X32 FILLER_360_2343 ();
 FILLCELL_X32 FILLER_360_2375 ();
 FILLCELL_X32 FILLER_360_2407 ();
 FILLCELL_X32 FILLER_360_2439 ();
 FILLCELL_X32 FILLER_360_2471 ();
 FILLCELL_X32 FILLER_360_2503 ();
 FILLCELL_X32 FILLER_360_2535 ();
 FILLCELL_X32 FILLER_360_2567 ();
 FILLCELL_X32 FILLER_360_2599 ();
 FILLCELL_X32 FILLER_360_2631 ();
 FILLCELL_X32 FILLER_360_2663 ();
 FILLCELL_X32 FILLER_360_2695 ();
 FILLCELL_X32 FILLER_360_2727 ();
 FILLCELL_X32 FILLER_360_2759 ();
 FILLCELL_X32 FILLER_360_2791 ();
 FILLCELL_X32 FILLER_360_2823 ();
 FILLCELL_X32 FILLER_360_2855 ();
 FILLCELL_X32 FILLER_360_2887 ();
 FILLCELL_X32 FILLER_360_2919 ();
 FILLCELL_X32 FILLER_360_2951 ();
 FILLCELL_X32 FILLER_360_2983 ();
 FILLCELL_X32 FILLER_360_3015 ();
 FILLCELL_X32 FILLER_360_3047 ();
 FILLCELL_X32 FILLER_360_3079 ();
 FILLCELL_X32 FILLER_360_3111 ();
 FILLCELL_X8 FILLER_360_3143 ();
 FILLCELL_X4 FILLER_360_3151 ();
 FILLCELL_X2 FILLER_360_3155 ();
 FILLCELL_X32 FILLER_360_3158 ();
 FILLCELL_X32 FILLER_360_3190 ();
 FILLCELL_X32 FILLER_360_3222 ();
 FILLCELL_X32 FILLER_360_3254 ();
 FILLCELL_X32 FILLER_360_3286 ();
 FILLCELL_X32 FILLER_360_3318 ();
 FILLCELL_X32 FILLER_360_3350 ();
 FILLCELL_X32 FILLER_360_3382 ();
 FILLCELL_X32 FILLER_360_3414 ();
 FILLCELL_X32 FILLER_360_3446 ();
 FILLCELL_X32 FILLER_360_3478 ();
 FILLCELL_X32 FILLER_360_3510 ();
 FILLCELL_X32 FILLER_360_3542 ();
 FILLCELL_X32 FILLER_360_3574 ();
 FILLCELL_X32 FILLER_360_3606 ();
 FILLCELL_X32 FILLER_360_3638 ();
 FILLCELL_X32 FILLER_360_3670 ();
 FILLCELL_X32 FILLER_360_3702 ();
 FILLCELL_X4 FILLER_360_3734 ();
 FILLCELL_X32 FILLER_361_1 ();
 FILLCELL_X32 FILLER_361_33 ();
 FILLCELL_X32 FILLER_361_65 ();
 FILLCELL_X32 FILLER_361_97 ();
 FILLCELL_X32 FILLER_361_129 ();
 FILLCELL_X32 FILLER_361_161 ();
 FILLCELL_X32 FILLER_361_193 ();
 FILLCELL_X32 FILLER_361_225 ();
 FILLCELL_X32 FILLER_361_257 ();
 FILLCELL_X32 FILLER_361_289 ();
 FILLCELL_X32 FILLER_361_321 ();
 FILLCELL_X32 FILLER_361_353 ();
 FILLCELL_X32 FILLER_361_385 ();
 FILLCELL_X32 FILLER_361_417 ();
 FILLCELL_X32 FILLER_361_449 ();
 FILLCELL_X32 FILLER_361_481 ();
 FILLCELL_X32 FILLER_361_513 ();
 FILLCELL_X32 FILLER_361_545 ();
 FILLCELL_X32 FILLER_361_577 ();
 FILLCELL_X32 FILLER_361_609 ();
 FILLCELL_X32 FILLER_361_641 ();
 FILLCELL_X32 FILLER_361_673 ();
 FILLCELL_X32 FILLER_361_705 ();
 FILLCELL_X32 FILLER_361_737 ();
 FILLCELL_X32 FILLER_361_769 ();
 FILLCELL_X32 FILLER_361_801 ();
 FILLCELL_X32 FILLER_361_833 ();
 FILLCELL_X32 FILLER_361_865 ();
 FILLCELL_X32 FILLER_361_897 ();
 FILLCELL_X32 FILLER_361_929 ();
 FILLCELL_X32 FILLER_361_961 ();
 FILLCELL_X32 FILLER_361_993 ();
 FILLCELL_X32 FILLER_361_1025 ();
 FILLCELL_X32 FILLER_361_1057 ();
 FILLCELL_X32 FILLER_361_1089 ();
 FILLCELL_X32 FILLER_361_1121 ();
 FILLCELL_X32 FILLER_361_1153 ();
 FILLCELL_X32 FILLER_361_1185 ();
 FILLCELL_X32 FILLER_361_1217 ();
 FILLCELL_X8 FILLER_361_1249 ();
 FILLCELL_X4 FILLER_361_1257 ();
 FILLCELL_X2 FILLER_361_1261 ();
 FILLCELL_X32 FILLER_361_1264 ();
 FILLCELL_X32 FILLER_361_1296 ();
 FILLCELL_X32 FILLER_361_1328 ();
 FILLCELL_X32 FILLER_361_1360 ();
 FILLCELL_X32 FILLER_361_1392 ();
 FILLCELL_X32 FILLER_361_1424 ();
 FILLCELL_X32 FILLER_361_1456 ();
 FILLCELL_X32 FILLER_361_1488 ();
 FILLCELL_X32 FILLER_361_1520 ();
 FILLCELL_X32 FILLER_361_1552 ();
 FILLCELL_X32 FILLER_361_1584 ();
 FILLCELL_X32 FILLER_361_1616 ();
 FILLCELL_X32 FILLER_361_1648 ();
 FILLCELL_X32 FILLER_361_1680 ();
 FILLCELL_X32 FILLER_361_1712 ();
 FILLCELL_X32 FILLER_361_1744 ();
 FILLCELL_X32 FILLER_361_1776 ();
 FILLCELL_X32 FILLER_361_1808 ();
 FILLCELL_X32 FILLER_361_1840 ();
 FILLCELL_X32 FILLER_361_1872 ();
 FILLCELL_X32 FILLER_361_1904 ();
 FILLCELL_X32 FILLER_361_1936 ();
 FILLCELL_X32 FILLER_361_1968 ();
 FILLCELL_X32 FILLER_361_2000 ();
 FILLCELL_X32 FILLER_361_2032 ();
 FILLCELL_X32 FILLER_361_2064 ();
 FILLCELL_X32 FILLER_361_2096 ();
 FILLCELL_X32 FILLER_361_2128 ();
 FILLCELL_X32 FILLER_361_2160 ();
 FILLCELL_X32 FILLER_361_2192 ();
 FILLCELL_X32 FILLER_361_2224 ();
 FILLCELL_X32 FILLER_361_2256 ();
 FILLCELL_X32 FILLER_361_2288 ();
 FILLCELL_X32 FILLER_361_2320 ();
 FILLCELL_X32 FILLER_361_2352 ();
 FILLCELL_X32 FILLER_361_2384 ();
 FILLCELL_X32 FILLER_361_2416 ();
 FILLCELL_X32 FILLER_361_2448 ();
 FILLCELL_X32 FILLER_361_2480 ();
 FILLCELL_X8 FILLER_361_2512 ();
 FILLCELL_X4 FILLER_361_2520 ();
 FILLCELL_X2 FILLER_361_2524 ();
 FILLCELL_X32 FILLER_361_2527 ();
 FILLCELL_X32 FILLER_361_2559 ();
 FILLCELL_X32 FILLER_361_2591 ();
 FILLCELL_X32 FILLER_361_2623 ();
 FILLCELL_X32 FILLER_361_2655 ();
 FILLCELL_X32 FILLER_361_2687 ();
 FILLCELL_X32 FILLER_361_2719 ();
 FILLCELL_X32 FILLER_361_2751 ();
 FILLCELL_X32 FILLER_361_2783 ();
 FILLCELL_X32 FILLER_361_2815 ();
 FILLCELL_X32 FILLER_361_2847 ();
 FILLCELL_X32 FILLER_361_2879 ();
 FILLCELL_X32 FILLER_361_2911 ();
 FILLCELL_X32 FILLER_361_2943 ();
 FILLCELL_X32 FILLER_361_2975 ();
 FILLCELL_X32 FILLER_361_3007 ();
 FILLCELL_X32 FILLER_361_3039 ();
 FILLCELL_X32 FILLER_361_3071 ();
 FILLCELL_X32 FILLER_361_3103 ();
 FILLCELL_X32 FILLER_361_3135 ();
 FILLCELL_X32 FILLER_361_3167 ();
 FILLCELL_X32 FILLER_361_3199 ();
 FILLCELL_X32 FILLER_361_3231 ();
 FILLCELL_X32 FILLER_361_3263 ();
 FILLCELL_X32 FILLER_361_3295 ();
 FILLCELL_X32 FILLER_361_3327 ();
 FILLCELL_X32 FILLER_361_3359 ();
 FILLCELL_X32 FILLER_361_3391 ();
 FILLCELL_X32 FILLER_361_3423 ();
 FILLCELL_X32 FILLER_361_3455 ();
 FILLCELL_X32 FILLER_361_3487 ();
 FILLCELL_X32 FILLER_361_3519 ();
 FILLCELL_X32 FILLER_361_3551 ();
 FILLCELL_X32 FILLER_361_3583 ();
 FILLCELL_X32 FILLER_361_3615 ();
 FILLCELL_X32 FILLER_361_3647 ();
 FILLCELL_X32 FILLER_361_3679 ();
 FILLCELL_X16 FILLER_361_3711 ();
 FILLCELL_X8 FILLER_361_3727 ();
 FILLCELL_X2 FILLER_361_3735 ();
 FILLCELL_X1 FILLER_361_3737 ();
 FILLCELL_X32 FILLER_362_1 ();
 FILLCELL_X32 FILLER_362_33 ();
 FILLCELL_X32 FILLER_362_65 ();
 FILLCELL_X32 FILLER_362_97 ();
 FILLCELL_X32 FILLER_362_129 ();
 FILLCELL_X32 FILLER_362_161 ();
 FILLCELL_X32 FILLER_362_193 ();
 FILLCELL_X32 FILLER_362_225 ();
 FILLCELL_X32 FILLER_362_257 ();
 FILLCELL_X32 FILLER_362_289 ();
 FILLCELL_X32 FILLER_362_321 ();
 FILLCELL_X32 FILLER_362_353 ();
 FILLCELL_X32 FILLER_362_385 ();
 FILLCELL_X32 FILLER_362_417 ();
 FILLCELL_X32 FILLER_362_449 ();
 FILLCELL_X32 FILLER_362_481 ();
 FILLCELL_X32 FILLER_362_513 ();
 FILLCELL_X32 FILLER_362_545 ();
 FILLCELL_X32 FILLER_362_577 ();
 FILLCELL_X16 FILLER_362_609 ();
 FILLCELL_X4 FILLER_362_625 ();
 FILLCELL_X2 FILLER_362_629 ();
 FILLCELL_X32 FILLER_362_632 ();
 FILLCELL_X32 FILLER_362_664 ();
 FILLCELL_X32 FILLER_362_696 ();
 FILLCELL_X32 FILLER_362_728 ();
 FILLCELL_X32 FILLER_362_760 ();
 FILLCELL_X32 FILLER_362_792 ();
 FILLCELL_X32 FILLER_362_824 ();
 FILLCELL_X32 FILLER_362_856 ();
 FILLCELL_X32 FILLER_362_888 ();
 FILLCELL_X32 FILLER_362_920 ();
 FILLCELL_X32 FILLER_362_952 ();
 FILLCELL_X32 FILLER_362_984 ();
 FILLCELL_X32 FILLER_362_1016 ();
 FILLCELL_X32 FILLER_362_1048 ();
 FILLCELL_X32 FILLER_362_1080 ();
 FILLCELL_X32 FILLER_362_1112 ();
 FILLCELL_X32 FILLER_362_1144 ();
 FILLCELL_X32 FILLER_362_1176 ();
 FILLCELL_X32 FILLER_362_1208 ();
 FILLCELL_X32 FILLER_362_1240 ();
 FILLCELL_X32 FILLER_362_1272 ();
 FILLCELL_X32 FILLER_362_1304 ();
 FILLCELL_X32 FILLER_362_1336 ();
 FILLCELL_X32 FILLER_362_1368 ();
 FILLCELL_X32 FILLER_362_1400 ();
 FILLCELL_X32 FILLER_362_1432 ();
 FILLCELL_X32 FILLER_362_1464 ();
 FILLCELL_X32 FILLER_362_1496 ();
 FILLCELL_X32 FILLER_362_1528 ();
 FILLCELL_X32 FILLER_362_1560 ();
 FILLCELL_X32 FILLER_362_1592 ();
 FILLCELL_X32 FILLER_362_1624 ();
 FILLCELL_X32 FILLER_362_1656 ();
 FILLCELL_X32 FILLER_362_1688 ();
 FILLCELL_X32 FILLER_362_1720 ();
 FILLCELL_X32 FILLER_362_1752 ();
 FILLCELL_X32 FILLER_362_1784 ();
 FILLCELL_X32 FILLER_362_1816 ();
 FILLCELL_X32 FILLER_362_1848 ();
 FILLCELL_X8 FILLER_362_1880 ();
 FILLCELL_X4 FILLER_362_1888 ();
 FILLCELL_X2 FILLER_362_1892 ();
 FILLCELL_X32 FILLER_362_1895 ();
 FILLCELL_X32 FILLER_362_1927 ();
 FILLCELL_X32 FILLER_362_1959 ();
 FILLCELL_X32 FILLER_362_1991 ();
 FILLCELL_X32 FILLER_362_2023 ();
 FILLCELL_X32 FILLER_362_2055 ();
 FILLCELL_X32 FILLER_362_2087 ();
 FILLCELL_X32 FILLER_362_2119 ();
 FILLCELL_X32 FILLER_362_2151 ();
 FILLCELL_X32 FILLER_362_2183 ();
 FILLCELL_X32 FILLER_362_2215 ();
 FILLCELL_X32 FILLER_362_2247 ();
 FILLCELL_X32 FILLER_362_2279 ();
 FILLCELL_X32 FILLER_362_2311 ();
 FILLCELL_X32 FILLER_362_2343 ();
 FILLCELL_X32 FILLER_362_2375 ();
 FILLCELL_X32 FILLER_362_2407 ();
 FILLCELL_X32 FILLER_362_2439 ();
 FILLCELL_X32 FILLER_362_2471 ();
 FILLCELL_X32 FILLER_362_2503 ();
 FILLCELL_X32 FILLER_362_2535 ();
 FILLCELL_X32 FILLER_362_2567 ();
 FILLCELL_X32 FILLER_362_2599 ();
 FILLCELL_X32 FILLER_362_2631 ();
 FILLCELL_X32 FILLER_362_2663 ();
 FILLCELL_X32 FILLER_362_2695 ();
 FILLCELL_X32 FILLER_362_2727 ();
 FILLCELL_X32 FILLER_362_2759 ();
 FILLCELL_X32 FILLER_362_2791 ();
 FILLCELL_X32 FILLER_362_2823 ();
 FILLCELL_X32 FILLER_362_2855 ();
 FILLCELL_X32 FILLER_362_2887 ();
 FILLCELL_X32 FILLER_362_2919 ();
 FILLCELL_X32 FILLER_362_2951 ();
 FILLCELL_X32 FILLER_362_2983 ();
 FILLCELL_X32 FILLER_362_3015 ();
 FILLCELL_X32 FILLER_362_3047 ();
 FILLCELL_X32 FILLER_362_3079 ();
 FILLCELL_X32 FILLER_362_3111 ();
 FILLCELL_X8 FILLER_362_3143 ();
 FILLCELL_X4 FILLER_362_3151 ();
 FILLCELL_X2 FILLER_362_3155 ();
 FILLCELL_X32 FILLER_362_3158 ();
 FILLCELL_X32 FILLER_362_3190 ();
 FILLCELL_X32 FILLER_362_3222 ();
 FILLCELL_X32 FILLER_362_3254 ();
 FILLCELL_X32 FILLER_362_3286 ();
 FILLCELL_X32 FILLER_362_3318 ();
 FILLCELL_X32 FILLER_362_3350 ();
 FILLCELL_X32 FILLER_362_3382 ();
 FILLCELL_X32 FILLER_362_3414 ();
 FILLCELL_X32 FILLER_362_3446 ();
 FILLCELL_X32 FILLER_362_3478 ();
 FILLCELL_X32 FILLER_362_3510 ();
 FILLCELL_X32 FILLER_362_3542 ();
 FILLCELL_X32 FILLER_362_3574 ();
 FILLCELL_X32 FILLER_362_3606 ();
 FILLCELL_X32 FILLER_362_3638 ();
 FILLCELL_X32 FILLER_362_3670 ();
 FILLCELL_X32 FILLER_362_3702 ();
 FILLCELL_X4 FILLER_362_3734 ();
 FILLCELL_X32 FILLER_363_1 ();
 FILLCELL_X32 FILLER_363_33 ();
 FILLCELL_X32 FILLER_363_65 ();
 FILLCELL_X32 FILLER_363_97 ();
 FILLCELL_X32 FILLER_363_129 ();
 FILLCELL_X32 FILLER_363_161 ();
 FILLCELL_X32 FILLER_363_193 ();
 FILLCELL_X32 FILLER_363_225 ();
 FILLCELL_X32 FILLER_363_257 ();
 FILLCELL_X32 FILLER_363_289 ();
 FILLCELL_X32 FILLER_363_321 ();
 FILLCELL_X32 FILLER_363_353 ();
 FILLCELL_X32 FILLER_363_385 ();
 FILLCELL_X32 FILLER_363_417 ();
 FILLCELL_X32 FILLER_363_449 ();
 FILLCELL_X32 FILLER_363_481 ();
 FILLCELL_X32 FILLER_363_513 ();
 FILLCELL_X32 FILLER_363_545 ();
 FILLCELL_X32 FILLER_363_577 ();
 FILLCELL_X32 FILLER_363_609 ();
 FILLCELL_X32 FILLER_363_641 ();
 FILLCELL_X32 FILLER_363_673 ();
 FILLCELL_X32 FILLER_363_705 ();
 FILLCELL_X32 FILLER_363_737 ();
 FILLCELL_X32 FILLER_363_769 ();
 FILLCELL_X32 FILLER_363_801 ();
 FILLCELL_X32 FILLER_363_833 ();
 FILLCELL_X32 FILLER_363_865 ();
 FILLCELL_X32 FILLER_363_897 ();
 FILLCELL_X32 FILLER_363_929 ();
 FILLCELL_X32 FILLER_363_961 ();
 FILLCELL_X32 FILLER_363_993 ();
 FILLCELL_X32 FILLER_363_1025 ();
 FILLCELL_X32 FILLER_363_1057 ();
 FILLCELL_X32 FILLER_363_1089 ();
 FILLCELL_X32 FILLER_363_1121 ();
 FILLCELL_X32 FILLER_363_1153 ();
 FILLCELL_X32 FILLER_363_1185 ();
 FILLCELL_X32 FILLER_363_1217 ();
 FILLCELL_X8 FILLER_363_1249 ();
 FILLCELL_X4 FILLER_363_1257 ();
 FILLCELL_X2 FILLER_363_1261 ();
 FILLCELL_X32 FILLER_363_1264 ();
 FILLCELL_X32 FILLER_363_1296 ();
 FILLCELL_X32 FILLER_363_1328 ();
 FILLCELL_X32 FILLER_363_1360 ();
 FILLCELL_X32 FILLER_363_1392 ();
 FILLCELL_X32 FILLER_363_1424 ();
 FILLCELL_X32 FILLER_363_1456 ();
 FILLCELL_X32 FILLER_363_1488 ();
 FILLCELL_X32 FILLER_363_1520 ();
 FILLCELL_X32 FILLER_363_1552 ();
 FILLCELL_X32 FILLER_363_1584 ();
 FILLCELL_X32 FILLER_363_1616 ();
 FILLCELL_X32 FILLER_363_1648 ();
 FILLCELL_X32 FILLER_363_1680 ();
 FILLCELL_X32 FILLER_363_1712 ();
 FILLCELL_X32 FILLER_363_1744 ();
 FILLCELL_X32 FILLER_363_1776 ();
 FILLCELL_X32 FILLER_363_1808 ();
 FILLCELL_X32 FILLER_363_1840 ();
 FILLCELL_X32 FILLER_363_1872 ();
 FILLCELL_X32 FILLER_363_1904 ();
 FILLCELL_X32 FILLER_363_1936 ();
 FILLCELL_X32 FILLER_363_1968 ();
 FILLCELL_X32 FILLER_363_2000 ();
 FILLCELL_X32 FILLER_363_2032 ();
 FILLCELL_X32 FILLER_363_2064 ();
 FILLCELL_X32 FILLER_363_2096 ();
 FILLCELL_X32 FILLER_363_2128 ();
 FILLCELL_X32 FILLER_363_2160 ();
 FILLCELL_X32 FILLER_363_2192 ();
 FILLCELL_X32 FILLER_363_2224 ();
 FILLCELL_X32 FILLER_363_2256 ();
 FILLCELL_X32 FILLER_363_2288 ();
 FILLCELL_X32 FILLER_363_2320 ();
 FILLCELL_X32 FILLER_363_2352 ();
 FILLCELL_X32 FILLER_363_2384 ();
 FILLCELL_X32 FILLER_363_2416 ();
 FILLCELL_X32 FILLER_363_2448 ();
 FILLCELL_X32 FILLER_363_2480 ();
 FILLCELL_X8 FILLER_363_2512 ();
 FILLCELL_X4 FILLER_363_2520 ();
 FILLCELL_X2 FILLER_363_2524 ();
 FILLCELL_X32 FILLER_363_2527 ();
 FILLCELL_X32 FILLER_363_2559 ();
 FILLCELL_X32 FILLER_363_2591 ();
 FILLCELL_X32 FILLER_363_2623 ();
 FILLCELL_X32 FILLER_363_2655 ();
 FILLCELL_X32 FILLER_363_2687 ();
 FILLCELL_X32 FILLER_363_2719 ();
 FILLCELL_X32 FILLER_363_2751 ();
 FILLCELL_X32 FILLER_363_2783 ();
 FILLCELL_X32 FILLER_363_2815 ();
 FILLCELL_X32 FILLER_363_2847 ();
 FILLCELL_X32 FILLER_363_2879 ();
 FILLCELL_X32 FILLER_363_2911 ();
 FILLCELL_X32 FILLER_363_2943 ();
 FILLCELL_X32 FILLER_363_2975 ();
 FILLCELL_X32 FILLER_363_3007 ();
 FILLCELL_X32 FILLER_363_3039 ();
 FILLCELL_X32 FILLER_363_3071 ();
 FILLCELL_X32 FILLER_363_3103 ();
 FILLCELL_X32 FILLER_363_3135 ();
 FILLCELL_X32 FILLER_363_3167 ();
 FILLCELL_X32 FILLER_363_3199 ();
 FILLCELL_X32 FILLER_363_3231 ();
 FILLCELL_X32 FILLER_363_3263 ();
 FILLCELL_X32 FILLER_363_3295 ();
 FILLCELL_X32 FILLER_363_3327 ();
 FILLCELL_X32 FILLER_363_3359 ();
 FILLCELL_X32 FILLER_363_3391 ();
 FILLCELL_X32 FILLER_363_3423 ();
 FILLCELL_X32 FILLER_363_3455 ();
 FILLCELL_X32 FILLER_363_3487 ();
 FILLCELL_X32 FILLER_363_3519 ();
 FILLCELL_X32 FILLER_363_3551 ();
 FILLCELL_X32 FILLER_363_3583 ();
 FILLCELL_X32 FILLER_363_3615 ();
 FILLCELL_X32 FILLER_363_3647 ();
 FILLCELL_X32 FILLER_363_3679 ();
 FILLCELL_X16 FILLER_363_3711 ();
 FILLCELL_X8 FILLER_363_3727 ();
 FILLCELL_X2 FILLER_363_3735 ();
 FILLCELL_X1 FILLER_363_3737 ();
 FILLCELL_X32 FILLER_364_1 ();
 FILLCELL_X32 FILLER_364_33 ();
 FILLCELL_X32 FILLER_364_65 ();
 FILLCELL_X32 FILLER_364_97 ();
 FILLCELL_X32 FILLER_364_129 ();
 FILLCELL_X32 FILLER_364_161 ();
 FILLCELL_X32 FILLER_364_193 ();
 FILLCELL_X32 FILLER_364_225 ();
 FILLCELL_X32 FILLER_364_257 ();
 FILLCELL_X32 FILLER_364_289 ();
 FILLCELL_X32 FILLER_364_321 ();
 FILLCELL_X32 FILLER_364_353 ();
 FILLCELL_X32 FILLER_364_385 ();
 FILLCELL_X32 FILLER_364_417 ();
 FILLCELL_X32 FILLER_364_449 ();
 FILLCELL_X32 FILLER_364_481 ();
 FILLCELL_X32 FILLER_364_513 ();
 FILLCELL_X32 FILLER_364_545 ();
 FILLCELL_X32 FILLER_364_577 ();
 FILLCELL_X16 FILLER_364_609 ();
 FILLCELL_X4 FILLER_364_625 ();
 FILLCELL_X2 FILLER_364_629 ();
 FILLCELL_X32 FILLER_364_632 ();
 FILLCELL_X32 FILLER_364_664 ();
 FILLCELL_X32 FILLER_364_696 ();
 FILLCELL_X32 FILLER_364_728 ();
 FILLCELL_X32 FILLER_364_760 ();
 FILLCELL_X32 FILLER_364_792 ();
 FILLCELL_X32 FILLER_364_824 ();
 FILLCELL_X32 FILLER_364_856 ();
 FILLCELL_X32 FILLER_364_888 ();
 FILLCELL_X32 FILLER_364_920 ();
 FILLCELL_X32 FILLER_364_952 ();
 FILLCELL_X32 FILLER_364_984 ();
 FILLCELL_X32 FILLER_364_1016 ();
 FILLCELL_X32 FILLER_364_1048 ();
 FILLCELL_X32 FILLER_364_1080 ();
 FILLCELL_X32 FILLER_364_1112 ();
 FILLCELL_X32 FILLER_364_1144 ();
 FILLCELL_X32 FILLER_364_1176 ();
 FILLCELL_X32 FILLER_364_1208 ();
 FILLCELL_X32 FILLER_364_1240 ();
 FILLCELL_X32 FILLER_364_1272 ();
 FILLCELL_X32 FILLER_364_1304 ();
 FILLCELL_X32 FILLER_364_1336 ();
 FILLCELL_X32 FILLER_364_1368 ();
 FILLCELL_X32 FILLER_364_1400 ();
 FILLCELL_X32 FILLER_364_1432 ();
 FILLCELL_X32 FILLER_364_1464 ();
 FILLCELL_X32 FILLER_364_1496 ();
 FILLCELL_X32 FILLER_364_1528 ();
 FILLCELL_X32 FILLER_364_1560 ();
 FILLCELL_X32 FILLER_364_1592 ();
 FILLCELL_X32 FILLER_364_1624 ();
 FILLCELL_X32 FILLER_364_1656 ();
 FILLCELL_X32 FILLER_364_1688 ();
 FILLCELL_X32 FILLER_364_1720 ();
 FILLCELL_X32 FILLER_364_1752 ();
 FILLCELL_X32 FILLER_364_1784 ();
 FILLCELL_X32 FILLER_364_1816 ();
 FILLCELL_X32 FILLER_364_1848 ();
 FILLCELL_X8 FILLER_364_1880 ();
 FILLCELL_X4 FILLER_364_1888 ();
 FILLCELL_X2 FILLER_364_1892 ();
 FILLCELL_X32 FILLER_364_1895 ();
 FILLCELL_X32 FILLER_364_1927 ();
 FILLCELL_X32 FILLER_364_1959 ();
 FILLCELL_X32 FILLER_364_1991 ();
 FILLCELL_X32 FILLER_364_2023 ();
 FILLCELL_X32 FILLER_364_2055 ();
 FILLCELL_X32 FILLER_364_2087 ();
 FILLCELL_X32 FILLER_364_2119 ();
 FILLCELL_X32 FILLER_364_2151 ();
 FILLCELL_X32 FILLER_364_2183 ();
 FILLCELL_X32 FILLER_364_2215 ();
 FILLCELL_X32 FILLER_364_2247 ();
 FILLCELL_X32 FILLER_364_2279 ();
 FILLCELL_X32 FILLER_364_2311 ();
 FILLCELL_X32 FILLER_364_2343 ();
 FILLCELL_X32 FILLER_364_2375 ();
 FILLCELL_X32 FILLER_364_2407 ();
 FILLCELL_X32 FILLER_364_2439 ();
 FILLCELL_X32 FILLER_364_2471 ();
 FILLCELL_X32 FILLER_364_2503 ();
 FILLCELL_X32 FILLER_364_2535 ();
 FILLCELL_X32 FILLER_364_2567 ();
 FILLCELL_X32 FILLER_364_2599 ();
 FILLCELL_X32 FILLER_364_2631 ();
 FILLCELL_X32 FILLER_364_2663 ();
 FILLCELL_X32 FILLER_364_2695 ();
 FILLCELL_X32 FILLER_364_2727 ();
 FILLCELL_X32 FILLER_364_2759 ();
 FILLCELL_X32 FILLER_364_2791 ();
 FILLCELL_X32 FILLER_364_2823 ();
 FILLCELL_X32 FILLER_364_2855 ();
 FILLCELL_X32 FILLER_364_2887 ();
 FILLCELL_X32 FILLER_364_2919 ();
 FILLCELL_X32 FILLER_364_2951 ();
 FILLCELL_X32 FILLER_364_2983 ();
 FILLCELL_X32 FILLER_364_3015 ();
 FILLCELL_X32 FILLER_364_3047 ();
 FILLCELL_X32 FILLER_364_3079 ();
 FILLCELL_X32 FILLER_364_3111 ();
 FILLCELL_X8 FILLER_364_3143 ();
 FILLCELL_X4 FILLER_364_3151 ();
 FILLCELL_X2 FILLER_364_3155 ();
 FILLCELL_X32 FILLER_364_3158 ();
 FILLCELL_X32 FILLER_364_3190 ();
 FILLCELL_X32 FILLER_364_3222 ();
 FILLCELL_X32 FILLER_364_3254 ();
 FILLCELL_X32 FILLER_364_3286 ();
 FILLCELL_X32 FILLER_364_3318 ();
 FILLCELL_X32 FILLER_364_3350 ();
 FILLCELL_X32 FILLER_364_3382 ();
 FILLCELL_X32 FILLER_364_3414 ();
 FILLCELL_X32 FILLER_364_3446 ();
 FILLCELL_X32 FILLER_364_3478 ();
 FILLCELL_X32 FILLER_364_3510 ();
 FILLCELL_X32 FILLER_364_3542 ();
 FILLCELL_X32 FILLER_364_3574 ();
 FILLCELL_X32 FILLER_364_3606 ();
 FILLCELL_X32 FILLER_364_3638 ();
 FILLCELL_X32 FILLER_364_3670 ();
 FILLCELL_X32 FILLER_364_3702 ();
 FILLCELL_X4 FILLER_364_3734 ();
 FILLCELL_X32 FILLER_365_1 ();
 FILLCELL_X32 FILLER_365_33 ();
 FILLCELL_X32 FILLER_365_65 ();
 FILLCELL_X32 FILLER_365_97 ();
 FILLCELL_X32 FILLER_365_129 ();
 FILLCELL_X32 FILLER_365_161 ();
 FILLCELL_X32 FILLER_365_193 ();
 FILLCELL_X32 FILLER_365_225 ();
 FILLCELL_X32 FILLER_365_257 ();
 FILLCELL_X32 FILLER_365_289 ();
 FILLCELL_X32 FILLER_365_321 ();
 FILLCELL_X32 FILLER_365_353 ();
 FILLCELL_X32 FILLER_365_385 ();
 FILLCELL_X32 FILLER_365_417 ();
 FILLCELL_X32 FILLER_365_449 ();
 FILLCELL_X32 FILLER_365_481 ();
 FILLCELL_X32 FILLER_365_513 ();
 FILLCELL_X32 FILLER_365_545 ();
 FILLCELL_X32 FILLER_365_577 ();
 FILLCELL_X32 FILLER_365_609 ();
 FILLCELL_X32 FILLER_365_641 ();
 FILLCELL_X32 FILLER_365_673 ();
 FILLCELL_X32 FILLER_365_705 ();
 FILLCELL_X32 FILLER_365_737 ();
 FILLCELL_X32 FILLER_365_769 ();
 FILLCELL_X32 FILLER_365_801 ();
 FILLCELL_X32 FILLER_365_833 ();
 FILLCELL_X32 FILLER_365_865 ();
 FILLCELL_X32 FILLER_365_897 ();
 FILLCELL_X32 FILLER_365_929 ();
 FILLCELL_X32 FILLER_365_961 ();
 FILLCELL_X32 FILLER_365_993 ();
 FILLCELL_X32 FILLER_365_1025 ();
 FILLCELL_X32 FILLER_365_1057 ();
 FILLCELL_X32 FILLER_365_1089 ();
 FILLCELL_X32 FILLER_365_1121 ();
 FILLCELL_X32 FILLER_365_1153 ();
 FILLCELL_X32 FILLER_365_1185 ();
 FILLCELL_X32 FILLER_365_1217 ();
 FILLCELL_X8 FILLER_365_1249 ();
 FILLCELL_X4 FILLER_365_1257 ();
 FILLCELL_X2 FILLER_365_1261 ();
 FILLCELL_X32 FILLER_365_1264 ();
 FILLCELL_X32 FILLER_365_1296 ();
 FILLCELL_X32 FILLER_365_1328 ();
 FILLCELL_X32 FILLER_365_1360 ();
 FILLCELL_X32 FILLER_365_1392 ();
 FILLCELL_X32 FILLER_365_1424 ();
 FILLCELL_X32 FILLER_365_1456 ();
 FILLCELL_X32 FILLER_365_1488 ();
 FILLCELL_X32 FILLER_365_1520 ();
 FILLCELL_X32 FILLER_365_1552 ();
 FILLCELL_X32 FILLER_365_1584 ();
 FILLCELL_X32 FILLER_365_1616 ();
 FILLCELL_X32 FILLER_365_1648 ();
 FILLCELL_X32 FILLER_365_1680 ();
 FILLCELL_X32 FILLER_365_1712 ();
 FILLCELL_X32 FILLER_365_1744 ();
 FILLCELL_X32 FILLER_365_1776 ();
 FILLCELL_X32 FILLER_365_1808 ();
 FILLCELL_X32 FILLER_365_1840 ();
 FILLCELL_X32 FILLER_365_1872 ();
 FILLCELL_X32 FILLER_365_1904 ();
 FILLCELL_X32 FILLER_365_1936 ();
 FILLCELL_X32 FILLER_365_1968 ();
 FILLCELL_X32 FILLER_365_2000 ();
 FILLCELL_X32 FILLER_365_2032 ();
 FILLCELL_X32 FILLER_365_2064 ();
 FILLCELL_X32 FILLER_365_2096 ();
 FILLCELL_X32 FILLER_365_2128 ();
 FILLCELL_X32 FILLER_365_2160 ();
 FILLCELL_X32 FILLER_365_2192 ();
 FILLCELL_X32 FILLER_365_2224 ();
 FILLCELL_X32 FILLER_365_2256 ();
 FILLCELL_X32 FILLER_365_2288 ();
 FILLCELL_X32 FILLER_365_2320 ();
 FILLCELL_X32 FILLER_365_2352 ();
 FILLCELL_X32 FILLER_365_2384 ();
 FILLCELL_X32 FILLER_365_2416 ();
 FILLCELL_X32 FILLER_365_2448 ();
 FILLCELL_X32 FILLER_365_2480 ();
 FILLCELL_X8 FILLER_365_2512 ();
 FILLCELL_X4 FILLER_365_2520 ();
 FILLCELL_X2 FILLER_365_2524 ();
 FILLCELL_X32 FILLER_365_2527 ();
 FILLCELL_X32 FILLER_365_2559 ();
 FILLCELL_X32 FILLER_365_2591 ();
 FILLCELL_X32 FILLER_365_2623 ();
 FILLCELL_X32 FILLER_365_2655 ();
 FILLCELL_X32 FILLER_365_2687 ();
 FILLCELL_X32 FILLER_365_2719 ();
 FILLCELL_X32 FILLER_365_2751 ();
 FILLCELL_X32 FILLER_365_2783 ();
 FILLCELL_X32 FILLER_365_2815 ();
 FILLCELL_X32 FILLER_365_2847 ();
 FILLCELL_X32 FILLER_365_2879 ();
 FILLCELL_X32 FILLER_365_2911 ();
 FILLCELL_X32 FILLER_365_2943 ();
 FILLCELL_X32 FILLER_365_2975 ();
 FILLCELL_X32 FILLER_365_3007 ();
 FILLCELL_X32 FILLER_365_3039 ();
 FILLCELL_X32 FILLER_365_3071 ();
 FILLCELL_X32 FILLER_365_3103 ();
 FILLCELL_X32 FILLER_365_3135 ();
 FILLCELL_X32 FILLER_365_3167 ();
 FILLCELL_X32 FILLER_365_3199 ();
 FILLCELL_X32 FILLER_365_3231 ();
 FILLCELL_X32 FILLER_365_3263 ();
 FILLCELL_X32 FILLER_365_3295 ();
 FILLCELL_X32 FILLER_365_3327 ();
 FILLCELL_X32 FILLER_365_3359 ();
 FILLCELL_X32 FILLER_365_3391 ();
 FILLCELL_X32 FILLER_365_3423 ();
 FILLCELL_X32 FILLER_365_3455 ();
 FILLCELL_X32 FILLER_365_3487 ();
 FILLCELL_X32 FILLER_365_3519 ();
 FILLCELL_X32 FILLER_365_3551 ();
 FILLCELL_X32 FILLER_365_3583 ();
 FILLCELL_X32 FILLER_365_3615 ();
 FILLCELL_X32 FILLER_365_3647 ();
 FILLCELL_X32 FILLER_365_3679 ();
 FILLCELL_X16 FILLER_365_3711 ();
 FILLCELL_X8 FILLER_365_3727 ();
 FILLCELL_X2 FILLER_365_3735 ();
 FILLCELL_X1 FILLER_365_3737 ();
 FILLCELL_X32 FILLER_366_1 ();
 FILLCELL_X32 FILLER_366_33 ();
 FILLCELL_X32 FILLER_366_65 ();
 FILLCELL_X32 FILLER_366_97 ();
 FILLCELL_X32 FILLER_366_129 ();
 FILLCELL_X32 FILLER_366_161 ();
 FILLCELL_X32 FILLER_366_193 ();
 FILLCELL_X32 FILLER_366_225 ();
 FILLCELL_X32 FILLER_366_257 ();
 FILLCELL_X32 FILLER_366_289 ();
 FILLCELL_X32 FILLER_366_321 ();
 FILLCELL_X32 FILLER_366_353 ();
 FILLCELL_X32 FILLER_366_385 ();
 FILLCELL_X32 FILLER_366_417 ();
 FILLCELL_X32 FILLER_366_449 ();
 FILLCELL_X32 FILLER_366_481 ();
 FILLCELL_X32 FILLER_366_513 ();
 FILLCELL_X32 FILLER_366_545 ();
 FILLCELL_X32 FILLER_366_577 ();
 FILLCELL_X16 FILLER_366_609 ();
 FILLCELL_X4 FILLER_366_625 ();
 FILLCELL_X2 FILLER_366_629 ();
 FILLCELL_X32 FILLER_366_632 ();
 FILLCELL_X32 FILLER_366_664 ();
 FILLCELL_X32 FILLER_366_696 ();
 FILLCELL_X32 FILLER_366_728 ();
 FILLCELL_X32 FILLER_366_760 ();
 FILLCELL_X32 FILLER_366_792 ();
 FILLCELL_X32 FILLER_366_824 ();
 FILLCELL_X32 FILLER_366_856 ();
 FILLCELL_X32 FILLER_366_888 ();
 FILLCELL_X32 FILLER_366_920 ();
 FILLCELL_X32 FILLER_366_952 ();
 FILLCELL_X32 FILLER_366_984 ();
 FILLCELL_X32 FILLER_366_1016 ();
 FILLCELL_X32 FILLER_366_1048 ();
 FILLCELL_X32 FILLER_366_1080 ();
 FILLCELL_X32 FILLER_366_1112 ();
 FILLCELL_X32 FILLER_366_1144 ();
 FILLCELL_X32 FILLER_366_1176 ();
 FILLCELL_X32 FILLER_366_1208 ();
 FILLCELL_X32 FILLER_366_1240 ();
 FILLCELL_X32 FILLER_366_1272 ();
 FILLCELL_X32 FILLER_366_1304 ();
 FILLCELL_X32 FILLER_366_1336 ();
 FILLCELL_X32 FILLER_366_1368 ();
 FILLCELL_X32 FILLER_366_1400 ();
 FILLCELL_X32 FILLER_366_1432 ();
 FILLCELL_X32 FILLER_366_1464 ();
 FILLCELL_X32 FILLER_366_1496 ();
 FILLCELL_X32 FILLER_366_1528 ();
 FILLCELL_X32 FILLER_366_1560 ();
 FILLCELL_X32 FILLER_366_1592 ();
 FILLCELL_X32 FILLER_366_1624 ();
 FILLCELL_X32 FILLER_366_1656 ();
 FILLCELL_X32 FILLER_366_1688 ();
 FILLCELL_X32 FILLER_366_1720 ();
 FILLCELL_X32 FILLER_366_1752 ();
 FILLCELL_X32 FILLER_366_1784 ();
 FILLCELL_X32 FILLER_366_1816 ();
 FILLCELL_X32 FILLER_366_1848 ();
 FILLCELL_X8 FILLER_366_1880 ();
 FILLCELL_X4 FILLER_366_1888 ();
 FILLCELL_X2 FILLER_366_1892 ();
 FILLCELL_X32 FILLER_366_1895 ();
 FILLCELL_X32 FILLER_366_1927 ();
 FILLCELL_X32 FILLER_366_1959 ();
 FILLCELL_X32 FILLER_366_1991 ();
 FILLCELL_X32 FILLER_366_2023 ();
 FILLCELL_X32 FILLER_366_2055 ();
 FILLCELL_X32 FILLER_366_2087 ();
 FILLCELL_X32 FILLER_366_2119 ();
 FILLCELL_X32 FILLER_366_2151 ();
 FILLCELL_X32 FILLER_366_2183 ();
 FILLCELL_X32 FILLER_366_2215 ();
 FILLCELL_X32 FILLER_366_2247 ();
 FILLCELL_X32 FILLER_366_2279 ();
 FILLCELL_X32 FILLER_366_2311 ();
 FILLCELL_X32 FILLER_366_2343 ();
 FILLCELL_X32 FILLER_366_2375 ();
 FILLCELL_X32 FILLER_366_2407 ();
 FILLCELL_X32 FILLER_366_2439 ();
 FILLCELL_X32 FILLER_366_2471 ();
 FILLCELL_X32 FILLER_366_2503 ();
 FILLCELL_X32 FILLER_366_2535 ();
 FILLCELL_X32 FILLER_366_2567 ();
 FILLCELL_X32 FILLER_366_2599 ();
 FILLCELL_X32 FILLER_366_2631 ();
 FILLCELL_X32 FILLER_366_2663 ();
 FILLCELL_X32 FILLER_366_2695 ();
 FILLCELL_X32 FILLER_366_2727 ();
 FILLCELL_X32 FILLER_366_2759 ();
 FILLCELL_X32 FILLER_366_2791 ();
 FILLCELL_X32 FILLER_366_2823 ();
 FILLCELL_X32 FILLER_366_2855 ();
 FILLCELL_X32 FILLER_366_2887 ();
 FILLCELL_X32 FILLER_366_2919 ();
 FILLCELL_X32 FILLER_366_2951 ();
 FILLCELL_X32 FILLER_366_2983 ();
 FILLCELL_X32 FILLER_366_3015 ();
 FILLCELL_X32 FILLER_366_3047 ();
 FILLCELL_X32 FILLER_366_3079 ();
 FILLCELL_X32 FILLER_366_3111 ();
 FILLCELL_X8 FILLER_366_3143 ();
 FILLCELL_X4 FILLER_366_3151 ();
 FILLCELL_X2 FILLER_366_3155 ();
 FILLCELL_X32 FILLER_366_3158 ();
 FILLCELL_X32 FILLER_366_3190 ();
 FILLCELL_X32 FILLER_366_3222 ();
 FILLCELL_X32 FILLER_366_3254 ();
 FILLCELL_X32 FILLER_366_3286 ();
 FILLCELL_X32 FILLER_366_3318 ();
 FILLCELL_X32 FILLER_366_3350 ();
 FILLCELL_X32 FILLER_366_3382 ();
 FILLCELL_X32 FILLER_366_3414 ();
 FILLCELL_X32 FILLER_366_3446 ();
 FILLCELL_X32 FILLER_366_3478 ();
 FILLCELL_X32 FILLER_366_3510 ();
 FILLCELL_X32 FILLER_366_3542 ();
 FILLCELL_X32 FILLER_366_3574 ();
 FILLCELL_X32 FILLER_366_3606 ();
 FILLCELL_X32 FILLER_366_3638 ();
 FILLCELL_X32 FILLER_366_3670 ();
 FILLCELL_X32 FILLER_366_3702 ();
 FILLCELL_X4 FILLER_366_3734 ();
 FILLCELL_X32 FILLER_367_1 ();
 FILLCELL_X32 FILLER_367_33 ();
 FILLCELL_X32 FILLER_367_65 ();
 FILLCELL_X32 FILLER_367_97 ();
 FILLCELL_X32 FILLER_367_129 ();
 FILLCELL_X32 FILLER_367_161 ();
 FILLCELL_X32 FILLER_367_193 ();
 FILLCELL_X32 FILLER_367_225 ();
 FILLCELL_X32 FILLER_367_257 ();
 FILLCELL_X32 FILLER_367_289 ();
 FILLCELL_X32 FILLER_367_321 ();
 FILLCELL_X32 FILLER_367_353 ();
 FILLCELL_X32 FILLER_367_385 ();
 FILLCELL_X32 FILLER_367_417 ();
 FILLCELL_X32 FILLER_367_449 ();
 FILLCELL_X32 FILLER_367_481 ();
 FILLCELL_X32 FILLER_367_513 ();
 FILLCELL_X32 FILLER_367_545 ();
 FILLCELL_X32 FILLER_367_577 ();
 FILLCELL_X32 FILLER_367_609 ();
 FILLCELL_X32 FILLER_367_641 ();
 FILLCELL_X32 FILLER_367_673 ();
 FILLCELL_X32 FILLER_367_705 ();
 FILLCELL_X32 FILLER_367_737 ();
 FILLCELL_X32 FILLER_367_769 ();
 FILLCELL_X32 FILLER_367_801 ();
 FILLCELL_X32 FILLER_367_833 ();
 FILLCELL_X32 FILLER_367_865 ();
 FILLCELL_X32 FILLER_367_897 ();
 FILLCELL_X32 FILLER_367_929 ();
 FILLCELL_X32 FILLER_367_961 ();
 FILLCELL_X32 FILLER_367_993 ();
 FILLCELL_X32 FILLER_367_1025 ();
 FILLCELL_X32 FILLER_367_1057 ();
 FILLCELL_X32 FILLER_367_1089 ();
 FILLCELL_X32 FILLER_367_1121 ();
 FILLCELL_X32 FILLER_367_1153 ();
 FILLCELL_X32 FILLER_367_1185 ();
 FILLCELL_X32 FILLER_367_1217 ();
 FILLCELL_X8 FILLER_367_1249 ();
 FILLCELL_X4 FILLER_367_1257 ();
 FILLCELL_X2 FILLER_367_1261 ();
 FILLCELL_X32 FILLER_367_1264 ();
 FILLCELL_X32 FILLER_367_1296 ();
 FILLCELL_X32 FILLER_367_1328 ();
 FILLCELL_X32 FILLER_367_1360 ();
 FILLCELL_X32 FILLER_367_1392 ();
 FILLCELL_X32 FILLER_367_1424 ();
 FILLCELL_X32 FILLER_367_1456 ();
 FILLCELL_X32 FILLER_367_1488 ();
 FILLCELL_X32 FILLER_367_1520 ();
 FILLCELL_X32 FILLER_367_1552 ();
 FILLCELL_X32 FILLER_367_1584 ();
 FILLCELL_X32 FILLER_367_1616 ();
 FILLCELL_X32 FILLER_367_1648 ();
 FILLCELL_X32 FILLER_367_1680 ();
 FILLCELL_X32 FILLER_367_1712 ();
 FILLCELL_X32 FILLER_367_1744 ();
 FILLCELL_X32 FILLER_367_1776 ();
 FILLCELL_X32 FILLER_367_1808 ();
 FILLCELL_X32 FILLER_367_1840 ();
 FILLCELL_X32 FILLER_367_1872 ();
 FILLCELL_X32 FILLER_367_1904 ();
 FILLCELL_X32 FILLER_367_1936 ();
 FILLCELL_X32 FILLER_367_1968 ();
 FILLCELL_X32 FILLER_367_2000 ();
 FILLCELL_X32 FILLER_367_2032 ();
 FILLCELL_X32 FILLER_367_2064 ();
 FILLCELL_X32 FILLER_367_2096 ();
 FILLCELL_X32 FILLER_367_2128 ();
 FILLCELL_X32 FILLER_367_2160 ();
 FILLCELL_X32 FILLER_367_2192 ();
 FILLCELL_X32 FILLER_367_2224 ();
 FILLCELL_X32 FILLER_367_2256 ();
 FILLCELL_X32 FILLER_367_2288 ();
 FILLCELL_X32 FILLER_367_2320 ();
 FILLCELL_X32 FILLER_367_2352 ();
 FILLCELL_X32 FILLER_367_2384 ();
 FILLCELL_X32 FILLER_367_2416 ();
 FILLCELL_X32 FILLER_367_2448 ();
 FILLCELL_X32 FILLER_367_2480 ();
 FILLCELL_X8 FILLER_367_2512 ();
 FILLCELL_X4 FILLER_367_2520 ();
 FILLCELL_X2 FILLER_367_2524 ();
 FILLCELL_X32 FILLER_367_2527 ();
 FILLCELL_X32 FILLER_367_2559 ();
 FILLCELL_X32 FILLER_367_2591 ();
 FILLCELL_X32 FILLER_367_2623 ();
 FILLCELL_X32 FILLER_367_2655 ();
 FILLCELL_X32 FILLER_367_2687 ();
 FILLCELL_X32 FILLER_367_2719 ();
 FILLCELL_X32 FILLER_367_2751 ();
 FILLCELL_X32 FILLER_367_2783 ();
 FILLCELL_X32 FILLER_367_2815 ();
 FILLCELL_X32 FILLER_367_2847 ();
 FILLCELL_X32 FILLER_367_2879 ();
 FILLCELL_X32 FILLER_367_2911 ();
 FILLCELL_X32 FILLER_367_2943 ();
 FILLCELL_X32 FILLER_367_2975 ();
 FILLCELL_X32 FILLER_367_3007 ();
 FILLCELL_X32 FILLER_367_3039 ();
 FILLCELL_X32 FILLER_367_3071 ();
 FILLCELL_X32 FILLER_367_3103 ();
 FILLCELL_X32 FILLER_367_3135 ();
 FILLCELL_X32 FILLER_367_3167 ();
 FILLCELL_X32 FILLER_367_3199 ();
 FILLCELL_X32 FILLER_367_3231 ();
 FILLCELL_X32 FILLER_367_3263 ();
 FILLCELL_X32 FILLER_367_3295 ();
 FILLCELL_X32 FILLER_367_3327 ();
 FILLCELL_X32 FILLER_367_3359 ();
 FILLCELL_X32 FILLER_367_3391 ();
 FILLCELL_X32 FILLER_367_3423 ();
 FILLCELL_X32 FILLER_367_3455 ();
 FILLCELL_X32 FILLER_367_3487 ();
 FILLCELL_X32 FILLER_367_3519 ();
 FILLCELL_X32 FILLER_367_3551 ();
 FILLCELL_X32 FILLER_367_3583 ();
 FILLCELL_X32 FILLER_367_3615 ();
 FILLCELL_X32 FILLER_367_3647 ();
 FILLCELL_X32 FILLER_367_3679 ();
 FILLCELL_X16 FILLER_367_3711 ();
 FILLCELL_X8 FILLER_367_3727 ();
 FILLCELL_X2 FILLER_367_3735 ();
 FILLCELL_X1 FILLER_367_3737 ();
 FILLCELL_X32 FILLER_368_1 ();
 FILLCELL_X32 FILLER_368_33 ();
 FILLCELL_X32 FILLER_368_65 ();
 FILLCELL_X32 FILLER_368_97 ();
 FILLCELL_X32 FILLER_368_129 ();
 FILLCELL_X32 FILLER_368_161 ();
 FILLCELL_X32 FILLER_368_193 ();
 FILLCELL_X32 FILLER_368_225 ();
 FILLCELL_X32 FILLER_368_257 ();
 FILLCELL_X32 FILLER_368_289 ();
 FILLCELL_X32 FILLER_368_321 ();
 FILLCELL_X32 FILLER_368_353 ();
 FILLCELL_X32 FILLER_368_385 ();
 FILLCELL_X32 FILLER_368_417 ();
 FILLCELL_X32 FILLER_368_449 ();
 FILLCELL_X32 FILLER_368_481 ();
 FILLCELL_X32 FILLER_368_513 ();
 FILLCELL_X32 FILLER_368_545 ();
 FILLCELL_X32 FILLER_368_577 ();
 FILLCELL_X16 FILLER_368_609 ();
 FILLCELL_X4 FILLER_368_625 ();
 FILLCELL_X2 FILLER_368_629 ();
 FILLCELL_X32 FILLER_368_632 ();
 FILLCELL_X32 FILLER_368_664 ();
 FILLCELL_X32 FILLER_368_696 ();
 FILLCELL_X32 FILLER_368_728 ();
 FILLCELL_X32 FILLER_368_760 ();
 FILLCELL_X32 FILLER_368_792 ();
 FILLCELL_X32 FILLER_368_824 ();
 FILLCELL_X32 FILLER_368_856 ();
 FILLCELL_X32 FILLER_368_888 ();
 FILLCELL_X32 FILLER_368_920 ();
 FILLCELL_X32 FILLER_368_952 ();
 FILLCELL_X32 FILLER_368_984 ();
 FILLCELL_X32 FILLER_368_1016 ();
 FILLCELL_X32 FILLER_368_1048 ();
 FILLCELL_X32 FILLER_368_1080 ();
 FILLCELL_X32 FILLER_368_1112 ();
 FILLCELL_X32 FILLER_368_1144 ();
 FILLCELL_X32 FILLER_368_1176 ();
 FILLCELL_X32 FILLER_368_1208 ();
 FILLCELL_X32 FILLER_368_1240 ();
 FILLCELL_X32 FILLER_368_1272 ();
 FILLCELL_X32 FILLER_368_1304 ();
 FILLCELL_X32 FILLER_368_1336 ();
 FILLCELL_X32 FILLER_368_1368 ();
 FILLCELL_X32 FILLER_368_1400 ();
 FILLCELL_X32 FILLER_368_1432 ();
 FILLCELL_X32 FILLER_368_1464 ();
 FILLCELL_X32 FILLER_368_1496 ();
 FILLCELL_X32 FILLER_368_1528 ();
 FILLCELL_X32 FILLER_368_1560 ();
 FILLCELL_X32 FILLER_368_1592 ();
 FILLCELL_X32 FILLER_368_1624 ();
 FILLCELL_X32 FILLER_368_1656 ();
 FILLCELL_X32 FILLER_368_1688 ();
 FILLCELL_X32 FILLER_368_1720 ();
 FILLCELL_X32 FILLER_368_1752 ();
 FILLCELL_X32 FILLER_368_1784 ();
 FILLCELL_X32 FILLER_368_1816 ();
 FILLCELL_X32 FILLER_368_1848 ();
 FILLCELL_X8 FILLER_368_1880 ();
 FILLCELL_X4 FILLER_368_1888 ();
 FILLCELL_X2 FILLER_368_1892 ();
 FILLCELL_X32 FILLER_368_1895 ();
 FILLCELL_X32 FILLER_368_1927 ();
 FILLCELL_X32 FILLER_368_1959 ();
 FILLCELL_X32 FILLER_368_1991 ();
 FILLCELL_X32 FILLER_368_2023 ();
 FILLCELL_X32 FILLER_368_2055 ();
 FILLCELL_X32 FILLER_368_2087 ();
 FILLCELL_X32 FILLER_368_2119 ();
 FILLCELL_X32 FILLER_368_2151 ();
 FILLCELL_X32 FILLER_368_2183 ();
 FILLCELL_X32 FILLER_368_2215 ();
 FILLCELL_X32 FILLER_368_2247 ();
 FILLCELL_X32 FILLER_368_2279 ();
 FILLCELL_X32 FILLER_368_2311 ();
 FILLCELL_X32 FILLER_368_2343 ();
 FILLCELL_X32 FILLER_368_2375 ();
 FILLCELL_X32 FILLER_368_2407 ();
 FILLCELL_X32 FILLER_368_2439 ();
 FILLCELL_X32 FILLER_368_2471 ();
 FILLCELL_X32 FILLER_368_2503 ();
 FILLCELL_X32 FILLER_368_2535 ();
 FILLCELL_X32 FILLER_368_2567 ();
 FILLCELL_X32 FILLER_368_2599 ();
 FILLCELL_X32 FILLER_368_2631 ();
 FILLCELL_X32 FILLER_368_2663 ();
 FILLCELL_X32 FILLER_368_2695 ();
 FILLCELL_X32 FILLER_368_2727 ();
 FILLCELL_X32 FILLER_368_2759 ();
 FILLCELL_X32 FILLER_368_2791 ();
 FILLCELL_X32 FILLER_368_2823 ();
 FILLCELL_X32 FILLER_368_2855 ();
 FILLCELL_X32 FILLER_368_2887 ();
 FILLCELL_X32 FILLER_368_2919 ();
 FILLCELL_X32 FILLER_368_2951 ();
 FILLCELL_X32 FILLER_368_2983 ();
 FILLCELL_X32 FILLER_368_3015 ();
 FILLCELL_X32 FILLER_368_3047 ();
 FILLCELL_X32 FILLER_368_3079 ();
 FILLCELL_X32 FILLER_368_3111 ();
 FILLCELL_X8 FILLER_368_3143 ();
 FILLCELL_X4 FILLER_368_3151 ();
 FILLCELL_X2 FILLER_368_3155 ();
 FILLCELL_X32 FILLER_368_3158 ();
 FILLCELL_X32 FILLER_368_3190 ();
 FILLCELL_X32 FILLER_368_3222 ();
 FILLCELL_X32 FILLER_368_3254 ();
 FILLCELL_X32 FILLER_368_3286 ();
 FILLCELL_X32 FILLER_368_3318 ();
 FILLCELL_X32 FILLER_368_3350 ();
 FILLCELL_X32 FILLER_368_3382 ();
 FILLCELL_X32 FILLER_368_3414 ();
 FILLCELL_X32 FILLER_368_3446 ();
 FILLCELL_X32 FILLER_368_3478 ();
 FILLCELL_X32 FILLER_368_3510 ();
 FILLCELL_X32 FILLER_368_3542 ();
 FILLCELL_X32 FILLER_368_3574 ();
 FILLCELL_X32 FILLER_368_3606 ();
 FILLCELL_X32 FILLER_368_3638 ();
 FILLCELL_X32 FILLER_368_3670 ();
 FILLCELL_X32 FILLER_368_3702 ();
 FILLCELL_X4 FILLER_368_3734 ();
 FILLCELL_X32 FILLER_369_1 ();
 FILLCELL_X32 FILLER_369_33 ();
 FILLCELL_X32 FILLER_369_65 ();
 FILLCELL_X32 FILLER_369_97 ();
 FILLCELL_X32 FILLER_369_129 ();
 FILLCELL_X32 FILLER_369_161 ();
 FILLCELL_X32 FILLER_369_193 ();
 FILLCELL_X32 FILLER_369_225 ();
 FILLCELL_X32 FILLER_369_257 ();
 FILLCELL_X32 FILLER_369_289 ();
 FILLCELL_X32 FILLER_369_321 ();
 FILLCELL_X32 FILLER_369_353 ();
 FILLCELL_X32 FILLER_369_385 ();
 FILLCELL_X32 FILLER_369_417 ();
 FILLCELL_X32 FILLER_369_449 ();
 FILLCELL_X32 FILLER_369_481 ();
 FILLCELL_X32 FILLER_369_513 ();
 FILLCELL_X32 FILLER_369_545 ();
 FILLCELL_X32 FILLER_369_577 ();
 FILLCELL_X32 FILLER_369_609 ();
 FILLCELL_X32 FILLER_369_641 ();
 FILLCELL_X32 FILLER_369_673 ();
 FILLCELL_X32 FILLER_369_705 ();
 FILLCELL_X32 FILLER_369_737 ();
 FILLCELL_X32 FILLER_369_769 ();
 FILLCELL_X32 FILLER_369_801 ();
 FILLCELL_X32 FILLER_369_833 ();
 FILLCELL_X32 FILLER_369_865 ();
 FILLCELL_X32 FILLER_369_897 ();
 FILLCELL_X32 FILLER_369_929 ();
 FILLCELL_X32 FILLER_369_961 ();
 FILLCELL_X32 FILLER_369_993 ();
 FILLCELL_X32 FILLER_369_1025 ();
 FILLCELL_X32 FILLER_369_1057 ();
 FILLCELL_X32 FILLER_369_1089 ();
 FILLCELL_X32 FILLER_369_1121 ();
 FILLCELL_X32 FILLER_369_1153 ();
 FILLCELL_X32 FILLER_369_1185 ();
 FILLCELL_X32 FILLER_369_1217 ();
 FILLCELL_X8 FILLER_369_1249 ();
 FILLCELL_X4 FILLER_369_1257 ();
 FILLCELL_X2 FILLER_369_1261 ();
 FILLCELL_X32 FILLER_369_1264 ();
 FILLCELL_X32 FILLER_369_1296 ();
 FILLCELL_X32 FILLER_369_1328 ();
 FILLCELL_X32 FILLER_369_1360 ();
 FILLCELL_X32 FILLER_369_1392 ();
 FILLCELL_X32 FILLER_369_1424 ();
 FILLCELL_X32 FILLER_369_1456 ();
 FILLCELL_X32 FILLER_369_1488 ();
 FILLCELL_X32 FILLER_369_1520 ();
 FILLCELL_X32 FILLER_369_1552 ();
 FILLCELL_X32 FILLER_369_1584 ();
 FILLCELL_X32 FILLER_369_1616 ();
 FILLCELL_X32 FILLER_369_1648 ();
 FILLCELL_X32 FILLER_369_1680 ();
 FILLCELL_X32 FILLER_369_1712 ();
 FILLCELL_X32 FILLER_369_1744 ();
 FILLCELL_X32 FILLER_369_1776 ();
 FILLCELL_X32 FILLER_369_1808 ();
 FILLCELL_X32 FILLER_369_1840 ();
 FILLCELL_X32 FILLER_369_1872 ();
 FILLCELL_X32 FILLER_369_1904 ();
 FILLCELL_X32 FILLER_369_1936 ();
 FILLCELL_X32 FILLER_369_1968 ();
 FILLCELL_X32 FILLER_369_2000 ();
 FILLCELL_X32 FILLER_369_2032 ();
 FILLCELL_X32 FILLER_369_2064 ();
 FILLCELL_X32 FILLER_369_2096 ();
 FILLCELL_X32 FILLER_369_2128 ();
 FILLCELL_X32 FILLER_369_2160 ();
 FILLCELL_X32 FILLER_369_2192 ();
 FILLCELL_X32 FILLER_369_2224 ();
 FILLCELL_X32 FILLER_369_2256 ();
 FILLCELL_X32 FILLER_369_2288 ();
 FILLCELL_X32 FILLER_369_2320 ();
 FILLCELL_X32 FILLER_369_2352 ();
 FILLCELL_X32 FILLER_369_2384 ();
 FILLCELL_X32 FILLER_369_2416 ();
 FILLCELL_X32 FILLER_369_2448 ();
 FILLCELL_X32 FILLER_369_2480 ();
 FILLCELL_X8 FILLER_369_2512 ();
 FILLCELL_X4 FILLER_369_2520 ();
 FILLCELL_X2 FILLER_369_2524 ();
 FILLCELL_X32 FILLER_369_2527 ();
 FILLCELL_X32 FILLER_369_2559 ();
 FILLCELL_X32 FILLER_369_2591 ();
 FILLCELL_X32 FILLER_369_2623 ();
 FILLCELL_X32 FILLER_369_2655 ();
 FILLCELL_X32 FILLER_369_2687 ();
 FILLCELL_X32 FILLER_369_2719 ();
 FILLCELL_X32 FILLER_369_2751 ();
 FILLCELL_X32 FILLER_369_2783 ();
 FILLCELL_X32 FILLER_369_2815 ();
 FILLCELL_X32 FILLER_369_2847 ();
 FILLCELL_X32 FILLER_369_2879 ();
 FILLCELL_X32 FILLER_369_2911 ();
 FILLCELL_X32 FILLER_369_2943 ();
 FILLCELL_X32 FILLER_369_2975 ();
 FILLCELL_X32 FILLER_369_3007 ();
 FILLCELL_X32 FILLER_369_3039 ();
 FILLCELL_X32 FILLER_369_3071 ();
 FILLCELL_X32 FILLER_369_3103 ();
 FILLCELL_X32 FILLER_369_3135 ();
 FILLCELL_X32 FILLER_369_3167 ();
 FILLCELL_X32 FILLER_369_3199 ();
 FILLCELL_X32 FILLER_369_3231 ();
 FILLCELL_X32 FILLER_369_3263 ();
 FILLCELL_X32 FILLER_369_3295 ();
 FILLCELL_X32 FILLER_369_3327 ();
 FILLCELL_X32 FILLER_369_3359 ();
 FILLCELL_X32 FILLER_369_3391 ();
 FILLCELL_X32 FILLER_369_3423 ();
 FILLCELL_X32 FILLER_369_3455 ();
 FILLCELL_X32 FILLER_369_3487 ();
 FILLCELL_X32 FILLER_369_3519 ();
 FILLCELL_X32 FILLER_369_3551 ();
 FILLCELL_X32 FILLER_369_3583 ();
 FILLCELL_X32 FILLER_369_3615 ();
 FILLCELL_X32 FILLER_369_3647 ();
 FILLCELL_X32 FILLER_369_3679 ();
 FILLCELL_X16 FILLER_369_3711 ();
 FILLCELL_X8 FILLER_369_3727 ();
 FILLCELL_X2 FILLER_369_3735 ();
 FILLCELL_X1 FILLER_369_3737 ();
 FILLCELL_X32 FILLER_370_1 ();
 FILLCELL_X32 FILLER_370_33 ();
 FILLCELL_X32 FILLER_370_65 ();
 FILLCELL_X32 FILLER_370_97 ();
 FILLCELL_X32 FILLER_370_129 ();
 FILLCELL_X32 FILLER_370_161 ();
 FILLCELL_X32 FILLER_370_193 ();
 FILLCELL_X32 FILLER_370_225 ();
 FILLCELL_X32 FILLER_370_257 ();
 FILLCELL_X32 FILLER_370_289 ();
 FILLCELL_X32 FILLER_370_321 ();
 FILLCELL_X32 FILLER_370_353 ();
 FILLCELL_X32 FILLER_370_385 ();
 FILLCELL_X32 FILLER_370_417 ();
 FILLCELL_X32 FILLER_370_449 ();
 FILLCELL_X32 FILLER_370_481 ();
 FILLCELL_X32 FILLER_370_513 ();
 FILLCELL_X32 FILLER_370_545 ();
 FILLCELL_X32 FILLER_370_577 ();
 FILLCELL_X16 FILLER_370_609 ();
 FILLCELL_X4 FILLER_370_625 ();
 FILLCELL_X2 FILLER_370_629 ();
 FILLCELL_X32 FILLER_370_632 ();
 FILLCELL_X32 FILLER_370_664 ();
 FILLCELL_X32 FILLER_370_696 ();
 FILLCELL_X32 FILLER_370_728 ();
 FILLCELL_X32 FILLER_370_760 ();
 FILLCELL_X32 FILLER_370_792 ();
 FILLCELL_X32 FILLER_370_824 ();
 FILLCELL_X32 FILLER_370_856 ();
 FILLCELL_X32 FILLER_370_888 ();
 FILLCELL_X32 FILLER_370_920 ();
 FILLCELL_X32 FILLER_370_952 ();
 FILLCELL_X32 FILLER_370_984 ();
 FILLCELL_X32 FILLER_370_1016 ();
 FILLCELL_X32 FILLER_370_1048 ();
 FILLCELL_X32 FILLER_370_1080 ();
 FILLCELL_X32 FILLER_370_1112 ();
 FILLCELL_X32 FILLER_370_1144 ();
 FILLCELL_X32 FILLER_370_1176 ();
 FILLCELL_X32 FILLER_370_1208 ();
 FILLCELL_X32 FILLER_370_1240 ();
 FILLCELL_X32 FILLER_370_1272 ();
 FILLCELL_X32 FILLER_370_1304 ();
 FILLCELL_X32 FILLER_370_1336 ();
 FILLCELL_X32 FILLER_370_1368 ();
 FILLCELL_X32 FILLER_370_1400 ();
 FILLCELL_X32 FILLER_370_1432 ();
 FILLCELL_X32 FILLER_370_1464 ();
 FILLCELL_X32 FILLER_370_1496 ();
 FILLCELL_X32 FILLER_370_1528 ();
 FILLCELL_X32 FILLER_370_1560 ();
 FILLCELL_X32 FILLER_370_1592 ();
 FILLCELL_X32 FILLER_370_1624 ();
 FILLCELL_X32 FILLER_370_1656 ();
 FILLCELL_X32 FILLER_370_1688 ();
 FILLCELL_X32 FILLER_370_1720 ();
 FILLCELL_X32 FILLER_370_1752 ();
 FILLCELL_X32 FILLER_370_1784 ();
 FILLCELL_X32 FILLER_370_1816 ();
 FILLCELL_X32 FILLER_370_1848 ();
 FILLCELL_X8 FILLER_370_1880 ();
 FILLCELL_X4 FILLER_370_1888 ();
 FILLCELL_X2 FILLER_370_1892 ();
 FILLCELL_X32 FILLER_370_1895 ();
 FILLCELL_X32 FILLER_370_1927 ();
 FILLCELL_X32 FILLER_370_1959 ();
 FILLCELL_X32 FILLER_370_1991 ();
 FILLCELL_X32 FILLER_370_2023 ();
 FILLCELL_X32 FILLER_370_2055 ();
 FILLCELL_X32 FILLER_370_2087 ();
 FILLCELL_X32 FILLER_370_2119 ();
 FILLCELL_X32 FILLER_370_2151 ();
 FILLCELL_X32 FILLER_370_2183 ();
 FILLCELL_X32 FILLER_370_2215 ();
 FILLCELL_X32 FILLER_370_2247 ();
 FILLCELL_X32 FILLER_370_2279 ();
 FILLCELL_X32 FILLER_370_2311 ();
 FILLCELL_X32 FILLER_370_2343 ();
 FILLCELL_X32 FILLER_370_2375 ();
 FILLCELL_X32 FILLER_370_2407 ();
 FILLCELL_X32 FILLER_370_2439 ();
 FILLCELL_X32 FILLER_370_2471 ();
 FILLCELL_X32 FILLER_370_2503 ();
 FILLCELL_X32 FILLER_370_2535 ();
 FILLCELL_X32 FILLER_370_2567 ();
 FILLCELL_X32 FILLER_370_2599 ();
 FILLCELL_X32 FILLER_370_2631 ();
 FILLCELL_X32 FILLER_370_2663 ();
 FILLCELL_X32 FILLER_370_2695 ();
 FILLCELL_X32 FILLER_370_2727 ();
 FILLCELL_X32 FILLER_370_2759 ();
 FILLCELL_X32 FILLER_370_2791 ();
 FILLCELL_X32 FILLER_370_2823 ();
 FILLCELL_X32 FILLER_370_2855 ();
 FILLCELL_X32 FILLER_370_2887 ();
 FILLCELL_X32 FILLER_370_2919 ();
 FILLCELL_X32 FILLER_370_2951 ();
 FILLCELL_X32 FILLER_370_2983 ();
 FILLCELL_X32 FILLER_370_3015 ();
 FILLCELL_X32 FILLER_370_3047 ();
 FILLCELL_X32 FILLER_370_3079 ();
 FILLCELL_X32 FILLER_370_3111 ();
 FILLCELL_X8 FILLER_370_3143 ();
 FILLCELL_X4 FILLER_370_3151 ();
 FILLCELL_X2 FILLER_370_3155 ();
 FILLCELL_X32 FILLER_370_3158 ();
 FILLCELL_X32 FILLER_370_3190 ();
 FILLCELL_X32 FILLER_370_3222 ();
 FILLCELL_X32 FILLER_370_3254 ();
 FILLCELL_X32 FILLER_370_3286 ();
 FILLCELL_X32 FILLER_370_3318 ();
 FILLCELL_X32 FILLER_370_3350 ();
 FILLCELL_X32 FILLER_370_3382 ();
 FILLCELL_X32 FILLER_370_3414 ();
 FILLCELL_X32 FILLER_370_3446 ();
 FILLCELL_X32 FILLER_370_3478 ();
 FILLCELL_X32 FILLER_370_3510 ();
 FILLCELL_X32 FILLER_370_3542 ();
 FILLCELL_X32 FILLER_370_3574 ();
 FILLCELL_X32 FILLER_370_3606 ();
 FILLCELL_X32 FILLER_370_3638 ();
 FILLCELL_X32 FILLER_370_3670 ();
 FILLCELL_X32 FILLER_370_3702 ();
 FILLCELL_X4 FILLER_370_3734 ();
 FILLCELL_X32 FILLER_371_1 ();
 FILLCELL_X32 FILLER_371_33 ();
 FILLCELL_X32 FILLER_371_65 ();
 FILLCELL_X32 FILLER_371_97 ();
 FILLCELL_X32 FILLER_371_129 ();
 FILLCELL_X32 FILLER_371_161 ();
 FILLCELL_X32 FILLER_371_193 ();
 FILLCELL_X32 FILLER_371_225 ();
 FILLCELL_X32 FILLER_371_257 ();
 FILLCELL_X32 FILLER_371_289 ();
 FILLCELL_X32 FILLER_371_321 ();
 FILLCELL_X32 FILLER_371_353 ();
 FILLCELL_X32 FILLER_371_385 ();
 FILLCELL_X32 FILLER_371_417 ();
 FILLCELL_X32 FILLER_371_449 ();
 FILLCELL_X32 FILLER_371_481 ();
 FILLCELL_X32 FILLER_371_513 ();
 FILLCELL_X32 FILLER_371_545 ();
 FILLCELL_X32 FILLER_371_577 ();
 FILLCELL_X32 FILLER_371_609 ();
 FILLCELL_X32 FILLER_371_641 ();
 FILLCELL_X32 FILLER_371_673 ();
 FILLCELL_X32 FILLER_371_705 ();
 FILLCELL_X32 FILLER_371_737 ();
 FILLCELL_X32 FILLER_371_769 ();
 FILLCELL_X32 FILLER_371_801 ();
 FILLCELL_X32 FILLER_371_833 ();
 FILLCELL_X32 FILLER_371_865 ();
 FILLCELL_X32 FILLER_371_897 ();
 FILLCELL_X32 FILLER_371_929 ();
 FILLCELL_X32 FILLER_371_961 ();
 FILLCELL_X32 FILLER_371_993 ();
 FILLCELL_X32 FILLER_371_1025 ();
 FILLCELL_X32 FILLER_371_1057 ();
 FILLCELL_X32 FILLER_371_1089 ();
 FILLCELL_X32 FILLER_371_1121 ();
 FILLCELL_X32 FILLER_371_1153 ();
 FILLCELL_X32 FILLER_371_1185 ();
 FILLCELL_X32 FILLER_371_1217 ();
 FILLCELL_X8 FILLER_371_1249 ();
 FILLCELL_X4 FILLER_371_1257 ();
 FILLCELL_X2 FILLER_371_1261 ();
 FILLCELL_X32 FILLER_371_1264 ();
 FILLCELL_X32 FILLER_371_1296 ();
 FILLCELL_X32 FILLER_371_1328 ();
 FILLCELL_X32 FILLER_371_1360 ();
 FILLCELL_X32 FILLER_371_1392 ();
 FILLCELL_X32 FILLER_371_1424 ();
 FILLCELL_X32 FILLER_371_1456 ();
 FILLCELL_X32 FILLER_371_1488 ();
 FILLCELL_X32 FILLER_371_1520 ();
 FILLCELL_X32 FILLER_371_1552 ();
 FILLCELL_X32 FILLER_371_1584 ();
 FILLCELL_X32 FILLER_371_1616 ();
 FILLCELL_X32 FILLER_371_1648 ();
 FILLCELL_X32 FILLER_371_1680 ();
 FILLCELL_X32 FILLER_371_1712 ();
 FILLCELL_X32 FILLER_371_1744 ();
 FILLCELL_X32 FILLER_371_1776 ();
 FILLCELL_X32 FILLER_371_1808 ();
 FILLCELL_X32 FILLER_371_1840 ();
 FILLCELL_X32 FILLER_371_1872 ();
 FILLCELL_X32 FILLER_371_1904 ();
 FILLCELL_X32 FILLER_371_1936 ();
 FILLCELL_X32 FILLER_371_1968 ();
 FILLCELL_X32 FILLER_371_2000 ();
 FILLCELL_X32 FILLER_371_2032 ();
 FILLCELL_X32 FILLER_371_2064 ();
 FILLCELL_X32 FILLER_371_2096 ();
 FILLCELL_X32 FILLER_371_2128 ();
 FILLCELL_X32 FILLER_371_2160 ();
 FILLCELL_X32 FILLER_371_2192 ();
 FILLCELL_X32 FILLER_371_2224 ();
 FILLCELL_X32 FILLER_371_2256 ();
 FILLCELL_X32 FILLER_371_2288 ();
 FILLCELL_X32 FILLER_371_2320 ();
 FILLCELL_X32 FILLER_371_2352 ();
 FILLCELL_X32 FILLER_371_2384 ();
 FILLCELL_X32 FILLER_371_2416 ();
 FILLCELL_X32 FILLER_371_2448 ();
 FILLCELL_X32 FILLER_371_2480 ();
 FILLCELL_X8 FILLER_371_2512 ();
 FILLCELL_X4 FILLER_371_2520 ();
 FILLCELL_X2 FILLER_371_2524 ();
 FILLCELL_X32 FILLER_371_2527 ();
 FILLCELL_X32 FILLER_371_2559 ();
 FILLCELL_X32 FILLER_371_2591 ();
 FILLCELL_X32 FILLER_371_2623 ();
 FILLCELL_X32 FILLER_371_2655 ();
 FILLCELL_X32 FILLER_371_2687 ();
 FILLCELL_X32 FILLER_371_2719 ();
 FILLCELL_X32 FILLER_371_2751 ();
 FILLCELL_X32 FILLER_371_2783 ();
 FILLCELL_X32 FILLER_371_2815 ();
 FILLCELL_X32 FILLER_371_2847 ();
 FILLCELL_X32 FILLER_371_2879 ();
 FILLCELL_X32 FILLER_371_2911 ();
 FILLCELL_X32 FILLER_371_2943 ();
 FILLCELL_X32 FILLER_371_2975 ();
 FILLCELL_X32 FILLER_371_3007 ();
 FILLCELL_X32 FILLER_371_3039 ();
 FILLCELL_X32 FILLER_371_3071 ();
 FILLCELL_X32 FILLER_371_3103 ();
 FILLCELL_X32 FILLER_371_3135 ();
 FILLCELL_X32 FILLER_371_3167 ();
 FILLCELL_X32 FILLER_371_3199 ();
 FILLCELL_X32 FILLER_371_3231 ();
 FILLCELL_X32 FILLER_371_3263 ();
 FILLCELL_X32 FILLER_371_3295 ();
 FILLCELL_X32 FILLER_371_3327 ();
 FILLCELL_X32 FILLER_371_3359 ();
 FILLCELL_X32 FILLER_371_3391 ();
 FILLCELL_X32 FILLER_371_3423 ();
 FILLCELL_X32 FILLER_371_3455 ();
 FILLCELL_X32 FILLER_371_3487 ();
 FILLCELL_X32 FILLER_371_3519 ();
 FILLCELL_X32 FILLER_371_3551 ();
 FILLCELL_X32 FILLER_371_3583 ();
 FILLCELL_X32 FILLER_371_3615 ();
 FILLCELL_X32 FILLER_371_3647 ();
 FILLCELL_X32 FILLER_371_3679 ();
 FILLCELL_X16 FILLER_371_3711 ();
 FILLCELL_X8 FILLER_371_3727 ();
 FILLCELL_X2 FILLER_371_3735 ();
 FILLCELL_X1 FILLER_371_3737 ();
 FILLCELL_X32 FILLER_372_1 ();
 FILLCELL_X32 FILLER_372_33 ();
 FILLCELL_X32 FILLER_372_65 ();
 FILLCELL_X32 FILLER_372_97 ();
 FILLCELL_X32 FILLER_372_129 ();
 FILLCELL_X32 FILLER_372_161 ();
 FILLCELL_X32 FILLER_372_193 ();
 FILLCELL_X32 FILLER_372_225 ();
 FILLCELL_X32 FILLER_372_257 ();
 FILLCELL_X32 FILLER_372_289 ();
 FILLCELL_X32 FILLER_372_321 ();
 FILLCELL_X32 FILLER_372_353 ();
 FILLCELL_X32 FILLER_372_385 ();
 FILLCELL_X32 FILLER_372_417 ();
 FILLCELL_X32 FILLER_372_449 ();
 FILLCELL_X32 FILLER_372_481 ();
 FILLCELL_X32 FILLER_372_513 ();
 FILLCELL_X32 FILLER_372_545 ();
 FILLCELL_X32 FILLER_372_577 ();
 FILLCELL_X16 FILLER_372_609 ();
 FILLCELL_X4 FILLER_372_625 ();
 FILLCELL_X2 FILLER_372_629 ();
 FILLCELL_X32 FILLER_372_632 ();
 FILLCELL_X32 FILLER_372_664 ();
 FILLCELL_X32 FILLER_372_696 ();
 FILLCELL_X32 FILLER_372_728 ();
 FILLCELL_X32 FILLER_372_760 ();
 FILLCELL_X32 FILLER_372_792 ();
 FILLCELL_X32 FILLER_372_824 ();
 FILLCELL_X32 FILLER_372_856 ();
 FILLCELL_X32 FILLER_372_888 ();
 FILLCELL_X32 FILLER_372_920 ();
 FILLCELL_X32 FILLER_372_952 ();
 FILLCELL_X32 FILLER_372_984 ();
 FILLCELL_X32 FILLER_372_1016 ();
 FILLCELL_X32 FILLER_372_1048 ();
 FILLCELL_X32 FILLER_372_1080 ();
 FILLCELL_X32 FILLER_372_1112 ();
 FILLCELL_X32 FILLER_372_1144 ();
 FILLCELL_X32 FILLER_372_1176 ();
 FILLCELL_X32 FILLER_372_1208 ();
 FILLCELL_X32 FILLER_372_1240 ();
 FILLCELL_X32 FILLER_372_1272 ();
 FILLCELL_X32 FILLER_372_1304 ();
 FILLCELL_X32 FILLER_372_1336 ();
 FILLCELL_X32 FILLER_372_1368 ();
 FILLCELL_X32 FILLER_372_1400 ();
 FILLCELL_X32 FILLER_372_1432 ();
 FILLCELL_X32 FILLER_372_1464 ();
 FILLCELL_X32 FILLER_372_1496 ();
 FILLCELL_X32 FILLER_372_1528 ();
 FILLCELL_X32 FILLER_372_1560 ();
 FILLCELL_X32 FILLER_372_1592 ();
 FILLCELL_X32 FILLER_372_1624 ();
 FILLCELL_X32 FILLER_372_1656 ();
 FILLCELL_X32 FILLER_372_1688 ();
 FILLCELL_X32 FILLER_372_1720 ();
 FILLCELL_X32 FILLER_372_1752 ();
 FILLCELL_X32 FILLER_372_1784 ();
 FILLCELL_X32 FILLER_372_1816 ();
 FILLCELL_X32 FILLER_372_1848 ();
 FILLCELL_X8 FILLER_372_1880 ();
 FILLCELL_X4 FILLER_372_1888 ();
 FILLCELL_X2 FILLER_372_1892 ();
 FILLCELL_X32 FILLER_372_1895 ();
 FILLCELL_X32 FILLER_372_1927 ();
 FILLCELL_X32 FILLER_372_1959 ();
 FILLCELL_X32 FILLER_372_1991 ();
 FILLCELL_X32 FILLER_372_2023 ();
 FILLCELL_X32 FILLER_372_2055 ();
 FILLCELL_X32 FILLER_372_2087 ();
 FILLCELL_X32 FILLER_372_2119 ();
 FILLCELL_X32 FILLER_372_2151 ();
 FILLCELL_X32 FILLER_372_2183 ();
 FILLCELL_X32 FILLER_372_2215 ();
 FILLCELL_X32 FILLER_372_2247 ();
 FILLCELL_X32 FILLER_372_2279 ();
 FILLCELL_X32 FILLER_372_2311 ();
 FILLCELL_X32 FILLER_372_2343 ();
 FILLCELL_X32 FILLER_372_2375 ();
 FILLCELL_X32 FILLER_372_2407 ();
 FILLCELL_X32 FILLER_372_2439 ();
 FILLCELL_X32 FILLER_372_2471 ();
 FILLCELL_X32 FILLER_372_2503 ();
 FILLCELL_X32 FILLER_372_2535 ();
 FILLCELL_X32 FILLER_372_2567 ();
 FILLCELL_X32 FILLER_372_2599 ();
 FILLCELL_X32 FILLER_372_2631 ();
 FILLCELL_X32 FILLER_372_2663 ();
 FILLCELL_X32 FILLER_372_2695 ();
 FILLCELL_X32 FILLER_372_2727 ();
 FILLCELL_X32 FILLER_372_2759 ();
 FILLCELL_X32 FILLER_372_2791 ();
 FILLCELL_X32 FILLER_372_2823 ();
 FILLCELL_X32 FILLER_372_2855 ();
 FILLCELL_X32 FILLER_372_2887 ();
 FILLCELL_X32 FILLER_372_2919 ();
 FILLCELL_X32 FILLER_372_2951 ();
 FILLCELL_X32 FILLER_372_2983 ();
 FILLCELL_X32 FILLER_372_3015 ();
 FILLCELL_X32 FILLER_372_3047 ();
 FILLCELL_X32 FILLER_372_3079 ();
 FILLCELL_X32 FILLER_372_3111 ();
 FILLCELL_X8 FILLER_372_3143 ();
 FILLCELL_X4 FILLER_372_3151 ();
 FILLCELL_X2 FILLER_372_3155 ();
 FILLCELL_X32 FILLER_372_3158 ();
 FILLCELL_X32 FILLER_372_3190 ();
 FILLCELL_X32 FILLER_372_3222 ();
 FILLCELL_X32 FILLER_372_3254 ();
 FILLCELL_X32 FILLER_372_3286 ();
 FILLCELL_X32 FILLER_372_3318 ();
 FILLCELL_X32 FILLER_372_3350 ();
 FILLCELL_X32 FILLER_372_3382 ();
 FILLCELL_X32 FILLER_372_3414 ();
 FILLCELL_X32 FILLER_372_3446 ();
 FILLCELL_X32 FILLER_372_3478 ();
 FILLCELL_X32 FILLER_372_3510 ();
 FILLCELL_X32 FILLER_372_3542 ();
 FILLCELL_X32 FILLER_372_3574 ();
 FILLCELL_X32 FILLER_372_3606 ();
 FILLCELL_X32 FILLER_372_3638 ();
 FILLCELL_X32 FILLER_372_3670 ();
 FILLCELL_X32 FILLER_372_3702 ();
 FILLCELL_X4 FILLER_372_3734 ();
 FILLCELL_X32 FILLER_373_1 ();
 FILLCELL_X32 FILLER_373_33 ();
 FILLCELL_X32 FILLER_373_65 ();
 FILLCELL_X32 FILLER_373_97 ();
 FILLCELL_X32 FILLER_373_129 ();
 FILLCELL_X32 FILLER_373_161 ();
 FILLCELL_X32 FILLER_373_193 ();
 FILLCELL_X32 FILLER_373_225 ();
 FILLCELL_X32 FILLER_373_257 ();
 FILLCELL_X32 FILLER_373_289 ();
 FILLCELL_X32 FILLER_373_321 ();
 FILLCELL_X32 FILLER_373_353 ();
 FILLCELL_X32 FILLER_373_385 ();
 FILLCELL_X32 FILLER_373_417 ();
 FILLCELL_X32 FILLER_373_449 ();
 FILLCELL_X32 FILLER_373_481 ();
 FILLCELL_X32 FILLER_373_513 ();
 FILLCELL_X32 FILLER_373_545 ();
 FILLCELL_X32 FILLER_373_577 ();
 FILLCELL_X32 FILLER_373_609 ();
 FILLCELL_X32 FILLER_373_641 ();
 FILLCELL_X32 FILLER_373_673 ();
 FILLCELL_X32 FILLER_373_705 ();
 FILLCELL_X32 FILLER_373_737 ();
 FILLCELL_X32 FILLER_373_769 ();
 FILLCELL_X32 FILLER_373_801 ();
 FILLCELL_X32 FILLER_373_833 ();
 FILLCELL_X32 FILLER_373_865 ();
 FILLCELL_X32 FILLER_373_897 ();
 FILLCELL_X32 FILLER_373_929 ();
 FILLCELL_X32 FILLER_373_961 ();
 FILLCELL_X32 FILLER_373_993 ();
 FILLCELL_X32 FILLER_373_1025 ();
 FILLCELL_X32 FILLER_373_1057 ();
 FILLCELL_X32 FILLER_373_1089 ();
 FILLCELL_X32 FILLER_373_1121 ();
 FILLCELL_X32 FILLER_373_1153 ();
 FILLCELL_X32 FILLER_373_1185 ();
 FILLCELL_X32 FILLER_373_1217 ();
 FILLCELL_X8 FILLER_373_1249 ();
 FILLCELL_X4 FILLER_373_1257 ();
 FILLCELL_X2 FILLER_373_1261 ();
 FILLCELL_X32 FILLER_373_1264 ();
 FILLCELL_X32 FILLER_373_1296 ();
 FILLCELL_X32 FILLER_373_1328 ();
 FILLCELL_X32 FILLER_373_1360 ();
 FILLCELL_X32 FILLER_373_1392 ();
 FILLCELL_X32 FILLER_373_1424 ();
 FILLCELL_X32 FILLER_373_1456 ();
 FILLCELL_X32 FILLER_373_1488 ();
 FILLCELL_X32 FILLER_373_1520 ();
 FILLCELL_X32 FILLER_373_1552 ();
 FILLCELL_X32 FILLER_373_1584 ();
 FILLCELL_X32 FILLER_373_1616 ();
 FILLCELL_X32 FILLER_373_1648 ();
 FILLCELL_X32 FILLER_373_1680 ();
 FILLCELL_X32 FILLER_373_1712 ();
 FILLCELL_X32 FILLER_373_1744 ();
 FILLCELL_X32 FILLER_373_1776 ();
 FILLCELL_X32 FILLER_373_1808 ();
 FILLCELL_X32 FILLER_373_1840 ();
 FILLCELL_X32 FILLER_373_1872 ();
 FILLCELL_X32 FILLER_373_1904 ();
 FILLCELL_X32 FILLER_373_1936 ();
 FILLCELL_X32 FILLER_373_1968 ();
 FILLCELL_X32 FILLER_373_2000 ();
 FILLCELL_X32 FILLER_373_2032 ();
 FILLCELL_X32 FILLER_373_2064 ();
 FILLCELL_X32 FILLER_373_2096 ();
 FILLCELL_X32 FILLER_373_2128 ();
 FILLCELL_X32 FILLER_373_2160 ();
 FILLCELL_X32 FILLER_373_2192 ();
 FILLCELL_X32 FILLER_373_2224 ();
 FILLCELL_X32 FILLER_373_2256 ();
 FILLCELL_X32 FILLER_373_2288 ();
 FILLCELL_X32 FILLER_373_2320 ();
 FILLCELL_X32 FILLER_373_2352 ();
 FILLCELL_X32 FILLER_373_2384 ();
 FILLCELL_X32 FILLER_373_2416 ();
 FILLCELL_X32 FILLER_373_2448 ();
 FILLCELL_X32 FILLER_373_2480 ();
 FILLCELL_X8 FILLER_373_2512 ();
 FILLCELL_X4 FILLER_373_2520 ();
 FILLCELL_X2 FILLER_373_2524 ();
 FILLCELL_X32 FILLER_373_2527 ();
 FILLCELL_X32 FILLER_373_2559 ();
 FILLCELL_X32 FILLER_373_2591 ();
 FILLCELL_X32 FILLER_373_2623 ();
 FILLCELL_X32 FILLER_373_2655 ();
 FILLCELL_X32 FILLER_373_2687 ();
 FILLCELL_X32 FILLER_373_2719 ();
 FILLCELL_X32 FILLER_373_2751 ();
 FILLCELL_X32 FILLER_373_2783 ();
 FILLCELL_X32 FILLER_373_2815 ();
 FILLCELL_X32 FILLER_373_2847 ();
 FILLCELL_X32 FILLER_373_2879 ();
 FILLCELL_X32 FILLER_373_2911 ();
 FILLCELL_X32 FILLER_373_2943 ();
 FILLCELL_X32 FILLER_373_2975 ();
 FILLCELL_X32 FILLER_373_3007 ();
 FILLCELL_X32 FILLER_373_3039 ();
 FILLCELL_X32 FILLER_373_3071 ();
 FILLCELL_X32 FILLER_373_3103 ();
 FILLCELL_X32 FILLER_373_3135 ();
 FILLCELL_X32 FILLER_373_3167 ();
 FILLCELL_X32 FILLER_373_3199 ();
 FILLCELL_X32 FILLER_373_3231 ();
 FILLCELL_X32 FILLER_373_3263 ();
 FILLCELL_X32 FILLER_373_3295 ();
 FILLCELL_X32 FILLER_373_3327 ();
 FILLCELL_X32 FILLER_373_3359 ();
 FILLCELL_X32 FILLER_373_3391 ();
 FILLCELL_X32 FILLER_373_3423 ();
 FILLCELL_X32 FILLER_373_3455 ();
 FILLCELL_X32 FILLER_373_3487 ();
 FILLCELL_X32 FILLER_373_3519 ();
 FILLCELL_X32 FILLER_373_3551 ();
 FILLCELL_X32 FILLER_373_3583 ();
 FILLCELL_X32 FILLER_373_3615 ();
 FILLCELL_X32 FILLER_373_3647 ();
 FILLCELL_X32 FILLER_373_3679 ();
 FILLCELL_X16 FILLER_373_3711 ();
 FILLCELL_X8 FILLER_373_3727 ();
 FILLCELL_X2 FILLER_373_3735 ();
 FILLCELL_X1 FILLER_373_3737 ();
 FILLCELL_X32 FILLER_374_1 ();
 FILLCELL_X32 FILLER_374_33 ();
 FILLCELL_X32 FILLER_374_65 ();
 FILLCELL_X32 FILLER_374_97 ();
 FILLCELL_X32 FILLER_374_129 ();
 FILLCELL_X32 FILLER_374_161 ();
 FILLCELL_X32 FILLER_374_193 ();
 FILLCELL_X32 FILLER_374_225 ();
 FILLCELL_X32 FILLER_374_257 ();
 FILLCELL_X32 FILLER_374_289 ();
 FILLCELL_X32 FILLER_374_321 ();
 FILLCELL_X32 FILLER_374_353 ();
 FILLCELL_X32 FILLER_374_385 ();
 FILLCELL_X32 FILLER_374_417 ();
 FILLCELL_X32 FILLER_374_449 ();
 FILLCELL_X32 FILLER_374_481 ();
 FILLCELL_X32 FILLER_374_513 ();
 FILLCELL_X32 FILLER_374_545 ();
 FILLCELL_X32 FILLER_374_577 ();
 FILLCELL_X16 FILLER_374_609 ();
 FILLCELL_X4 FILLER_374_625 ();
 FILLCELL_X2 FILLER_374_629 ();
 FILLCELL_X32 FILLER_374_632 ();
 FILLCELL_X32 FILLER_374_664 ();
 FILLCELL_X32 FILLER_374_696 ();
 FILLCELL_X32 FILLER_374_728 ();
 FILLCELL_X32 FILLER_374_760 ();
 FILLCELL_X32 FILLER_374_792 ();
 FILLCELL_X32 FILLER_374_824 ();
 FILLCELL_X32 FILLER_374_856 ();
 FILLCELL_X32 FILLER_374_888 ();
 FILLCELL_X32 FILLER_374_920 ();
 FILLCELL_X32 FILLER_374_952 ();
 FILLCELL_X32 FILLER_374_984 ();
 FILLCELL_X32 FILLER_374_1016 ();
 FILLCELL_X32 FILLER_374_1048 ();
 FILLCELL_X32 FILLER_374_1080 ();
 FILLCELL_X32 FILLER_374_1112 ();
 FILLCELL_X32 FILLER_374_1144 ();
 FILLCELL_X32 FILLER_374_1176 ();
 FILLCELL_X32 FILLER_374_1208 ();
 FILLCELL_X32 FILLER_374_1240 ();
 FILLCELL_X32 FILLER_374_1272 ();
 FILLCELL_X32 FILLER_374_1304 ();
 FILLCELL_X32 FILLER_374_1336 ();
 FILLCELL_X32 FILLER_374_1368 ();
 FILLCELL_X32 FILLER_374_1400 ();
 FILLCELL_X32 FILLER_374_1432 ();
 FILLCELL_X32 FILLER_374_1464 ();
 FILLCELL_X32 FILLER_374_1496 ();
 FILLCELL_X32 FILLER_374_1528 ();
 FILLCELL_X32 FILLER_374_1560 ();
 FILLCELL_X32 FILLER_374_1592 ();
 FILLCELL_X32 FILLER_374_1624 ();
 FILLCELL_X32 FILLER_374_1656 ();
 FILLCELL_X32 FILLER_374_1688 ();
 FILLCELL_X32 FILLER_374_1720 ();
 FILLCELL_X32 FILLER_374_1752 ();
 FILLCELL_X32 FILLER_374_1784 ();
 FILLCELL_X32 FILLER_374_1816 ();
 FILLCELL_X32 FILLER_374_1848 ();
 FILLCELL_X8 FILLER_374_1880 ();
 FILLCELL_X4 FILLER_374_1888 ();
 FILLCELL_X2 FILLER_374_1892 ();
 FILLCELL_X32 FILLER_374_1895 ();
 FILLCELL_X32 FILLER_374_1927 ();
 FILLCELL_X32 FILLER_374_1959 ();
 FILLCELL_X32 FILLER_374_1991 ();
 FILLCELL_X32 FILLER_374_2023 ();
 FILLCELL_X32 FILLER_374_2055 ();
 FILLCELL_X32 FILLER_374_2087 ();
 FILLCELL_X32 FILLER_374_2119 ();
 FILLCELL_X32 FILLER_374_2151 ();
 FILLCELL_X32 FILLER_374_2183 ();
 FILLCELL_X32 FILLER_374_2215 ();
 FILLCELL_X32 FILLER_374_2247 ();
 FILLCELL_X32 FILLER_374_2279 ();
 FILLCELL_X32 FILLER_374_2311 ();
 FILLCELL_X32 FILLER_374_2343 ();
 FILLCELL_X32 FILLER_374_2375 ();
 FILLCELL_X32 FILLER_374_2407 ();
 FILLCELL_X32 FILLER_374_2439 ();
 FILLCELL_X32 FILLER_374_2471 ();
 FILLCELL_X32 FILLER_374_2503 ();
 FILLCELL_X32 FILLER_374_2535 ();
 FILLCELL_X32 FILLER_374_2567 ();
 FILLCELL_X32 FILLER_374_2599 ();
 FILLCELL_X32 FILLER_374_2631 ();
 FILLCELL_X32 FILLER_374_2663 ();
 FILLCELL_X32 FILLER_374_2695 ();
 FILLCELL_X32 FILLER_374_2727 ();
 FILLCELL_X32 FILLER_374_2759 ();
 FILLCELL_X32 FILLER_374_2791 ();
 FILLCELL_X32 FILLER_374_2823 ();
 FILLCELL_X32 FILLER_374_2855 ();
 FILLCELL_X32 FILLER_374_2887 ();
 FILLCELL_X32 FILLER_374_2919 ();
 FILLCELL_X32 FILLER_374_2951 ();
 FILLCELL_X32 FILLER_374_2983 ();
 FILLCELL_X32 FILLER_374_3015 ();
 FILLCELL_X32 FILLER_374_3047 ();
 FILLCELL_X32 FILLER_374_3079 ();
 FILLCELL_X32 FILLER_374_3111 ();
 FILLCELL_X8 FILLER_374_3143 ();
 FILLCELL_X4 FILLER_374_3151 ();
 FILLCELL_X2 FILLER_374_3155 ();
 FILLCELL_X32 FILLER_374_3158 ();
 FILLCELL_X32 FILLER_374_3190 ();
 FILLCELL_X32 FILLER_374_3222 ();
 FILLCELL_X32 FILLER_374_3254 ();
 FILLCELL_X32 FILLER_374_3286 ();
 FILLCELL_X32 FILLER_374_3318 ();
 FILLCELL_X32 FILLER_374_3350 ();
 FILLCELL_X32 FILLER_374_3382 ();
 FILLCELL_X32 FILLER_374_3414 ();
 FILLCELL_X32 FILLER_374_3446 ();
 FILLCELL_X32 FILLER_374_3478 ();
 FILLCELL_X32 FILLER_374_3510 ();
 FILLCELL_X32 FILLER_374_3542 ();
 FILLCELL_X32 FILLER_374_3574 ();
 FILLCELL_X32 FILLER_374_3606 ();
 FILLCELL_X32 FILLER_374_3638 ();
 FILLCELL_X32 FILLER_374_3670 ();
 FILLCELL_X32 FILLER_374_3702 ();
 FILLCELL_X4 FILLER_374_3734 ();
 FILLCELL_X32 FILLER_375_1 ();
 FILLCELL_X32 FILLER_375_33 ();
 FILLCELL_X32 FILLER_375_65 ();
 FILLCELL_X32 FILLER_375_97 ();
 FILLCELL_X32 FILLER_375_129 ();
 FILLCELL_X32 FILLER_375_161 ();
 FILLCELL_X32 FILLER_375_193 ();
 FILLCELL_X32 FILLER_375_225 ();
 FILLCELL_X32 FILLER_375_257 ();
 FILLCELL_X32 FILLER_375_289 ();
 FILLCELL_X32 FILLER_375_321 ();
 FILLCELL_X32 FILLER_375_353 ();
 FILLCELL_X32 FILLER_375_385 ();
 FILLCELL_X32 FILLER_375_417 ();
 FILLCELL_X32 FILLER_375_449 ();
 FILLCELL_X32 FILLER_375_481 ();
 FILLCELL_X32 FILLER_375_513 ();
 FILLCELL_X32 FILLER_375_545 ();
 FILLCELL_X32 FILLER_375_577 ();
 FILLCELL_X32 FILLER_375_609 ();
 FILLCELL_X32 FILLER_375_641 ();
 FILLCELL_X32 FILLER_375_673 ();
 FILLCELL_X32 FILLER_375_705 ();
 FILLCELL_X32 FILLER_375_737 ();
 FILLCELL_X32 FILLER_375_769 ();
 FILLCELL_X32 FILLER_375_801 ();
 FILLCELL_X32 FILLER_375_833 ();
 FILLCELL_X32 FILLER_375_865 ();
 FILLCELL_X32 FILLER_375_897 ();
 FILLCELL_X32 FILLER_375_929 ();
 FILLCELL_X32 FILLER_375_961 ();
 FILLCELL_X32 FILLER_375_993 ();
 FILLCELL_X32 FILLER_375_1025 ();
 FILLCELL_X32 FILLER_375_1057 ();
 FILLCELL_X32 FILLER_375_1089 ();
 FILLCELL_X32 FILLER_375_1121 ();
 FILLCELL_X32 FILLER_375_1153 ();
 FILLCELL_X32 FILLER_375_1185 ();
 FILLCELL_X32 FILLER_375_1217 ();
 FILLCELL_X8 FILLER_375_1249 ();
 FILLCELL_X4 FILLER_375_1257 ();
 FILLCELL_X2 FILLER_375_1261 ();
 FILLCELL_X32 FILLER_375_1264 ();
 FILLCELL_X32 FILLER_375_1296 ();
 FILLCELL_X32 FILLER_375_1328 ();
 FILLCELL_X32 FILLER_375_1360 ();
 FILLCELL_X32 FILLER_375_1392 ();
 FILLCELL_X32 FILLER_375_1424 ();
 FILLCELL_X32 FILLER_375_1456 ();
 FILLCELL_X32 FILLER_375_1488 ();
 FILLCELL_X32 FILLER_375_1520 ();
 FILLCELL_X32 FILLER_375_1552 ();
 FILLCELL_X32 FILLER_375_1584 ();
 FILLCELL_X32 FILLER_375_1616 ();
 FILLCELL_X32 FILLER_375_1648 ();
 FILLCELL_X32 FILLER_375_1680 ();
 FILLCELL_X32 FILLER_375_1712 ();
 FILLCELL_X32 FILLER_375_1744 ();
 FILLCELL_X32 FILLER_375_1776 ();
 FILLCELL_X32 FILLER_375_1808 ();
 FILLCELL_X32 FILLER_375_1840 ();
 FILLCELL_X32 FILLER_375_1872 ();
 FILLCELL_X32 FILLER_375_1904 ();
 FILLCELL_X32 FILLER_375_1936 ();
 FILLCELL_X32 FILLER_375_1968 ();
 FILLCELL_X32 FILLER_375_2000 ();
 FILLCELL_X32 FILLER_375_2032 ();
 FILLCELL_X32 FILLER_375_2064 ();
 FILLCELL_X32 FILLER_375_2096 ();
 FILLCELL_X32 FILLER_375_2128 ();
 FILLCELL_X32 FILLER_375_2160 ();
 FILLCELL_X32 FILLER_375_2192 ();
 FILLCELL_X32 FILLER_375_2224 ();
 FILLCELL_X32 FILLER_375_2256 ();
 FILLCELL_X32 FILLER_375_2288 ();
 FILLCELL_X32 FILLER_375_2320 ();
 FILLCELL_X32 FILLER_375_2352 ();
 FILLCELL_X32 FILLER_375_2384 ();
 FILLCELL_X32 FILLER_375_2416 ();
 FILLCELL_X32 FILLER_375_2448 ();
 FILLCELL_X32 FILLER_375_2480 ();
 FILLCELL_X8 FILLER_375_2512 ();
 FILLCELL_X4 FILLER_375_2520 ();
 FILLCELL_X2 FILLER_375_2524 ();
 FILLCELL_X32 FILLER_375_2527 ();
 FILLCELL_X32 FILLER_375_2559 ();
 FILLCELL_X32 FILLER_375_2591 ();
 FILLCELL_X32 FILLER_375_2623 ();
 FILLCELL_X32 FILLER_375_2655 ();
 FILLCELL_X32 FILLER_375_2687 ();
 FILLCELL_X32 FILLER_375_2719 ();
 FILLCELL_X32 FILLER_375_2751 ();
 FILLCELL_X32 FILLER_375_2783 ();
 FILLCELL_X32 FILLER_375_2815 ();
 FILLCELL_X32 FILLER_375_2847 ();
 FILLCELL_X32 FILLER_375_2879 ();
 FILLCELL_X32 FILLER_375_2911 ();
 FILLCELL_X32 FILLER_375_2943 ();
 FILLCELL_X32 FILLER_375_2975 ();
 FILLCELL_X32 FILLER_375_3007 ();
 FILLCELL_X32 FILLER_375_3039 ();
 FILLCELL_X32 FILLER_375_3071 ();
 FILLCELL_X32 FILLER_375_3103 ();
 FILLCELL_X32 FILLER_375_3135 ();
 FILLCELL_X32 FILLER_375_3167 ();
 FILLCELL_X32 FILLER_375_3199 ();
 FILLCELL_X32 FILLER_375_3231 ();
 FILLCELL_X32 FILLER_375_3263 ();
 FILLCELL_X32 FILLER_375_3295 ();
 FILLCELL_X32 FILLER_375_3327 ();
 FILLCELL_X32 FILLER_375_3359 ();
 FILLCELL_X32 FILLER_375_3391 ();
 FILLCELL_X32 FILLER_375_3423 ();
 FILLCELL_X32 FILLER_375_3455 ();
 FILLCELL_X32 FILLER_375_3487 ();
 FILLCELL_X32 FILLER_375_3519 ();
 FILLCELL_X32 FILLER_375_3551 ();
 FILLCELL_X32 FILLER_375_3583 ();
 FILLCELL_X32 FILLER_375_3615 ();
 FILLCELL_X32 FILLER_375_3647 ();
 FILLCELL_X32 FILLER_375_3679 ();
 FILLCELL_X16 FILLER_375_3711 ();
 FILLCELL_X8 FILLER_375_3727 ();
 FILLCELL_X2 FILLER_375_3735 ();
 FILLCELL_X1 FILLER_375_3737 ();
 FILLCELL_X32 FILLER_376_1 ();
 FILLCELL_X32 FILLER_376_33 ();
 FILLCELL_X32 FILLER_376_65 ();
 FILLCELL_X32 FILLER_376_97 ();
 FILLCELL_X32 FILLER_376_129 ();
 FILLCELL_X32 FILLER_376_161 ();
 FILLCELL_X32 FILLER_376_193 ();
 FILLCELL_X32 FILLER_376_225 ();
 FILLCELL_X32 FILLER_376_257 ();
 FILLCELL_X32 FILLER_376_289 ();
 FILLCELL_X32 FILLER_376_321 ();
 FILLCELL_X32 FILLER_376_353 ();
 FILLCELL_X32 FILLER_376_385 ();
 FILLCELL_X32 FILLER_376_417 ();
 FILLCELL_X32 FILLER_376_449 ();
 FILLCELL_X32 FILLER_376_481 ();
 FILLCELL_X32 FILLER_376_513 ();
 FILLCELL_X32 FILLER_376_545 ();
 FILLCELL_X32 FILLER_376_577 ();
 FILLCELL_X16 FILLER_376_609 ();
 FILLCELL_X4 FILLER_376_625 ();
 FILLCELL_X2 FILLER_376_629 ();
 FILLCELL_X32 FILLER_376_632 ();
 FILLCELL_X32 FILLER_376_664 ();
 FILLCELL_X32 FILLER_376_696 ();
 FILLCELL_X32 FILLER_376_728 ();
 FILLCELL_X32 FILLER_376_760 ();
 FILLCELL_X32 FILLER_376_792 ();
 FILLCELL_X32 FILLER_376_824 ();
 FILLCELL_X32 FILLER_376_856 ();
 FILLCELL_X32 FILLER_376_888 ();
 FILLCELL_X32 FILLER_376_920 ();
 FILLCELL_X32 FILLER_376_952 ();
 FILLCELL_X32 FILLER_376_984 ();
 FILLCELL_X32 FILLER_376_1016 ();
 FILLCELL_X32 FILLER_376_1048 ();
 FILLCELL_X32 FILLER_376_1080 ();
 FILLCELL_X32 FILLER_376_1112 ();
 FILLCELL_X32 FILLER_376_1144 ();
 FILLCELL_X32 FILLER_376_1176 ();
 FILLCELL_X32 FILLER_376_1208 ();
 FILLCELL_X32 FILLER_376_1240 ();
 FILLCELL_X32 FILLER_376_1272 ();
 FILLCELL_X32 FILLER_376_1304 ();
 FILLCELL_X32 FILLER_376_1336 ();
 FILLCELL_X32 FILLER_376_1368 ();
 FILLCELL_X32 FILLER_376_1400 ();
 FILLCELL_X32 FILLER_376_1432 ();
 FILLCELL_X32 FILLER_376_1464 ();
 FILLCELL_X32 FILLER_376_1496 ();
 FILLCELL_X32 FILLER_376_1528 ();
 FILLCELL_X32 FILLER_376_1560 ();
 FILLCELL_X32 FILLER_376_1592 ();
 FILLCELL_X32 FILLER_376_1624 ();
 FILLCELL_X32 FILLER_376_1656 ();
 FILLCELL_X32 FILLER_376_1688 ();
 FILLCELL_X32 FILLER_376_1720 ();
 FILLCELL_X32 FILLER_376_1752 ();
 FILLCELL_X32 FILLER_376_1784 ();
 FILLCELL_X32 FILLER_376_1816 ();
 FILLCELL_X32 FILLER_376_1848 ();
 FILLCELL_X8 FILLER_376_1880 ();
 FILLCELL_X4 FILLER_376_1888 ();
 FILLCELL_X2 FILLER_376_1892 ();
 FILLCELL_X32 FILLER_376_1895 ();
 FILLCELL_X32 FILLER_376_1927 ();
 FILLCELL_X32 FILLER_376_1959 ();
 FILLCELL_X32 FILLER_376_1991 ();
 FILLCELL_X32 FILLER_376_2023 ();
 FILLCELL_X32 FILLER_376_2055 ();
 FILLCELL_X32 FILLER_376_2087 ();
 FILLCELL_X32 FILLER_376_2119 ();
 FILLCELL_X32 FILLER_376_2151 ();
 FILLCELL_X32 FILLER_376_2183 ();
 FILLCELL_X32 FILLER_376_2215 ();
 FILLCELL_X32 FILLER_376_2247 ();
 FILLCELL_X32 FILLER_376_2279 ();
 FILLCELL_X32 FILLER_376_2311 ();
 FILLCELL_X32 FILLER_376_2343 ();
 FILLCELL_X32 FILLER_376_2375 ();
 FILLCELL_X32 FILLER_376_2407 ();
 FILLCELL_X32 FILLER_376_2439 ();
 FILLCELL_X32 FILLER_376_2471 ();
 FILLCELL_X32 FILLER_376_2503 ();
 FILLCELL_X32 FILLER_376_2535 ();
 FILLCELL_X32 FILLER_376_2567 ();
 FILLCELL_X32 FILLER_376_2599 ();
 FILLCELL_X32 FILLER_376_2631 ();
 FILLCELL_X32 FILLER_376_2663 ();
 FILLCELL_X32 FILLER_376_2695 ();
 FILLCELL_X32 FILLER_376_2727 ();
 FILLCELL_X32 FILLER_376_2759 ();
 FILLCELL_X32 FILLER_376_2791 ();
 FILLCELL_X32 FILLER_376_2823 ();
 FILLCELL_X32 FILLER_376_2855 ();
 FILLCELL_X32 FILLER_376_2887 ();
 FILLCELL_X32 FILLER_376_2919 ();
 FILLCELL_X32 FILLER_376_2951 ();
 FILLCELL_X32 FILLER_376_2983 ();
 FILLCELL_X32 FILLER_376_3015 ();
 FILLCELL_X32 FILLER_376_3047 ();
 FILLCELL_X32 FILLER_376_3079 ();
 FILLCELL_X32 FILLER_376_3111 ();
 FILLCELL_X8 FILLER_376_3143 ();
 FILLCELL_X4 FILLER_376_3151 ();
 FILLCELL_X2 FILLER_376_3155 ();
 FILLCELL_X32 FILLER_376_3158 ();
 FILLCELL_X32 FILLER_376_3190 ();
 FILLCELL_X32 FILLER_376_3222 ();
 FILLCELL_X32 FILLER_376_3254 ();
 FILLCELL_X32 FILLER_376_3286 ();
 FILLCELL_X32 FILLER_376_3318 ();
 FILLCELL_X32 FILLER_376_3350 ();
 FILLCELL_X32 FILLER_376_3382 ();
 FILLCELL_X32 FILLER_376_3414 ();
 FILLCELL_X32 FILLER_376_3446 ();
 FILLCELL_X32 FILLER_376_3478 ();
 FILLCELL_X32 FILLER_376_3510 ();
 FILLCELL_X32 FILLER_376_3542 ();
 FILLCELL_X32 FILLER_376_3574 ();
 FILLCELL_X32 FILLER_376_3606 ();
 FILLCELL_X32 FILLER_376_3638 ();
 FILLCELL_X32 FILLER_376_3670 ();
 FILLCELL_X32 FILLER_376_3702 ();
 FILLCELL_X4 FILLER_376_3734 ();
 FILLCELL_X32 FILLER_377_1 ();
 FILLCELL_X32 FILLER_377_33 ();
 FILLCELL_X32 FILLER_377_65 ();
 FILLCELL_X32 FILLER_377_97 ();
 FILLCELL_X32 FILLER_377_129 ();
 FILLCELL_X32 FILLER_377_161 ();
 FILLCELL_X32 FILLER_377_193 ();
 FILLCELL_X32 FILLER_377_225 ();
 FILLCELL_X32 FILLER_377_257 ();
 FILLCELL_X32 FILLER_377_289 ();
 FILLCELL_X32 FILLER_377_321 ();
 FILLCELL_X32 FILLER_377_353 ();
 FILLCELL_X32 FILLER_377_385 ();
 FILLCELL_X32 FILLER_377_417 ();
 FILLCELL_X32 FILLER_377_449 ();
 FILLCELL_X32 FILLER_377_481 ();
 FILLCELL_X32 FILLER_377_513 ();
 FILLCELL_X32 FILLER_377_545 ();
 FILLCELL_X32 FILLER_377_577 ();
 FILLCELL_X32 FILLER_377_609 ();
 FILLCELL_X32 FILLER_377_641 ();
 FILLCELL_X32 FILLER_377_673 ();
 FILLCELL_X32 FILLER_377_705 ();
 FILLCELL_X32 FILLER_377_737 ();
 FILLCELL_X32 FILLER_377_769 ();
 FILLCELL_X32 FILLER_377_801 ();
 FILLCELL_X32 FILLER_377_833 ();
 FILLCELL_X32 FILLER_377_865 ();
 FILLCELL_X32 FILLER_377_897 ();
 FILLCELL_X32 FILLER_377_929 ();
 FILLCELL_X32 FILLER_377_961 ();
 FILLCELL_X32 FILLER_377_993 ();
 FILLCELL_X32 FILLER_377_1025 ();
 FILLCELL_X32 FILLER_377_1057 ();
 FILLCELL_X32 FILLER_377_1089 ();
 FILLCELL_X32 FILLER_377_1121 ();
 FILLCELL_X32 FILLER_377_1153 ();
 FILLCELL_X32 FILLER_377_1185 ();
 FILLCELL_X32 FILLER_377_1217 ();
 FILLCELL_X8 FILLER_377_1249 ();
 FILLCELL_X4 FILLER_377_1257 ();
 FILLCELL_X2 FILLER_377_1261 ();
 FILLCELL_X32 FILLER_377_1264 ();
 FILLCELL_X32 FILLER_377_1296 ();
 FILLCELL_X32 FILLER_377_1328 ();
 FILLCELL_X32 FILLER_377_1360 ();
 FILLCELL_X32 FILLER_377_1392 ();
 FILLCELL_X32 FILLER_377_1424 ();
 FILLCELL_X32 FILLER_377_1456 ();
 FILLCELL_X32 FILLER_377_1488 ();
 FILLCELL_X32 FILLER_377_1520 ();
 FILLCELL_X32 FILLER_377_1552 ();
 FILLCELL_X32 FILLER_377_1584 ();
 FILLCELL_X32 FILLER_377_1616 ();
 FILLCELL_X32 FILLER_377_1648 ();
 FILLCELL_X32 FILLER_377_1680 ();
 FILLCELL_X32 FILLER_377_1712 ();
 FILLCELL_X32 FILLER_377_1744 ();
 FILLCELL_X32 FILLER_377_1776 ();
 FILLCELL_X32 FILLER_377_1808 ();
 FILLCELL_X32 FILLER_377_1840 ();
 FILLCELL_X32 FILLER_377_1872 ();
 FILLCELL_X32 FILLER_377_1904 ();
 FILLCELL_X32 FILLER_377_1936 ();
 FILLCELL_X32 FILLER_377_1968 ();
 FILLCELL_X32 FILLER_377_2000 ();
 FILLCELL_X32 FILLER_377_2032 ();
 FILLCELL_X32 FILLER_377_2064 ();
 FILLCELL_X32 FILLER_377_2096 ();
 FILLCELL_X32 FILLER_377_2128 ();
 FILLCELL_X32 FILLER_377_2160 ();
 FILLCELL_X32 FILLER_377_2192 ();
 FILLCELL_X32 FILLER_377_2224 ();
 FILLCELL_X32 FILLER_377_2256 ();
 FILLCELL_X32 FILLER_377_2288 ();
 FILLCELL_X32 FILLER_377_2320 ();
 FILLCELL_X32 FILLER_377_2352 ();
 FILLCELL_X32 FILLER_377_2384 ();
 FILLCELL_X32 FILLER_377_2416 ();
 FILLCELL_X32 FILLER_377_2448 ();
 FILLCELL_X32 FILLER_377_2480 ();
 FILLCELL_X8 FILLER_377_2512 ();
 FILLCELL_X4 FILLER_377_2520 ();
 FILLCELL_X2 FILLER_377_2524 ();
 FILLCELL_X32 FILLER_377_2527 ();
 FILLCELL_X32 FILLER_377_2559 ();
 FILLCELL_X32 FILLER_377_2591 ();
 FILLCELL_X32 FILLER_377_2623 ();
 FILLCELL_X32 FILLER_377_2655 ();
 FILLCELL_X32 FILLER_377_2687 ();
 FILLCELL_X32 FILLER_377_2719 ();
 FILLCELL_X32 FILLER_377_2751 ();
 FILLCELL_X32 FILLER_377_2783 ();
 FILLCELL_X32 FILLER_377_2815 ();
 FILLCELL_X32 FILLER_377_2847 ();
 FILLCELL_X32 FILLER_377_2879 ();
 FILLCELL_X32 FILLER_377_2911 ();
 FILLCELL_X32 FILLER_377_2943 ();
 FILLCELL_X32 FILLER_377_2975 ();
 FILLCELL_X32 FILLER_377_3007 ();
 FILLCELL_X32 FILLER_377_3039 ();
 FILLCELL_X32 FILLER_377_3071 ();
 FILLCELL_X32 FILLER_377_3103 ();
 FILLCELL_X32 FILLER_377_3135 ();
 FILLCELL_X32 FILLER_377_3167 ();
 FILLCELL_X32 FILLER_377_3199 ();
 FILLCELL_X32 FILLER_377_3231 ();
 FILLCELL_X32 FILLER_377_3263 ();
 FILLCELL_X32 FILLER_377_3295 ();
 FILLCELL_X32 FILLER_377_3327 ();
 FILLCELL_X32 FILLER_377_3359 ();
 FILLCELL_X32 FILLER_377_3391 ();
 FILLCELL_X32 FILLER_377_3423 ();
 FILLCELL_X32 FILLER_377_3455 ();
 FILLCELL_X32 FILLER_377_3487 ();
 FILLCELL_X32 FILLER_377_3519 ();
 FILLCELL_X32 FILLER_377_3551 ();
 FILLCELL_X32 FILLER_377_3583 ();
 FILLCELL_X32 FILLER_377_3615 ();
 FILLCELL_X32 FILLER_377_3647 ();
 FILLCELL_X32 FILLER_377_3679 ();
 FILLCELL_X16 FILLER_377_3711 ();
 FILLCELL_X8 FILLER_377_3727 ();
 FILLCELL_X2 FILLER_377_3735 ();
 FILLCELL_X1 FILLER_377_3737 ();
 FILLCELL_X32 FILLER_378_1 ();
 FILLCELL_X32 FILLER_378_33 ();
 FILLCELL_X32 FILLER_378_65 ();
 FILLCELL_X32 FILLER_378_97 ();
 FILLCELL_X32 FILLER_378_129 ();
 FILLCELL_X32 FILLER_378_161 ();
 FILLCELL_X32 FILLER_378_193 ();
 FILLCELL_X32 FILLER_378_225 ();
 FILLCELL_X32 FILLER_378_257 ();
 FILLCELL_X32 FILLER_378_289 ();
 FILLCELL_X32 FILLER_378_321 ();
 FILLCELL_X32 FILLER_378_353 ();
 FILLCELL_X32 FILLER_378_385 ();
 FILLCELL_X32 FILLER_378_417 ();
 FILLCELL_X32 FILLER_378_449 ();
 FILLCELL_X32 FILLER_378_481 ();
 FILLCELL_X32 FILLER_378_513 ();
 FILLCELL_X32 FILLER_378_545 ();
 FILLCELL_X32 FILLER_378_577 ();
 FILLCELL_X16 FILLER_378_609 ();
 FILLCELL_X4 FILLER_378_625 ();
 FILLCELL_X2 FILLER_378_629 ();
 FILLCELL_X32 FILLER_378_632 ();
 FILLCELL_X32 FILLER_378_664 ();
 FILLCELL_X32 FILLER_378_696 ();
 FILLCELL_X32 FILLER_378_728 ();
 FILLCELL_X32 FILLER_378_760 ();
 FILLCELL_X32 FILLER_378_792 ();
 FILLCELL_X32 FILLER_378_824 ();
 FILLCELL_X32 FILLER_378_856 ();
 FILLCELL_X32 FILLER_378_888 ();
 FILLCELL_X32 FILLER_378_920 ();
 FILLCELL_X32 FILLER_378_952 ();
 FILLCELL_X32 FILLER_378_984 ();
 FILLCELL_X32 FILLER_378_1016 ();
 FILLCELL_X32 FILLER_378_1048 ();
 FILLCELL_X32 FILLER_378_1080 ();
 FILLCELL_X32 FILLER_378_1112 ();
 FILLCELL_X32 FILLER_378_1144 ();
 FILLCELL_X32 FILLER_378_1176 ();
 FILLCELL_X32 FILLER_378_1208 ();
 FILLCELL_X32 FILLER_378_1240 ();
 FILLCELL_X32 FILLER_378_1272 ();
 FILLCELL_X32 FILLER_378_1304 ();
 FILLCELL_X32 FILLER_378_1336 ();
 FILLCELL_X32 FILLER_378_1368 ();
 FILLCELL_X32 FILLER_378_1400 ();
 FILLCELL_X32 FILLER_378_1432 ();
 FILLCELL_X32 FILLER_378_1464 ();
 FILLCELL_X32 FILLER_378_1496 ();
 FILLCELL_X32 FILLER_378_1528 ();
 FILLCELL_X32 FILLER_378_1560 ();
 FILLCELL_X32 FILLER_378_1592 ();
 FILLCELL_X32 FILLER_378_1624 ();
 FILLCELL_X32 FILLER_378_1656 ();
 FILLCELL_X32 FILLER_378_1688 ();
 FILLCELL_X32 FILLER_378_1720 ();
 FILLCELL_X32 FILLER_378_1752 ();
 FILLCELL_X32 FILLER_378_1784 ();
 FILLCELL_X32 FILLER_378_1816 ();
 FILLCELL_X32 FILLER_378_1848 ();
 FILLCELL_X8 FILLER_378_1880 ();
 FILLCELL_X4 FILLER_378_1888 ();
 FILLCELL_X2 FILLER_378_1892 ();
 FILLCELL_X32 FILLER_378_1895 ();
 FILLCELL_X32 FILLER_378_1927 ();
 FILLCELL_X32 FILLER_378_1959 ();
 FILLCELL_X32 FILLER_378_1991 ();
 FILLCELL_X32 FILLER_378_2023 ();
 FILLCELL_X32 FILLER_378_2055 ();
 FILLCELL_X32 FILLER_378_2087 ();
 FILLCELL_X32 FILLER_378_2119 ();
 FILLCELL_X32 FILLER_378_2151 ();
 FILLCELL_X32 FILLER_378_2183 ();
 FILLCELL_X32 FILLER_378_2215 ();
 FILLCELL_X32 FILLER_378_2247 ();
 FILLCELL_X32 FILLER_378_2279 ();
 FILLCELL_X32 FILLER_378_2311 ();
 FILLCELL_X32 FILLER_378_2343 ();
 FILLCELL_X32 FILLER_378_2375 ();
 FILLCELL_X32 FILLER_378_2407 ();
 FILLCELL_X32 FILLER_378_2439 ();
 FILLCELL_X32 FILLER_378_2471 ();
 FILLCELL_X32 FILLER_378_2503 ();
 FILLCELL_X32 FILLER_378_2535 ();
 FILLCELL_X32 FILLER_378_2567 ();
 FILLCELL_X32 FILLER_378_2599 ();
 FILLCELL_X32 FILLER_378_2631 ();
 FILLCELL_X32 FILLER_378_2663 ();
 FILLCELL_X32 FILLER_378_2695 ();
 FILLCELL_X32 FILLER_378_2727 ();
 FILLCELL_X32 FILLER_378_2759 ();
 FILLCELL_X32 FILLER_378_2791 ();
 FILLCELL_X32 FILLER_378_2823 ();
 FILLCELL_X32 FILLER_378_2855 ();
 FILLCELL_X32 FILLER_378_2887 ();
 FILLCELL_X32 FILLER_378_2919 ();
 FILLCELL_X32 FILLER_378_2951 ();
 FILLCELL_X32 FILLER_378_2983 ();
 FILLCELL_X32 FILLER_378_3015 ();
 FILLCELL_X32 FILLER_378_3047 ();
 FILLCELL_X32 FILLER_378_3079 ();
 FILLCELL_X32 FILLER_378_3111 ();
 FILLCELL_X8 FILLER_378_3143 ();
 FILLCELL_X4 FILLER_378_3151 ();
 FILLCELL_X2 FILLER_378_3155 ();
 FILLCELL_X32 FILLER_378_3158 ();
 FILLCELL_X32 FILLER_378_3190 ();
 FILLCELL_X32 FILLER_378_3222 ();
 FILLCELL_X32 FILLER_378_3254 ();
 FILLCELL_X32 FILLER_378_3286 ();
 FILLCELL_X32 FILLER_378_3318 ();
 FILLCELL_X32 FILLER_378_3350 ();
 FILLCELL_X32 FILLER_378_3382 ();
 FILLCELL_X32 FILLER_378_3414 ();
 FILLCELL_X32 FILLER_378_3446 ();
 FILLCELL_X32 FILLER_378_3478 ();
 FILLCELL_X32 FILLER_378_3510 ();
 FILLCELL_X32 FILLER_378_3542 ();
 FILLCELL_X32 FILLER_378_3574 ();
 FILLCELL_X32 FILLER_378_3606 ();
 FILLCELL_X32 FILLER_378_3638 ();
 FILLCELL_X32 FILLER_378_3670 ();
 FILLCELL_X32 FILLER_378_3702 ();
 FILLCELL_X4 FILLER_378_3734 ();
 FILLCELL_X32 FILLER_379_1 ();
 FILLCELL_X32 FILLER_379_33 ();
 FILLCELL_X32 FILLER_379_65 ();
 FILLCELL_X32 FILLER_379_97 ();
 FILLCELL_X32 FILLER_379_129 ();
 FILLCELL_X32 FILLER_379_161 ();
 FILLCELL_X32 FILLER_379_193 ();
 FILLCELL_X32 FILLER_379_225 ();
 FILLCELL_X32 FILLER_379_257 ();
 FILLCELL_X32 FILLER_379_289 ();
 FILLCELL_X32 FILLER_379_321 ();
 FILLCELL_X32 FILLER_379_353 ();
 FILLCELL_X32 FILLER_379_385 ();
 FILLCELL_X32 FILLER_379_417 ();
 FILLCELL_X32 FILLER_379_449 ();
 FILLCELL_X32 FILLER_379_481 ();
 FILLCELL_X32 FILLER_379_513 ();
 FILLCELL_X32 FILLER_379_545 ();
 FILLCELL_X32 FILLER_379_577 ();
 FILLCELL_X32 FILLER_379_609 ();
 FILLCELL_X32 FILLER_379_641 ();
 FILLCELL_X32 FILLER_379_673 ();
 FILLCELL_X32 FILLER_379_705 ();
 FILLCELL_X32 FILLER_379_737 ();
 FILLCELL_X32 FILLER_379_769 ();
 FILLCELL_X32 FILLER_379_801 ();
 FILLCELL_X32 FILLER_379_833 ();
 FILLCELL_X32 FILLER_379_865 ();
 FILLCELL_X32 FILLER_379_897 ();
 FILLCELL_X32 FILLER_379_929 ();
 FILLCELL_X32 FILLER_379_961 ();
 FILLCELL_X32 FILLER_379_993 ();
 FILLCELL_X32 FILLER_379_1025 ();
 FILLCELL_X32 FILLER_379_1057 ();
 FILLCELL_X32 FILLER_379_1089 ();
 FILLCELL_X32 FILLER_379_1121 ();
 FILLCELL_X32 FILLER_379_1153 ();
 FILLCELL_X32 FILLER_379_1185 ();
 FILLCELL_X32 FILLER_379_1217 ();
 FILLCELL_X8 FILLER_379_1249 ();
 FILLCELL_X4 FILLER_379_1257 ();
 FILLCELL_X2 FILLER_379_1261 ();
 FILLCELL_X32 FILLER_379_1264 ();
 FILLCELL_X32 FILLER_379_1296 ();
 FILLCELL_X32 FILLER_379_1328 ();
 FILLCELL_X32 FILLER_379_1360 ();
 FILLCELL_X32 FILLER_379_1392 ();
 FILLCELL_X32 FILLER_379_1424 ();
 FILLCELL_X32 FILLER_379_1456 ();
 FILLCELL_X32 FILLER_379_1488 ();
 FILLCELL_X32 FILLER_379_1520 ();
 FILLCELL_X32 FILLER_379_1552 ();
 FILLCELL_X32 FILLER_379_1584 ();
 FILLCELL_X32 FILLER_379_1616 ();
 FILLCELL_X32 FILLER_379_1648 ();
 FILLCELL_X32 FILLER_379_1680 ();
 FILLCELL_X32 FILLER_379_1712 ();
 FILLCELL_X32 FILLER_379_1744 ();
 FILLCELL_X32 FILLER_379_1776 ();
 FILLCELL_X32 FILLER_379_1808 ();
 FILLCELL_X32 FILLER_379_1840 ();
 FILLCELL_X32 FILLER_379_1872 ();
 FILLCELL_X32 FILLER_379_1904 ();
 FILLCELL_X32 FILLER_379_1936 ();
 FILLCELL_X32 FILLER_379_1968 ();
 FILLCELL_X32 FILLER_379_2000 ();
 FILLCELL_X32 FILLER_379_2032 ();
 FILLCELL_X32 FILLER_379_2064 ();
 FILLCELL_X32 FILLER_379_2096 ();
 FILLCELL_X32 FILLER_379_2128 ();
 FILLCELL_X32 FILLER_379_2160 ();
 FILLCELL_X32 FILLER_379_2192 ();
 FILLCELL_X32 FILLER_379_2224 ();
 FILLCELL_X32 FILLER_379_2256 ();
 FILLCELL_X32 FILLER_379_2288 ();
 FILLCELL_X32 FILLER_379_2320 ();
 FILLCELL_X32 FILLER_379_2352 ();
 FILLCELL_X32 FILLER_379_2384 ();
 FILLCELL_X32 FILLER_379_2416 ();
 FILLCELL_X32 FILLER_379_2448 ();
 FILLCELL_X32 FILLER_379_2480 ();
 FILLCELL_X8 FILLER_379_2512 ();
 FILLCELL_X4 FILLER_379_2520 ();
 FILLCELL_X2 FILLER_379_2524 ();
 FILLCELL_X32 FILLER_379_2527 ();
 FILLCELL_X32 FILLER_379_2559 ();
 FILLCELL_X32 FILLER_379_2591 ();
 FILLCELL_X32 FILLER_379_2623 ();
 FILLCELL_X32 FILLER_379_2655 ();
 FILLCELL_X32 FILLER_379_2687 ();
 FILLCELL_X32 FILLER_379_2719 ();
 FILLCELL_X32 FILLER_379_2751 ();
 FILLCELL_X32 FILLER_379_2783 ();
 FILLCELL_X32 FILLER_379_2815 ();
 FILLCELL_X32 FILLER_379_2847 ();
 FILLCELL_X32 FILLER_379_2879 ();
 FILLCELL_X32 FILLER_379_2911 ();
 FILLCELL_X32 FILLER_379_2943 ();
 FILLCELL_X32 FILLER_379_2975 ();
 FILLCELL_X32 FILLER_379_3007 ();
 FILLCELL_X32 FILLER_379_3039 ();
 FILLCELL_X32 FILLER_379_3071 ();
 FILLCELL_X32 FILLER_379_3103 ();
 FILLCELL_X32 FILLER_379_3135 ();
 FILLCELL_X32 FILLER_379_3167 ();
 FILLCELL_X32 FILLER_379_3199 ();
 FILLCELL_X32 FILLER_379_3231 ();
 FILLCELL_X32 FILLER_379_3263 ();
 FILLCELL_X32 FILLER_379_3295 ();
 FILLCELL_X32 FILLER_379_3327 ();
 FILLCELL_X32 FILLER_379_3359 ();
 FILLCELL_X32 FILLER_379_3391 ();
 FILLCELL_X32 FILLER_379_3423 ();
 FILLCELL_X32 FILLER_379_3455 ();
 FILLCELL_X32 FILLER_379_3487 ();
 FILLCELL_X32 FILLER_379_3519 ();
 FILLCELL_X32 FILLER_379_3551 ();
 FILLCELL_X32 FILLER_379_3583 ();
 FILLCELL_X32 FILLER_379_3615 ();
 FILLCELL_X32 FILLER_379_3647 ();
 FILLCELL_X32 FILLER_379_3679 ();
 FILLCELL_X16 FILLER_379_3711 ();
 FILLCELL_X8 FILLER_379_3727 ();
 FILLCELL_X2 FILLER_379_3735 ();
 FILLCELL_X1 FILLER_379_3737 ();
 FILLCELL_X32 FILLER_380_1 ();
 FILLCELL_X32 FILLER_380_33 ();
 FILLCELL_X32 FILLER_380_65 ();
 FILLCELL_X32 FILLER_380_97 ();
 FILLCELL_X32 FILLER_380_129 ();
 FILLCELL_X32 FILLER_380_161 ();
 FILLCELL_X32 FILLER_380_193 ();
 FILLCELL_X32 FILLER_380_225 ();
 FILLCELL_X32 FILLER_380_257 ();
 FILLCELL_X32 FILLER_380_289 ();
 FILLCELL_X32 FILLER_380_321 ();
 FILLCELL_X32 FILLER_380_353 ();
 FILLCELL_X32 FILLER_380_385 ();
 FILLCELL_X32 FILLER_380_417 ();
 FILLCELL_X32 FILLER_380_449 ();
 FILLCELL_X32 FILLER_380_481 ();
 FILLCELL_X32 FILLER_380_513 ();
 FILLCELL_X32 FILLER_380_545 ();
 FILLCELL_X32 FILLER_380_577 ();
 FILLCELL_X16 FILLER_380_609 ();
 FILLCELL_X4 FILLER_380_625 ();
 FILLCELL_X2 FILLER_380_629 ();
 FILLCELL_X32 FILLER_380_632 ();
 FILLCELL_X32 FILLER_380_664 ();
 FILLCELL_X32 FILLER_380_696 ();
 FILLCELL_X32 FILLER_380_728 ();
 FILLCELL_X32 FILLER_380_760 ();
 FILLCELL_X32 FILLER_380_792 ();
 FILLCELL_X32 FILLER_380_824 ();
 FILLCELL_X32 FILLER_380_856 ();
 FILLCELL_X32 FILLER_380_888 ();
 FILLCELL_X32 FILLER_380_920 ();
 FILLCELL_X32 FILLER_380_952 ();
 FILLCELL_X32 FILLER_380_984 ();
 FILLCELL_X32 FILLER_380_1016 ();
 FILLCELL_X32 FILLER_380_1048 ();
 FILLCELL_X32 FILLER_380_1080 ();
 FILLCELL_X32 FILLER_380_1112 ();
 FILLCELL_X32 FILLER_380_1144 ();
 FILLCELL_X32 FILLER_380_1176 ();
 FILLCELL_X32 FILLER_380_1208 ();
 FILLCELL_X32 FILLER_380_1240 ();
 FILLCELL_X32 FILLER_380_1272 ();
 FILLCELL_X32 FILLER_380_1304 ();
 FILLCELL_X32 FILLER_380_1336 ();
 FILLCELL_X32 FILLER_380_1368 ();
 FILLCELL_X32 FILLER_380_1400 ();
 FILLCELL_X32 FILLER_380_1432 ();
 FILLCELL_X32 FILLER_380_1464 ();
 FILLCELL_X32 FILLER_380_1496 ();
 FILLCELL_X32 FILLER_380_1528 ();
 FILLCELL_X32 FILLER_380_1560 ();
 FILLCELL_X32 FILLER_380_1592 ();
 FILLCELL_X32 FILLER_380_1624 ();
 FILLCELL_X32 FILLER_380_1656 ();
 FILLCELL_X32 FILLER_380_1688 ();
 FILLCELL_X32 FILLER_380_1720 ();
 FILLCELL_X32 FILLER_380_1752 ();
 FILLCELL_X32 FILLER_380_1784 ();
 FILLCELL_X32 FILLER_380_1816 ();
 FILLCELL_X32 FILLER_380_1848 ();
 FILLCELL_X8 FILLER_380_1880 ();
 FILLCELL_X4 FILLER_380_1888 ();
 FILLCELL_X2 FILLER_380_1892 ();
 FILLCELL_X32 FILLER_380_1895 ();
 FILLCELL_X32 FILLER_380_1927 ();
 FILLCELL_X32 FILLER_380_1959 ();
 FILLCELL_X32 FILLER_380_1991 ();
 FILLCELL_X32 FILLER_380_2023 ();
 FILLCELL_X32 FILLER_380_2055 ();
 FILLCELL_X32 FILLER_380_2087 ();
 FILLCELL_X32 FILLER_380_2119 ();
 FILLCELL_X32 FILLER_380_2151 ();
 FILLCELL_X32 FILLER_380_2183 ();
 FILLCELL_X32 FILLER_380_2215 ();
 FILLCELL_X32 FILLER_380_2247 ();
 FILLCELL_X32 FILLER_380_2279 ();
 FILLCELL_X32 FILLER_380_2311 ();
 FILLCELL_X32 FILLER_380_2343 ();
 FILLCELL_X32 FILLER_380_2375 ();
 FILLCELL_X32 FILLER_380_2407 ();
 FILLCELL_X32 FILLER_380_2439 ();
 FILLCELL_X32 FILLER_380_2471 ();
 FILLCELL_X32 FILLER_380_2503 ();
 FILLCELL_X32 FILLER_380_2535 ();
 FILLCELL_X32 FILLER_380_2567 ();
 FILLCELL_X32 FILLER_380_2599 ();
 FILLCELL_X32 FILLER_380_2631 ();
 FILLCELL_X32 FILLER_380_2663 ();
 FILLCELL_X32 FILLER_380_2695 ();
 FILLCELL_X32 FILLER_380_2727 ();
 FILLCELL_X32 FILLER_380_2759 ();
 FILLCELL_X32 FILLER_380_2791 ();
 FILLCELL_X32 FILLER_380_2823 ();
 FILLCELL_X32 FILLER_380_2855 ();
 FILLCELL_X32 FILLER_380_2887 ();
 FILLCELL_X32 FILLER_380_2919 ();
 FILLCELL_X32 FILLER_380_2951 ();
 FILLCELL_X32 FILLER_380_2983 ();
 FILLCELL_X32 FILLER_380_3015 ();
 FILLCELL_X32 FILLER_380_3047 ();
 FILLCELL_X32 FILLER_380_3079 ();
 FILLCELL_X32 FILLER_380_3111 ();
 FILLCELL_X8 FILLER_380_3143 ();
 FILLCELL_X4 FILLER_380_3151 ();
 FILLCELL_X2 FILLER_380_3155 ();
 FILLCELL_X32 FILLER_380_3158 ();
 FILLCELL_X32 FILLER_380_3190 ();
 FILLCELL_X32 FILLER_380_3222 ();
 FILLCELL_X32 FILLER_380_3254 ();
 FILLCELL_X32 FILLER_380_3286 ();
 FILLCELL_X32 FILLER_380_3318 ();
 FILLCELL_X32 FILLER_380_3350 ();
 FILLCELL_X32 FILLER_380_3382 ();
 FILLCELL_X32 FILLER_380_3414 ();
 FILLCELL_X32 FILLER_380_3446 ();
 FILLCELL_X32 FILLER_380_3478 ();
 FILLCELL_X32 FILLER_380_3510 ();
 FILLCELL_X32 FILLER_380_3542 ();
 FILLCELL_X32 FILLER_380_3574 ();
 FILLCELL_X32 FILLER_380_3606 ();
 FILLCELL_X32 FILLER_380_3638 ();
 FILLCELL_X32 FILLER_380_3670 ();
 FILLCELL_X32 FILLER_380_3702 ();
 FILLCELL_X4 FILLER_380_3734 ();
 FILLCELL_X32 FILLER_381_1 ();
 FILLCELL_X32 FILLER_381_33 ();
 FILLCELL_X32 FILLER_381_65 ();
 FILLCELL_X32 FILLER_381_97 ();
 FILLCELL_X32 FILLER_381_129 ();
 FILLCELL_X32 FILLER_381_161 ();
 FILLCELL_X32 FILLER_381_193 ();
 FILLCELL_X32 FILLER_381_225 ();
 FILLCELL_X32 FILLER_381_257 ();
 FILLCELL_X32 FILLER_381_289 ();
 FILLCELL_X32 FILLER_381_321 ();
 FILLCELL_X32 FILLER_381_353 ();
 FILLCELL_X32 FILLER_381_385 ();
 FILLCELL_X32 FILLER_381_417 ();
 FILLCELL_X32 FILLER_381_449 ();
 FILLCELL_X32 FILLER_381_481 ();
 FILLCELL_X32 FILLER_381_513 ();
 FILLCELL_X32 FILLER_381_545 ();
 FILLCELL_X32 FILLER_381_577 ();
 FILLCELL_X32 FILLER_381_609 ();
 FILLCELL_X32 FILLER_381_641 ();
 FILLCELL_X32 FILLER_381_673 ();
 FILLCELL_X32 FILLER_381_705 ();
 FILLCELL_X32 FILLER_381_737 ();
 FILLCELL_X32 FILLER_381_769 ();
 FILLCELL_X32 FILLER_381_801 ();
 FILLCELL_X32 FILLER_381_833 ();
 FILLCELL_X32 FILLER_381_865 ();
 FILLCELL_X32 FILLER_381_897 ();
 FILLCELL_X32 FILLER_381_929 ();
 FILLCELL_X32 FILLER_381_961 ();
 FILLCELL_X32 FILLER_381_993 ();
 FILLCELL_X32 FILLER_381_1025 ();
 FILLCELL_X32 FILLER_381_1057 ();
 FILLCELL_X32 FILLER_381_1089 ();
 FILLCELL_X32 FILLER_381_1121 ();
 FILLCELL_X32 FILLER_381_1153 ();
 FILLCELL_X32 FILLER_381_1185 ();
 FILLCELL_X32 FILLER_381_1217 ();
 FILLCELL_X8 FILLER_381_1249 ();
 FILLCELL_X4 FILLER_381_1257 ();
 FILLCELL_X2 FILLER_381_1261 ();
 FILLCELL_X32 FILLER_381_1264 ();
 FILLCELL_X32 FILLER_381_1296 ();
 FILLCELL_X32 FILLER_381_1328 ();
 FILLCELL_X32 FILLER_381_1360 ();
 FILLCELL_X32 FILLER_381_1392 ();
 FILLCELL_X32 FILLER_381_1424 ();
 FILLCELL_X32 FILLER_381_1456 ();
 FILLCELL_X32 FILLER_381_1488 ();
 FILLCELL_X32 FILLER_381_1520 ();
 FILLCELL_X32 FILLER_381_1552 ();
 FILLCELL_X32 FILLER_381_1584 ();
 FILLCELL_X32 FILLER_381_1616 ();
 FILLCELL_X32 FILLER_381_1648 ();
 FILLCELL_X32 FILLER_381_1680 ();
 FILLCELL_X32 FILLER_381_1712 ();
 FILLCELL_X32 FILLER_381_1744 ();
 FILLCELL_X32 FILLER_381_1776 ();
 FILLCELL_X32 FILLER_381_1808 ();
 FILLCELL_X32 FILLER_381_1840 ();
 FILLCELL_X32 FILLER_381_1872 ();
 FILLCELL_X32 FILLER_381_1904 ();
 FILLCELL_X32 FILLER_381_1936 ();
 FILLCELL_X32 FILLER_381_1968 ();
 FILLCELL_X32 FILLER_381_2000 ();
 FILLCELL_X32 FILLER_381_2032 ();
 FILLCELL_X32 FILLER_381_2064 ();
 FILLCELL_X32 FILLER_381_2096 ();
 FILLCELL_X32 FILLER_381_2128 ();
 FILLCELL_X32 FILLER_381_2160 ();
 FILLCELL_X32 FILLER_381_2192 ();
 FILLCELL_X32 FILLER_381_2224 ();
 FILLCELL_X32 FILLER_381_2256 ();
 FILLCELL_X32 FILLER_381_2288 ();
 FILLCELL_X32 FILLER_381_2320 ();
 FILLCELL_X32 FILLER_381_2352 ();
 FILLCELL_X32 FILLER_381_2384 ();
 FILLCELL_X32 FILLER_381_2416 ();
 FILLCELL_X32 FILLER_381_2448 ();
 FILLCELL_X32 FILLER_381_2480 ();
 FILLCELL_X8 FILLER_381_2512 ();
 FILLCELL_X4 FILLER_381_2520 ();
 FILLCELL_X2 FILLER_381_2524 ();
 FILLCELL_X32 FILLER_381_2527 ();
 FILLCELL_X32 FILLER_381_2559 ();
 FILLCELL_X32 FILLER_381_2591 ();
 FILLCELL_X32 FILLER_381_2623 ();
 FILLCELL_X32 FILLER_381_2655 ();
 FILLCELL_X32 FILLER_381_2687 ();
 FILLCELL_X32 FILLER_381_2719 ();
 FILLCELL_X32 FILLER_381_2751 ();
 FILLCELL_X32 FILLER_381_2783 ();
 FILLCELL_X32 FILLER_381_2815 ();
 FILLCELL_X32 FILLER_381_2847 ();
 FILLCELL_X32 FILLER_381_2879 ();
 FILLCELL_X32 FILLER_381_2911 ();
 FILLCELL_X32 FILLER_381_2943 ();
 FILLCELL_X32 FILLER_381_2975 ();
 FILLCELL_X32 FILLER_381_3007 ();
 FILLCELL_X32 FILLER_381_3039 ();
 FILLCELL_X32 FILLER_381_3071 ();
 FILLCELL_X32 FILLER_381_3103 ();
 FILLCELL_X32 FILLER_381_3135 ();
 FILLCELL_X32 FILLER_381_3167 ();
 FILLCELL_X32 FILLER_381_3199 ();
 FILLCELL_X32 FILLER_381_3231 ();
 FILLCELL_X32 FILLER_381_3263 ();
 FILLCELL_X32 FILLER_381_3295 ();
 FILLCELL_X32 FILLER_381_3327 ();
 FILLCELL_X32 FILLER_381_3359 ();
 FILLCELL_X32 FILLER_381_3391 ();
 FILLCELL_X32 FILLER_381_3423 ();
 FILLCELL_X32 FILLER_381_3455 ();
 FILLCELL_X32 FILLER_381_3487 ();
 FILLCELL_X32 FILLER_381_3519 ();
 FILLCELL_X32 FILLER_381_3551 ();
 FILLCELL_X32 FILLER_381_3583 ();
 FILLCELL_X32 FILLER_381_3615 ();
 FILLCELL_X32 FILLER_381_3647 ();
 FILLCELL_X32 FILLER_381_3679 ();
 FILLCELL_X16 FILLER_381_3711 ();
 FILLCELL_X8 FILLER_381_3727 ();
 FILLCELL_X2 FILLER_381_3735 ();
 FILLCELL_X1 FILLER_381_3737 ();
 FILLCELL_X32 FILLER_382_1 ();
 FILLCELL_X32 FILLER_382_33 ();
 FILLCELL_X32 FILLER_382_65 ();
 FILLCELL_X32 FILLER_382_97 ();
 FILLCELL_X32 FILLER_382_129 ();
 FILLCELL_X32 FILLER_382_161 ();
 FILLCELL_X32 FILLER_382_193 ();
 FILLCELL_X32 FILLER_382_225 ();
 FILLCELL_X32 FILLER_382_257 ();
 FILLCELL_X32 FILLER_382_289 ();
 FILLCELL_X32 FILLER_382_321 ();
 FILLCELL_X32 FILLER_382_353 ();
 FILLCELL_X32 FILLER_382_385 ();
 FILLCELL_X32 FILLER_382_417 ();
 FILLCELL_X32 FILLER_382_449 ();
 FILLCELL_X32 FILLER_382_481 ();
 FILLCELL_X32 FILLER_382_513 ();
 FILLCELL_X32 FILLER_382_545 ();
 FILLCELL_X32 FILLER_382_577 ();
 FILLCELL_X16 FILLER_382_609 ();
 FILLCELL_X4 FILLER_382_625 ();
 FILLCELL_X2 FILLER_382_629 ();
 FILLCELL_X32 FILLER_382_632 ();
 FILLCELL_X32 FILLER_382_664 ();
 FILLCELL_X32 FILLER_382_696 ();
 FILLCELL_X32 FILLER_382_728 ();
 FILLCELL_X32 FILLER_382_760 ();
 FILLCELL_X32 FILLER_382_792 ();
 FILLCELL_X32 FILLER_382_824 ();
 FILLCELL_X32 FILLER_382_856 ();
 FILLCELL_X32 FILLER_382_888 ();
 FILLCELL_X32 FILLER_382_920 ();
 FILLCELL_X32 FILLER_382_952 ();
 FILLCELL_X32 FILLER_382_984 ();
 FILLCELL_X32 FILLER_382_1016 ();
 FILLCELL_X32 FILLER_382_1048 ();
 FILLCELL_X32 FILLER_382_1080 ();
 FILLCELL_X32 FILLER_382_1112 ();
 FILLCELL_X32 FILLER_382_1144 ();
 FILLCELL_X32 FILLER_382_1176 ();
 FILLCELL_X32 FILLER_382_1208 ();
 FILLCELL_X32 FILLER_382_1240 ();
 FILLCELL_X32 FILLER_382_1272 ();
 FILLCELL_X32 FILLER_382_1304 ();
 FILLCELL_X32 FILLER_382_1336 ();
 FILLCELL_X32 FILLER_382_1368 ();
 FILLCELL_X32 FILLER_382_1400 ();
 FILLCELL_X32 FILLER_382_1432 ();
 FILLCELL_X32 FILLER_382_1464 ();
 FILLCELL_X32 FILLER_382_1496 ();
 FILLCELL_X32 FILLER_382_1528 ();
 FILLCELL_X32 FILLER_382_1560 ();
 FILLCELL_X32 FILLER_382_1592 ();
 FILLCELL_X32 FILLER_382_1624 ();
 FILLCELL_X32 FILLER_382_1656 ();
 FILLCELL_X32 FILLER_382_1688 ();
 FILLCELL_X32 FILLER_382_1720 ();
 FILLCELL_X32 FILLER_382_1752 ();
 FILLCELL_X32 FILLER_382_1784 ();
 FILLCELL_X32 FILLER_382_1816 ();
 FILLCELL_X32 FILLER_382_1848 ();
 FILLCELL_X8 FILLER_382_1880 ();
 FILLCELL_X4 FILLER_382_1888 ();
 FILLCELL_X2 FILLER_382_1892 ();
 FILLCELL_X32 FILLER_382_1895 ();
 FILLCELL_X32 FILLER_382_1927 ();
 FILLCELL_X32 FILLER_382_1959 ();
 FILLCELL_X32 FILLER_382_1991 ();
 FILLCELL_X32 FILLER_382_2023 ();
 FILLCELL_X32 FILLER_382_2055 ();
 FILLCELL_X32 FILLER_382_2087 ();
 FILLCELL_X32 FILLER_382_2119 ();
 FILLCELL_X32 FILLER_382_2151 ();
 FILLCELL_X32 FILLER_382_2183 ();
 FILLCELL_X32 FILLER_382_2215 ();
 FILLCELL_X32 FILLER_382_2247 ();
 FILLCELL_X32 FILLER_382_2279 ();
 FILLCELL_X32 FILLER_382_2311 ();
 FILLCELL_X32 FILLER_382_2343 ();
 FILLCELL_X32 FILLER_382_2375 ();
 FILLCELL_X32 FILLER_382_2407 ();
 FILLCELL_X32 FILLER_382_2439 ();
 FILLCELL_X32 FILLER_382_2471 ();
 FILLCELL_X32 FILLER_382_2503 ();
 FILLCELL_X32 FILLER_382_2535 ();
 FILLCELL_X32 FILLER_382_2567 ();
 FILLCELL_X32 FILLER_382_2599 ();
 FILLCELL_X32 FILLER_382_2631 ();
 FILLCELL_X32 FILLER_382_2663 ();
 FILLCELL_X32 FILLER_382_2695 ();
 FILLCELL_X32 FILLER_382_2727 ();
 FILLCELL_X32 FILLER_382_2759 ();
 FILLCELL_X32 FILLER_382_2791 ();
 FILLCELL_X32 FILLER_382_2823 ();
 FILLCELL_X32 FILLER_382_2855 ();
 FILLCELL_X32 FILLER_382_2887 ();
 FILLCELL_X32 FILLER_382_2919 ();
 FILLCELL_X32 FILLER_382_2951 ();
 FILLCELL_X32 FILLER_382_2983 ();
 FILLCELL_X32 FILLER_382_3015 ();
 FILLCELL_X32 FILLER_382_3047 ();
 FILLCELL_X32 FILLER_382_3079 ();
 FILLCELL_X32 FILLER_382_3111 ();
 FILLCELL_X8 FILLER_382_3143 ();
 FILLCELL_X4 FILLER_382_3151 ();
 FILLCELL_X2 FILLER_382_3155 ();
 FILLCELL_X32 FILLER_382_3158 ();
 FILLCELL_X32 FILLER_382_3190 ();
 FILLCELL_X32 FILLER_382_3222 ();
 FILLCELL_X32 FILLER_382_3254 ();
 FILLCELL_X32 FILLER_382_3286 ();
 FILLCELL_X32 FILLER_382_3318 ();
 FILLCELL_X32 FILLER_382_3350 ();
 FILLCELL_X32 FILLER_382_3382 ();
 FILLCELL_X32 FILLER_382_3414 ();
 FILLCELL_X32 FILLER_382_3446 ();
 FILLCELL_X32 FILLER_382_3478 ();
 FILLCELL_X32 FILLER_382_3510 ();
 FILLCELL_X32 FILLER_382_3542 ();
 FILLCELL_X32 FILLER_382_3574 ();
 FILLCELL_X32 FILLER_382_3606 ();
 FILLCELL_X32 FILLER_382_3638 ();
 FILLCELL_X32 FILLER_382_3670 ();
 FILLCELL_X32 FILLER_382_3702 ();
 FILLCELL_X4 FILLER_382_3734 ();
 FILLCELL_X32 FILLER_383_1 ();
 FILLCELL_X32 FILLER_383_33 ();
 FILLCELL_X32 FILLER_383_65 ();
 FILLCELL_X32 FILLER_383_97 ();
 FILLCELL_X32 FILLER_383_129 ();
 FILLCELL_X32 FILLER_383_161 ();
 FILLCELL_X32 FILLER_383_193 ();
 FILLCELL_X32 FILLER_383_225 ();
 FILLCELL_X32 FILLER_383_257 ();
 FILLCELL_X32 FILLER_383_289 ();
 FILLCELL_X32 FILLER_383_321 ();
 FILLCELL_X32 FILLER_383_353 ();
 FILLCELL_X32 FILLER_383_385 ();
 FILLCELL_X32 FILLER_383_417 ();
 FILLCELL_X32 FILLER_383_449 ();
 FILLCELL_X32 FILLER_383_481 ();
 FILLCELL_X32 FILLER_383_513 ();
 FILLCELL_X32 FILLER_383_545 ();
 FILLCELL_X32 FILLER_383_577 ();
 FILLCELL_X32 FILLER_383_609 ();
 FILLCELL_X32 FILLER_383_641 ();
 FILLCELL_X32 FILLER_383_673 ();
 FILLCELL_X32 FILLER_383_705 ();
 FILLCELL_X32 FILLER_383_737 ();
 FILLCELL_X32 FILLER_383_769 ();
 FILLCELL_X32 FILLER_383_801 ();
 FILLCELL_X32 FILLER_383_833 ();
 FILLCELL_X32 FILLER_383_865 ();
 FILLCELL_X32 FILLER_383_897 ();
 FILLCELL_X32 FILLER_383_929 ();
 FILLCELL_X32 FILLER_383_961 ();
 FILLCELL_X32 FILLER_383_993 ();
 FILLCELL_X32 FILLER_383_1025 ();
 FILLCELL_X32 FILLER_383_1057 ();
 FILLCELL_X32 FILLER_383_1089 ();
 FILLCELL_X32 FILLER_383_1121 ();
 FILLCELL_X32 FILLER_383_1153 ();
 FILLCELL_X32 FILLER_383_1185 ();
 FILLCELL_X32 FILLER_383_1217 ();
 FILLCELL_X8 FILLER_383_1249 ();
 FILLCELL_X4 FILLER_383_1257 ();
 FILLCELL_X2 FILLER_383_1261 ();
 FILLCELL_X32 FILLER_383_1264 ();
 FILLCELL_X32 FILLER_383_1296 ();
 FILLCELL_X32 FILLER_383_1328 ();
 FILLCELL_X32 FILLER_383_1360 ();
 FILLCELL_X32 FILLER_383_1392 ();
 FILLCELL_X32 FILLER_383_1424 ();
 FILLCELL_X32 FILLER_383_1456 ();
 FILLCELL_X32 FILLER_383_1488 ();
 FILLCELL_X32 FILLER_383_1520 ();
 FILLCELL_X32 FILLER_383_1552 ();
 FILLCELL_X32 FILLER_383_1584 ();
 FILLCELL_X32 FILLER_383_1616 ();
 FILLCELL_X32 FILLER_383_1648 ();
 FILLCELL_X32 FILLER_383_1680 ();
 FILLCELL_X32 FILLER_383_1712 ();
 FILLCELL_X32 FILLER_383_1744 ();
 FILLCELL_X32 FILLER_383_1776 ();
 FILLCELL_X32 FILLER_383_1808 ();
 FILLCELL_X32 FILLER_383_1840 ();
 FILLCELL_X32 FILLER_383_1872 ();
 FILLCELL_X32 FILLER_383_1904 ();
 FILLCELL_X32 FILLER_383_1936 ();
 FILLCELL_X32 FILLER_383_1968 ();
 FILLCELL_X32 FILLER_383_2000 ();
 FILLCELL_X32 FILLER_383_2032 ();
 FILLCELL_X32 FILLER_383_2064 ();
 FILLCELL_X32 FILLER_383_2096 ();
 FILLCELL_X32 FILLER_383_2128 ();
 FILLCELL_X32 FILLER_383_2160 ();
 FILLCELL_X32 FILLER_383_2192 ();
 FILLCELL_X32 FILLER_383_2224 ();
 FILLCELL_X32 FILLER_383_2256 ();
 FILLCELL_X32 FILLER_383_2288 ();
 FILLCELL_X32 FILLER_383_2320 ();
 FILLCELL_X32 FILLER_383_2352 ();
 FILLCELL_X32 FILLER_383_2384 ();
 FILLCELL_X32 FILLER_383_2416 ();
 FILLCELL_X32 FILLER_383_2448 ();
 FILLCELL_X32 FILLER_383_2480 ();
 FILLCELL_X8 FILLER_383_2512 ();
 FILLCELL_X4 FILLER_383_2520 ();
 FILLCELL_X2 FILLER_383_2524 ();
 FILLCELL_X32 FILLER_383_2527 ();
 FILLCELL_X32 FILLER_383_2559 ();
 FILLCELL_X32 FILLER_383_2591 ();
 FILLCELL_X32 FILLER_383_2623 ();
 FILLCELL_X32 FILLER_383_2655 ();
 FILLCELL_X32 FILLER_383_2687 ();
 FILLCELL_X32 FILLER_383_2719 ();
 FILLCELL_X32 FILLER_383_2751 ();
 FILLCELL_X32 FILLER_383_2783 ();
 FILLCELL_X32 FILLER_383_2815 ();
 FILLCELL_X32 FILLER_383_2847 ();
 FILLCELL_X32 FILLER_383_2879 ();
 FILLCELL_X32 FILLER_383_2911 ();
 FILLCELL_X32 FILLER_383_2943 ();
 FILLCELL_X32 FILLER_383_2975 ();
 FILLCELL_X32 FILLER_383_3007 ();
 FILLCELL_X32 FILLER_383_3039 ();
 FILLCELL_X32 FILLER_383_3071 ();
 FILLCELL_X32 FILLER_383_3103 ();
 FILLCELL_X32 FILLER_383_3135 ();
 FILLCELL_X32 FILLER_383_3167 ();
 FILLCELL_X32 FILLER_383_3199 ();
 FILLCELL_X32 FILLER_383_3231 ();
 FILLCELL_X32 FILLER_383_3263 ();
 FILLCELL_X32 FILLER_383_3295 ();
 FILLCELL_X32 FILLER_383_3327 ();
 FILLCELL_X32 FILLER_383_3359 ();
 FILLCELL_X32 FILLER_383_3391 ();
 FILLCELL_X32 FILLER_383_3423 ();
 FILLCELL_X32 FILLER_383_3455 ();
 FILLCELL_X32 FILLER_383_3487 ();
 FILLCELL_X32 FILLER_383_3519 ();
 FILLCELL_X32 FILLER_383_3551 ();
 FILLCELL_X32 FILLER_383_3583 ();
 FILLCELL_X32 FILLER_383_3615 ();
 FILLCELL_X32 FILLER_383_3647 ();
 FILLCELL_X32 FILLER_383_3679 ();
 FILLCELL_X16 FILLER_383_3711 ();
 FILLCELL_X8 FILLER_383_3727 ();
 FILLCELL_X2 FILLER_383_3735 ();
 FILLCELL_X1 FILLER_383_3737 ();
 FILLCELL_X32 FILLER_384_1 ();
 FILLCELL_X32 FILLER_384_33 ();
 FILLCELL_X32 FILLER_384_65 ();
 FILLCELL_X32 FILLER_384_97 ();
 FILLCELL_X32 FILLER_384_129 ();
 FILLCELL_X32 FILLER_384_161 ();
 FILLCELL_X32 FILLER_384_193 ();
 FILLCELL_X32 FILLER_384_225 ();
 FILLCELL_X32 FILLER_384_257 ();
 FILLCELL_X32 FILLER_384_289 ();
 FILLCELL_X32 FILLER_384_321 ();
 FILLCELL_X32 FILLER_384_353 ();
 FILLCELL_X32 FILLER_384_385 ();
 FILLCELL_X32 FILLER_384_417 ();
 FILLCELL_X32 FILLER_384_449 ();
 FILLCELL_X32 FILLER_384_481 ();
 FILLCELL_X32 FILLER_384_513 ();
 FILLCELL_X32 FILLER_384_545 ();
 FILLCELL_X32 FILLER_384_577 ();
 FILLCELL_X16 FILLER_384_609 ();
 FILLCELL_X4 FILLER_384_625 ();
 FILLCELL_X2 FILLER_384_629 ();
 FILLCELL_X32 FILLER_384_632 ();
 FILLCELL_X32 FILLER_384_664 ();
 FILLCELL_X32 FILLER_384_696 ();
 FILLCELL_X32 FILLER_384_728 ();
 FILLCELL_X32 FILLER_384_760 ();
 FILLCELL_X32 FILLER_384_792 ();
 FILLCELL_X32 FILLER_384_824 ();
 FILLCELL_X32 FILLER_384_856 ();
 FILLCELL_X32 FILLER_384_888 ();
 FILLCELL_X32 FILLER_384_920 ();
 FILLCELL_X32 FILLER_384_952 ();
 FILLCELL_X32 FILLER_384_984 ();
 FILLCELL_X32 FILLER_384_1016 ();
 FILLCELL_X32 FILLER_384_1048 ();
 FILLCELL_X32 FILLER_384_1080 ();
 FILLCELL_X32 FILLER_384_1112 ();
 FILLCELL_X32 FILLER_384_1144 ();
 FILLCELL_X32 FILLER_384_1176 ();
 FILLCELL_X32 FILLER_384_1208 ();
 FILLCELL_X32 FILLER_384_1240 ();
 FILLCELL_X32 FILLER_384_1272 ();
 FILLCELL_X32 FILLER_384_1304 ();
 FILLCELL_X32 FILLER_384_1336 ();
 FILLCELL_X32 FILLER_384_1368 ();
 FILLCELL_X32 FILLER_384_1400 ();
 FILLCELL_X32 FILLER_384_1432 ();
 FILLCELL_X32 FILLER_384_1464 ();
 FILLCELL_X32 FILLER_384_1496 ();
 FILLCELL_X32 FILLER_384_1528 ();
 FILLCELL_X32 FILLER_384_1560 ();
 FILLCELL_X32 FILLER_384_1592 ();
 FILLCELL_X32 FILLER_384_1624 ();
 FILLCELL_X32 FILLER_384_1656 ();
 FILLCELL_X32 FILLER_384_1688 ();
 FILLCELL_X32 FILLER_384_1720 ();
 FILLCELL_X32 FILLER_384_1752 ();
 FILLCELL_X32 FILLER_384_1784 ();
 FILLCELL_X32 FILLER_384_1816 ();
 FILLCELL_X32 FILLER_384_1848 ();
 FILLCELL_X8 FILLER_384_1880 ();
 FILLCELL_X4 FILLER_384_1888 ();
 FILLCELL_X2 FILLER_384_1892 ();
 FILLCELL_X32 FILLER_384_1895 ();
 FILLCELL_X32 FILLER_384_1927 ();
 FILLCELL_X32 FILLER_384_1959 ();
 FILLCELL_X32 FILLER_384_1991 ();
 FILLCELL_X32 FILLER_384_2023 ();
 FILLCELL_X32 FILLER_384_2055 ();
 FILLCELL_X32 FILLER_384_2087 ();
 FILLCELL_X32 FILLER_384_2119 ();
 FILLCELL_X32 FILLER_384_2151 ();
 FILLCELL_X32 FILLER_384_2183 ();
 FILLCELL_X32 FILLER_384_2215 ();
 FILLCELL_X32 FILLER_384_2247 ();
 FILLCELL_X32 FILLER_384_2279 ();
 FILLCELL_X32 FILLER_384_2311 ();
 FILLCELL_X32 FILLER_384_2343 ();
 FILLCELL_X32 FILLER_384_2375 ();
 FILLCELL_X32 FILLER_384_2407 ();
 FILLCELL_X32 FILLER_384_2439 ();
 FILLCELL_X32 FILLER_384_2471 ();
 FILLCELL_X32 FILLER_384_2503 ();
 FILLCELL_X32 FILLER_384_2535 ();
 FILLCELL_X32 FILLER_384_2567 ();
 FILLCELL_X32 FILLER_384_2599 ();
 FILLCELL_X32 FILLER_384_2631 ();
 FILLCELL_X32 FILLER_384_2663 ();
 FILLCELL_X32 FILLER_384_2695 ();
 FILLCELL_X32 FILLER_384_2727 ();
 FILLCELL_X32 FILLER_384_2759 ();
 FILLCELL_X32 FILLER_384_2791 ();
 FILLCELL_X32 FILLER_384_2823 ();
 FILLCELL_X32 FILLER_384_2855 ();
 FILLCELL_X32 FILLER_384_2887 ();
 FILLCELL_X32 FILLER_384_2919 ();
 FILLCELL_X32 FILLER_384_2951 ();
 FILLCELL_X32 FILLER_384_2983 ();
 FILLCELL_X32 FILLER_384_3015 ();
 FILLCELL_X32 FILLER_384_3047 ();
 FILLCELL_X32 FILLER_384_3079 ();
 FILLCELL_X32 FILLER_384_3111 ();
 FILLCELL_X8 FILLER_384_3143 ();
 FILLCELL_X4 FILLER_384_3151 ();
 FILLCELL_X2 FILLER_384_3155 ();
 FILLCELL_X32 FILLER_384_3158 ();
 FILLCELL_X32 FILLER_384_3190 ();
 FILLCELL_X32 FILLER_384_3222 ();
 FILLCELL_X32 FILLER_384_3254 ();
 FILLCELL_X32 FILLER_384_3286 ();
 FILLCELL_X32 FILLER_384_3318 ();
 FILLCELL_X32 FILLER_384_3350 ();
 FILLCELL_X32 FILLER_384_3382 ();
 FILLCELL_X32 FILLER_384_3414 ();
 FILLCELL_X32 FILLER_384_3446 ();
 FILLCELL_X32 FILLER_384_3478 ();
 FILLCELL_X32 FILLER_384_3510 ();
 FILLCELL_X32 FILLER_384_3542 ();
 FILLCELL_X32 FILLER_384_3574 ();
 FILLCELL_X32 FILLER_384_3606 ();
 FILLCELL_X32 FILLER_384_3638 ();
 FILLCELL_X32 FILLER_384_3670 ();
 FILLCELL_X32 FILLER_384_3702 ();
 FILLCELL_X4 FILLER_384_3734 ();
 FILLCELL_X32 FILLER_385_1 ();
 FILLCELL_X32 FILLER_385_33 ();
 FILLCELL_X32 FILLER_385_65 ();
 FILLCELL_X32 FILLER_385_97 ();
 FILLCELL_X32 FILLER_385_129 ();
 FILLCELL_X32 FILLER_385_161 ();
 FILLCELL_X32 FILLER_385_193 ();
 FILLCELL_X32 FILLER_385_225 ();
 FILLCELL_X32 FILLER_385_257 ();
 FILLCELL_X32 FILLER_385_289 ();
 FILLCELL_X32 FILLER_385_321 ();
 FILLCELL_X32 FILLER_385_353 ();
 FILLCELL_X32 FILLER_385_385 ();
 FILLCELL_X32 FILLER_385_417 ();
 FILLCELL_X32 FILLER_385_449 ();
 FILLCELL_X32 FILLER_385_481 ();
 FILLCELL_X32 FILLER_385_513 ();
 FILLCELL_X32 FILLER_385_545 ();
 FILLCELL_X32 FILLER_385_577 ();
 FILLCELL_X32 FILLER_385_609 ();
 FILLCELL_X32 FILLER_385_641 ();
 FILLCELL_X32 FILLER_385_673 ();
 FILLCELL_X32 FILLER_385_705 ();
 FILLCELL_X32 FILLER_385_737 ();
 FILLCELL_X32 FILLER_385_769 ();
 FILLCELL_X32 FILLER_385_801 ();
 FILLCELL_X32 FILLER_385_833 ();
 FILLCELL_X32 FILLER_385_865 ();
 FILLCELL_X32 FILLER_385_897 ();
 FILLCELL_X32 FILLER_385_929 ();
 FILLCELL_X32 FILLER_385_961 ();
 FILLCELL_X32 FILLER_385_993 ();
 FILLCELL_X32 FILLER_385_1025 ();
 FILLCELL_X32 FILLER_385_1057 ();
 FILLCELL_X32 FILLER_385_1089 ();
 FILLCELL_X32 FILLER_385_1121 ();
 FILLCELL_X32 FILLER_385_1153 ();
 FILLCELL_X32 FILLER_385_1185 ();
 FILLCELL_X32 FILLER_385_1217 ();
 FILLCELL_X8 FILLER_385_1249 ();
 FILLCELL_X4 FILLER_385_1257 ();
 FILLCELL_X2 FILLER_385_1261 ();
 FILLCELL_X32 FILLER_385_1264 ();
 FILLCELL_X32 FILLER_385_1296 ();
 FILLCELL_X32 FILLER_385_1328 ();
 FILLCELL_X32 FILLER_385_1360 ();
 FILLCELL_X32 FILLER_385_1392 ();
 FILLCELL_X32 FILLER_385_1424 ();
 FILLCELL_X32 FILLER_385_1456 ();
 FILLCELL_X32 FILLER_385_1488 ();
 FILLCELL_X32 FILLER_385_1520 ();
 FILLCELL_X32 FILLER_385_1552 ();
 FILLCELL_X32 FILLER_385_1584 ();
 FILLCELL_X32 FILLER_385_1616 ();
 FILLCELL_X32 FILLER_385_1648 ();
 FILLCELL_X32 FILLER_385_1680 ();
 FILLCELL_X32 FILLER_385_1712 ();
 FILLCELL_X32 FILLER_385_1744 ();
 FILLCELL_X32 FILLER_385_1776 ();
 FILLCELL_X32 FILLER_385_1808 ();
 FILLCELL_X32 FILLER_385_1840 ();
 FILLCELL_X32 FILLER_385_1872 ();
 FILLCELL_X32 FILLER_385_1904 ();
 FILLCELL_X32 FILLER_385_1936 ();
 FILLCELL_X32 FILLER_385_1968 ();
 FILLCELL_X32 FILLER_385_2000 ();
 FILLCELL_X32 FILLER_385_2032 ();
 FILLCELL_X32 FILLER_385_2064 ();
 FILLCELL_X32 FILLER_385_2096 ();
 FILLCELL_X32 FILLER_385_2128 ();
 FILLCELL_X32 FILLER_385_2160 ();
 FILLCELL_X32 FILLER_385_2192 ();
 FILLCELL_X32 FILLER_385_2224 ();
 FILLCELL_X32 FILLER_385_2256 ();
 FILLCELL_X32 FILLER_385_2288 ();
 FILLCELL_X32 FILLER_385_2320 ();
 FILLCELL_X32 FILLER_385_2352 ();
 FILLCELL_X32 FILLER_385_2384 ();
 FILLCELL_X32 FILLER_385_2416 ();
 FILLCELL_X32 FILLER_385_2448 ();
 FILLCELL_X32 FILLER_385_2480 ();
 FILLCELL_X8 FILLER_385_2512 ();
 FILLCELL_X4 FILLER_385_2520 ();
 FILLCELL_X2 FILLER_385_2524 ();
 FILLCELL_X32 FILLER_385_2527 ();
 FILLCELL_X32 FILLER_385_2559 ();
 FILLCELL_X32 FILLER_385_2591 ();
 FILLCELL_X32 FILLER_385_2623 ();
 FILLCELL_X32 FILLER_385_2655 ();
 FILLCELL_X32 FILLER_385_2687 ();
 FILLCELL_X32 FILLER_385_2719 ();
 FILLCELL_X32 FILLER_385_2751 ();
 FILLCELL_X32 FILLER_385_2783 ();
 FILLCELL_X32 FILLER_385_2815 ();
 FILLCELL_X32 FILLER_385_2847 ();
 FILLCELL_X32 FILLER_385_2879 ();
 FILLCELL_X32 FILLER_385_2911 ();
 FILLCELL_X32 FILLER_385_2943 ();
 FILLCELL_X32 FILLER_385_2975 ();
 FILLCELL_X32 FILLER_385_3007 ();
 FILLCELL_X32 FILLER_385_3039 ();
 FILLCELL_X32 FILLER_385_3071 ();
 FILLCELL_X32 FILLER_385_3103 ();
 FILLCELL_X32 FILLER_385_3135 ();
 FILLCELL_X32 FILLER_385_3167 ();
 FILLCELL_X32 FILLER_385_3199 ();
 FILLCELL_X32 FILLER_385_3231 ();
 FILLCELL_X32 FILLER_385_3263 ();
 FILLCELL_X32 FILLER_385_3295 ();
 FILLCELL_X32 FILLER_385_3327 ();
 FILLCELL_X32 FILLER_385_3359 ();
 FILLCELL_X32 FILLER_385_3391 ();
 FILLCELL_X32 FILLER_385_3423 ();
 FILLCELL_X32 FILLER_385_3455 ();
 FILLCELL_X32 FILLER_385_3487 ();
 FILLCELL_X32 FILLER_385_3519 ();
 FILLCELL_X32 FILLER_385_3551 ();
 FILLCELL_X32 FILLER_385_3583 ();
 FILLCELL_X32 FILLER_385_3615 ();
 FILLCELL_X32 FILLER_385_3647 ();
 FILLCELL_X32 FILLER_385_3679 ();
 FILLCELL_X16 FILLER_385_3711 ();
 FILLCELL_X8 FILLER_385_3727 ();
 FILLCELL_X2 FILLER_385_3735 ();
 FILLCELL_X1 FILLER_385_3737 ();
 FILLCELL_X32 FILLER_386_1 ();
 FILLCELL_X32 FILLER_386_33 ();
 FILLCELL_X32 FILLER_386_65 ();
 FILLCELL_X32 FILLER_386_97 ();
 FILLCELL_X32 FILLER_386_129 ();
 FILLCELL_X32 FILLER_386_161 ();
 FILLCELL_X32 FILLER_386_193 ();
 FILLCELL_X32 FILLER_386_225 ();
 FILLCELL_X32 FILLER_386_257 ();
 FILLCELL_X32 FILLER_386_289 ();
 FILLCELL_X32 FILLER_386_321 ();
 FILLCELL_X32 FILLER_386_353 ();
 FILLCELL_X32 FILLER_386_385 ();
 FILLCELL_X32 FILLER_386_417 ();
 FILLCELL_X32 FILLER_386_449 ();
 FILLCELL_X32 FILLER_386_481 ();
 FILLCELL_X32 FILLER_386_513 ();
 FILLCELL_X32 FILLER_386_545 ();
 FILLCELL_X32 FILLER_386_577 ();
 FILLCELL_X16 FILLER_386_609 ();
 FILLCELL_X4 FILLER_386_625 ();
 FILLCELL_X2 FILLER_386_629 ();
 FILLCELL_X32 FILLER_386_632 ();
 FILLCELL_X32 FILLER_386_664 ();
 FILLCELL_X32 FILLER_386_696 ();
 FILLCELL_X32 FILLER_386_728 ();
 FILLCELL_X32 FILLER_386_760 ();
 FILLCELL_X32 FILLER_386_792 ();
 FILLCELL_X32 FILLER_386_824 ();
 FILLCELL_X32 FILLER_386_856 ();
 FILLCELL_X32 FILLER_386_888 ();
 FILLCELL_X32 FILLER_386_920 ();
 FILLCELL_X32 FILLER_386_952 ();
 FILLCELL_X32 FILLER_386_984 ();
 FILLCELL_X32 FILLER_386_1016 ();
 FILLCELL_X32 FILLER_386_1048 ();
 FILLCELL_X32 FILLER_386_1080 ();
 FILLCELL_X32 FILLER_386_1112 ();
 FILLCELL_X32 FILLER_386_1144 ();
 FILLCELL_X32 FILLER_386_1176 ();
 FILLCELL_X32 FILLER_386_1208 ();
 FILLCELL_X32 FILLER_386_1240 ();
 FILLCELL_X32 FILLER_386_1272 ();
 FILLCELL_X32 FILLER_386_1304 ();
 FILLCELL_X32 FILLER_386_1336 ();
 FILLCELL_X32 FILLER_386_1368 ();
 FILLCELL_X32 FILLER_386_1400 ();
 FILLCELL_X32 FILLER_386_1432 ();
 FILLCELL_X32 FILLER_386_1464 ();
 FILLCELL_X32 FILLER_386_1496 ();
 FILLCELL_X32 FILLER_386_1528 ();
 FILLCELL_X32 FILLER_386_1560 ();
 FILLCELL_X32 FILLER_386_1592 ();
 FILLCELL_X32 FILLER_386_1624 ();
 FILLCELL_X32 FILLER_386_1656 ();
 FILLCELL_X32 FILLER_386_1688 ();
 FILLCELL_X32 FILLER_386_1720 ();
 FILLCELL_X32 FILLER_386_1752 ();
 FILLCELL_X32 FILLER_386_1784 ();
 FILLCELL_X32 FILLER_386_1816 ();
 FILLCELL_X32 FILLER_386_1848 ();
 FILLCELL_X8 FILLER_386_1880 ();
 FILLCELL_X4 FILLER_386_1888 ();
 FILLCELL_X2 FILLER_386_1892 ();
 FILLCELL_X32 FILLER_386_1895 ();
 FILLCELL_X32 FILLER_386_1927 ();
 FILLCELL_X32 FILLER_386_1959 ();
 FILLCELL_X32 FILLER_386_1991 ();
 FILLCELL_X32 FILLER_386_2023 ();
 FILLCELL_X32 FILLER_386_2055 ();
 FILLCELL_X32 FILLER_386_2087 ();
 FILLCELL_X32 FILLER_386_2119 ();
 FILLCELL_X32 FILLER_386_2151 ();
 FILLCELL_X32 FILLER_386_2183 ();
 FILLCELL_X32 FILLER_386_2215 ();
 FILLCELL_X32 FILLER_386_2247 ();
 FILLCELL_X32 FILLER_386_2279 ();
 FILLCELL_X32 FILLER_386_2311 ();
 FILLCELL_X32 FILLER_386_2343 ();
 FILLCELL_X32 FILLER_386_2375 ();
 FILLCELL_X32 FILLER_386_2407 ();
 FILLCELL_X32 FILLER_386_2439 ();
 FILLCELL_X32 FILLER_386_2471 ();
 FILLCELL_X32 FILLER_386_2503 ();
 FILLCELL_X32 FILLER_386_2535 ();
 FILLCELL_X32 FILLER_386_2567 ();
 FILLCELL_X32 FILLER_386_2599 ();
 FILLCELL_X32 FILLER_386_2631 ();
 FILLCELL_X32 FILLER_386_2663 ();
 FILLCELL_X32 FILLER_386_2695 ();
 FILLCELL_X32 FILLER_386_2727 ();
 FILLCELL_X32 FILLER_386_2759 ();
 FILLCELL_X32 FILLER_386_2791 ();
 FILLCELL_X32 FILLER_386_2823 ();
 FILLCELL_X32 FILLER_386_2855 ();
 FILLCELL_X32 FILLER_386_2887 ();
 FILLCELL_X32 FILLER_386_2919 ();
 FILLCELL_X32 FILLER_386_2951 ();
 FILLCELL_X32 FILLER_386_2983 ();
 FILLCELL_X32 FILLER_386_3015 ();
 FILLCELL_X32 FILLER_386_3047 ();
 FILLCELL_X32 FILLER_386_3079 ();
 FILLCELL_X32 FILLER_386_3111 ();
 FILLCELL_X8 FILLER_386_3143 ();
 FILLCELL_X4 FILLER_386_3151 ();
 FILLCELL_X2 FILLER_386_3155 ();
 FILLCELL_X32 FILLER_386_3158 ();
 FILLCELL_X32 FILLER_386_3190 ();
 FILLCELL_X32 FILLER_386_3222 ();
 FILLCELL_X32 FILLER_386_3254 ();
 FILLCELL_X32 FILLER_386_3286 ();
 FILLCELL_X32 FILLER_386_3318 ();
 FILLCELL_X32 FILLER_386_3350 ();
 FILLCELL_X32 FILLER_386_3382 ();
 FILLCELL_X32 FILLER_386_3414 ();
 FILLCELL_X32 FILLER_386_3446 ();
 FILLCELL_X32 FILLER_386_3478 ();
 FILLCELL_X32 FILLER_386_3510 ();
 FILLCELL_X32 FILLER_386_3542 ();
 FILLCELL_X32 FILLER_386_3574 ();
 FILLCELL_X32 FILLER_386_3606 ();
 FILLCELL_X32 FILLER_386_3638 ();
 FILLCELL_X32 FILLER_386_3670 ();
 FILLCELL_X32 FILLER_386_3702 ();
 FILLCELL_X4 FILLER_386_3734 ();
 FILLCELL_X32 FILLER_387_1 ();
 FILLCELL_X32 FILLER_387_33 ();
 FILLCELL_X32 FILLER_387_65 ();
 FILLCELL_X32 FILLER_387_97 ();
 FILLCELL_X32 FILLER_387_129 ();
 FILLCELL_X32 FILLER_387_161 ();
 FILLCELL_X32 FILLER_387_193 ();
 FILLCELL_X32 FILLER_387_225 ();
 FILLCELL_X32 FILLER_387_257 ();
 FILLCELL_X32 FILLER_387_289 ();
 FILLCELL_X32 FILLER_387_321 ();
 FILLCELL_X32 FILLER_387_353 ();
 FILLCELL_X32 FILLER_387_385 ();
 FILLCELL_X32 FILLER_387_417 ();
 FILLCELL_X32 FILLER_387_449 ();
 FILLCELL_X32 FILLER_387_481 ();
 FILLCELL_X32 FILLER_387_513 ();
 FILLCELL_X32 FILLER_387_545 ();
 FILLCELL_X32 FILLER_387_577 ();
 FILLCELL_X32 FILLER_387_609 ();
 FILLCELL_X32 FILLER_387_641 ();
 FILLCELL_X32 FILLER_387_673 ();
 FILLCELL_X32 FILLER_387_705 ();
 FILLCELL_X32 FILLER_387_737 ();
 FILLCELL_X32 FILLER_387_769 ();
 FILLCELL_X32 FILLER_387_801 ();
 FILLCELL_X32 FILLER_387_833 ();
 FILLCELL_X32 FILLER_387_865 ();
 FILLCELL_X32 FILLER_387_897 ();
 FILLCELL_X32 FILLER_387_929 ();
 FILLCELL_X32 FILLER_387_961 ();
 FILLCELL_X32 FILLER_387_993 ();
 FILLCELL_X32 FILLER_387_1025 ();
 FILLCELL_X32 FILLER_387_1057 ();
 FILLCELL_X32 FILLER_387_1089 ();
 FILLCELL_X32 FILLER_387_1121 ();
 FILLCELL_X32 FILLER_387_1153 ();
 FILLCELL_X32 FILLER_387_1185 ();
 FILLCELL_X32 FILLER_387_1217 ();
 FILLCELL_X8 FILLER_387_1249 ();
 FILLCELL_X4 FILLER_387_1257 ();
 FILLCELL_X2 FILLER_387_1261 ();
 FILLCELL_X32 FILLER_387_1264 ();
 FILLCELL_X32 FILLER_387_1296 ();
 FILLCELL_X32 FILLER_387_1328 ();
 FILLCELL_X32 FILLER_387_1360 ();
 FILLCELL_X32 FILLER_387_1392 ();
 FILLCELL_X32 FILLER_387_1424 ();
 FILLCELL_X32 FILLER_387_1456 ();
 FILLCELL_X32 FILLER_387_1488 ();
 FILLCELL_X32 FILLER_387_1520 ();
 FILLCELL_X32 FILLER_387_1552 ();
 FILLCELL_X32 FILLER_387_1584 ();
 FILLCELL_X32 FILLER_387_1616 ();
 FILLCELL_X32 FILLER_387_1648 ();
 FILLCELL_X32 FILLER_387_1680 ();
 FILLCELL_X32 FILLER_387_1712 ();
 FILLCELL_X32 FILLER_387_1744 ();
 FILLCELL_X32 FILLER_387_1776 ();
 FILLCELL_X32 FILLER_387_1808 ();
 FILLCELL_X32 FILLER_387_1840 ();
 FILLCELL_X32 FILLER_387_1872 ();
 FILLCELL_X32 FILLER_387_1904 ();
 FILLCELL_X32 FILLER_387_1936 ();
 FILLCELL_X32 FILLER_387_1968 ();
 FILLCELL_X32 FILLER_387_2000 ();
 FILLCELL_X32 FILLER_387_2032 ();
 FILLCELL_X32 FILLER_387_2064 ();
 FILLCELL_X32 FILLER_387_2096 ();
 FILLCELL_X32 FILLER_387_2128 ();
 FILLCELL_X32 FILLER_387_2160 ();
 FILLCELL_X32 FILLER_387_2192 ();
 FILLCELL_X32 FILLER_387_2224 ();
 FILLCELL_X32 FILLER_387_2256 ();
 FILLCELL_X32 FILLER_387_2288 ();
 FILLCELL_X32 FILLER_387_2320 ();
 FILLCELL_X32 FILLER_387_2352 ();
 FILLCELL_X32 FILLER_387_2384 ();
 FILLCELL_X32 FILLER_387_2416 ();
 FILLCELL_X32 FILLER_387_2448 ();
 FILLCELL_X32 FILLER_387_2480 ();
 FILLCELL_X8 FILLER_387_2512 ();
 FILLCELL_X4 FILLER_387_2520 ();
 FILLCELL_X2 FILLER_387_2524 ();
 FILLCELL_X32 FILLER_387_2527 ();
 FILLCELL_X32 FILLER_387_2559 ();
 FILLCELL_X32 FILLER_387_2591 ();
 FILLCELL_X32 FILLER_387_2623 ();
 FILLCELL_X32 FILLER_387_2655 ();
 FILLCELL_X32 FILLER_387_2687 ();
 FILLCELL_X32 FILLER_387_2719 ();
 FILLCELL_X32 FILLER_387_2751 ();
 FILLCELL_X32 FILLER_387_2783 ();
 FILLCELL_X32 FILLER_387_2815 ();
 FILLCELL_X32 FILLER_387_2847 ();
 FILLCELL_X32 FILLER_387_2879 ();
 FILLCELL_X32 FILLER_387_2911 ();
 FILLCELL_X32 FILLER_387_2943 ();
 FILLCELL_X32 FILLER_387_2975 ();
 FILLCELL_X32 FILLER_387_3007 ();
 FILLCELL_X32 FILLER_387_3039 ();
 FILLCELL_X32 FILLER_387_3071 ();
 FILLCELL_X32 FILLER_387_3103 ();
 FILLCELL_X32 FILLER_387_3135 ();
 FILLCELL_X32 FILLER_387_3167 ();
 FILLCELL_X32 FILLER_387_3199 ();
 FILLCELL_X32 FILLER_387_3231 ();
 FILLCELL_X32 FILLER_387_3263 ();
 FILLCELL_X32 FILLER_387_3295 ();
 FILLCELL_X32 FILLER_387_3327 ();
 FILLCELL_X32 FILLER_387_3359 ();
 FILLCELL_X32 FILLER_387_3391 ();
 FILLCELL_X32 FILLER_387_3423 ();
 FILLCELL_X32 FILLER_387_3455 ();
 FILLCELL_X32 FILLER_387_3487 ();
 FILLCELL_X32 FILLER_387_3519 ();
 FILLCELL_X32 FILLER_387_3551 ();
 FILLCELL_X32 FILLER_387_3583 ();
 FILLCELL_X32 FILLER_387_3615 ();
 FILLCELL_X32 FILLER_387_3647 ();
 FILLCELL_X32 FILLER_387_3679 ();
 FILLCELL_X16 FILLER_387_3711 ();
 FILLCELL_X8 FILLER_387_3727 ();
 FILLCELL_X2 FILLER_387_3735 ();
 FILLCELL_X1 FILLER_387_3737 ();
 FILLCELL_X32 FILLER_388_1 ();
 FILLCELL_X32 FILLER_388_33 ();
 FILLCELL_X32 FILLER_388_65 ();
 FILLCELL_X32 FILLER_388_97 ();
 FILLCELL_X32 FILLER_388_129 ();
 FILLCELL_X32 FILLER_388_161 ();
 FILLCELL_X32 FILLER_388_193 ();
 FILLCELL_X32 FILLER_388_225 ();
 FILLCELL_X32 FILLER_388_257 ();
 FILLCELL_X32 FILLER_388_289 ();
 FILLCELL_X32 FILLER_388_321 ();
 FILLCELL_X32 FILLER_388_353 ();
 FILLCELL_X32 FILLER_388_385 ();
 FILLCELL_X32 FILLER_388_417 ();
 FILLCELL_X32 FILLER_388_449 ();
 FILLCELL_X32 FILLER_388_481 ();
 FILLCELL_X32 FILLER_388_513 ();
 FILLCELL_X32 FILLER_388_545 ();
 FILLCELL_X32 FILLER_388_577 ();
 FILLCELL_X16 FILLER_388_609 ();
 FILLCELL_X4 FILLER_388_625 ();
 FILLCELL_X2 FILLER_388_629 ();
 FILLCELL_X32 FILLER_388_632 ();
 FILLCELL_X32 FILLER_388_664 ();
 FILLCELL_X32 FILLER_388_696 ();
 FILLCELL_X32 FILLER_388_728 ();
 FILLCELL_X32 FILLER_388_760 ();
 FILLCELL_X32 FILLER_388_792 ();
 FILLCELL_X32 FILLER_388_824 ();
 FILLCELL_X32 FILLER_388_856 ();
 FILLCELL_X32 FILLER_388_888 ();
 FILLCELL_X32 FILLER_388_920 ();
 FILLCELL_X32 FILLER_388_952 ();
 FILLCELL_X32 FILLER_388_984 ();
 FILLCELL_X32 FILLER_388_1016 ();
 FILLCELL_X32 FILLER_388_1048 ();
 FILLCELL_X32 FILLER_388_1080 ();
 FILLCELL_X32 FILLER_388_1112 ();
 FILLCELL_X32 FILLER_388_1144 ();
 FILLCELL_X32 FILLER_388_1176 ();
 FILLCELL_X32 FILLER_388_1208 ();
 FILLCELL_X32 FILLER_388_1240 ();
 FILLCELL_X32 FILLER_388_1272 ();
 FILLCELL_X32 FILLER_388_1304 ();
 FILLCELL_X32 FILLER_388_1336 ();
 FILLCELL_X32 FILLER_388_1368 ();
 FILLCELL_X32 FILLER_388_1400 ();
 FILLCELL_X32 FILLER_388_1432 ();
 FILLCELL_X32 FILLER_388_1464 ();
 FILLCELL_X32 FILLER_388_1496 ();
 FILLCELL_X32 FILLER_388_1528 ();
 FILLCELL_X32 FILLER_388_1560 ();
 FILLCELL_X32 FILLER_388_1592 ();
 FILLCELL_X32 FILLER_388_1624 ();
 FILLCELL_X32 FILLER_388_1656 ();
 FILLCELL_X32 FILLER_388_1688 ();
 FILLCELL_X32 FILLER_388_1720 ();
 FILLCELL_X32 FILLER_388_1752 ();
 FILLCELL_X32 FILLER_388_1784 ();
 FILLCELL_X32 FILLER_388_1816 ();
 FILLCELL_X32 FILLER_388_1848 ();
 FILLCELL_X8 FILLER_388_1880 ();
 FILLCELL_X4 FILLER_388_1888 ();
 FILLCELL_X2 FILLER_388_1892 ();
 FILLCELL_X32 FILLER_388_1895 ();
 FILLCELL_X32 FILLER_388_1927 ();
 FILLCELL_X32 FILLER_388_1959 ();
 FILLCELL_X32 FILLER_388_1991 ();
 FILLCELL_X32 FILLER_388_2023 ();
 FILLCELL_X32 FILLER_388_2055 ();
 FILLCELL_X32 FILLER_388_2087 ();
 FILLCELL_X32 FILLER_388_2119 ();
 FILLCELL_X32 FILLER_388_2151 ();
 FILLCELL_X32 FILLER_388_2183 ();
 FILLCELL_X32 FILLER_388_2215 ();
 FILLCELL_X32 FILLER_388_2247 ();
 FILLCELL_X32 FILLER_388_2279 ();
 FILLCELL_X32 FILLER_388_2311 ();
 FILLCELL_X32 FILLER_388_2343 ();
 FILLCELL_X32 FILLER_388_2375 ();
 FILLCELL_X32 FILLER_388_2407 ();
 FILLCELL_X32 FILLER_388_2439 ();
 FILLCELL_X32 FILLER_388_2471 ();
 FILLCELL_X32 FILLER_388_2503 ();
 FILLCELL_X32 FILLER_388_2535 ();
 FILLCELL_X32 FILLER_388_2567 ();
 FILLCELL_X32 FILLER_388_2599 ();
 FILLCELL_X32 FILLER_388_2631 ();
 FILLCELL_X32 FILLER_388_2663 ();
 FILLCELL_X32 FILLER_388_2695 ();
 FILLCELL_X32 FILLER_388_2727 ();
 FILLCELL_X32 FILLER_388_2759 ();
 FILLCELL_X32 FILLER_388_2791 ();
 FILLCELL_X32 FILLER_388_2823 ();
 FILLCELL_X32 FILLER_388_2855 ();
 FILLCELL_X32 FILLER_388_2887 ();
 FILLCELL_X32 FILLER_388_2919 ();
 FILLCELL_X32 FILLER_388_2951 ();
 FILLCELL_X32 FILLER_388_2983 ();
 FILLCELL_X32 FILLER_388_3015 ();
 FILLCELL_X32 FILLER_388_3047 ();
 FILLCELL_X32 FILLER_388_3079 ();
 FILLCELL_X32 FILLER_388_3111 ();
 FILLCELL_X8 FILLER_388_3143 ();
 FILLCELL_X4 FILLER_388_3151 ();
 FILLCELL_X2 FILLER_388_3155 ();
 FILLCELL_X32 FILLER_388_3158 ();
 FILLCELL_X32 FILLER_388_3190 ();
 FILLCELL_X32 FILLER_388_3222 ();
 FILLCELL_X32 FILLER_388_3254 ();
 FILLCELL_X32 FILLER_388_3286 ();
 FILLCELL_X32 FILLER_388_3318 ();
 FILLCELL_X32 FILLER_388_3350 ();
 FILLCELL_X32 FILLER_388_3382 ();
 FILLCELL_X32 FILLER_388_3414 ();
 FILLCELL_X32 FILLER_388_3446 ();
 FILLCELL_X32 FILLER_388_3478 ();
 FILLCELL_X32 FILLER_388_3510 ();
 FILLCELL_X32 FILLER_388_3542 ();
 FILLCELL_X32 FILLER_388_3574 ();
 FILLCELL_X32 FILLER_388_3606 ();
 FILLCELL_X32 FILLER_388_3638 ();
 FILLCELL_X32 FILLER_388_3670 ();
 FILLCELL_X32 FILLER_388_3702 ();
 FILLCELL_X4 FILLER_388_3734 ();
 FILLCELL_X32 FILLER_389_1 ();
 FILLCELL_X32 FILLER_389_33 ();
 FILLCELL_X32 FILLER_389_65 ();
 FILLCELL_X32 FILLER_389_97 ();
 FILLCELL_X32 FILLER_389_129 ();
 FILLCELL_X32 FILLER_389_161 ();
 FILLCELL_X32 FILLER_389_193 ();
 FILLCELL_X32 FILLER_389_225 ();
 FILLCELL_X32 FILLER_389_257 ();
 FILLCELL_X32 FILLER_389_289 ();
 FILLCELL_X32 FILLER_389_321 ();
 FILLCELL_X32 FILLER_389_353 ();
 FILLCELL_X32 FILLER_389_385 ();
 FILLCELL_X32 FILLER_389_417 ();
 FILLCELL_X32 FILLER_389_449 ();
 FILLCELL_X32 FILLER_389_481 ();
 FILLCELL_X32 FILLER_389_513 ();
 FILLCELL_X32 FILLER_389_545 ();
 FILLCELL_X32 FILLER_389_577 ();
 FILLCELL_X32 FILLER_389_609 ();
 FILLCELL_X32 FILLER_389_641 ();
 FILLCELL_X32 FILLER_389_673 ();
 FILLCELL_X32 FILLER_389_705 ();
 FILLCELL_X32 FILLER_389_737 ();
 FILLCELL_X32 FILLER_389_769 ();
 FILLCELL_X32 FILLER_389_801 ();
 FILLCELL_X32 FILLER_389_833 ();
 FILLCELL_X32 FILLER_389_865 ();
 FILLCELL_X32 FILLER_389_897 ();
 FILLCELL_X32 FILLER_389_929 ();
 FILLCELL_X32 FILLER_389_961 ();
 FILLCELL_X32 FILLER_389_993 ();
 FILLCELL_X32 FILLER_389_1025 ();
 FILLCELL_X32 FILLER_389_1057 ();
 FILLCELL_X32 FILLER_389_1089 ();
 FILLCELL_X32 FILLER_389_1121 ();
 FILLCELL_X32 FILLER_389_1153 ();
 FILLCELL_X32 FILLER_389_1185 ();
 FILLCELL_X32 FILLER_389_1217 ();
 FILLCELL_X8 FILLER_389_1249 ();
 FILLCELL_X4 FILLER_389_1257 ();
 FILLCELL_X2 FILLER_389_1261 ();
 FILLCELL_X32 FILLER_389_1264 ();
 FILLCELL_X32 FILLER_389_1296 ();
 FILLCELL_X32 FILLER_389_1328 ();
 FILLCELL_X32 FILLER_389_1360 ();
 FILLCELL_X32 FILLER_389_1392 ();
 FILLCELL_X32 FILLER_389_1424 ();
 FILLCELL_X32 FILLER_389_1456 ();
 FILLCELL_X32 FILLER_389_1488 ();
 FILLCELL_X32 FILLER_389_1520 ();
 FILLCELL_X32 FILLER_389_1552 ();
 FILLCELL_X32 FILLER_389_1584 ();
 FILLCELL_X32 FILLER_389_1616 ();
 FILLCELL_X32 FILLER_389_1648 ();
 FILLCELL_X32 FILLER_389_1680 ();
 FILLCELL_X32 FILLER_389_1712 ();
 FILLCELL_X32 FILLER_389_1744 ();
 FILLCELL_X32 FILLER_389_1776 ();
 FILLCELL_X32 FILLER_389_1808 ();
 FILLCELL_X32 FILLER_389_1840 ();
 FILLCELL_X32 FILLER_389_1872 ();
 FILLCELL_X32 FILLER_389_1904 ();
 FILLCELL_X32 FILLER_389_1936 ();
 FILLCELL_X32 FILLER_389_1968 ();
 FILLCELL_X32 FILLER_389_2000 ();
 FILLCELL_X32 FILLER_389_2032 ();
 FILLCELL_X32 FILLER_389_2064 ();
 FILLCELL_X32 FILLER_389_2096 ();
 FILLCELL_X32 FILLER_389_2128 ();
 FILLCELL_X32 FILLER_389_2160 ();
 FILLCELL_X32 FILLER_389_2192 ();
 FILLCELL_X32 FILLER_389_2224 ();
 FILLCELL_X32 FILLER_389_2256 ();
 FILLCELL_X32 FILLER_389_2288 ();
 FILLCELL_X32 FILLER_389_2320 ();
 FILLCELL_X32 FILLER_389_2352 ();
 FILLCELL_X32 FILLER_389_2384 ();
 FILLCELL_X32 FILLER_389_2416 ();
 FILLCELL_X32 FILLER_389_2448 ();
 FILLCELL_X32 FILLER_389_2480 ();
 FILLCELL_X8 FILLER_389_2512 ();
 FILLCELL_X4 FILLER_389_2520 ();
 FILLCELL_X2 FILLER_389_2524 ();
 FILLCELL_X32 FILLER_389_2527 ();
 FILLCELL_X32 FILLER_389_2559 ();
 FILLCELL_X32 FILLER_389_2591 ();
 FILLCELL_X32 FILLER_389_2623 ();
 FILLCELL_X32 FILLER_389_2655 ();
 FILLCELL_X32 FILLER_389_2687 ();
 FILLCELL_X32 FILLER_389_2719 ();
 FILLCELL_X32 FILLER_389_2751 ();
 FILLCELL_X32 FILLER_389_2783 ();
 FILLCELL_X32 FILLER_389_2815 ();
 FILLCELL_X32 FILLER_389_2847 ();
 FILLCELL_X32 FILLER_389_2879 ();
 FILLCELL_X32 FILLER_389_2911 ();
 FILLCELL_X32 FILLER_389_2943 ();
 FILLCELL_X32 FILLER_389_2975 ();
 FILLCELL_X32 FILLER_389_3007 ();
 FILLCELL_X32 FILLER_389_3039 ();
 FILLCELL_X32 FILLER_389_3071 ();
 FILLCELL_X32 FILLER_389_3103 ();
 FILLCELL_X32 FILLER_389_3135 ();
 FILLCELL_X32 FILLER_389_3167 ();
 FILLCELL_X32 FILLER_389_3199 ();
 FILLCELL_X32 FILLER_389_3231 ();
 FILLCELL_X32 FILLER_389_3263 ();
 FILLCELL_X32 FILLER_389_3295 ();
 FILLCELL_X32 FILLER_389_3327 ();
 FILLCELL_X32 FILLER_389_3359 ();
 FILLCELL_X32 FILLER_389_3391 ();
 FILLCELL_X32 FILLER_389_3423 ();
 FILLCELL_X32 FILLER_389_3455 ();
 FILLCELL_X32 FILLER_389_3487 ();
 FILLCELL_X32 FILLER_389_3519 ();
 FILLCELL_X32 FILLER_389_3551 ();
 FILLCELL_X32 FILLER_389_3583 ();
 FILLCELL_X32 FILLER_389_3615 ();
 FILLCELL_X32 FILLER_389_3647 ();
 FILLCELL_X32 FILLER_389_3679 ();
 FILLCELL_X16 FILLER_389_3711 ();
 FILLCELL_X8 FILLER_389_3727 ();
 FILLCELL_X2 FILLER_389_3735 ();
 FILLCELL_X1 FILLER_389_3737 ();
 FILLCELL_X32 FILLER_390_1 ();
 FILLCELL_X32 FILLER_390_33 ();
 FILLCELL_X32 FILLER_390_65 ();
 FILLCELL_X32 FILLER_390_97 ();
 FILLCELL_X32 FILLER_390_129 ();
 FILLCELL_X32 FILLER_390_161 ();
 FILLCELL_X32 FILLER_390_193 ();
 FILLCELL_X32 FILLER_390_225 ();
 FILLCELL_X32 FILLER_390_257 ();
 FILLCELL_X32 FILLER_390_289 ();
 FILLCELL_X32 FILLER_390_321 ();
 FILLCELL_X32 FILLER_390_353 ();
 FILLCELL_X32 FILLER_390_385 ();
 FILLCELL_X32 FILLER_390_417 ();
 FILLCELL_X32 FILLER_390_449 ();
 FILLCELL_X32 FILLER_390_481 ();
 FILLCELL_X32 FILLER_390_513 ();
 FILLCELL_X32 FILLER_390_545 ();
 FILLCELL_X32 FILLER_390_577 ();
 FILLCELL_X16 FILLER_390_609 ();
 FILLCELL_X4 FILLER_390_625 ();
 FILLCELL_X2 FILLER_390_629 ();
 FILLCELL_X32 FILLER_390_632 ();
 FILLCELL_X32 FILLER_390_664 ();
 FILLCELL_X32 FILLER_390_696 ();
 FILLCELL_X32 FILLER_390_728 ();
 FILLCELL_X32 FILLER_390_760 ();
 FILLCELL_X32 FILLER_390_792 ();
 FILLCELL_X32 FILLER_390_824 ();
 FILLCELL_X32 FILLER_390_856 ();
 FILLCELL_X32 FILLER_390_888 ();
 FILLCELL_X32 FILLER_390_920 ();
 FILLCELL_X32 FILLER_390_952 ();
 FILLCELL_X32 FILLER_390_984 ();
 FILLCELL_X32 FILLER_390_1016 ();
 FILLCELL_X32 FILLER_390_1048 ();
 FILLCELL_X32 FILLER_390_1080 ();
 FILLCELL_X32 FILLER_390_1112 ();
 FILLCELL_X32 FILLER_390_1144 ();
 FILLCELL_X32 FILLER_390_1176 ();
 FILLCELL_X32 FILLER_390_1208 ();
 FILLCELL_X32 FILLER_390_1240 ();
 FILLCELL_X32 FILLER_390_1272 ();
 FILLCELL_X32 FILLER_390_1304 ();
 FILLCELL_X32 FILLER_390_1336 ();
 FILLCELL_X32 FILLER_390_1368 ();
 FILLCELL_X32 FILLER_390_1400 ();
 FILLCELL_X32 FILLER_390_1432 ();
 FILLCELL_X32 FILLER_390_1464 ();
 FILLCELL_X32 FILLER_390_1496 ();
 FILLCELL_X32 FILLER_390_1528 ();
 FILLCELL_X32 FILLER_390_1560 ();
 FILLCELL_X32 FILLER_390_1592 ();
 FILLCELL_X32 FILLER_390_1624 ();
 FILLCELL_X32 FILLER_390_1656 ();
 FILLCELL_X32 FILLER_390_1688 ();
 FILLCELL_X32 FILLER_390_1720 ();
 FILLCELL_X32 FILLER_390_1752 ();
 FILLCELL_X32 FILLER_390_1784 ();
 FILLCELL_X32 FILLER_390_1816 ();
 FILLCELL_X32 FILLER_390_1848 ();
 FILLCELL_X8 FILLER_390_1880 ();
 FILLCELL_X4 FILLER_390_1888 ();
 FILLCELL_X2 FILLER_390_1892 ();
 FILLCELL_X32 FILLER_390_1895 ();
 FILLCELL_X32 FILLER_390_1927 ();
 FILLCELL_X32 FILLER_390_1959 ();
 FILLCELL_X32 FILLER_390_1991 ();
 FILLCELL_X32 FILLER_390_2023 ();
 FILLCELL_X32 FILLER_390_2055 ();
 FILLCELL_X32 FILLER_390_2087 ();
 FILLCELL_X32 FILLER_390_2119 ();
 FILLCELL_X32 FILLER_390_2151 ();
 FILLCELL_X32 FILLER_390_2183 ();
 FILLCELL_X32 FILLER_390_2215 ();
 FILLCELL_X32 FILLER_390_2247 ();
 FILLCELL_X32 FILLER_390_2279 ();
 FILLCELL_X32 FILLER_390_2311 ();
 FILLCELL_X32 FILLER_390_2343 ();
 FILLCELL_X32 FILLER_390_2375 ();
 FILLCELL_X32 FILLER_390_2407 ();
 FILLCELL_X32 FILLER_390_2439 ();
 FILLCELL_X32 FILLER_390_2471 ();
 FILLCELL_X32 FILLER_390_2503 ();
 FILLCELL_X32 FILLER_390_2535 ();
 FILLCELL_X32 FILLER_390_2567 ();
 FILLCELL_X32 FILLER_390_2599 ();
 FILLCELL_X32 FILLER_390_2631 ();
 FILLCELL_X32 FILLER_390_2663 ();
 FILLCELL_X32 FILLER_390_2695 ();
 FILLCELL_X32 FILLER_390_2727 ();
 FILLCELL_X32 FILLER_390_2759 ();
 FILLCELL_X32 FILLER_390_2791 ();
 FILLCELL_X32 FILLER_390_2823 ();
 FILLCELL_X32 FILLER_390_2855 ();
 FILLCELL_X32 FILLER_390_2887 ();
 FILLCELL_X32 FILLER_390_2919 ();
 FILLCELL_X32 FILLER_390_2951 ();
 FILLCELL_X32 FILLER_390_2983 ();
 FILLCELL_X32 FILLER_390_3015 ();
 FILLCELL_X32 FILLER_390_3047 ();
 FILLCELL_X32 FILLER_390_3079 ();
 FILLCELL_X32 FILLER_390_3111 ();
 FILLCELL_X8 FILLER_390_3143 ();
 FILLCELL_X4 FILLER_390_3151 ();
 FILLCELL_X2 FILLER_390_3155 ();
 FILLCELL_X32 FILLER_390_3158 ();
 FILLCELL_X32 FILLER_390_3190 ();
 FILLCELL_X32 FILLER_390_3222 ();
 FILLCELL_X32 FILLER_390_3254 ();
 FILLCELL_X32 FILLER_390_3286 ();
 FILLCELL_X32 FILLER_390_3318 ();
 FILLCELL_X32 FILLER_390_3350 ();
 FILLCELL_X32 FILLER_390_3382 ();
 FILLCELL_X32 FILLER_390_3414 ();
 FILLCELL_X32 FILLER_390_3446 ();
 FILLCELL_X32 FILLER_390_3478 ();
 FILLCELL_X32 FILLER_390_3510 ();
 FILLCELL_X32 FILLER_390_3542 ();
 FILLCELL_X32 FILLER_390_3574 ();
 FILLCELL_X32 FILLER_390_3606 ();
 FILLCELL_X32 FILLER_390_3638 ();
 FILLCELL_X32 FILLER_390_3670 ();
 FILLCELL_X32 FILLER_390_3702 ();
 FILLCELL_X4 FILLER_390_3734 ();
 FILLCELL_X32 FILLER_391_1 ();
 FILLCELL_X32 FILLER_391_33 ();
 FILLCELL_X32 FILLER_391_65 ();
 FILLCELL_X32 FILLER_391_97 ();
 FILLCELL_X32 FILLER_391_129 ();
 FILLCELL_X32 FILLER_391_161 ();
 FILLCELL_X32 FILLER_391_193 ();
 FILLCELL_X32 FILLER_391_225 ();
 FILLCELL_X32 FILLER_391_257 ();
 FILLCELL_X32 FILLER_391_289 ();
 FILLCELL_X32 FILLER_391_321 ();
 FILLCELL_X32 FILLER_391_353 ();
 FILLCELL_X32 FILLER_391_385 ();
 FILLCELL_X32 FILLER_391_417 ();
 FILLCELL_X32 FILLER_391_449 ();
 FILLCELL_X32 FILLER_391_481 ();
 FILLCELL_X32 FILLER_391_513 ();
 FILLCELL_X32 FILLER_391_545 ();
 FILLCELL_X32 FILLER_391_577 ();
 FILLCELL_X32 FILLER_391_609 ();
 FILLCELL_X32 FILLER_391_641 ();
 FILLCELL_X32 FILLER_391_673 ();
 FILLCELL_X32 FILLER_391_705 ();
 FILLCELL_X32 FILLER_391_737 ();
 FILLCELL_X32 FILLER_391_769 ();
 FILLCELL_X32 FILLER_391_801 ();
 FILLCELL_X32 FILLER_391_833 ();
 FILLCELL_X32 FILLER_391_865 ();
 FILLCELL_X32 FILLER_391_897 ();
 FILLCELL_X32 FILLER_391_929 ();
 FILLCELL_X32 FILLER_391_961 ();
 FILLCELL_X32 FILLER_391_993 ();
 FILLCELL_X32 FILLER_391_1025 ();
 FILLCELL_X32 FILLER_391_1057 ();
 FILLCELL_X32 FILLER_391_1089 ();
 FILLCELL_X32 FILLER_391_1121 ();
 FILLCELL_X32 FILLER_391_1153 ();
 FILLCELL_X32 FILLER_391_1185 ();
 FILLCELL_X32 FILLER_391_1217 ();
 FILLCELL_X8 FILLER_391_1249 ();
 FILLCELL_X4 FILLER_391_1257 ();
 FILLCELL_X2 FILLER_391_1261 ();
 FILLCELL_X32 FILLER_391_1264 ();
 FILLCELL_X32 FILLER_391_1296 ();
 FILLCELL_X32 FILLER_391_1328 ();
 FILLCELL_X32 FILLER_391_1360 ();
 FILLCELL_X32 FILLER_391_1392 ();
 FILLCELL_X32 FILLER_391_1424 ();
 FILLCELL_X32 FILLER_391_1456 ();
 FILLCELL_X32 FILLER_391_1488 ();
 FILLCELL_X32 FILLER_391_1520 ();
 FILLCELL_X32 FILLER_391_1552 ();
 FILLCELL_X32 FILLER_391_1584 ();
 FILLCELL_X32 FILLER_391_1616 ();
 FILLCELL_X32 FILLER_391_1648 ();
 FILLCELL_X32 FILLER_391_1680 ();
 FILLCELL_X32 FILLER_391_1712 ();
 FILLCELL_X32 FILLER_391_1744 ();
 FILLCELL_X32 FILLER_391_1776 ();
 FILLCELL_X32 FILLER_391_1808 ();
 FILLCELL_X32 FILLER_391_1840 ();
 FILLCELL_X32 FILLER_391_1872 ();
 FILLCELL_X32 FILLER_391_1904 ();
 FILLCELL_X32 FILLER_391_1936 ();
 FILLCELL_X32 FILLER_391_1968 ();
 FILLCELL_X32 FILLER_391_2000 ();
 FILLCELL_X32 FILLER_391_2032 ();
 FILLCELL_X32 FILLER_391_2064 ();
 FILLCELL_X32 FILLER_391_2096 ();
 FILLCELL_X32 FILLER_391_2128 ();
 FILLCELL_X32 FILLER_391_2160 ();
 FILLCELL_X32 FILLER_391_2192 ();
 FILLCELL_X32 FILLER_391_2224 ();
 FILLCELL_X32 FILLER_391_2256 ();
 FILLCELL_X32 FILLER_391_2288 ();
 FILLCELL_X32 FILLER_391_2320 ();
 FILLCELL_X32 FILLER_391_2352 ();
 FILLCELL_X32 FILLER_391_2384 ();
 FILLCELL_X32 FILLER_391_2416 ();
 FILLCELL_X32 FILLER_391_2448 ();
 FILLCELL_X32 FILLER_391_2480 ();
 FILLCELL_X8 FILLER_391_2512 ();
 FILLCELL_X4 FILLER_391_2520 ();
 FILLCELL_X2 FILLER_391_2524 ();
 FILLCELL_X32 FILLER_391_2527 ();
 FILLCELL_X32 FILLER_391_2559 ();
 FILLCELL_X32 FILLER_391_2591 ();
 FILLCELL_X32 FILLER_391_2623 ();
 FILLCELL_X32 FILLER_391_2655 ();
 FILLCELL_X32 FILLER_391_2687 ();
 FILLCELL_X32 FILLER_391_2719 ();
 FILLCELL_X32 FILLER_391_2751 ();
 FILLCELL_X32 FILLER_391_2783 ();
 FILLCELL_X32 FILLER_391_2815 ();
 FILLCELL_X32 FILLER_391_2847 ();
 FILLCELL_X32 FILLER_391_2879 ();
 FILLCELL_X32 FILLER_391_2911 ();
 FILLCELL_X32 FILLER_391_2943 ();
 FILLCELL_X32 FILLER_391_2975 ();
 FILLCELL_X32 FILLER_391_3007 ();
 FILLCELL_X32 FILLER_391_3039 ();
 FILLCELL_X32 FILLER_391_3071 ();
 FILLCELL_X32 FILLER_391_3103 ();
 FILLCELL_X32 FILLER_391_3135 ();
 FILLCELL_X32 FILLER_391_3167 ();
 FILLCELL_X32 FILLER_391_3199 ();
 FILLCELL_X32 FILLER_391_3231 ();
 FILLCELL_X32 FILLER_391_3263 ();
 FILLCELL_X32 FILLER_391_3295 ();
 FILLCELL_X32 FILLER_391_3327 ();
 FILLCELL_X32 FILLER_391_3359 ();
 FILLCELL_X32 FILLER_391_3391 ();
 FILLCELL_X32 FILLER_391_3423 ();
 FILLCELL_X32 FILLER_391_3455 ();
 FILLCELL_X32 FILLER_391_3487 ();
 FILLCELL_X32 FILLER_391_3519 ();
 FILLCELL_X32 FILLER_391_3551 ();
 FILLCELL_X32 FILLER_391_3583 ();
 FILLCELL_X32 FILLER_391_3615 ();
 FILLCELL_X32 FILLER_391_3647 ();
 FILLCELL_X32 FILLER_391_3679 ();
 FILLCELL_X16 FILLER_391_3711 ();
 FILLCELL_X8 FILLER_391_3727 ();
 FILLCELL_X2 FILLER_391_3735 ();
 FILLCELL_X1 FILLER_391_3737 ();
 FILLCELL_X32 FILLER_392_1 ();
 FILLCELL_X32 FILLER_392_33 ();
 FILLCELL_X32 FILLER_392_65 ();
 FILLCELL_X32 FILLER_392_97 ();
 FILLCELL_X32 FILLER_392_129 ();
 FILLCELL_X32 FILLER_392_161 ();
 FILLCELL_X32 FILLER_392_193 ();
 FILLCELL_X32 FILLER_392_225 ();
 FILLCELL_X32 FILLER_392_257 ();
 FILLCELL_X32 FILLER_392_289 ();
 FILLCELL_X32 FILLER_392_321 ();
 FILLCELL_X32 FILLER_392_353 ();
 FILLCELL_X32 FILLER_392_385 ();
 FILLCELL_X32 FILLER_392_417 ();
 FILLCELL_X32 FILLER_392_449 ();
 FILLCELL_X32 FILLER_392_481 ();
 FILLCELL_X32 FILLER_392_513 ();
 FILLCELL_X32 FILLER_392_545 ();
 FILLCELL_X32 FILLER_392_577 ();
 FILLCELL_X16 FILLER_392_609 ();
 FILLCELL_X4 FILLER_392_625 ();
 FILLCELL_X2 FILLER_392_629 ();
 FILLCELL_X32 FILLER_392_632 ();
 FILLCELL_X32 FILLER_392_664 ();
 FILLCELL_X32 FILLER_392_696 ();
 FILLCELL_X32 FILLER_392_728 ();
 FILLCELL_X32 FILLER_392_760 ();
 FILLCELL_X32 FILLER_392_792 ();
 FILLCELL_X32 FILLER_392_824 ();
 FILLCELL_X32 FILLER_392_856 ();
 FILLCELL_X32 FILLER_392_888 ();
 FILLCELL_X32 FILLER_392_920 ();
 FILLCELL_X32 FILLER_392_952 ();
 FILLCELL_X32 FILLER_392_984 ();
 FILLCELL_X32 FILLER_392_1016 ();
 FILLCELL_X32 FILLER_392_1048 ();
 FILLCELL_X32 FILLER_392_1080 ();
 FILLCELL_X32 FILLER_392_1112 ();
 FILLCELL_X32 FILLER_392_1144 ();
 FILLCELL_X32 FILLER_392_1176 ();
 FILLCELL_X32 FILLER_392_1208 ();
 FILLCELL_X32 FILLER_392_1240 ();
 FILLCELL_X32 FILLER_392_1272 ();
 FILLCELL_X32 FILLER_392_1304 ();
 FILLCELL_X32 FILLER_392_1336 ();
 FILLCELL_X32 FILLER_392_1368 ();
 FILLCELL_X32 FILLER_392_1400 ();
 FILLCELL_X32 FILLER_392_1432 ();
 FILLCELL_X32 FILLER_392_1464 ();
 FILLCELL_X32 FILLER_392_1496 ();
 FILLCELL_X32 FILLER_392_1528 ();
 FILLCELL_X32 FILLER_392_1560 ();
 FILLCELL_X32 FILLER_392_1592 ();
 FILLCELL_X32 FILLER_392_1624 ();
 FILLCELL_X32 FILLER_392_1656 ();
 FILLCELL_X32 FILLER_392_1688 ();
 FILLCELL_X32 FILLER_392_1720 ();
 FILLCELL_X32 FILLER_392_1752 ();
 FILLCELL_X32 FILLER_392_1784 ();
 FILLCELL_X32 FILLER_392_1816 ();
 FILLCELL_X32 FILLER_392_1848 ();
 FILLCELL_X8 FILLER_392_1880 ();
 FILLCELL_X4 FILLER_392_1888 ();
 FILLCELL_X2 FILLER_392_1892 ();
 FILLCELL_X32 FILLER_392_1895 ();
 FILLCELL_X32 FILLER_392_1927 ();
 FILLCELL_X32 FILLER_392_1959 ();
 FILLCELL_X32 FILLER_392_1991 ();
 FILLCELL_X32 FILLER_392_2023 ();
 FILLCELL_X32 FILLER_392_2055 ();
 FILLCELL_X32 FILLER_392_2087 ();
 FILLCELL_X32 FILLER_392_2119 ();
 FILLCELL_X32 FILLER_392_2151 ();
 FILLCELL_X32 FILLER_392_2183 ();
 FILLCELL_X32 FILLER_392_2215 ();
 FILLCELL_X32 FILLER_392_2247 ();
 FILLCELL_X32 FILLER_392_2279 ();
 FILLCELL_X32 FILLER_392_2311 ();
 FILLCELL_X32 FILLER_392_2343 ();
 FILLCELL_X32 FILLER_392_2375 ();
 FILLCELL_X32 FILLER_392_2407 ();
 FILLCELL_X32 FILLER_392_2439 ();
 FILLCELL_X32 FILLER_392_2471 ();
 FILLCELL_X32 FILLER_392_2503 ();
 FILLCELL_X32 FILLER_392_2535 ();
 FILLCELL_X32 FILLER_392_2567 ();
 FILLCELL_X32 FILLER_392_2599 ();
 FILLCELL_X32 FILLER_392_2631 ();
 FILLCELL_X32 FILLER_392_2663 ();
 FILLCELL_X32 FILLER_392_2695 ();
 FILLCELL_X32 FILLER_392_2727 ();
 FILLCELL_X32 FILLER_392_2759 ();
 FILLCELL_X32 FILLER_392_2791 ();
 FILLCELL_X32 FILLER_392_2823 ();
 FILLCELL_X32 FILLER_392_2855 ();
 FILLCELL_X32 FILLER_392_2887 ();
 FILLCELL_X32 FILLER_392_2919 ();
 FILLCELL_X32 FILLER_392_2951 ();
 FILLCELL_X32 FILLER_392_2983 ();
 FILLCELL_X32 FILLER_392_3015 ();
 FILLCELL_X32 FILLER_392_3047 ();
 FILLCELL_X32 FILLER_392_3079 ();
 FILLCELL_X32 FILLER_392_3111 ();
 FILLCELL_X8 FILLER_392_3143 ();
 FILLCELL_X4 FILLER_392_3151 ();
 FILLCELL_X2 FILLER_392_3155 ();
 FILLCELL_X32 FILLER_392_3158 ();
 FILLCELL_X32 FILLER_392_3190 ();
 FILLCELL_X32 FILLER_392_3222 ();
 FILLCELL_X32 FILLER_392_3254 ();
 FILLCELL_X32 FILLER_392_3286 ();
 FILLCELL_X32 FILLER_392_3318 ();
 FILLCELL_X32 FILLER_392_3350 ();
 FILLCELL_X32 FILLER_392_3382 ();
 FILLCELL_X32 FILLER_392_3414 ();
 FILLCELL_X32 FILLER_392_3446 ();
 FILLCELL_X32 FILLER_392_3478 ();
 FILLCELL_X32 FILLER_392_3510 ();
 FILLCELL_X32 FILLER_392_3542 ();
 FILLCELL_X32 FILLER_392_3574 ();
 FILLCELL_X32 FILLER_392_3606 ();
 FILLCELL_X32 FILLER_392_3638 ();
 FILLCELL_X32 FILLER_392_3670 ();
 FILLCELL_X32 FILLER_392_3702 ();
 FILLCELL_X4 FILLER_392_3734 ();
 FILLCELL_X32 FILLER_393_1 ();
 FILLCELL_X32 FILLER_393_33 ();
 FILLCELL_X32 FILLER_393_65 ();
 FILLCELL_X32 FILLER_393_97 ();
 FILLCELL_X32 FILLER_393_129 ();
 FILLCELL_X32 FILLER_393_161 ();
 FILLCELL_X32 FILLER_393_193 ();
 FILLCELL_X32 FILLER_393_225 ();
 FILLCELL_X32 FILLER_393_257 ();
 FILLCELL_X32 FILLER_393_289 ();
 FILLCELL_X32 FILLER_393_321 ();
 FILLCELL_X32 FILLER_393_353 ();
 FILLCELL_X32 FILLER_393_385 ();
 FILLCELL_X32 FILLER_393_417 ();
 FILLCELL_X32 FILLER_393_449 ();
 FILLCELL_X32 FILLER_393_481 ();
 FILLCELL_X32 FILLER_393_513 ();
 FILLCELL_X32 FILLER_393_545 ();
 FILLCELL_X32 FILLER_393_577 ();
 FILLCELL_X32 FILLER_393_609 ();
 FILLCELL_X32 FILLER_393_641 ();
 FILLCELL_X32 FILLER_393_673 ();
 FILLCELL_X32 FILLER_393_705 ();
 FILLCELL_X32 FILLER_393_737 ();
 FILLCELL_X32 FILLER_393_769 ();
 FILLCELL_X32 FILLER_393_801 ();
 FILLCELL_X32 FILLER_393_833 ();
 FILLCELL_X32 FILLER_393_865 ();
 FILLCELL_X32 FILLER_393_897 ();
 FILLCELL_X32 FILLER_393_929 ();
 FILLCELL_X32 FILLER_393_961 ();
 FILLCELL_X32 FILLER_393_993 ();
 FILLCELL_X32 FILLER_393_1025 ();
 FILLCELL_X32 FILLER_393_1057 ();
 FILLCELL_X32 FILLER_393_1089 ();
 FILLCELL_X32 FILLER_393_1121 ();
 FILLCELL_X32 FILLER_393_1153 ();
 FILLCELL_X32 FILLER_393_1185 ();
 FILLCELL_X32 FILLER_393_1217 ();
 FILLCELL_X8 FILLER_393_1249 ();
 FILLCELL_X4 FILLER_393_1257 ();
 FILLCELL_X2 FILLER_393_1261 ();
 FILLCELL_X32 FILLER_393_1264 ();
 FILLCELL_X32 FILLER_393_1296 ();
 FILLCELL_X32 FILLER_393_1328 ();
 FILLCELL_X32 FILLER_393_1360 ();
 FILLCELL_X32 FILLER_393_1392 ();
 FILLCELL_X32 FILLER_393_1424 ();
 FILLCELL_X32 FILLER_393_1456 ();
 FILLCELL_X32 FILLER_393_1488 ();
 FILLCELL_X32 FILLER_393_1520 ();
 FILLCELL_X32 FILLER_393_1552 ();
 FILLCELL_X32 FILLER_393_1584 ();
 FILLCELL_X32 FILLER_393_1616 ();
 FILLCELL_X32 FILLER_393_1648 ();
 FILLCELL_X32 FILLER_393_1680 ();
 FILLCELL_X32 FILLER_393_1712 ();
 FILLCELL_X32 FILLER_393_1744 ();
 FILLCELL_X32 FILLER_393_1776 ();
 FILLCELL_X32 FILLER_393_1808 ();
 FILLCELL_X32 FILLER_393_1840 ();
 FILLCELL_X32 FILLER_393_1872 ();
 FILLCELL_X32 FILLER_393_1904 ();
 FILLCELL_X32 FILLER_393_1936 ();
 FILLCELL_X32 FILLER_393_1968 ();
 FILLCELL_X32 FILLER_393_2000 ();
 FILLCELL_X32 FILLER_393_2032 ();
 FILLCELL_X32 FILLER_393_2064 ();
 FILLCELL_X32 FILLER_393_2096 ();
 FILLCELL_X32 FILLER_393_2128 ();
 FILLCELL_X32 FILLER_393_2160 ();
 FILLCELL_X32 FILLER_393_2192 ();
 FILLCELL_X32 FILLER_393_2224 ();
 FILLCELL_X32 FILLER_393_2256 ();
 FILLCELL_X32 FILLER_393_2288 ();
 FILLCELL_X32 FILLER_393_2320 ();
 FILLCELL_X32 FILLER_393_2352 ();
 FILLCELL_X32 FILLER_393_2384 ();
 FILLCELL_X32 FILLER_393_2416 ();
 FILLCELL_X32 FILLER_393_2448 ();
 FILLCELL_X32 FILLER_393_2480 ();
 FILLCELL_X8 FILLER_393_2512 ();
 FILLCELL_X4 FILLER_393_2520 ();
 FILLCELL_X2 FILLER_393_2524 ();
 FILLCELL_X32 FILLER_393_2527 ();
 FILLCELL_X32 FILLER_393_2559 ();
 FILLCELL_X32 FILLER_393_2591 ();
 FILLCELL_X32 FILLER_393_2623 ();
 FILLCELL_X32 FILLER_393_2655 ();
 FILLCELL_X32 FILLER_393_2687 ();
 FILLCELL_X32 FILLER_393_2719 ();
 FILLCELL_X32 FILLER_393_2751 ();
 FILLCELL_X32 FILLER_393_2783 ();
 FILLCELL_X32 FILLER_393_2815 ();
 FILLCELL_X32 FILLER_393_2847 ();
 FILLCELL_X32 FILLER_393_2879 ();
 FILLCELL_X32 FILLER_393_2911 ();
 FILLCELL_X32 FILLER_393_2943 ();
 FILLCELL_X32 FILLER_393_2975 ();
 FILLCELL_X32 FILLER_393_3007 ();
 FILLCELL_X32 FILLER_393_3039 ();
 FILLCELL_X32 FILLER_393_3071 ();
 FILLCELL_X32 FILLER_393_3103 ();
 FILLCELL_X32 FILLER_393_3135 ();
 FILLCELL_X32 FILLER_393_3167 ();
 FILLCELL_X32 FILLER_393_3199 ();
 FILLCELL_X32 FILLER_393_3231 ();
 FILLCELL_X32 FILLER_393_3263 ();
 FILLCELL_X32 FILLER_393_3295 ();
 FILLCELL_X32 FILLER_393_3327 ();
 FILLCELL_X32 FILLER_393_3359 ();
 FILLCELL_X32 FILLER_393_3391 ();
 FILLCELL_X32 FILLER_393_3423 ();
 FILLCELL_X32 FILLER_393_3455 ();
 FILLCELL_X32 FILLER_393_3487 ();
 FILLCELL_X32 FILLER_393_3519 ();
 FILLCELL_X32 FILLER_393_3551 ();
 FILLCELL_X32 FILLER_393_3583 ();
 FILLCELL_X32 FILLER_393_3615 ();
 FILLCELL_X32 FILLER_393_3647 ();
 FILLCELL_X32 FILLER_393_3679 ();
 FILLCELL_X16 FILLER_393_3711 ();
 FILLCELL_X8 FILLER_393_3727 ();
 FILLCELL_X2 FILLER_393_3735 ();
 FILLCELL_X1 FILLER_393_3737 ();
 FILLCELL_X32 FILLER_394_1 ();
 FILLCELL_X32 FILLER_394_33 ();
 FILLCELL_X32 FILLER_394_65 ();
 FILLCELL_X32 FILLER_394_97 ();
 FILLCELL_X32 FILLER_394_129 ();
 FILLCELL_X32 FILLER_394_161 ();
 FILLCELL_X32 FILLER_394_193 ();
 FILLCELL_X32 FILLER_394_225 ();
 FILLCELL_X32 FILLER_394_257 ();
 FILLCELL_X32 FILLER_394_289 ();
 FILLCELL_X32 FILLER_394_321 ();
 FILLCELL_X32 FILLER_394_353 ();
 FILLCELL_X32 FILLER_394_385 ();
 FILLCELL_X32 FILLER_394_417 ();
 FILLCELL_X32 FILLER_394_449 ();
 FILLCELL_X32 FILLER_394_481 ();
 FILLCELL_X32 FILLER_394_513 ();
 FILLCELL_X32 FILLER_394_545 ();
 FILLCELL_X32 FILLER_394_577 ();
 FILLCELL_X16 FILLER_394_609 ();
 FILLCELL_X4 FILLER_394_625 ();
 FILLCELL_X2 FILLER_394_629 ();
 FILLCELL_X32 FILLER_394_632 ();
 FILLCELL_X32 FILLER_394_664 ();
 FILLCELL_X32 FILLER_394_696 ();
 FILLCELL_X32 FILLER_394_728 ();
 FILLCELL_X32 FILLER_394_760 ();
 FILLCELL_X32 FILLER_394_792 ();
 FILLCELL_X32 FILLER_394_824 ();
 FILLCELL_X32 FILLER_394_856 ();
 FILLCELL_X32 FILLER_394_888 ();
 FILLCELL_X32 FILLER_394_920 ();
 FILLCELL_X32 FILLER_394_952 ();
 FILLCELL_X32 FILLER_394_984 ();
 FILLCELL_X32 FILLER_394_1016 ();
 FILLCELL_X32 FILLER_394_1048 ();
 FILLCELL_X32 FILLER_394_1080 ();
 FILLCELL_X32 FILLER_394_1112 ();
 FILLCELL_X32 FILLER_394_1144 ();
 FILLCELL_X32 FILLER_394_1176 ();
 FILLCELL_X32 FILLER_394_1208 ();
 FILLCELL_X32 FILLER_394_1240 ();
 FILLCELL_X32 FILLER_394_1272 ();
 FILLCELL_X32 FILLER_394_1304 ();
 FILLCELL_X32 FILLER_394_1336 ();
 FILLCELL_X32 FILLER_394_1368 ();
 FILLCELL_X32 FILLER_394_1400 ();
 FILLCELL_X32 FILLER_394_1432 ();
 FILLCELL_X32 FILLER_394_1464 ();
 FILLCELL_X32 FILLER_394_1496 ();
 FILLCELL_X32 FILLER_394_1528 ();
 FILLCELL_X32 FILLER_394_1560 ();
 FILLCELL_X32 FILLER_394_1592 ();
 FILLCELL_X32 FILLER_394_1624 ();
 FILLCELL_X32 FILLER_394_1656 ();
 FILLCELL_X32 FILLER_394_1688 ();
 FILLCELL_X32 FILLER_394_1720 ();
 FILLCELL_X32 FILLER_394_1752 ();
 FILLCELL_X32 FILLER_394_1784 ();
 FILLCELL_X32 FILLER_394_1816 ();
 FILLCELL_X32 FILLER_394_1848 ();
 FILLCELL_X8 FILLER_394_1880 ();
 FILLCELL_X4 FILLER_394_1888 ();
 FILLCELL_X2 FILLER_394_1892 ();
 FILLCELL_X32 FILLER_394_1895 ();
 FILLCELL_X32 FILLER_394_1927 ();
 FILLCELL_X32 FILLER_394_1959 ();
 FILLCELL_X32 FILLER_394_1991 ();
 FILLCELL_X32 FILLER_394_2023 ();
 FILLCELL_X32 FILLER_394_2055 ();
 FILLCELL_X32 FILLER_394_2087 ();
 FILLCELL_X32 FILLER_394_2119 ();
 FILLCELL_X32 FILLER_394_2151 ();
 FILLCELL_X32 FILLER_394_2183 ();
 FILLCELL_X32 FILLER_394_2215 ();
 FILLCELL_X32 FILLER_394_2247 ();
 FILLCELL_X32 FILLER_394_2279 ();
 FILLCELL_X32 FILLER_394_2311 ();
 FILLCELL_X32 FILLER_394_2343 ();
 FILLCELL_X32 FILLER_394_2375 ();
 FILLCELL_X32 FILLER_394_2407 ();
 FILLCELL_X32 FILLER_394_2439 ();
 FILLCELL_X32 FILLER_394_2471 ();
 FILLCELL_X32 FILLER_394_2503 ();
 FILLCELL_X32 FILLER_394_2535 ();
 FILLCELL_X32 FILLER_394_2567 ();
 FILLCELL_X32 FILLER_394_2599 ();
 FILLCELL_X32 FILLER_394_2631 ();
 FILLCELL_X32 FILLER_394_2663 ();
 FILLCELL_X32 FILLER_394_2695 ();
 FILLCELL_X32 FILLER_394_2727 ();
 FILLCELL_X32 FILLER_394_2759 ();
 FILLCELL_X32 FILLER_394_2791 ();
 FILLCELL_X32 FILLER_394_2823 ();
 FILLCELL_X32 FILLER_394_2855 ();
 FILLCELL_X32 FILLER_394_2887 ();
 FILLCELL_X32 FILLER_394_2919 ();
 FILLCELL_X32 FILLER_394_2951 ();
 FILLCELL_X32 FILLER_394_2983 ();
 FILLCELL_X32 FILLER_394_3015 ();
 FILLCELL_X32 FILLER_394_3047 ();
 FILLCELL_X32 FILLER_394_3079 ();
 FILLCELL_X32 FILLER_394_3111 ();
 FILLCELL_X8 FILLER_394_3143 ();
 FILLCELL_X4 FILLER_394_3151 ();
 FILLCELL_X2 FILLER_394_3155 ();
 FILLCELL_X32 FILLER_394_3158 ();
 FILLCELL_X32 FILLER_394_3190 ();
 FILLCELL_X32 FILLER_394_3222 ();
 FILLCELL_X32 FILLER_394_3254 ();
 FILLCELL_X32 FILLER_394_3286 ();
 FILLCELL_X32 FILLER_394_3318 ();
 FILLCELL_X32 FILLER_394_3350 ();
 FILLCELL_X32 FILLER_394_3382 ();
 FILLCELL_X32 FILLER_394_3414 ();
 FILLCELL_X32 FILLER_394_3446 ();
 FILLCELL_X32 FILLER_394_3478 ();
 FILLCELL_X32 FILLER_394_3510 ();
 FILLCELL_X32 FILLER_394_3542 ();
 FILLCELL_X32 FILLER_394_3574 ();
 FILLCELL_X32 FILLER_394_3606 ();
 FILLCELL_X32 FILLER_394_3638 ();
 FILLCELL_X32 FILLER_394_3670 ();
 FILLCELL_X32 FILLER_394_3702 ();
 FILLCELL_X4 FILLER_394_3734 ();
 FILLCELL_X32 FILLER_395_1 ();
 FILLCELL_X32 FILLER_395_33 ();
 FILLCELL_X32 FILLER_395_65 ();
 FILLCELL_X32 FILLER_395_97 ();
 FILLCELL_X32 FILLER_395_129 ();
 FILLCELL_X32 FILLER_395_161 ();
 FILLCELL_X32 FILLER_395_193 ();
 FILLCELL_X32 FILLER_395_225 ();
 FILLCELL_X32 FILLER_395_257 ();
 FILLCELL_X32 FILLER_395_289 ();
 FILLCELL_X32 FILLER_395_321 ();
 FILLCELL_X32 FILLER_395_353 ();
 FILLCELL_X32 FILLER_395_385 ();
 FILLCELL_X32 FILLER_395_417 ();
 FILLCELL_X32 FILLER_395_449 ();
 FILLCELL_X32 FILLER_395_481 ();
 FILLCELL_X32 FILLER_395_513 ();
 FILLCELL_X32 FILLER_395_545 ();
 FILLCELL_X32 FILLER_395_577 ();
 FILLCELL_X32 FILLER_395_609 ();
 FILLCELL_X32 FILLER_395_641 ();
 FILLCELL_X32 FILLER_395_673 ();
 FILLCELL_X32 FILLER_395_705 ();
 FILLCELL_X32 FILLER_395_737 ();
 FILLCELL_X32 FILLER_395_769 ();
 FILLCELL_X32 FILLER_395_801 ();
 FILLCELL_X32 FILLER_395_833 ();
 FILLCELL_X32 FILLER_395_865 ();
 FILLCELL_X32 FILLER_395_897 ();
 FILLCELL_X32 FILLER_395_929 ();
 FILLCELL_X32 FILLER_395_961 ();
 FILLCELL_X32 FILLER_395_993 ();
 FILLCELL_X32 FILLER_395_1025 ();
 FILLCELL_X32 FILLER_395_1057 ();
 FILLCELL_X32 FILLER_395_1089 ();
 FILLCELL_X32 FILLER_395_1121 ();
 FILLCELL_X32 FILLER_395_1153 ();
 FILLCELL_X32 FILLER_395_1185 ();
 FILLCELL_X32 FILLER_395_1217 ();
 FILLCELL_X8 FILLER_395_1249 ();
 FILLCELL_X4 FILLER_395_1257 ();
 FILLCELL_X2 FILLER_395_1261 ();
 FILLCELL_X32 FILLER_395_1264 ();
 FILLCELL_X32 FILLER_395_1296 ();
 FILLCELL_X32 FILLER_395_1328 ();
 FILLCELL_X32 FILLER_395_1360 ();
 FILLCELL_X32 FILLER_395_1392 ();
 FILLCELL_X32 FILLER_395_1424 ();
 FILLCELL_X32 FILLER_395_1456 ();
 FILLCELL_X32 FILLER_395_1488 ();
 FILLCELL_X32 FILLER_395_1520 ();
 FILLCELL_X32 FILLER_395_1552 ();
 FILLCELL_X32 FILLER_395_1584 ();
 FILLCELL_X32 FILLER_395_1616 ();
 FILLCELL_X32 FILLER_395_1648 ();
 FILLCELL_X32 FILLER_395_1680 ();
 FILLCELL_X32 FILLER_395_1712 ();
 FILLCELL_X32 FILLER_395_1744 ();
 FILLCELL_X32 FILLER_395_1776 ();
 FILLCELL_X32 FILLER_395_1808 ();
 FILLCELL_X32 FILLER_395_1840 ();
 FILLCELL_X32 FILLER_395_1872 ();
 FILLCELL_X32 FILLER_395_1904 ();
 FILLCELL_X32 FILLER_395_1936 ();
 FILLCELL_X32 FILLER_395_1968 ();
 FILLCELL_X32 FILLER_395_2000 ();
 FILLCELL_X32 FILLER_395_2032 ();
 FILLCELL_X32 FILLER_395_2064 ();
 FILLCELL_X32 FILLER_395_2096 ();
 FILLCELL_X32 FILLER_395_2128 ();
 FILLCELL_X32 FILLER_395_2160 ();
 FILLCELL_X32 FILLER_395_2192 ();
 FILLCELL_X32 FILLER_395_2224 ();
 FILLCELL_X32 FILLER_395_2256 ();
 FILLCELL_X32 FILLER_395_2288 ();
 FILLCELL_X32 FILLER_395_2320 ();
 FILLCELL_X32 FILLER_395_2352 ();
 FILLCELL_X32 FILLER_395_2384 ();
 FILLCELL_X32 FILLER_395_2416 ();
 FILLCELL_X32 FILLER_395_2448 ();
 FILLCELL_X32 FILLER_395_2480 ();
 FILLCELL_X8 FILLER_395_2512 ();
 FILLCELL_X4 FILLER_395_2520 ();
 FILLCELL_X2 FILLER_395_2524 ();
 FILLCELL_X32 FILLER_395_2527 ();
 FILLCELL_X32 FILLER_395_2559 ();
 FILLCELL_X32 FILLER_395_2591 ();
 FILLCELL_X32 FILLER_395_2623 ();
 FILLCELL_X32 FILLER_395_2655 ();
 FILLCELL_X32 FILLER_395_2687 ();
 FILLCELL_X32 FILLER_395_2719 ();
 FILLCELL_X32 FILLER_395_2751 ();
 FILLCELL_X32 FILLER_395_2783 ();
 FILLCELL_X32 FILLER_395_2815 ();
 FILLCELL_X32 FILLER_395_2847 ();
 FILLCELL_X32 FILLER_395_2879 ();
 FILLCELL_X32 FILLER_395_2911 ();
 FILLCELL_X32 FILLER_395_2943 ();
 FILLCELL_X32 FILLER_395_2975 ();
 FILLCELL_X32 FILLER_395_3007 ();
 FILLCELL_X32 FILLER_395_3039 ();
 FILLCELL_X32 FILLER_395_3071 ();
 FILLCELL_X32 FILLER_395_3103 ();
 FILLCELL_X32 FILLER_395_3135 ();
 FILLCELL_X32 FILLER_395_3167 ();
 FILLCELL_X32 FILLER_395_3199 ();
 FILLCELL_X32 FILLER_395_3231 ();
 FILLCELL_X32 FILLER_395_3263 ();
 FILLCELL_X32 FILLER_395_3295 ();
 FILLCELL_X32 FILLER_395_3327 ();
 FILLCELL_X32 FILLER_395_3359 ();
 FILLCELL_X32 FILLER_395_3391 ();
 FILLCELL_X32 FILLER_395_3423 ();
 FILLCELL_X32 FILLER_395_3455 ();
 FILLCELL_X32 FILLER_395_3487 ();
 FILLCELL_X32 FILLER_395_3519 ();
 FILLCELL_X32 FILLER_395_3551 ();
 FILLCELL_X32 FILLER_395_3583 ();
 FILLCELL_X32 FILLER_395_3615 ();
 FILLCELL_X32 FILLER_395_3647 ();
 FILLCELL_X32 FILLER_395_3679 ();
 FILLCELL_X16 FILLER_395_3711 ();
 FILLCELL_X8 FILLER_395_3727 ();
 FILLCELL_X2 FILLER_395_3735 ();
 FILLCELL_X1 FILLER_395_3737 ();
 FILLCELL_X32 FILLER_396_1 ();
 FILLCELL_X32 FILLER_396_33 ();
 FILLCELL_X32 FILLER_396_65 ();
 FILLCELL_X32 FILLER_396_97 ();
 FILLCELL_X32 FILLER_396_129 ();
 FILLCELL_X32 FILLER_396_161 ();
 FILLCELL_X32 FILLER_396_193 ();
 FILLCELL_X32 FILLER_396_225 ();
 FILLCELL_X32 FILLER_396_257 ();
 FILLCELL_X32 FILLER_396_289 ();
 FILLCELL_X32 FILLER_396_321 ();
 FILLCELL_X32 FILLER_396_353 ();
 FILLCELL_X32 FILLER_396_385 ();
 FILLCELL_X32 FILLER_396_417 ();
 FILLCELL_X32 FILLER_396_449 ();
 FILLCELL_X32 FILLER_396_481 ();
 FILLCELL_X32 FILLER_396_513 ();
 FILLCELL_X32 FILLER_396_545 ();
 FILLCELL_X32 FILLER_396_577 ();
 FILLCELL_X16 FILLER_396_609 ();
 FILLCELL_X4 FILLER_396_625 ();
 FILLCELL_X2 FILLER_396_629 ();
 FILLCELL_X32 FILLER_396_632 ();
 FILLCELL_X32 FILLER_396_664 ();
 FILLCELL_X32 FILLER_396_696 ();
 FILLCELL_X32 FILLER_396_728 ();
 FILLCELL_X32 FILLER_396_760 ();
 FILLCELL_X32 FILLER_396_792 ();
 FILLCELL_X32 FILLER_396_824 ();
 FILLCELL_X32 FILLER_396_856 ();
 FILLCELL_X32 FILLER_396_888 ();
 FILLCELL_X32 FILLER_396_920 ();
 FILLCELL_X32 FILLER_396_952 ();
 FILLCELL_X32 FILLER_396_984 ();
 FILLCELL_X32 FILLER_396_1016 ();
 FILLCELL_X32 FILLER_396_1048 ();
 FILLCELL_X32 FILLER_396_1080 ();
 FILLCELL_X32 FILLER_396_1112 ();
 FILLCELL_X32 FILLER_396_1144 ();
 FILLCELL_X32 FILLER_396_1176 ();
 FILLCELL_X32 FILLER_396_1208 ();
 FILLCELL_X32 FILLER_396_1240 ();
 FILLCELL_X32 FILLER_396_1272 ();
 FILLCELL_X32 FILLER_396_1304 ();
 FILLCELL_X32 FILLER_396_1336 ();
 FILLCELL_X32 FILLER_396_1368 ();
 FILLCELL_X32 FILLER_396_1400 ();
 FILLCELL_X32 FILLER_396_1432 ();
 FILLCELL_X32 FILLER_396_1464 ();
 FILLCELL_X32 FILLER_396_1496 ();
 FILLCELL_X32 FILLER_396_1528 ();
 FILLCELL_X32 FILLER_396_1560 ();
 FILLCELL_X32 FILLER_396_1592 ();
 FILLCELL_X32 FILLER_396_1624 ();
 FILLCELL_X32 FILLER_396_1656 ();
 FILLCELL_X32 FILLER_396_1688 ();
 FILLCELL_X32 FILLER_396_1720 ();
 FILLCELL_X32 FILLER_396_1752 ();
 FILLCELL_X32 FILLER_396_1784 ();
 FILLCELL_X32 FILLER_396_1816 ();
 FILLCELL_X32 FILLER_396_1848 ();
 FILLCELL_X8 FILLER_396_1880 ();
 FILLCELL_X4 FILLER_396_1888 ();
 FILLCELL_X2 FILLER_396_1892 ();
 FILLCELL_X32 FILLER_396_1895 ();
 FILLCELL_X32 FILLER_396_1927 ();
 FILLCELL_X32 FILLER_396_1959 ();
 FILLCELL_X32 FILLER_396_1991 ();
 FILLCELL_X32 FILLER_396_2023 ();
 FILLCELL_X32 FILLER_396_2055 ();
 FILLCELL_X32 FILLER_396_2087 ();
 FILLCELL_X32 FILLER_396_2119 ();
 FILLCELL_X32 FILLER_396_2151 ();
 FILLCELL_X32 FILLER_396_2183 ();
 FILLCELL_X32 FILLER_396_2215 ();
 FILLCELL_X32 FILLER_396_2247 ();
 FILLCELL_X32 FILLER_396_2279 ();
 FILLCELL_X32 FILLER_396_2311 ();
 FILLCELL_X32 FILLER_396_2343 ();
 FILLCELL_X32 FILLER_396_2375 ();
 FILLCELL_X32 FILLER_396_2407 ();
 FILLCELL_X32 FILLER_396_2439 ();
 FILLCELL_X32 FILLER_396_2471 ();
 FILLCELL_X32 FILLER_396_2503 ();
 FILLCELL_X32 FILLER_396_2535 ();
 FILLCELL_X32 FILLER_396_2567 ();
 FILLCELL_X32 FILLER_396_2599 ();
 FILLCELL_X32 FILLER_396_2631 ();
 FILLCELL_X32 FILLER_396_2663 ();
 FILLCELL_X32 FILLER_396_2695 ();
 FILLCELL_X32 FILLER_396_2727 ();
 FILLCELL_X32 FILLER_396_2759 ();
 FILLCELL_X32 FILLER_396_2791 ();
 FILLCELL_X32 FILLER_396_2823 ();
 FILLCELL_X32 FILLER_396_2855 ();
 FILLCELL_X32 FILLER_396_2887 ();
 FILLCELL_X32 FILLER_396_2919 ();
 FILLCELL_X32 FILLER_396_2951 ();
 FILLCELL_X32 FILLER_396_2983 ();
 FILLCELL_X32 FILLER_396_3015 ();
 FILLCELL_X32 FILLER_396_3047 ();
 FILLCELL_X32 FILLER_396_3079 ();
 FILLCELL_X32 FILLER_396_3111 ();
 FILLCELL_X8 FILLER_396_3143 ();
 FILLCELL_X4 FILLER_396_3151 ();
 FILLCELL_X2 FILLER_396_3155 ();
 FILLCELL_X32 FILLER_396_3158 ();
 FILLCELL_X32 FILLER_396_3190 ();
 FILLCELL_X32 FILLER_396_3222 ();
 FILLCELL_X32 FILLER_396_3254 ();
 FILLCELL_X32 FILLER_396_3286 ();
 FILLCELL_X32 FILLER_396_3318 ();
 FILLCELL_X32 FILLER_396_3350 ();
 FILLCELL_X32 FILLER_396_3382 ();
 FILLCELL_X32 FILLER_396_3414 ();
 FILLCELL_X32 FILLER_396_3446 ();
 FILLCELL_X32 FILLER_396_3478 ();
 FILLCELL_X32 FILLER_396_3510 ();
 FILLCELL_X32 FILLER_396_3542 ();
 FILLCELL_X32 FILLER_396_3574 ();
 FILLCELL_X32 FILLER_396_3606 ();
 FILLCELL_X32 FILLER_396_3638 ();
 FILLCELL_X32 FILLER_396_3670 ();
 FILLCELL_X32 FILLER_396_3702 ();
 FILLCELL_X4 FILLER_396_3734 ();
 FILLCELL_X32 FILLER_397_1 ();
 FILLCELL_X32 FILLER_397_33 ();
 FILLCELL_X32 FILLER_397_65 ();
 FILLCELL_X32 FILLER_397_97 ();
 FILLCELL_X32 FILLER_397_129 ();
 FILLCELL_X32 FILLER_397_161 ();
 FILLCELL_X32 FILLER_397_193 ();
 FILLCELL_X32 FILLER_397_225 ();
 FILLCELL_X32 FILLER_397_257 ();
 FILLCELL_X32 FILLER_397_289 ();
 FILLCELL_X32 FILLER_397_321 ();
 FILLCELL_X32 FILLER_397_353 ();
 FILLCELL_X32 FILLER_397_385 ();
 FILLCELL_X32 FILLER_397_417 ();
 FILLCELL_X32 FILLER_397_449 ();
 FILLCELL_X32 FILLER_397_481 ();
 FILLCELL_X32 FILLER_397_513 ();
 FILLCELL_X32 FILLER_397_545 ();
 FILLCELL_X32 FILLER_397_577 ();
 FILLCELL_X32 FILLER_397_609 ();
 FILLCELL_X32 FILLER_397_641 ();
 FILLCELL_X32 FILLER_397_673 ();
 FILLCELL_X32 FILLER_397_705 ();
 FILLCELL_X32 FILLER_397_737 ();
 FILLCELL_X32 FILLER_397_769 ();
 FILLCELL_X32 FILLER_397_801 ();
 FILLCELL_X32 FILLER_397_833 ();
 FILLCELL_X32 FILLER_397_865 ();
 FILLCELL_X32 FILLER_397_897 ();
 FILLCELL_X32 FILLER_397_929 ();
 FILLCELL_X32 FILLER_397_961 ();
 FILLCELL_X32 FILLER_397_993 ();
 FILLCELL_X32 FILLER_397_1025 ();
 FILLCELL_X32 FILLER_397_1057 ();
 FILLCELL_X32 FILLER_397_1089 ();
 FILLCELL_X32 FILLER_397_1121 ();
 FILLCELL_X32 FILLER_397_1153 ();
 FILLCELL_X32 FILLER_397_1185 ();
 FILLCELL_X32 FILLER_397_1217 ();
 FILLCELL_X8 FILLER_397_1249 ();
 FILLCELL_X4 FILLER_397_1257 ();
 FILLCELL_X2 FILLER_397_1261 ();
 FILLCELL_X32 FILLER_397_1264 ();
 FILLCELL_X32 FILLER_397_1296 ();
 FILLCELL_X32 FILLER_397_1328 ();
 FILLCELL_X32 FILLER_397_1360 ();
 FILLCELL_X32 FILLER_397_1392 ();
 FILLCELL_X32 FILLER_397_1424 ();
 FILLCELL_X32 FILLER_397_1456 ();
 FILLCELL_X32 FILLER_397_1488 ();
 FILLCELL_X32 FILLER_397_1520 ();
 FILLCELL_X32 FILLER_397_1552 ();
 FILLCELL_X32 FILLER_397_1584 ();
 FILLCELL_X32 FILLER_397_1616 ();
 FILLCELL_X32 FILLER_397_1648 ();
 FILLCELL_X32 FILLER_397_1680 ();
 FILLCELL_X32 FILLER_397_1712 ();
 FILLCELL_X32 FILLER_397_1744 ();
 FILLCELL_X32 FILLER_397_1776 ();
 FILLCELL_X32 FILLER_397_1808 ();
 FILLCELL_X32 FILLER_397_1840 ();
 FILLCELL_X32 FILLER_397_1872 ();
 FILLCELL_X32 FILLER_397_1904 ();
 FILLCELL_X32 FILLER_397_1936 ();
 FILLCELL_X32 FILLER_397_1968 ();
 FILLCELL_X32 FILLER_397_2000 ();
 FILLCELL_X32 FILLER_397_2032 ();
 FILLCELL_X32 FILLER_397_2064 ();
 FILLCELL_X32 FILLER_397_2096 ();
 FILLCELL_X32 FILLER_397_2128 ();
 FILLCELL_X32 FILLER_397_2160 ();
 FILLCELL_X32 FILLER_397_2192 ();
 FILLCELL_X32 FILLER_397_2224 ();
 FILLCELL_X32 FILLER_397_2256 ();
 FILLCELL_X32 FILLER_397_2288 ();
 FILLCELL_X32 FILLER_397_2320 ();
 FILLCELL_X32 FILLER_397_2352 ();
 FILLCELL_X32 FILLER_397_2384 ();
 FILLCELL_X32 FILLER_397_2416 ();
 FILLCELL_X32 FILLER_397_2448 ();
 FILLCELL_X32 FILLER_397_2480 ();
 FILLCELL_X8 FILLER_397_2512 ();
 FILLCELL_X4 FILLER_397_2520 ();
 FILLCELL_X2 FILLER_397_2524 ();
 FILLCELL_X32 FILLER_397_2527 ();
 FILLCELL_X32 FILLER_397_2559 ();
 FILLCELL_X32 FILLER_397_2591 ();
 FILLCELL_X32 FILLER_397_2623 ();
 FILLCELL_X32 FILLER_397_2655 ();
 FILLCELL_X32 FILLER_397_2687 ();
 FILLCELL_X32 FILLER_397_2719 ();
 FILLCELL_X32 FILLER_397_2751 ();
 FILLCELL_X32 FILLER_397_2783 ();
 FILLCELL_X32 FILLER_397_2815 ();
 FILLCELL_X32 FILLER_397_2847 ();
 FILLCELL_X32 FILLER_397_2879 ();
 FILLCELL_X32 FILLER_397_2911 ();
 FILLCELL_X32 FILLER_397_2943 ();
 FILLCELL_X32 FILLER_397_2975 ();
 FILLCELL_X32 FILLER_397_3007 ();
 FILLCELL_X32 FILLER_397_3039 ();
 FILLCELL_X32 FILLER_397_3071 ();
 FILLCELL_X32 FILLER_397_3103 ();
 FILLCELL_X32 FILLER_397_3135 ();
 FILLCELL_X32 FILLER_397_3167 ();
 FILLCELL_X32 FILLER_397_3199 ();
 FILLCELL_X32 FILLER_397_3231 ();
 FILLCELL_X32 FILLER_397_3263 ();
 FILLCELL_X32 FILLER_397_3295 ();
 FILLCELL_X32 FILLER_397_3327 ();
 FILLCELL_X32 FILLER_397_3359 ();
 FILLCELL_X32 FILLER_397_3391 ();
 FILLCELL_X32 FILLER_397_3423 ();
 FILLCELL_X32 FILLER_397_3455 ();
 FILLCELL_X32 FILLER_397_3487 ();
 FILLCELL_X32 FILLER_397_3519 ();
 FILLCELL_X32 FILLER_397_3551 ();
 FILLCELL_X32 FILLER_397_3583 ();
 FILLCELL_X32 FILLER_397_3615 ();
 FILLCELL_X32 FILLER_397_3647 ();
 FILLCELL_X32 FILLER_397_3679 ();
 FILLCELL_X16 FILLER_397_3711 ();
 FILLCELL_X8 FILLER_397_3727 ();
 FILLCELL_X2 FILLER_397_3735 ();
 FILLCELL_X1 FILLER_397_3737 ();
 FILLCELL_X32 FILLER_398_1 ();
 FILLCELL_X32 FILLER_398_33 ();
 FILLCELL_X32 FILLER_398_65 ();
 FILLCELL_X32 FILLER_398_97 ();
 FILLCELL_X32 FILLER_398_129 ();
 FILLCELL_X32 FILLER_398_161 ();
 FILLCELL_X32 FILLER_398_193 ();
 FILLCELL_X32 FILLER_398_225 ();
 FILLCELL_X32 FILLER_398_257 ();
 FILLCELL_X32 FILLER_398_289 ();
 FILLCELL_X32 FILLER_398_321 ();
 FILLCELL_X32 FILLER_398_353 ();
 FILLCELL_X32 FILLER_398_385 ();
 FILLCELL_X32 FILLER_398_417 ();
 FILLCELL_X32 FILLER_398_449 ();
 FILLCELL_X32 FILLER_398_481 ();
 FILLCELL_X32 FILLER_398_513 ();
 FILLCELL_X32 FILLER_398_545 ();
 FILLCELL_X32 FILLER_398_577 ();
 FILLCELL_X16 FILLER_398_609 ();
 FILLCELL_X4 FILLER_398_625 ();
 FILLCELL_X2 FILLER_398_629 ();
 FILLCELL_X32 FILLER_398_632 ();
 FILLCELL_X32 FILLER_398_664 ();
 FILLCELL_X32 FILLER_398_696 ();
 FILLCELL_X32 FILLER_398_728 ();
 FILLCELL_X32 FILLER_398_760 ();
 FILLCELL_X32 FILLER_398_792 ();
 FILLCELL_X32 FILLER_398_824 ();
 FILLCELL_X32 FILLER_398_856 ();
 FILLCELL_X32 FILLER_398_888 ();
 FILLCELL_X32 FILLER_398_920 ();
 FILLCELL_X32 FILLER_398_952 ();
 FILLCELL_X32 FILLER_398_984 ();
 FILLCELL_X32 FILLER_398_1016 ();
 FILLCELL_X32 FILLER_398_1048 ();
 FILLCELL_X32 FILLER_398_1080 ();
 FILLCELL_X32 FILLER_398_1112 ();
 FILLCELL_X32 FILLER_398_1144 ();
 FILLCELL_X32 FILLER_398_1176 ();
 FILLCELL_X32 FILLER_398_1208 ();
 FILLCELL_X32 FILLER_398_1240 ();
 FILLCELL_X32 FILLER_398_1272 ();
 FILLCELL_X32 FILLER_398_1304 ();
 FILLCELL_X32 FILLER_398_1336 ();
 FILLCELL_X32 FILLER_398_1368 ();
 FILLCELL_X32 FILLER_398_1400 ();
 FILLCELL_X32 FILLER_398_1432 ();
 FILLCELL_X32 FILLER_398_1464 ();
 FILLCELL_X32 FILLER_398_1496 ();
 FILLCELL_X32 FILLER_398_1528 ();
 FILLCELL_X32 FILLER_398_1560 ();
 FILLCELL_X32 FILLER_398_1592 ();
 FILLCELL_X32 FILLER_398_1624 ();
 FILLCELL_X32 FILLER_398_1656 ();
 FILLCELL_X32 FILLER_398_1688 ();
 FILLCELL_X32 FILLER_398_1720 ();
 FILLCELL_X32 FILLER_398_1752 ();
 FILLCELL_X32 FILLER_398_1784 ();
 FILLCELL_X32 FILLER_398_1816 ();
 FILLCELL_X32 FILLER_398_1848 ();
 FILLCELL_X8 FILLER_398_1880 ();
 FILLCELL_X4 FILLER_398_1888 ();
 FILLCELL_X2 FILLER_398_1892 ();
 FILLCELL_X32 FILLER_398_1895 ();
 FILLCELL_X32 FILLER_398_1927 ();
 FILLCELL_X32 FILLER_398_1959 ();
 FILLCELL_X32 FILLER_398_1991 ();
 FILLCELL_X32 FILLER_398_2023 ();
 FILLCELL_X32 FILLER_398_2055 ();
 FILLCELL_X32 FILLER_398_2087 ();
 FILLCELL_X32 FILLER_398_2119 ();
 FILLCELL_X32 FILLER_398_2151 ();
 FILLCELL_X32 FILLER_398_2183 ();
 FILLCELL_X32 FILLER_398_2215 ();
 FILLCELL_X32 FILLER_398_2247 ();
 FILLCELL_X32 FILLER_398_2279 ();
 FILLCELL_X32 FILLER_398_2311 ();
 FILLCELL_X32 FILLER_398_2343 ();
 FILLCELL_X32 FILLER_398_2375 ();
 FILLCELL_X32 FILLER_398_2407 ();
 FILLCELL_X32 FILLER_398_2439 ();
 FILLCELL_X32 FILLER_398_2471 ();
 FILLCELL_X32 FILLER_398_2503 ();
 FILLCELL_X32 FILLER_398_2535 ();
 FILLCELL_X32 FILLER_398_2567 ();
 FILLCELL_X32 FILLER_398_2599 ();
 FILLCELL_X32 FILLER_398_2631 ();
 FILLCELL_X32 FILLER_398_2663 ();
 FILLCELL_X32 FILLER_398_2695 ();
 FILLCELL_X32 FILLER_398_2727 ();
 FILLCELL_X32 FILLER_398_2759 ();
 FILLCELL_X32 FILLER_398_2791 ();
 FILLCELL_X32 FILLER_398_2823 ();
 FILLCELL_X32 FILLER_398_2855 ();
 FILLCELL_X32 FILLER_398_2887 ();
 FILLCELL_X32 FILLER_398_2919 ();
 FILLCELL_X32 FILLER_398_2951 ();
 FILLCELL_X32 FILLER_398_2983 ();
 FILLCELL_X32 FILLER_398_3015 ();
 FILLCELL_X32 FILLER_398_3047 ();
 FILLCELL_X32 FILLER_398_3079 ();
 FILLCELL_X32 FILLER_398_3111 ();
 FILLCELL_X8 FILLER_398_3143 ();
 FILLCELL_X4 FILLER_398_3151 ();
 FILLCELL_X2 FILLER_398_3155 ();
 FILLCELL_X32 FILLER_398_3158 ();
 FILLCELL_X32 FILLER_398_3190 ();
 FILLCELL_X32 FILLER_398_3222 ();
 FILLCELL_X32 FILLER_398_3254 ();
 FILLCELL_X32 FILLER_398_3286 ();
 FILLCELL_X32 FILLER_398_3318 ();
 FILLCELL_X32 FILLER_398_3350 ();
 FILLCELL_X32 FILLER_398_3382 ();
 FILLCELL_X32 FILLER_398_3414 ();
 FILLCELL_X32 FILLER_398_3446 ();
 FILLCELL_X32 FILLER_398_3478 ();
 FILLCELL_X32 FILLER_398_3510 ();
 FILLCELL_X32 FILLER_398_3542 ();
 FILLCELL_X32 FILLER_398_3574 ();
 FILLCELL_X32 FILLER_398_3606 ();
 FILLCELL_X32 FILLER_398_3638 ();
 FILLCELL_X32 FILLER_398_3670 ();
 FILLCELL_X32 FILLER_398_3702 ();
 FILLCELL_X4 FILLER_398_3734 ();
 FILLCELL_X32 FILLER_399_1 ();
 FILLCELL_X32 FILLER_399_33 ();
 FILLCELL_X32 FILLER_399_65 ();
 FILLCELL_X32 FILLER_399_97 ();
 FILLCELL_X32 FILLER_399_129 ();
 FILLCELL_X32 FILLER_399_161 ();
 FILLCELL_X32 FILLER_399_193 ();
 FILLCELL_X32 FILLER_399_225 ();
 FILLCELL_X32 FILLER_399_257 ();
 FILLCELL_X32 FILLER_399_289 ();
 FILLCELL_X32 FILLER_399_321 ();
 FILLCELL_X32 FILLER_399_353 ();
 FILLCELL_X32 FILLER_399_385 ();
 FILLCELL_X32 FILLER_399_417 ();
 FILLCELL_X32 FILLER_399_449 ();
 FILLCELL_X32 FILLER_399_481 ();
 FILLCELL_X32 FILLER_399_513 ();
 FILLCELL_X32 FILLER_399_545 ();
 FILLCELL_X32 FILLER_399_577 ();
 FILLCELL_X32 FILLER_399_609 ();
 FILLCELL_X32 FILLER_399_641 ();
 FILLCELL_X32 FILLER_399_673 ();
 FILLCELL_X32 FILLER_399_705 ();
 FILLCELL_X32 FILLER_399_737 ();
 FILLCELL_X32 FILLER_399_769 ();
 FILLCELL_X32 FILLER_399_801 ();
 FILLCELL_X32 FILLER_399_833 ();
 FILLCELL_X32 FILLER_399_865 ();
 FILLCELL_X32 FILLER_399_897 ();
 FILLCELL_X32 FILLER_399_929 ();
 FILLCELL_X32 FILLER_399_961 ();
 FILLCELL_X32 FILLER_399_993 ();
 FILLCELL_X32 FILLER_399_1025 ();
 FILLCELL_X32 FILLER_399_1057 ();
 FILLCELL_X32 FILLER_399_1089 ();
 FILLCELL_X32 FILLER_399_1121 ();
 FILLCELL_X32 FILLER_399_1153 ();
 FILLCELL_X32 FILLER_399_1185 ();
 FILLCELL_X32 FILLER_399_1217 ();
 FILLCELL_X8 FILLER_399_1249 ();
 FILLCELL_X4 FILLER_399_1257 ();
 FILLCELL_X2 FILLER_399_1261 ();
 FILLCELL_X32 FILLER_399_1264 ();
 FILLCELL_X32 FILLER_399_1296 ();
 FILLCELL_X32 FILLER_399_1328 ();
 FILLCELL_X32 FILLER_399_1360 ();
 FILLCELL_X32 FILLER_399_1392 ();
 FILLCELL_X32 FILLER_399_1424 ();
 FILLCELL_X32 FILLER_399_1456 ();
 FILLCELL_X32 FILLER_399_1488 ();
 FILLCELL_X32 FILLER_399_1520 ();
 FILLCELL_X32 FILLER_399_1552 ();
 FILLCELL_X32 FILLER_399_1584 ();
 FILLCELL_X32 FILLER_399_1616 ();
 FILLCELL_X32 FILLER_399_1648 ();
 FILLCELL_X32 FILLER_399_1680 ();
 FILLCELL_X32 FILLER_399_1712 ();
 FILLCELL_X32 FILLER_399_1744 ();
 FILLCELL_X32 FILLER_399_1776 ();
 FILLCELL_X32 FILLER_399_1808 ();
 FILLCELL_X32 FILLER_399_1840 ();
 FILLCELL_X32 FILLER_399_1872 ();
 FILLCELL_X32 FILLER_399_1904 ();
 FILLCELL_X32 FILLER_399_1936 ();
 FILLCELL_X32 FILLER_399_1968 ();
 FILLCELL_X32 FILLER_399_2000 ();
 FILLCELL_X32 FILLER_399_2032 ();
 FILLCELL_X32 FILLER_399_2064 ();
 FILLCELL_X32 FILLER_399_2096 ();
 FILLCELL_X32 FILLER_399_2128 ();
 FILLCELL_X32 FILLER_399_2160 ();
 FILLCELL_X32 FILLER_399_2192 ();
 FILLCELL_X32 FILLER_399_2224 ();
 FILLCELL_X32 FILLER_399_2256 ();
 FILLCELL_X32 FILLER_399_2288 ();
 FILLCELL_X32 FILLER_399_2320 ();
 FILLCELL_X32 FILLER_399_2352 ();
 FILLCELL_X32 FILLER_399_2384 ();
 FILLCELL_X32 FILLER_399_2416 ();
 FILLCELL_X32 FILLER_399_2448 ();
 FILLCELL_X32 FILLER_399_2480 ();
 FILLCELL_X8 FILLER_399_2512 ();
 FILLCELL_X4 FILLER_399_2520 ();
 FILLCELL_X2 FILLER_399_2524 ();
 FILLCELL_X32 FILLER_399_2527 ();
 FILLCELL_X32 FILLER_399_2559 ();
 FILLCELL_X32 FILLER_399_2591 ();
 FILLCELL_X32 FILLER_399_2623 ();
 FILLCELL_X32 FILLER_399_2655 ();
 FILLCELL_X32 FILLER_399_2687 ();
 FILLCELL_X32 FILLER_399_2719 ();
 FILLCELL_X32 FILLER_399_2751 ();
 FILLCELL_X32 FILLER_399_2783 ();
 FILLCELL_X32 FILLER_399_2815 ();
 FILLCELL_X32 FILLER_399_2847 ();
 FILLCELL_X32 FILLER_399_2879 ();
 FILLCELL_X32 FILLER_399_2911 ();
 FILLCELL_X32 FILLER_399_2943 ();
 FILLCELL_X32 FILLER_399_2975 ();
 FILLCELL_X32 FILLER_399_3007 ();
 FILLCELL_X32 FILLER_399_3039 ();
 FILLCELL_X32 FILLER_399_3071 ();
 FILLCELL_X32 FILLER_399_3103 ();
 FILLCELL_X32 FILLER_399_3135 ();
 FILLCELL_X32 FILLER_399_3167 ();
 FILLCELL_X32 FILLER_399_3199 ();
 FILLCELL_X32 FILLER_399_3231 ();
 FILLCELL_X32 FILLER_399_3263 ();
 FILLCELL_X32 FILLER_399_3295 ();
 FILLCELL_X32 FILLER_399_3327 ();
 FILLCELL_X32 FILLER_399_3359 ();
 FILLCELL_X32 FILLER_399_3391 ();
 FILLCELL_X32 FILLER_399_3423 ();
 FILLCELL_X32 FILLER_399_3455 ();
 FILLCELL_X32 FILLER_399_3487 ();
 FILLCELL_X32 FILLER_399_3519 ();
 FILLCELL_X32 FILLER_399_3551 ();
 FILLCELL_X32 FILLER_399_3583 ();
 FILLCELL_X32 FILLER_399_3615 ();
 FILLCELL_X32 FILLER_399_3647 ();
 FILLCELL_X32 FILLER_399_3679 ();
 FILLCELL_X16 FILLER_399_3711 ();
 FILLCELL_X8 FILLER_399_3727 ();
 FILLCELL_X2 FILLER_399_3735 ();
 FILLCELL_X1 FILLER_399_3737 ();
 FILLCELL_X32 FILLER_400_1 ();
 FILLCELL_X32 FILLER_400_33 ();
 FILLCELL_X32 FILLER_400_65 ();
 FILLCELL_X32 FILLER_400_97 ();
 FILLCELL_X32 FILLER_400_129 ();
 FILLCELL_X32 FILLER_400_161 ();
 FILLCELL_X32 FILLER_400_193 ();
 FILLCELL_X32 FILLER_400_225 ();
 FILLCELL_X32 FILLER_400_257 ();
 FILLCELL_X32 FILLER_400_289 ();
 FILLCELL_X32 FILLER_400_321 ();
 FILLCELL_X32 FILLER_400_353 ();
 FILLCELL_X32 FILLER_400_385 ();
 FILLCELL_X32 FILLER_400_417 ();
 FILLCELL_X32 FILLER_400_449 ();
 FILLCELL_X32 FILLER_400_481 ();
 FILLCELL_X32 FILLER_400_513 ();
 FILLCELL_X32 FILLER_400_545 ();
 FILLCELL_X32 FILLER_400_577 ();
 FILLCELL_X16 FILLER_400_609 ();
 FILLCELL_X4 FILLER_400_625 ();
 FILLCELL_X2 FILLER_400_629 ();
 FILLCELL_X32 FILLER_400_632 ();
 FILLCELL_X32 FILLER_400_664 ();
 FILLCELL_X32 FILLER_400_696 ();
 FILLCELL_X32 FILLER_400_728 ();
 FILLCELL_X32 FILLER_400_760 ();
 FILLCELL_X32 FILLER_400_792 ();
 FILLCELL_X32 FILLER_400_824 ();
 FILLCELL_X32 FILLER_400_856 ();
 FILLCELL_X32 FILLER_400_888 ();
 FILLCELL_X32 FILLER_400_920 ();
 FILLCELL_X32 FILLER_400_952 ();
 FILLCELL_X32 FILLER_400_984 ();
 FILLCELL_X32 FILLER_400_1016 ();
 FILLCELL_X32 FILLER_400_1048 ();
 FILLCELL_X32 FILLER_400_1080 ();
 FILLCELL_X32 FILLER_400_1112 ();
 FILLCELL_X32 FILLER_400_1144 ();
 FILLCELL_X32 FILLER_400_1176 ();
 FILLCELL_X32 FILLER_400_1208 ();
 FILLCELL_X32 FILLER_400_1240 ();
 FILLCELL_X32 FILLER_400_1272 ();
 FILLCELL_X32 FILLER_400_1304 ();
 FILLCELL_X32 FILLER_400_1336 ();
 FILLCELL_X32 FILLER_400_1368 ();
 FILLCELL_X32 FILLER_400_1400 ();
 FILLCELL_X32 FILLER_400_1432 ();
 FILLCELL_X32 FILLER_400_1464 ();
 FILLCELL_X32 FILLER_400_1496 ();
 FILLCELL_X32 FILLER_400_1528 ();
 FILLCELL_X32 FILLER_400_1560 ();
 FILLCELL_X32 FILLER_400_1592 ();
 FILLCELL_X32 FILLER_400_1624 ();
 FILLCELL_X32 FILLER_400_1656 ();
 FILLCELL_X32 FILLER_400_1688 ();
 FILLCELL_X32 FILLER_400_1720 ();
 FILLCELL_X32 FILLER_400_1752 ();
 FILLCELL_X32 FILLER_400_1784 ();
 FILLCELL_X32 FILLER_400_1816 ();
 FILLCELL_X32 FILLER_400_1848 ();
 FILLCELL_X8 FILLER_400_1880 ();
 FILLCELL_X4 FILLER_400_1888 ();
 FILLCELL_X2 FILLER_400_1892 ();
 FILLCELL_X32 FILLER_400_1895 ();
 FILLCELL_X32 FILLER_400_1927 ();
 FILLCELL_X32 FILLER_400_1959 ();
 FILLCELL_X32 FILLER_400_1991 ();
 FILLCELL_X32 FILLER_400_2023 ();
 FILLCELL_X32 FILLER_400_2055 ();
 FILLCELL_X32 FILLER_400_2087 ();
 FILLCELL_X32 FILLER_400_2119 ();
 FILLCELL_X32 FILLER_400_2151 ();
 FILLCELL_X32 FILLER_400_2183 ();
 FILLCELL_X32 FILLER_400_2215 ();
 FILLCELL_X32 FILLER_400_2247 ();
 FILLCELL_X32 FILLER_400_2279 ();
 FILLCELL_X32 FILLER_400_2311 ();
 FILLCELL_X32 FILLER_400_2343 ();
 FILLCELL_X32 FILLER_400_2375 ();
 FILLCELL_X32 FILLER_400_2407 ();
 FILLCELL_X32 FILLER_400_2439 ();
 FILLCELL_X32 FILLER_400_2471 ();
 FILLCELL_X32 FILLER_400_2503 ();
 FILLCELL_X32 FILLER_400_2535 ();
 FILLCELL_X32 FILLER_400_2567 ();
 FILLCELL_X32 FILLER_400_2599 ();
 FILLCELL_X32 FILLER_400_2631 ();
 FILLCELL_X32 FILLER_400_2663 ();
 FILLCELL_X32 FILLER_400_2695 ();
 FILLCELL_X32 FILLER_400_2727 ();
 FILLCELL_X32 FILLER_400_2759 ();
 FILLCELL_X32 FILLER_400_2791 ();
 FILLCELL_X32 FILLER_400_2823 ();
 FILLCELL_X32 FILLER_400_2855 ();
 FILLCELL_X32 FILLER_400_2887 ();
 FILLCELL_X32 FILLER_400_2919 ();
 FILLCELL_X32 FILLER_400_2951 ();
 FILLCELL_X32 FILLER_400_2983 ();
 FILLCELL_X32 FILLER_400_3015 ();
 FILLCELL_X32 FILLER_400_3047 ();
 FILLCELL_X32 FILLER_400_3079 ();
 FILLCELL_X32 FILLER_400_3111 ();
 FILLCELL_X8 FILLER_400_3143 ();
 FILLCELL_X4 FILLER_400_3151 ();
 FILLCELL_X2 FILLER_400_3155 ();
 FILLCELL_X32 FILLER_400_3158 ();
 FILLCELL_X32 FILLER_400_3190 ();
 FILLCELL_X32 FILLER_400_3222 ();
 FILLCELL_X32 FILLER_400_3254 ();
 FILLCELL_X32 FILLER_400_3286 ();
 FILLCELL_X32 FILLER_400_3318 ();
 FILLCELL_X32 FILLER_400_3350 ();
 FILLCELL_X32 FILLER_400_3382 ();
 FILLCELL_X32 FILLER_400_3414 ();
 FILLCELL_X32 FILLER_400_3446 ();
 FILLCELL_X32 FILLER_400_3478 ();
 FILLCELL_X32 FILLER_400_3510 ();
 FILLCELL_X32 FILLER_400_3542 ();
 FILLCELL_X32 FILLER_400_3574 ();
 FILLCELL_X32 FILLER_400_3606 ();
 FILLCELL_X32 FILLER_400_3638 ();
 FILLCELL_X32 FILLER_400_3670 ();
 FILLCELL_X32 FILLER_400_3702 ();
 FILLCELL_X4 FILLER_400_3734 ();
 FILLCELL_X32 FILLER_401_1 ();
 FILLCELL_X32 FILLER_401_33 ();
 FILLCELL_X32 FILLER_401_65 ();
 FILLCELL_X32 FILLER_401_97 ();
 FILLCELL_X32 FILLER_401_129 ();
 FILLCELL_X32 FILLER_401_161 ();
 FILLCELL_X32 FILLER_401_193 ();
 FILLCELL_X32 FILLER_401_225 ();
 FILLCELL_X32 FILLER_401_257 ();
 FILLCELL_X32 FILLER_401_289 ();
 FILLCELL_X32 FILLER_401_321 ();
 FILLCELL_X32 FILLER_401_353 ();
 FILLCELL_X32 FILLER_401_385 ();
 FILLCELL_X32 FILLER_401_417 ();
 FILLCELL_X32 FILLER_401_449 ();
 FILLCELL_X32 FILLER_401_481 ();
 FILLCELL_X32 FILLER_401_513 ();
 FILLCELL_X32 FILLER_401_545 ();
 FILLCELL_X32 FILLER_401_577 ();
 FILLCELL_X32 FILLER_401_609 ();
 FILLCELL_X32 FILLER_401_641 ();
 FILLCELL_X32 FILLER_401_673 ();
 FILLCELL_X32 FILLER_401_705 ();
 FILLCELL_X32 FILLER_401_737 ();
 FILLCELL_X32 FILLER_401_769 ();
 FILLCELL_X32 FILLER_401_801 ();
 FILLCELL_X32 FILLER_401_833 ();
 FILLCELL_X32 FILLER_401_865 ();
 FILLCELL_X32 FILLER_401_897 ();
 FILLCELL_X32 FILLER_401_929 ();
 FILLCELL_X32 FILLER_401_961 ();
 FILLCELL_X32 FILLER_401_993 ();
 FILLCELL_X32 FILLER_401_1025 ();
 FILLCELL_X32 FILLER_401_1057 ();
 FILLCELL_X32 FILLER_401_1089 ();
 FILLCELL_X32 FILLER_401_1121 ();
 FILLCELL_X32 FILLER_401_1153 ();
 FILLCELL_X32 FILLER_401_1185 ();
 FILLCELL_X32 FILLER_401_1217 ();
 FILLCELL_X8 FILLER_401_1249 ();
 FILLCELL_X4 FILLER_401_1257 ();
 FILLCELL_X2 FILLER_401_1261 ();
 FILLCELL_X32 FILLER_401_1264 ();
 FILLCELL_X32 FILLER_401_1296 ();
 FILLCELL_X32 FILLER_401_1328 ();
 FILLCELL_X32 FILLER_401_1360 ();
 FILLCELL_X32 FILLER_401_1392 ();
 FILLCELL_X32 FILLER_401_1424 ();
 FILLCELL_X32 FILLER_401_1456 ();
 FILLCELL_X32 FILLER_401_1488 ();
 FILLCELL_X32 FILLER_401_1520 ();
 FILLCELL_X32 FILLER_401_1552 ();
 FILLCELL_X32 FILLER_401_1584 ();
 FILLCELL_X32 FILLER_401_1616 ();
 FILLCELL_X32 FILLER_401_1648 ();
 FILLCELL_X32 FILLER_401_1680 ();
 FILLCELL_X32 FILLER_401_1712 ();
 FILLCELL_X32 FILLER_401_1744 ();
 FILLCELL_X32 FILLER_401_1776 ();
 FILLCELL_X32 FILLER_401_1808 ();
 FILLCELL_X32 FILLER_401_1840 ();
 FILLCELL_X32 FILLER_401_1872 ();
 FILLCELL_X32 FILLER_401_1904 ();
 FILLCELL_X32 FILLER_401_1936 ();
 FILLCELL_X32 FILLER_401_1968 ();
 FILLCELL_X32 FILLER_401_2000 ();
 FILLCELL_X32 FILLER_401_2032 ();
 FILLCELL_X32 FILLER_401_2064 ();
 FILLCELL_X32 FILLER_401_2096 ();
 FILLCELL_X32 FILLER_401_2128 ();
 FILLCELL_X32 FILLER_401_2160 ();
 FILLCELL_X32 FILLER_401_2192 ();
 FILLCELL_X32 FILLER_401_2224 ();
 FILLCELL_X32 FILLER_401_2256 ();
 FILLCELL_X32 FILLER_401_2288 ();
 FILLCELL_X32 FILLER_401_2320 ();
 FILLCELL_X32 FILLER_401_2352 ();
 FILLCELL_X32 FILLER_401_2384 ();
 FILLCELL_X32 FILLER_401_2416 ();
 FILLCELL_X32 FILLER_401_2448 ();
 FILLCELL_X32 FILLER_401_2480 ();
 FILLCELL_X8 FILLER_401_2512 ();
 FILLCELL_X4 FILLER_401_2520 ();
 FILLCELL_X2 FILLER_401_2524 ();
 FILLCELL_X32 FILLER_401_2527 ();
 FILLCELL_X32 FILLER_401_2559 ();
 FILLCELL_X32 FILLER_401_2591 ();
 FILLCELL_X32 FILLER_401_2623 ();
 FILLCELL_X32 FILLER_401_2655 ();
 FILLCELL_X32 FILLER_401_2687 ();
 FILLCELL_X32 FILLER_401_2719 ();
 FILLCELL_X32 FILLER_401_2751 ();
 FILLCELL_X32 FILLER_401_2783 ();
 FILLCELL_X32 FILLER_401_2815 ();
 FILLCELL_X32 FILLER_401_2847 ();
 FILLCELL_X32 FILLER_401_2879 ();
 FILLCELL_X32 FILLER_401_2911 ();
 FILLCELL_X32 FILLER_401_2943 ();
 FILLCELL_X32 FILLER_401_2975 ();
 FILLCELL_X32 FILLER_401_3007 ();
 FILLCELL_X32 FILLER_401_3039 ();
 FILLCELL_X32 FILLER_401_3071 ();
 FILLCELL_X32 FILLER_401_3103 ();
 FILLCELL_X32 FILLER_401_3135 ();
 FILLCELL_X32 FILLER_401_3167 ();
 FILLCELL_X32 FILLER_401_3199 ();
 FILLCELL_X32 FILLER_401_3231 ();
 FILLCELL_X32 FILLER_401_3263 ();
 FILLCELL_X32 FILLER_401_3295 ();
 FILLCELL_X32 FILLER_401_3327 ();
 FILLCELL_X32 FILLER_401_3359 ();
 FILLCELL_X32 FILLER_401_3391 ();
 FILLCELL_X32 FILLER_401_3423 ();
 FILLCELL_X32 FILLER_401_3455 ();
 FILLCELL_X32 FILLER_401_3487 ();
 FILLCELL_X32 FILLER_401_3519 ();
 FILLCELL_X32 FILLER_401_3551 ();
 FILLCELL_X32 FILLER_401_3583 ();
 FILLCELL_X32 FILLER_401_3615 ();
 FILLCELL_X32 FILLER_401_3647 ();
 FILLCELL_X32 FILLER_401_3679 ();
 FILLCELL_X16 FILLER_401_3711 ();
 FILLCELL_X8 FILLER_401_3727 ();
 FILLCELL_X2 FILLER_401_3735 ();
 FILLCELL_X1 FILLER_401_3737 ();
 FILLCELL_X32 FILLER_402_1 ();
 FILLCELL_X32 FILLER_402_33 ();
 FILLCELL_X32 FILLER_402_65 ();
 FILLCELL_X32 FILLER_402_97 ();
 FILLCELL_X32 FILLER_402_129 ();
 FILLCELL_X32 FILLER_402_161 ();
 FILLCELL_X32 FILLER_402_193 ();
 FILLCELL_X32 FILLER_402_225 ();
 FILLCELL_X32 FILLER_402_257 ();
 FILLCELL_X32 FILLER_402_289 ();
 FILLCELL_X32 FILLER_402_321 ();
 FILLCELL_X32 FILLER_402_353 ();
 FILLCELL_X32 FILLER_402_385 ();
 FILLCELL_X32 FILLER_402_417 ();
 FILLCELL_X32 FILLER_402_449 ();
 FILLCELL_X32 FILLER_402_481 ();
 FILLCELL_X32 FILLER_402_513 ();
 FILLCELL_X32 FILLER_402_545 ();
 FILLCELL_X32 FILLER_402_577 ();
 FILLCELL_X16 FILLER_402_609 ();
 FILLCELL_X4 FILLER_402_625 ();
 FILLCELL_X2 FILLER_402_629 ();
 FILLCELL_X32 FILLER_402_632 ();
 FILLCELL_X32 FILLER_402_664 ();
 FILLCELL_X32 FILLER_402_696 ();
 FILLCELL_X32 FILLER_402_728 ();
 FILLCELL_X32 FILLER_402_760 ();
 FILLCELL_X32 FILLER_402_792 ();
 FILLCELL_X32 FILLER_402_824 ();
 FILLCELL_X32 FILLER_402_856 ();
 FILLCELL_X32 FILLER_402_888 ();
 FILLCELL_X32 FILLER_402_920 ();
 FILLCELL_X32 FILLER_402_952 ();
 FILLCELL_X32 FILLER_402_984 ();
 FILLCELL_X32 FILLER_402_1016 ();
 FILLCELL_X32 FILLER_402_1048 ();
 FILLCELL_X32 FILLER_402_1080 ();
 FILLCELL_X32 FILLER_402_1112 ();
 FILLCELL_X32 FILLER_402_1144 ();
 FILLCELL_X32 FILLER_402_1176 ();
 FILLCELL_X32 FILLER_402_1208 ();
 FILLCELL_X32 FILLER_402_1240 ();
 FILLCELL_X32 FILLER_402_1272 ();
 FILLCELL_X32 FILLER_402_1304 ();
 FILLCELL_X32 FILLER_402_1336 ();
 FILLCELL_X32 FILLER_402_1368 ();
 FILLCELL_X32 FILLER_402_1400 ();
 FILLCELL_X32 FILLER_402_1432 ();
 FILLCELL_X32 FILLER_402_1464 ();
 FILLCELL_X32 FILLER_402_1496 ();
 FILLCELL_X32 FILLER_402_1528 ();
 FILLCELL_X32 FILLER_402_1560 ();
 FILLCELL_X32 FILLER_402_1592 ();
 FILLCELL_X32 FILLER_402_1624 ();
 FILLCELL_X32 FILLER_402_1656 ();
 FILLCELL_X32 FILLER_402_1688 ();
 FILLCELL_X32 FILLER_402_1720 ();
 FILLCELL_X32 FILLER_402_1752 ();
 FILLCELL_X32 FILLER_402_1784 ();
 FILLCELL_X32 FILLER_402_1816 ();
 FILLCELL_X32 FILLER_402_1848 ();
 FILLCELL_X8 FILLER_402_1880 ();
 FILLCELL_X4 FILLER_402_1888 ();
 FILLCELL_X2 FILLER_402_1892 ();
 FILLCELL_X32 FILLER_402_1895 ();
 FILLCELL_X32 FILLER_402_1927 ();
 FILLCELL_X32 FILLER_402_1959 ();
 FILLCELL_X32 FILLER_402_1991 ();
 FILLCELL_X32 FILLER_402_2023 ();
 FILLCELL_X32 FILLER_402_2055 ();
 FILLCELL_X32 FILLER_402_2087 ();
 FILLCELL_X32 FILLER_402_2119 ();
 FILLCELL_X32 FILLER_402_2151 ();
 FILLCELL_X32 FILLER_402_2183 ();
 FILLCELL_X32 FILLER_402_2215 ();
 FILLCELL_X32 FILLER_402_2247 ();
 FILLCELL_X32 FILLER_402_2279 ();
 FILLCELL_X32 FILLER_402_2311 ();
 FILLCELL_X32 FILLER_402_2343 ();
 FILLCELL_X32 FILLER_402_2375 ();
 FILLCELL_X32 FILLER_402_2407 ();
 FILLCELL_X32 FILLER_402_2439 ();
 FILLCELL_X32 FILLER_402_2471 ();
 FILLCELL_X32 FILLER_402_2503 ();
 FILLCELL_X32 FILLER_402_2535 ();
 FILLCELL_X32 FILLER_402_2567 ();
 FILLCELL_X32 FILLER_402_2599 ();
 FILLCELL_X32 FILLER_402_2631 ();
 FILLCELL_X32 FILLER_402_2663 ();
 FILLCELL_X32 FILLER_402_2695 ();
 FILLCELL_X32 FILLER_402_2727 ();
 FILLCELL_X32 FILLER_402_2759 ();
 FILLCELL_X32 FILLER_402_2791 ();
 FILLCELL_X32 FILLER_402_2823 ();
 FILLCELL_X32 FILLER_402_2855 ();
 FILLCELL_X32 FILLER_402_2887 ();
 FILLCELL_X32 FILLER_402_2919 ();
 FILLCELL_X32 FILLER_402_2951 ();
 FILLCELL_X32 FILLER_402_2983 ();
 FILLCELL_X32 FILLER_402_3015 ();
 FILLCELL_X32 FILLER_402_3047 ();
 FILLCELL_X32 FILLER_402_3079 ();
 FILLCELL_X32 FILLER_402_3111 ();
 FILLCELL_X8 FILLER_402_3143 ();
 FILLCELL_X4 FILLER_402_3151 ();
 FILLCELL_X2 FILLER_402_3155 ();
 FILLCELL_X32 FILLER_402_3158 ();
 FILLCELL_X32 FILLER_402_3190 ();
 FILLCELL_X32 FILLER_402_3222 ();
 FILLCELL_X32 FILLER_402_3254 ();
 FILLCELL_X32 FILLER_402_3286 ();
 FILLCELL_X32 FILLER_402_3318 ();
 FILLCELL_X32 FILLER_402_3350 ();
 FILLCELL_X32 FILLER_402_3382 ();
 FILLCELL_X32 FILLER_402_3414 ();
 FILLCELL_X32 FILLER_402_3446 ();
 FILLCELL_X32 FILLER_402_3478 ();
 FILLCELL_X32 FILLER_402_3510 ();
 FILLCELL_X32 FILLER_402_3542 ();
 FILLCELL_X32 FILLER_402_3574 ();
 FILLCELL_X32 FILLER_402_3606 ();
 FILLCELL_X32 FILLER_402_3638 ();
 FILLCELL_X32 FILLER_402_3670 ();
 FILLCELL_X32 FILLER_402_3702 ();
 FILLCELL_X4 FILLER_402_3734 ();
 FILLCELL_X32 FILLER_403_1 ();
 FILLCELL_X32 FILLER_403_33 ();
 FILLCELL_X32 FILLER_403_65 ();
 FILLCELL_X32 FILLER_403_97 ();
 FILLCELL_X32 FILLER_403_129 ();
 FILLCELL_X32 FILLER_403_161 ();
 FILLCELL_X32 FILLER_403_193 ();
 FILLCELL_X32 FILLER_403_225 ();
 FILLCELL_X32 FILLER_403_257 ();
 FILLCELL_X32 FILLER_403_289 ();
 FILLCELL_X32 FILLER_403_321 ();
 FILLCELL_X32 FILLER_403_353 ();
 FILLCELL_X32 FILLER_403_385 ();
 FILLCELL_X32 FILLER_403_417 ();
 FILLCELL_X32 FILLER_403_449 ();
 FILLCELL_X32 FILLER_403_481 ();
 FILLCELL_X32 FILLER_403_513 ();
 FILLCELL_X32 FILLER_403_545 ();
 FILLCELL_X32 FILLER_403_577 ();
 FILLCELL_X32 FILLER_403_609 ();
 FILLCELL_X32 FILLER_403_641 ();
 FILLCELL_X32 FILLER_403_673 ();
 FILLCELL_X32 FILLER_403_705 ();
 FILLCELL_X32 FILLER_403_737 ();
 FILLCELL_X32 FILLER_403_769 ();
 FILLCELL_X32 FILLER_403_801 ();
 FILLCELL_X32 FILLER_403_833 ();
 FILLCELL_X32 FILLER_403_865 ();
 FILLCELL_X32 FILLER_403_897 ();
 FILLCELL_X32 FILLER_403_929 ();
 FILLCELL_X32 FILLER_403_961 ();
 FILLCELL_X32 FILLER_403_993 ();
 FILLCELL_X32 FILLER_403_1025 ();
 FILLCELL_X32 FILLER_403_1057 ();
 FILLCELL_X32 FILLER_403_1089 ();
 FILLCELL_X32 FILLER_403_1121 ();
 FILLCELL_X32 FILLER_403_1153 ();
 FILLCELL_X32 FILLER_403_1185 ();
 FILLCELL_X32 FILLER_403_1217 ();
 FILLCELL_X8 FILLER_403_1249 ();
 FILLCELL_X4 FILLER_403_1257 ();
 FILLCELL_X2 FILLER_403_1261 ();
 FILLCELL_X32 FILLER_403_1264 ();
 FILLCELL_X32 FILLER_403_1296 ();
 FILLCELL_X32 FILLER_403_1328 ();
 FILLCELL_X32 FILLER_403_1360 ();
 FILLCELL_X32 FILLER_403_1392 ();
 FILLCELL_X32 FILLER_403_1424 ();
 FILLCELL_X32 FILLER_403_1456 ();
 FILLCELL_X32 FILLER_403_1488 ();
 FILLCELL_X32 FILLER_403_1520 ();
 FILLCELL_X32 FILLER_403_1552 ();
 FILLCELL_X32 FILLER_403_1584 ();
 FILLCELL_X32 FILLER_403_1616 ();
 FILLCELL_X32 FILLER_403_1648 ();
 FILLCELL_X32 FILLER_403_1680 ();
 FILLCELL_X32 FILLER_403_1712 ();
 FILLCELL_X32 FILLER_403_1744 ();
 FILLCELL_X32 FILLER_403_1776 ();
 FILLCELL_X32 FILLER_403_1808 ();
 FILLCELL_X32 FILLER_403_1840 ();
 FILLCELL_X32 FILLER_403_1872 ();
 FILLCELL_X32 FILLER_403_1904 ();
 FILLCELL_X32 FILLER_403_1936 ();
 FILLCELL_X32 FILLER_403_1968 ();
 FILLCELL_X32 FILLER_403_2000 ();
 FILLCELL_X32 FILLER_403_2032 ();
 FILLCELL_X32 FILLER_403_2064 ();
 FILLCELL_X32 FILLER_403_2096 ();
 FILLCELL_X32 FILLER_403_2128 ();
 FILLCELL_X32 FILLER_403_2160 ();
 FILLCELL_X32 FILLER_403_2192 ();
 FILLCELL_X32 FILLER_403_2224 ();
 FILLCELL_X32 FILLER_403_2256 ();
 FILLCELL_X32 FILLER_403_2288 ();
 FILLCELL_X32 FILLER_403_2320 ();
 FILLCELL_X32 FILLER_403_2352 ();
 FILLCELL_X32 FILLER_403_2384 ();
 FILLCELL_X32 FILLER_403_2416 ();
 FILLCELL_X32 FILLER_403_2448 ();
 FILLCELL_X32 FILLER_403_2480 ();
 FILLCELL_X8 FILLER_403_2512 ();
 FILLCELL_X4 FILLER_403_2520 ();
 FILLCELL_X2 FILLER_403_2524 ();
 FILLCELL_X32 FILLER_403_2527 ();
 FILLCELL_X32 FILLER_403_2559 ();
 FILLCELL_X32 FILLER_403_2591 ();
 FILLCELL_X32 FILLER_403_2623 ();
 FILLCELL_X32 FILLER_403_2655 ();
 FILLCELL_X32 FILLER_403_2687 ();
 FILLCELL_X32 FILLER_403_2719 ();
 FILLCELL_X32 FILLER_403_2751 ();
 FILLCELL_X32 FILLER_403_2783 ();
 FILLCELL_X32 FILLER_403_2815 ();
 FILLCELL_X32 FILLER_403_2847 ();
 FILLCELL_X32 FILLER_403_2879 ();
 FILLCELL_X32 FILLER_403_2911 ();
 FILLCELL_X32 FILLER_403_2943 ();
 FILLCELL_X32 FILLER_403_2975 ();
 FILLCELL_X32 FILLER_403_3007 ();
 FILLCELL_X32 FILLER_403_3039 ();
 FILLCELL_X32 FILLER_403_3071 ();
 FILLCELL_X32 FILLER_403_3103 ();
 FILLCELL_X32 FILLER_403_3135 ();
 FILLCELL_X32 FILLER_403_3167 ();
 FILLCELL_X32 FILLER_403_3199 ();
 FILLCELL_X32 FILLER_403_3231 ();
 FILLCELL_X32 FILLER_403_3263 ();
 FILLCELL_X32 FILLER_403_3295 ();
 FILLCELL_X32 FILLER_403_3327 ();
 FILLCELL_X32 FILLER_403_3359 ();
 FILLCELL_X32 FILLER_403_3391 ();
 FILLCELL_X32 FILLER_403_3423 ();
 FILLCELL_X32 FILLER_403_3455 ();
 FILLCELL_X32 FILLER_403_3487 ();
 FILLCELL_X32 FILLER_403_3519 ();
 FILLCELL_X32 FILLER_403_3551 ();
 FILLCELL_X32 FILLER_403_3583 ();
 FILLCELL_X32 FILLER_403_3615 ();
 FILLCELL_X32 FILLER_403_3647 ();
 FILLCELL_X32 FILLER_403_3679 ();
 FILLCELL_X16 FILLER_403_3711 ();
 FILLCELL_X8 FILLER_403_3727 ();
 FILLCELL_X2 FILLER_403_3735 ();
 FILLCELL_X1 FILLER_403_3737 ();
 FILLCELL_X32 FILLER_404_1 ();
 FILLCELL_X32 FILLER_404_33 ();
 FILLCELL_X32 FILLER_404_65 ();
 FILLCELL_X32 FILLER_404_97 ();
 FILLCELL_X32 FILLER_404_129 ();
 FILLCELL_X32 FILLER_404_161 ();
 FILLCELL_X32 FILLER_404_193 ();
 FILLCELL_X32 FILLER_404_225 ();
 FILLCELL_X32 FILLER_404_257 ();
 FILLCELL_X32 FILLER_404_289 ();
 FILLCELL_X32 FILLER_404_321 ();
 FILLCELL_X32 FILLER_404_353 ();
 FILLCELL_X32 FILLER_404_385 ();
 FILLCELL_X32 FILLER_404_417 ();
 FILLCELL_X32 FILLER_404_449 ();
 FILLCELL_X32 FILLER_404_481 ();
 FILLCELL_X32 FILLER_404_513 ();
 FILLCELL_X32 FILLER_404_545 ();
 FILLCELL_X32 FILLER_404_577 ();
 FILLCELL_X16 FILLER_404_609 ();
 FILLCELL_X4 FILLER_404_625 ();
 FILLCELL_X2 FILLER_404_629 ();
 FILLCELL_X32 FILLER_404_632 ();
 FILLCELL_X32 FILLER_404_664 ();
 FILLCELL_X32 FILLER_404_696 ();
 FILLCELL_X32 FILLER_404_728 ();
 FILLCELL_X32 FILLER_404_760 ();
 FILLCELL_X32 FILLER_404_792 ();
 FILLCELL_X32 FILLER_404_824 ();
 FILLCELL_X32 FILLER_404_856 ();
 FILLCELL_X32 FILLER_404_888 ();
 FILLCELL_X32 FILLER_404_920 ();
 FILLCELL_X32 FILLER_404_952 ();
 FILLCELL_X32 FILLER_404_984 ();
 FILLCELL_X32 FILLER_404_1016 ();
 FILLCELL_X32 FILLER_404_1048 ();
 FILLCELL_X32 FILLER_404_1080 ();
 FILLCELL_X32 FILLER_404_1112 ();
 FILLCELL_X32 FILLER_404_1144 ();
 FILLCELL_X32 FILLER_404_1176 ();
 FILLCELL_X32 FILLER_404_1208 ();
 FILLCELL_X32 FILLER_404_1240 ();
 FILLCELL_X32 FILLER_404_1272 ();
 FILLCELL_X32 FILLER_404_1304 ();
 FILLCELL_X32 FILLER_404_1336 ();
 FILLCELL_X32 FILLER_404_1368 ();
 FILLCELL_X32 FILLER_404_1400 ();
 FILLCELL_X32 FILLER_404_1432 ();
 FILLCELL_X32 FILLER_404_1464 ();
 FILLCELL_X32 FILLER_404_1496 ();
 FILLCELL_X32 FILLER_404_1528 ();
 FILLCELL_X32 FILLER_404_1560 ();
 FILLCELL_X32 FILLER_404_1592 ();
 FILLCELL_X32 FILLER_404_1624 ();
 FILLCELL_X32 FILLER_404_1656 ();
 FILLCELL_X32 FILLER_404_1688 ();
 FILLCELL_X32 FILLER_404_1720 ();
 FILLCELL_X32 FILLER_404_1752 ();
 FILLCELL_X32 FILLER_404_1784 ();
 FILLCELL_X32 FILLER_404_1816 ();
 FILLCELL_X32 FILLER_404_1848 ();
 FILLCELL_X8 FILLER_404_1880 ();
 FILLCELL_X4 FILLER_404_1888 ();
 FILLCELL_X2 FILLER_404_1892 ();
 FILLCELL_X32 FILLER_404_1895 ();
 FILLCELL_X32 FILLER_404_1927 ();
 FILLCELL_X32 FILLER_404_1959 ();
 FILLCELL_X32 FILLER_404_1991 ();
 FILLCELL_X32 FILLER_404_2023 ();
 FILLCELL_X32 FILLER_404_2055 ();
 FILLCELL_X32 FILLER_404_2087 ();
 FILLCELL_X32 FILLER_404_2119 ();
 FILLCELL_X32 FILLER_404_2151 ();
 FILLCELL_X32 FILLER_404_2183 ();
 FILLCELL_X32 FILLER_404_2215 ();
 FILLCELL_X32 FILLER_404_2247 ();
 FILLCELL_X32 FILLER_404_2279 ();
 FILLCELL_X32 FILLER_404_2311 ();
 FILLCELL_X32 FILLER_404_2343 ();
 FILLCELL_X32 FILLER_404_2375 ();
 FILLCELL_X32 FILLER_404_2407 ();
 FILLCELL_X32 FILLER_404_2439 ();
 FILLCELL_X32 FILLER_404_2471 ();
 FILLCELL_X32 FILLER_404_2503 ();
 FILLCELL_X32 FILLER_404_2535 ();
 FILLCELL_X32 FILLER_404_2567 ();
 FILLCELL_X32 FILLER_404_2599 ();
 FILLCELL_X32 FILLER_404_2631 ();
 FILLCELL_X32 FILLER_404_2663 ();
 FILLCELL_X32 FILLER_404_2695 ();
 FILLCELL_X32 FILLER_404_2727 ();
 FILLCELL_X32 FILLER_404_2759 ();
 FILLCELL_X32 FILLER_404_2791 ();
 FILLCELL_X32 FILLER_404_2823 ();
 FILLCELL_X32 FILLER_404_2855 ();
 FILLCELL_X32 FILLER_404_2887 ();
 FILLCELL_X32 FILLER_404_2919 ();
 FILLCELL_X32 FILLER_404_2951 ();
 FILLCELL_X32 FILLER_404_2983 ();
 FILLCELL_X32 FILLER_404_3015 ();
 FILLCELL_X32 FILLER_404_3047 ();
 FILLCELL_X32 FILLER_404_3079 ();
 FILLCELL_X32 FILLER_404_3111 ();
 FILLCELL_X8 FILLER_404_3143 ();
 FILLCELL_X4 FILLER_404_3151 ();
 FILLCELL_X2 FILLER_404_3155 ();
 FILLCELL_X32 FILLER_404_3158 ();
 FILLCELL_X32 FILLER_404_3190 ();
 FILLCELL_X32 FILLER_404_3222 ();
 FILLCELL_X32 FILLER_404_3254 ();
 FILLCELL_X32 FILLER_404_3286 ();
 FILLCELL_X32 FILLER_404_3318 ();
 FILLCELL_X32 FILLER_404_3350 ();
 FILLCELL_X32 FILLER_404_3382 ();
 FILLCELL_X32 FILLER_404_3414 ();
 FILLCELL_X32 FILLER_404_3446 ();
 FILLCELL_X32 FILLER_404_3478 ();
 FILLCELL_X32 FILLER_404_3510 ();
 FILLCELL_X32 FILLER_404_3542 ();
 FILLCELL_X32 FILLER_404_3574 ();
 FILLCELL_X32 FILLER_404_3606 ();
 FILLCELL_X32 FILLER_404_3638 ();
 FILLCELL_X32 FILLER_404_3670 ();
 FILLCELL_X32 FILLER_404_3702 ();
 FILLCELL_X4 FILLER_404_3734 ();
 FILLCELL_X32 FILLER_405_1 ();
 FILLCELL_X32 FILLER_405_33 ();
 FILLCELL_X32 FILLER_405_65 ();
 FILLCELL_X32 FILLER_405_97 ();
 FILLCELL_X32 FILLER_405_129 ();
 FILLCELL_X32 FILLER_405_161 ();
 FILLCELL_X32 FILLER_405_193 ();
 FILLCELL_X32 FILLER_405_225 ();
 FILLCELL_X32 FILLER_405_257 ();
 FILLCELL_X32 FILLER_405_289 ();
 FILLCELL_X32 FILLER_405_321 ();
 FILLCELL_X32 FILLER_405_353 ();
 FILLCELL_X32 FILLER_405_385 ();
 FILLCELL_X32 FILLER_405_417 ();
 FILLCELL_X32 FILLER_405_449 ();
 FILLCELL_X32 FILLER_405_481 ();
 FILLCELL_X32 FILLER_405_513 ();
 FILLCELL_X32 FILLER_405_545 ();
 FILLCELL_X32 FILLER_405_577 ();
 FILLCELL_X32 FILLER_405_609 ();
 FILLCELL_X32 FILLER_405_641 ();
 FILLCELL_X32 FILLER_405_673 ();
 FILLCELL_X32 FILLER_405_705 ();
 FILLCELL_X32 FILLER_405_737 ();
 FILLCELL_X32 FILLER_405_769 ();
 FILLCELL_X32 FILLER_405_801 ();
 FILLCELL_X32 FILLER_405_833 ();
 FILLCELL_X32 FILLER_405_865 ();
 FILLCELL_X32 FILLER_405_897 ();
 FILLCELL_X32 FILLER_405_929 ();
 FILLCELL_X32 FILLER_405_961 ();
 FILLCELL_X32 FILLER_405_993 ();
 FILLCELL_X32 FILLER_405_1025 ();
 FILLCELL_X32 FILLER_405_1057 ();
 FILLCELL_X32 FILLER_405_1089 ();
 FILLCELL_X32 FILLER_405_1121 ();
 FILLCELL_X32 FILLER_405_1153 ();
 FILLCELL_X32 FILLER_405_1185 ();
 FILLCELL_X32 FILLER_405_1217 ();
 FILLCELL_X8 FILLER_405_1249 ();
 FILLCELL_X4 FILLER_405_1257 ();
 FILLCELL_X2 FILLER_405_1261 ();
 FILLCELL_X32 FILLER_405_1264 ();
 FILLCELL_X32 FILLER_405_1296 ();
 FILLCELL_X32 FILLER_405_1328 ();
 FILLCELL_X32 FILLER_405_1360 ();
 FILLCELL_X32 FILLER_405_1392 ();
 FILLCELL_X32 FILLER_405_1424 ();
 FILLCELL_X32 FILLER_405_1456 ();
 FILLCELL_X32 FILLER_405_1488 ();
 FILLCELL_X32 FILLER_405_1520 ();
 FILLCELL_X32 FILLER_405_1552 ();
 FILLCELL_X32 FILLER_405_1584 ();
 FILLCELL_X32 FILLER_405_1616 ();
 FILLCELL_X32 FILLER_405_1648 ();
 FILLCELL_X32 FILLER_405_1680 ();
 FILLCELL_X32 FILLER_405_1712 ();
 FILLCELL_X32 FILLER_405_1744 ();
 FILLCELL_X32 FILLER_405_1776 ();
 FILLCELL_X32 FILLER_405_1808 ();
 FILLCELL_X32 FILLER_405_1840 ();
 FILLCELL_X32 FILLER_405_1872 ();
 FILLCELL_X32 FILLER_405_1904 ();
 FILLCELL_X32 FILLER_405_1936 ();
 FILLCELL_X32 FILLER_405_1968 ();
 FILLCELL_X32 FILLER_405_2000 ();
 FILLCELL_X32 FILLER_405_2032 ();
 FILLCELL_X32 FILLER_405_2064 ();
 FILLCELL_X32 FILLER_405_2096 ();
 FILLCELL_X32 FILLER_405_2128 ();
 FILLCELL_X32 FILLER_405_2160 ();
 FILLCELL_X32 FILLER_405_2192 ();
 FILLCELL_X32 FILLER_405_2224 ();
 FILLCELL_X32 FILLER_405_2256 ();
 FILLCELL_X32 FILLER_405_2288 ();
 FILLCELL_X32 FILLER_405_2320 ();
 FILLCELL_X32 FILLER_405_2352 ();
 FILLCELL_X32 FILLER_405_2384 ();
 FILLCELL_X32 FILLER_405_2416 ();
 FILLCELL_X32 FILLER_405_2448 ();
 FILLCELL_X32 FILLER_405_2480 ();
 FILLCELL_X8 FILLER_405_2512 ();
 FILLCELL_X4 FILLER_405_2520 ();
 FILLCELL_X2 FILLER_405_2524 ();
 FILLCELL_X32 FILLER_405_2527 ();
 FILLCELL_X32 FILLER_405_2559 ();
 FILLCELL_X32 FILLER_405_2591 ();
 FILLCELL_X32 FILLER_405_2623 ();
 FILLCELL_X32 FILLER_405_2655 ();
 FILLCELL_X32 FILLER_405_2687 ();
 FILLCELL_X32 FILLER_405_2719 ();
 FILLCELL_X32 FILLER_405_2751 ();
 FILLCELL_X32 FILLER_405_2783 ();
 FILLCELL_X32 FILLER_405_2815 ();
 FILLCELL_X32 FILLER_405_2847 ();
 FILLCELL_X32 FILLER_405_2879 ();
 FILLCELL_X32 FILLER_405_2911 ();
 FILLCELL_X32 FILLER_405_2943 ();
 FILLCELL_X32 FILLER_405_2975 ();
 FILLCELL_X32 FILLER_405_3007 ();
 FILLCELL_X32 FILLER_405_3039 ();
 FILLCELL_X32 FILLER_405_3071 ();
 FILLCELL_X32 FILLER_405_3103 ();
 FILLCELL_X32 FILLER_405_3135 ();
 FILLCELL_X32 FILLER_405_3167 ();
 FILLCELL_X32 FILLER_405_3199 ();
 FILLCELL_X32 FILLER_405_3231 ();
 FILLCELL_X32 FILLER_405_3263 ();
 FILLCELL_X32 FILLER_405_3295 ();
 FILLCELL_X32 FILLER_405_3327 ();
 FILLCELL_X32 FILLER_405_3359 ();
 FILLCELL_X32 FILLER_405_3391 ();
 FILLCELL_X32 FILLER_405_3423 ();
 FILLCELL_X32 FILLER_405_3455 ();
 FILLCELL_X32 FILLER_405_3487 ();
 FILLCELL_X32 FILLER_405_3519 ();
 FILLCELL_X32 FILLER_405_3551 ();
 FILLCELL_X32 FILLER_405_3583 ();
 FILLCELL_X32 FILLER_405_3615 ();
 FILLCELL_X32 FILLER_405_3647 ();
 FILLCELL_X32 FILLER_405_3679 ();
 FILLCELL_X16 FILLER_405_3711 ();
 FILLCELL_X8 FILLER_405_3727 ();
 FILLCELL_X2 FILLER_405_3735 ();
 FILLCELL_X1 FILLER_405_3737 ();
 FILLCELL_X32 FILLER_406_1 ();
 FILLCELL_X32 FILLER_406_33 ();
 FILLCELL_X32 FILLER_406_65 ();
 FILLCELL_X32 FILLER_406_97 ();
 FILLCELL_X32 FILLER_406_129 ();
 FILLCELL_X32 FILLER_406_161 ();
 FILLCELL_X32 FILLER_406_193 ();
 FILLCELL_X32 FILLER_406_225 ();
 FILLCELL_X32 FILLER_406_257 ();
 FILLCELL_X32 FILLER_406_289 ();
 FILLCELL_X32 FILLER_406_321 ();
 FILLCELL_X32 FILLER_406_353 ();
 FILLCELL_X32 FILLER_406_385 ();
 FILLCELL_X32 FILLER_406_417 ();
 FILLCELL_X32 FILLER_406_449 ();
 FILLCELL_X32 FILLER_406_481 ();
 FILLCELL_X32 FILLER_406_513 ();
 FILLCELL_X32 FILLER_406_545 ();
 FILLCELL_X32 FILLER_406_577 ();
 FILLCELL_X16 FILLER_406_609 ();
 FILLCELL_X4 FILLER_406_625 ();
 FILLCELL_X2 FILLER_406_629 ();
 FILLCELL_X32 FILLER_406_632 ();
 FILLCELL_X32 FILLER_406_664 ();
 FILLCELL_X32 FILLER_406_696 ();
 FILLCELL_X32 FILLER_406_728 ();
 FILLCELL_X32 FILLER_406_760 ();
 FILLCELL_X32 FILLER_406_792 ();
 FILLCELL_X32 FILLER_406_824 ();
 FILLCELL_X32 FILLER_406_856 ();
 FILLCELL_X32 FILLER_406_888 ();
 FILLCELL_X32 FILLER_406_920 ();
 FILLCELL_X32 FILLER_406_952 ();
 FILLCELL_X32 FILLER_406_984 ();
 FILLCELL_X32 FILLER_406_1016 ();
 FILLCELL_X32 FILLER_406_1048 ();
 FILLCELL_X32 FILLER_406_1080 ();
 FILLCELL_X32 FILLER_406_1112 ();
 FILLCELL_X32 FILLER_406_1144 ();
 FILLCELL_X32 FILLER_406_1176 ();
 FILLCELL_X32 FILLER_406_1208 ();
 FILLCELL_X32 FILLER_406_1240 ();
 FILLCELL_X32 FILLER_406_1272 ();
 FILLCELL_X32 FILLER_406_1304 ();
 FILLCELL_X32 FILLER_406_1336 ();
 FILLCELL_X32 FILLER_406_1368 ();
 FILLCELL_X32 FILLER_406_1400 ();
 FILLCELL_X32 FILLER_406_1432 ();
 FILLCELL_X32 FILLER_406_1464 ();
 FILLCELL_X32 FILLER_406_1496 ();
 FILLCELL_X32 FILLER_406_1528 ();
 FILLCELL_X32 FILLER_406_1560 ();
 FILLCELL_X32 FILLER_406_1592 ();
 FILLCELL_X32 FILLER_406_1624 ();
 FILLCELL_X32 FILLER_406_1656 ();
 FILLCELL_X32 FILLER_406_1688 ();
 FILLCELL_X32 FILLER_406_1720 ();
 FILLCELL_X32 FILLER_406_1752 ();
 FILLCELL_X32 FILLER_406_1784 ();
 FILLCELL_X32 FILLER_406_1816 ();
 FILLCELL_X32 FILLER_406_1848 ();
 FILLCELL_X8 FILLER_406_1880 ();
 FILLCELL_X4 FILLER_406_1888 ();
 FILLCELL_X2 FILLER_406_1892 ();
 FILLCELL_X32 FILLER_406_1895 ();
 FILLCELL_X32 FILLER_406_1927 ();
 FILLCELL_X32 FILLER_406_1959 ();
 FILLCELL_X32 FILLER_406_1991 ();
 FILLCELL_X32 FILLER_406_2023 ();
 FILLCELL_X32 FILLER_406_2055 ();
 FILLCELL_X32 FILLER_406_2087 ();
 FILLCELL_X32 FILLER_406_2119 ();
 FILLCELL_X32 FILLER_406_2151 ();
 FILLCELL_X32 FILLER_406_2183 ();
 FILLCELL_X32 FILLER_406_2215 ();
 FILLCELL_X32 FILLER_406_2247 ();
 FILLCELL_X32 FILLER_406_2279 ();
 FILLCELL_X32 FILLER_406_2311 ();
 FILLCELL_X32 FILLER_406_2343 ();
 FILLCELL_X32 FILLER_406_2375 ();
 FILLCELL_X32 FILLER_406_2407 ();
 FILLCELL_X32 FILLER_406_2439 ();
 FILLCELL_X32 FILLER_406_2471 ();
 FILLCELL_X32 FILLER_406_2503 ();
 FILLCELL_X32 FILLER_406_2535 ();
 FILLCELL_X32 FILLER_406_2567 ();
 FILLCELL_X32 FILLER_406_2599 ();
 FILLCELL_X32 FILLER_406_2631 ();
 FILLCELL_X32 FILLER_406_2663 ();
 FILLCELL_X32 FILLER_406_2695 ();
 FILLCELL_X32 FILLER_406_2727 ();
 FILLCELL_X32 FILLER_406_2759 ();
 FILLCELL_X32 FILLER_406_2791 ();
 FILLCELL_X32 FILLER_406_2823 ();
 FILLCELL_X32 FILLER_406_2855 ();
 FILLCELL_X32 FILLER_406_2887 ();
 FILLCELL_X32 FILLER_406_2919 ();
 FILLCELL_X32 FILLER_406_2951 ();
 FILLCELL_X32 FILLER_406_2983 ();
 FILLCELL_X32 FILLER_406_3015 ();
 FILLCELL_X32 FILLER_406_3047 ();
 FILLCELL_X32 FILLER_406_3079 ();
 FILLCELL_X32 FILLER_406_3111 ();
 FILLCELL_X8 FILLER_406_3143 ();
 FILLCELL_X4 FILLER_406_3151 ();
 FILLCELL_X2 FILLER_406_3155 ();
 FILLCELL_X32 FILLER_406_3158 ();
 FILLCELL_X32 FILLER_406_3190 ();
 FILLCELL_X32 FILLER_406_3222 ();
 FILLCELL_X32 FILLER_406_3254 ();
 FILLCELL_X32 FILLER_406_3286 ();
 FILLCELL_X32 FILLER_406_3318 ();
 FILLCELL_X32 FILLER_406_3350 ();
 FILLCELL_X32 FILLER_406_3382 ();
 FILLCELL_X32 FILLER_406_3414 ();
 FILLCELL_X32 FILLER_406_3446 ();
 FILLCELL_X32 FILLER_406_3478 ();
 FILLCELL_X32 FILLER_406_3510 ();
 FILLCELL_X32 FILLER_406_3542 ();
 FILLCELL_X32 FILLER_406_3574 ();
 FILLCELL_X32 FILLER_406_3606 ();
 FILLCELL_X32 FILLER_406_3638 ();
 FILLCELL_X32 FILLER_406_3670 ();
 FILLCELL_X32 FILLER_406_3702 ();
 FILLCELL_X4 FILLER_406_3734 ();
 FILLCELL_X32 FILLER_407_1 ();
 FILLCELL_X32 FILLER_407_33 ();
 FILLCELL_X32 FILLER_407_65 ();
 FILLCELL_X32 FILLER_407_97 ();
 FILLCELL_X32 FILLER_407_129 ();
 FILLCELL_X32 FILLER_407_161 ();
 FILLCELL_X32 FILLER_407_193 ();
 FILLCELL_X32 FILLER_407_225 ();
 FILLCELL_X32 FILLER_407_257 ();
 FILLCELL_X32 FILLER_407_289 ();
 FILLCELL_X32 FILLER_407_321 ();
 FILLCELL_X32 FILLER_407_353 ();
 FILLCELL_X32 FILLER_407_385 ();
 FILLCELL_X32 FILLER_407_417 ();
 FILLCELL_X32 FILLER_407_449 ();
 FILLCELL_X32 FILLER_407_481 ();
 FILLCELL_X32 FILLER_407_513 ();
 FILLCELL_X32 FILLER_407_545 ();
 FILLCELL_X32 FILLER_407_577 ();
 FILLCELL_X32 FILLER_407_609 ();
 FILLCELL_X32 FILLER_407_641 ();
 FILLCELL_X32 FILLER_407_673 ();
 FILLCELL_X32 FILLER_407_705 ();
 FILLCELL_X32 FILLER_407_737 ();
 FILLCELL_X32 FILLER_407_769 ();
 FILLCELL_X32 FILLER_407_801 ();
 FILLCELL_X32 FILLER_407_833 ();
 FILLCELL_X32 FILLER_407_865 ();
 FILLCELL_X32 FILLER_407_897 ();
 FILLCELL_X32 FILLER_407_929 ();
 FILLCELL_X32 FILLER_407_961 ();
 FILLCELL_X32 FILLER_407_993 ();
 FILLCELL_X32 FILLER_407_1025 ();
 FILLCELL_X32 FILLER_407_1057 ();
 FILLCELL_X32 FILLER_407_1089 ();
 FILLCELL_X32 FILLER_407_1121 ();
 FILLCELL_X32 FILLER_407_1153 ();
 FILLCELL_X32 FILLER_407_1185 ();
 FILLCELL_X32 FILLER_407_1217 ();
 FILLCELL_X8 FILLER_407_1249 ();
 FILLCELL_X4 FILLER_407_1257 ();
 FILLCELL_X2 FILLER_407_1261 ();
 FILLCELL_X32 FILLER_407_1264 ();
 FILLCELL_X32 FILLER_407_1296 ();
 FILLCELL_X32 FILLER_407_1328 ();
 FILLCELL_X32 FILLER_407_1360 ();
 FILLCELL_X32 FILLER_407_1392 ();
 FILLCELL_X32 FILLER_407_1424 ();
 FILLCELL_X32 FILLER_407_1456 ();
 FILLCELL_X32 FILLER_407_1488 ();
 FILLCELL_X32 FILLER_407_1520 ();
 FILLCELL_X32 FILLER_407_1552 ();
 FILLCELL_X32 FILLER_407_1584 ();
 FILLCELL_X32 FILLER_407_1616 ();
 FILLCELL_X32 FILLER_407_1648 ();
 FILLCELL_X32 FILLER_407_1680 ();
 FILLCELL_X32 FILLER_407_1712 ();
 FILLCELL_X32 FILLER_407_1744 ();
 FILLCELL_X32 FILLER_407_1776 ();
 FILLCELL_X32 FILLER_407_1808 ();
 FILLCELL_X32 FILLER_407_1840 ();
 FILLCELL_X32 FILLER_407_1872 ();
 FILLCELL_X32 FILLER_407_1904 ();
 FILLCELL_X32 FILLER_407_1936 ();
 FILLCELL_X32 FILLER_407_1968 ();
 FILLCELL_X32 FILLER_407_2000 ();
 FILLCELL_X32 FILLER_407_2032 ();
 FILLCELL_X32 FILLER_407_2064 ();
 FILLCELL_X32 FILLER_407_2096 ();
 FILLCELL_X32 FILLER_407_2128 ();
 FILLCELL_X32 FILLER_407_2160 ();
 FILLCELL_X32 FILLER_407_2192 ();
 FILLCELL_X32 FILLER_407_2224 ();
 FILLCELL_X32 FILLER_407_2256 ();
 FILLCELL_X32 FILLER_407_2288 ();
 FILLCELL_X32 FILLER_407_2320 ();
 FILLCELL_X32 FILLER_407_2352 ();
 FILLCELL_X32 FILLER_407_2384 ();
 FILLCELL_X32 FILLER_407_2416 ();
 FILLCELL_X32 FILLER_407_2448 ();
 FILLCELL_X32 FILLER_407_2480 ();
 FILLCELL_X8 FILLER_407_2512 ();
 FILLCELL_X4 FILLER_407_2520 ();
 FILLCELL_X2 FILLER_407_2524 ();
 FILLCELL_X32 FILLER_407_2527 ();
 FILLCELL_X32 FILLER_407_2559 ();
 FILLCELL_X32 FILLER_407_2591 ();
 FILLCELL_X32 FILLER_407_2623 ();
 FILLCELL_X32 FILLER_407_2655 ();
 FILLCELL_X32 FILLER_407_2687 ();
 FILLCELL_X32 FILLER_407_2719 ();
 FILLCELL_X32 FILLER_407_2751 ();
 FILLCELL_X32 FILLER_407_2783 ();
 FILLCELL_X32 FILLER_407_2815 ();
 FILLCELL_X32 FILLER_407_2847 ();
 FILLCELL_X32 FILLER_407_2879 ();
 FILLCELL_X32 FILLER_407_2911 ();
 FILLCELL_X32 FILLER_407_2943 ();
 FILLCELL_X32 FILLER_407_2975 ();
 FILLCELL_X32 FILLER_407_3007 ();
 FILLCELL_X32 FILLER_407_3039 ();
 FILLCELL_X32 FILLER_407_3071 ();
 FILLCELL_X32 FILLER_407_3103 ();
 FILLCELL_X32 FILLER_407_3135 ();
 FILLCELL_X32 FILLER_407_3167 ();
 FILLCELL_X32 FILLER_407_3199 ();
 FILLCELL_X32 FILLER_407_3231 ();
 FILLCELL_X32 FILLER_407_3263 ();
 FILLCELL_X32 FILLER_407_3295 ();
 FILLCELL_X32 FILLER_407_3327 ();
 FILLCELL_X32 FILLER_407_3359 ();
 FILLCELL_X32 FILLER_407_3391 ();
 FILLCELL_X32 FILLER_407_3423 ();
 FILLCELL_X32 FILLER_407_3455 ();
 FILLCELL_X32 FILLER_407_3487 ();
 FILLCELL_X32 FILLER_407_3519 ();
 FILLCELL_X32 FILLER_407_3551 ();
 FILLCELL_X32 FILLER_407_3583 ();
 FILLCELL_X32 FILLER_407_3615 ();
 FILLCELL_X32 FILLER_407_3647 ();
 FILLCELL_X32 FILLER_407_3679 ();
 FILLCELL_X16 FILLER_407_3711 ();
 FILLCELL_X8 FILLER_407_3727 ();
 FILLCELL_X2 FILLER_407_3735 ();
 FILLCELL_X1 FILLER_407_3737 ();
 FILLCELL_X32 FILLER_408_1 ();
 FILLCELL_X32 FILLER_408_33 ();
 FILLCELL_X32 FILLER_408_65 ();
 FILLCELL_X32 FILLER_408_97 ();
 FILLCELL_X32 FILLER_408_129 ();
 FILLCELL_X32 FILLER_408_161 ();
 FILLCELL_X32 FILLER_408_193 ();
 FILLCELL_X32 FILLER_408_225 ();
 FILLCELL_X32 FILLER_408_257 ();
 FILLCELL_X32 FILLER_408_289 ();
 FILLCELL_X32 FILLER_408_321 ();
 FILLCELL_X32 FILLER_408_353 ();
 FILLCELL_X32 FILLER_408_385 ();
 FILLCELL_X32 FILLER_408_417 ();
 FILLCELL_X32 FILLER_408_449 ();
 FILLCELL_X32 FILLER_408_481 ();
 FILLCELL_X32 FILLER_408_513 ();
 FILLCELL_X32 FILLER_408_545 ();
 FILLCELL_X32 FILLER_408_577 ();
 FILLCELL_X16 FILLER_408_609 ();
 FILLCELL_X4 FILLER_408_625 ();
 FILLCELL_X2 FILLER_408_629 ();
 FILLCELL_X32 FILLER_408_632 ();
 FILLCELL_X32 FILLER_408_664 ();
 FILLCELL_X32 FILLER_408_696 ();
 FILLCELL_X32 FILLER_408_728 ();
 FILLCELL_X32 FILLER_408_760 ();
 FILLCELL_X32 FILLER_408_792 ();
 FILLCELL_X32 FILLER_408_824 ();
 FILLCELL_X32 FILLER_408_856 ();
 FILLCELL_X32 FILLER_408_888 ();
 FILLCELL_X32 FILLER_408_920 ();
 FILLCELL_X32 FILLER_408_952 ();
 FILLCELL_X32 FILLER_408_984 ();
 FILLCELL_X32 FILLER_408_1016 ();
 FILLCELL_X32 FILLER_408_1048 ();
 FILLCELL_X32 FILLER_408_1080 ();
 FILLCELL_X32 FILLER_408_1112 ();
 FILLCELL_X32 FILLER_408_1144 ();
 FILLCELL_X32 FILLER_408_1176 ();
 FILLCELL_X32 FILLER_408_1208 ();
 FILLCELL_X32 FILLER_408_1240 ();
 FILLCELL_X32 FILLER_408_1272 ();
 FILLCELL_X32 FILLER_408_1304 ();
 FILLCELL_X32 FILLER_408_1336 ();
 FILLCELL_X32 FILLER_408_1368 ();
 FILLCELL_X32 FILLER_408_1400 ();
 FILLCELL_X32 FILLER_408_1432 ();
 FILLCELL_X32 FILLER_408_1464 ();
 FILLCELL_X32 FILLER_408_1496 ();
 FILLCELL_X32 FILLER_408_1528 ();
 FILLCELL_X32 FILLER_408_1560 ();
 FILLCELL_X32 FILLER_408_1592 ();
 FILLCELL_X32 FILLER_408_1624 ();
 FILLCELL_X32 FILLER_408_1656 ();
 FILLCELL_X32 FILLER_408_1688 ();
 FILLCELL_X32 FILLER_408_1720 ();
 FILLCELL_X32 FILLER_408_1752 ();
 FILLCELL_X32 FILLER_408_1784 ();
 FILLCELL_X32 FILLER_408_1816 ();
 FILLCELL_X32 FILLER_408_1848 ();
 FILLCELL_X8 FILLER_408_1880 ();
 FILLCELL_X4 FILLER_408_1888 ();
 FILLCELL_X2 FILLER_408_1892 ();
 FILLCELL_X32 FILLER_408_1895 ();
 FILLCELL_X32 FILLER_408_1927 ();
 FILLCELL_X32 FILLER_408_1959 ();
 FILLCELL_X32 FILLER_408_1991 ();
 FILLCELL_X32 FILLER_408_2023 ();
 FILLCELL_X32 FILLER_408_2055 ();
 FILLCELL_X32 FILLER_408_2087 ();
 FILLCELL_X32 FILLER_408_2119 ();
 FILLCELL_X32 FILLER_408_2151 ();
 FILLCELL_X32 FILLER_408_2183 ();
 FILLCELL_X32 FILLER_408_2215 ();
 FILLCELL_X32 FILLER_408_2247 ();
 FILLCELL_X32 FILLER_408_2279 ();
 FILLCELL_X32 FILLER_408_2311 ();
 FILLCELL_X32 FILLER_408_2343 ();
 FILLCELL_X32 FILLER_408_2375 ();
 FILLCELL_X32 FILLER_408_2407 ();
 FILLCELL_X32 FILLER_408_2439 ();
 FILLCELL_X32 FILLER_408_2471 ();
 FILLCELL_X32 FILLER_408_2503 ();
 FILLCELL_X32 FILLER_408_2535 ();
 FILLCELL_X32 FILLER_408_2567 ();
 FILLCELL_X32 FILLER_408_2599 ();
 FILLCELL_X32 FILLER_408_2631 ();
 FILLCELL_X32 FILLER_408_2663 ();
 FILLCELL_X32 FILLER_408_2695 ();
 FILLCELL_X32 FILLER_408_2727 ();
 FILLCELL_X32 FILLER_408_2759 ();
 FILLCELL_X32 FILLER_408_2791 ();
 FILLCELL_X32 FILLER_408_2823 ();
 FILLCELL_X32 FILLER_408_2855 ();
 FILLCELL_X32 FILLER_408_2887 ();
 FILLCELL_X32 FILLER_408_2919 ();
 FILLCELL_X32 FILLER_408_2951 ();
 FILLCELL_X32 FILLER_408_2983 ();
 FILLCELL_X32 FILLER_408_3015 ();
 FILLCELL_X32 FILLER_408_3047 ();
 FILLCELL_X32 FILLER_408_3079 ();
 FILLCELL_X32 FILLER_408_3111 ();
 FILLCELL_X8 FILLER_408_3143 ();
 FILLCELL_X4 FILLER_408_3151 ();
 FILLCELL_X2 FILLER_408_3155 ();
 FILLCELL_X32 FILLER_408_3158 ();
 FILLCELL_X32 FILLER_408_3190 ();
 FILLCELL_X32 FILLER_408_3222 ();
 FILLCELL_X32 FILLER_408_3254 ();
 FILLCELL_X32 FILLER_408_3286 ();
 FILLCELL_X32 FILLER_408_3318 ();
 FILLCELL_X32 FILLER_408_3350 ();
 FILLCELL_X32 FILLER_408_3382 ();
 FILLCELL_X32 FILLER_408_3414 ();
 FILLCELL_X32 FILLER_408_3446 ();
 FILLCELL_X32 FILLER_408_3478 ();
 FILLCELL_X32 FILLER_408_3510 ();
 FILLCELL_X32 FILLER_408_3542 ();
 FILLCELL_X32 FILLER_408_3574 ();
 FILLCELL_X32 FILLER_408_3606 ();
 FILLCELL_X32 FILLER_408_3638 ();
 FILLCELL_X32 FILLER_408_3670 ();
 FILLCELL_X32 FILLER_408_3702 ();
 FILLCELL_X4 FILLER_408_3734 ();
 FILLCELL_X32 FILLER_409_1 ();
 FILLCELL_X32 FILLER_409_33 ();
 FILLCELL_X32 FILLER_409_65 ();
 FILLCELL_X32 FILLER_409_97 ();
 FILLCELL_X32 FILLER_409_129 ();
 FILLCELL_X32 FILLER_409_161 ();
 FILLCELL_X32 FILLER_409_193 ();
 FILLCELL_X32 FILLER_409_225 ();
 FILLCELL_X32 FILLER_409_257 ();
 FILLCELL_X32 FILLER_409_289 ();
 FILLCELL_X32 FILLER_409_321 ();
 FILLCELL_X32 FILLER_409_353 ();
 FILLCELL_X32 FILLER_409_385 ();
 FILLCELL_X32 FILLER_409_417 ();
 FILLCELL_X32 FILLER_409_449 ();
 FILLCELL_X32 FILLER_409_481 ();
 FILLCELL_X32 FILLER_409_513 ();
 FILLCELL_X32 FILLER_409_545 ();
 FILLCELL_X32 FILLER_409_577 ();
 FILLCELL_X32 FILLER_409_609 ();
 FILLCELL_X32 FILLER_409_641 ();
 FILLCELL_X32 FILLER_409_673 ();
 FILLCELL_X32 FILLER_409_705 ();
 FILLCELL_X32 FILLER_409_737 ();
 FILLCELL_X32 FILLER_409_769 ();
 FILLCELL_X32 FILLER_409_801 ();
 FILLCELL_X32 FILLER_409_833 ();
 FILLCELL_X32 FILLER_409_865 ();
 FILLCELL_X32 FILLER_409_897 ();
 FILLCELL_X32 FILLER_409_929 ();
 FILLCELL_X32 FILLER_409_961 ();
 FILLCELL_X32 FILLER_409_993 ();
 FILLCELL_X32 FILLER_409_1025 ();
 FILLCELL_X32 FILLER_409_1057 ();
 FILLCELL_X32 FILLER_409_1089 ();
 FILLCELL_X32 FILLER_409_1121 ();
 FILLCELL_X32 FILLER_409_1153 ();
 FILLCELL_X32 FILLER_409_1185 ();
 FILLCELL_X32 FILLER_409_1217 ();
 FILLCELL_X8 FILLER_409_1249 ();
 FILLCELL_X4 FILLER_409_1257 ();
 FILLCELL_X2 FILLER_409_1261 ();
 FILLCELL_X32 FILLER_409_1264 ();
 FILLCELL_X32 FILLER_409_1296 ();
 FILLCELL_X32 FILLER_409_1328 ();
 FILLCELL_X32 FILLER_409_1360 ();
 FILLCELL_X32 FILLER_409_1392 ();
 FILLCELL_X32 FILLER_409_1424 ();
 FILLCELL_X32 FILLER_409_1456 ();
 FILLCELL_X32 FILLER_409_1488 ();
 FILLCELL_X32 FILLER_409_1520 ();
 FILLCELL_X32 FILLER_409_1552 ();
 FILLCELL_X32 FILLER_409_1584 ();
 FILLCELL_X32 FILLER_409_1616 ();
 FILLCELL_X32 FILLER_409_1648 ();
 FILLCELL_X32 FILLER_409_1680 ();
 FILLCELL_X32 FILLER_409_1712 ();
 FILLCELL_X32 FILLER_409_1744 ();
 FILLCELL_X32 FILLER_409_1776 ();
 FILLCELL_X32 FILLER_409_1808 ();
 FILLCELL_X32 FILLER_409_1840 ();
 FILLCELL_X32 FILLER_409_1872 ();
 FILLCELL_X32 FILLER_409_1904 ();
 FILLCELL_X32 FILLER_409_1936 ();
 FILLCELL_X32 FILLER_409_1968 ();
 FILLCELL_X32 FILLER_409_2000 ();
 FILLCELL_X32 FILLER_409_2032 ();
 FILLCELL_X32 FILLER_409_2064 ();
 FILLCELL_X32 FILLER_409_2096 ();
 FILLCELL_X32 FILLER_409_2128 ();
 FILLCELL_X32 FILLER_409_2160 ();
 FILLCELL_X32 FILLER_409_2192 ();
 FILLCELL_X32 FILLER_409_2224 ();
 FILLCELL_X32 FILLER_409_2256 ();
 FILLCELL_X32 FILLER_409_2288 ();
 FILLCELL_X32 FILLER_409_2320 ();
 FILLCELL_X32 FILLER_409_2352 ();
 FILLCELL_X32 FILLER_409_2384 ();
 FILLCELL_X32 FILLER_409_2416 ();
 FILLCELL_X32 FILLER_409_2448 ();
 FILLCELL_X32 FILLER_409_2480 ();
 FILLCELL_X8 FILLER_409_2512 ();
 FILLCELL_X4 FILLER_409_2520 ();
 FILLCELL_X2 FILLER_409_2524 ();
 FILLCELL_X32 FILLER_409_2527 ();
 FILLCELL_X32 FILLER_409_2559 ();
 FILLCELL_X32 FILLER_409_2591 ();
 FILLCELL_X32 FILLER_409_2623 ();
 FILLCELL_X32 FILLER_409_2655 ();
 FILLCELL_X32 FILLER_409_2687 ();
 FILLCELL_X32 FILLER_409_2719 ();
 FILLCELL_X32 FILLER_409_2751 ();
 FILLCELL_X32 FILLER_409_2783 ();
 FILLCELL_X32 FILLER_409_2815 ();
 FILLCELL_X32 FILLER_409_2847 ();
 FILLCELL_X32 FILLER_409_2879 ();
 FILLCELL_X32 FILLER_409_2911 ();
 FILLCELL_X32 FILLER_409_2943 ();
 FILLCELL_X32 FILLER_409_2975 ();
 FILLCELL_X32 FILLER_409_3007 ();
 FILLCELL_X32 FILLER_409_3039 ();
 FILLCELL_X32 FILLER_409_3071 ();
 FILLCELL_X32 FILLER_409_3103 ();
 FILLCELL_X32 FILLER_409_3135 ();
 FILLCELL_X32 FILLER_409_3167 ();
 FILLCELL_X32 FILLER_409_3199 ();
 FILLCELL_X32 FILLER_409_3231 ();
 FILLCELL_X32 FILLER_409_3263 ();
 FILLCELL_X32 FILLER_409_3295 ();
 FILLCELL_X32 FILLER_409_3327 ();
 FILLCELL_X32 FILLER_409_3359 ();
 FILLCELL_X32 FILLER_409_3391 ();
 FILLCELL_X32 FILLER_409_3423 ();
 FILLCELL_X32 FILLER_409_3455 ();
 FILLCELL_X32 FILLER_409_3487 ();
 FILLCELL_X32 FILLER_409_3519 ();
 FILLCELL_X32 FILLER_409_3551 ();
 FILLCELL_X32 FILLER_409_3583 ();
 FILLCELL_X32 FILLER_409_3615 ();
 FILLCELL_X32 FILLER_409_3647 ();
 FILLCELL_X32 FILLER_409_3679 ();
 FILLCELL_X16 FILLER_409_3711 ();
 FILLCELL_X8 FILLER_409_3727 ();
 FILLCELL_X2 FILLER_409_3735 ();
 FILLCELL_X1 FILLER_409_3737 ();
 FILLCELL_X32 FILLER_410_1 ();
 FILLCELL_X32 FILLER_410_33 ();
 FILLCELL_X32 FILLER_410_65 ();
 FILLCELL_X32 FILLER_410_97 ();
 FILLCELL_X32 FILLER_410_129 ();
 FILLCELL_X32 FILLER_410_161 ();
 FILLCELL_X32 FILLER_410_193 ();
 FILLCELL_X32 FILLER_410_225 ();
 FILLCELL_X32 FILLER_410_257 ();
 FILLCELL_X32 FILLER_410_289 ();
 FILLCELL_X32 FILLER_410_321 ();
 FILLCELL_X32 FILLER_410_353 ();
 FILLCELL_X32 FILLER_410_385 ();
 FILLCELL_X32 FILLER_410_417 ();
 FILLCELL_X32 FILLER_410_449 ();
 FILLCELL_X32 FILLER_410_481 ();
 FILLCELL_X32 FILLER_410_513 ();
 FILLCELL_X32 FILLER_410_545 ();
 FILLCELL_X32 FILLER_410_577 ();
 FILLCELL_X16 FILLER_410_609 ();
 FILLCELL_X4 FILLER_410_625 ();
 FILLCELL_X2 FILLER_410_629 ();
 FILLCELL_X32 FILLER_410_632 ();
 FILLCELL_X32 FILLER_410_664 ();
 FILLCELL_X32 FILLER_410_696 ();
 FILLCELL_X32 FILLER_410_728 ();
 FILLCELL_X32 FILLER_410_760 ();
 FILLCELL_X32 FILLER_410_792 ();
 FILLCELL_X32 FILLER_410_824 ();
 FILLCELL_X32 FILLER_410_856 ();
 FILLCELL_X32 FILLER_410_888 ();
 FILLCELL_X32 FILLER_410_920 ();
 FILLCELL_X32 FILLER_410_952 ();
 FILLCELL_X32 FILLER_410_984 ();
 FILLCELL_X32 FILLER_410_1016 ();
 FILLCELL_X32 FILLER_410_1048 ();
 FILLCELL_X32 FILLER_410_1080 ();
 FILLCELL_X32 FILLER_410_1112 ();
 FILLCELL_X32 FILLER_410_1144 ();
 FILLCELL_X32 FILLER_410_1176 ();
 FILLCELL_X32 FILLER_410_1208 ();
 FILLCELL_X32 FILLER_410_1240 ();
 FILLCELL_X32 FILLER_410_1272 ();
 FILLCELL_X32 FILLER_410_1304 ();
 FILLCELL_X32 FILLER_410_1336 ();
 FILLCELL_X32 FILLER_410_1368 ();
 FILLCELL_X32 FILLER_410_1400 ();
 FILLCELL_X32 FILLER_410_1432 ();
 FILLCELL_X32 FILLER_410_1464 ();
 FILLCELL_X32 FILLER_410_1496 ();
 FILLCELL_X32 FILLER_410_1528 ();
 FILLCELL_X32 FILLER_410_1560 ();
 FILLCELL_X32 FILLER_410_1592 ();
 FILLCELL_X32 FILLER_410_1624 ();
 FILLCELL_X32 FILLER_410_1656 ();
 FILLCELL_X32 FILLER_410_1688 ();
 FILLCELL_X32 FILLER_410_1720 ();
 FILLCELL_X32 FILLER_410_1752 ();
 FILLCELL_X32 FILLER_410_1784 ();
 FILLCELL_X32 FILLER_410_1816 ();
 FILLCELL_X32 FILLER_410_1848 ();
 FILLCELL_X8 FILLER_410_1880 ();
 FILLCELL_X4 FILLER_410_1888 ();
 FILLCELL_X2 FILLER_410_1892 ();
 FILLCELL_X32 FILLER_410_1895 ();
 FILLCELL_X32 FILLER_410_1927 ();
 FILLCELL_X32 FILLER_410_1959 ();
 FILLCELL_X32 FILLER_410_1991 ();
 FILLCELL_X32 FILLER_410_2023 ();
 FILLCELL_X32 FILLER_410_2055 ();
 FILLCELL_X32 FILLER_410_2087 ();
 FILLCELL_X32 FILLER_410_2119 ();
 FILLCELL_X32 FILLER_410_2151 ();
 FILLCELL_X32 FILLER_410_2183 ();
 FILLCELL_X32 FILLER_410_2215 ();
 FILLCELL_X32 FILLER_410_2247 ();
 FILLCELL_X32 FILLER_410_2279 ();
 FILLCELL_X32 FILLER_410_2311 ();
 FILLCELL_X32 FILLER_410_2343 ();
 FILLCELL_X32 FILLER_410_2375 ();
 FILLCELL_X32 FILLER_410_2407 ();
 FILLCELL_X32 FILLER_410_2439 ();
 FILLCELL_X32 FILLER_410_2471 ();
 FILLCELL_X32 FILLER_410_2503 ();
 FILLCELL_X32 FILLER_410_2535 ();
 FILLCELL_X32 FILLER_410_2567 ();
 FILLCELL_X32 FILLER_410_2599 ();
 FILLCELL_X32 FILLER_410_2631 ();
 FILLCELL_X32 FILLER_410_2663 ();
 FILLCELL_X32 FILLER_410_2695 ();
 FILLCELL_X32 FILLER_410_2727 ();
 FILLCELL_X32 FILLER_410_2759 ();
 FILLCELL_X32 FILLER_410_2791 ();
 FILLCELL_X32 FILLER_410_2823 ();
 FILLCELL_X32 FILLER_410_2855 ();
 FILLCELL_X32 FILLER_410_2887 ();
 FILLCELL_X32 FILLER_410_2919 ();
 FILLCELL_X32 FILLER_410_2951 ();
 FILLCELL_X32 FILLER_410_2983 ();
 FILLCELL_X32 FILLER_410_3015 ();
 FILLCELL_X32 FILLER_410_3047 ();
 FILLCELL_X32 FILLER_410_3079 ();
 FILLCELL_X32 FILLER_410_3111 ();
 FILLCELL_X8 FILLER_410_3143 ();
 FILLCELL_X4 FILLER_410_3151 ();
 FILLCELL_X2 FILLER_410_3155 ();
 FILLCELL_X32 FILLER_410_3158 ();
 FILLCELL_X32 FILLER_410_3190 ();
 FILLCELL_X32 FILLER_410_3222 ();
 FILLCELL_X32 FILLER_410_3254 ();
 FILLCELL_X32 FILLER_410_3286 ();
 FILLCELL_X32 FILLER_410_3318 ();
 FILLCELL_X32 FILLER_410_3350 ();
 FILLCELL_X32 FILLER_410_3382 ();
 FILLCELL_X32 FILLER_410_3414 ();
 FILLCELL_X32 FILLER_410_3446 ();
 FILLCELL_X32 FILLER_410_3478 ();
 FILLCELL_X32 FILLER_410_3510 ();
 FILLCELL_X32 FILLER_410_3542 ();
 FILLCELL_X32 FILLER_410_3574 ();
 FILLCELL_X32 FILLER_410_3606 ();
 FILLCELL_X32 FILLER_410_3638 ();
 FILLCELL_X32 FILLER_410_3670 ();
 FILLCELL_X32 FILLER_410_3702 ();
 FILLCELL_X4 FILLER_410_3734 ();
 FILLCELL_X32 FILLER_411_1 ();
 FILLCELL_X32 FILLER_411_33 ();
 FILLCELL_X32 FILLER_411_65 ();
 FILLCELL_X32 FILLER_411_97 ();
 FILLCELL_X32 FILLER_411_129 ();
 FILLCELL_X32 FILLER_411_161 ();
 FILLCELL_X32 FILLER_411_193 ();
 FILLCELL_X32 FILLER_411_225 ();
 FILLCELL_X32 FILLER_411_257 ();
 FILLCELL_X32 FILLER_411_289 ();
 FILLCELL_X32 FILLER_411_321 ();
 FILLCELL_X32 FILLER_411_353 ();
 FILLCELL_X32 FILLER_411_385 ();
 FILLCELL_X32 FILLER_411_417 ();
 FILLCELL_X32 FILLER_411_449 ();
 FILLCELL_X32 FILLER_411_481 ();
 FILLCELL_X32 FILLER_411_513 ();
 FILLCELL_X32 FILLER_411_545 ();
 FILLCELL_X32 FILLER_411_577 ();
 FILLCELL_X32 FILLER_411_609 ();
 FILLCELL_X32 FILLER_411_641 ();
 FILLCELL_X32 FILLER_411_673 ();
 FILLCELL_X32 FILLER_411_705 ();
 FILLCELL_X32 FILLER_411_737 ();
 FILLCELL_X32 FILLER_411_769 ();
 FILLCELL_X32 FILLER_411_801 ();
 FILLCELL_X32 FILLER_411_833 ();
 FILLCELL_X32 FILLER_411_865 ();
 FILLCELL_X32 FILLER_411_897 ();
 FILLCELL_X32 FILLER_411_929 ();
 FILLCELL_X32 FILLER_411_961 ();
 FILLCELL_X32 FILLER_411_993 ();
 FILLCELL_X32 FILLER_411_1025 ();
 FILLCELL_X32 FILLER_411_1057 ();
 FILLCELL_X32 FILLER_411_1089 ();
 FILLCELL_X32 FILLER_411_1121 ();
 FILLCELL_X32 FILLER_411_1153 ();
 FILLCELL_X32 FILLER_411_1185 ();
 FILLCELL_X32 FILLER_411_1217 ();
 FILLCELL_X8 FILLER_411_1249 ();
 FILLCELL_X4 FILLER_411_1257 ();
 FILLCELL_X2 FILLER_411_1261 ();
 FILLCELL_X32 FILLER_411_1264 ();
 FILLCELL_X32 FILLER_411_1296 ();
 FILLCELL_X32 FILLER_411_1328 ();
 FILLCELL_X32 FILLER_411_1360 ();
 FILLCELL_X32 FILLER_411_1392 ();
 FILLCELL_X32 FILLER_411_1424 ();
 FILLCELL_X32 FILLER_411_1456 ();
 FILLCELL_X32 FILLER_411_1488 ();
 FILLCELL_X32 FILLER_411_1520 ();
 FILLCELL_X32 FILLER_411_1552 ();
 FILLCELL_X32 FILLER_411_1584 ();
 FILLCELL_X32 FILLER_411_1616 ();
 FILLCELL_X32 FILLER_411_1648 ();
 FILLCELL_X32 FILLER_411_1680 ();
 FILLCELL_X32 FILLER_411_1712 ();
 FILLCELL_X32 FILLER_411_1744 ();
 FILLCELL_X32 FILLER_411_1776 ();
 FILLCELL_X32 FILLER_411_1808 ();
 FILLCELL_X32 FILLER_411_1840 ();
 FILLCELL_X32 FILLER_411_1872 ();
 FILLCELL_X32 FILLER_411_1904 ();
 FILLCELL_X32 FILLER_411_1936 ();
 FILLCELL_X32 FILLER_411_1968 ();
 FILLCELL_X32 FILLER_411_2000 ();
 FILLCELL_X32 FILLER_411_2032 ();
 FILLCELL_X32 FILLER_411_2064 ();
 FILLCELL_X32 FILLER_411_2096 ();
 FILLCELL_X32 FILLER_411_2128 ();
 FILLCELL_X32 FILLER_411_2160 ();
 FILLCELL_X32 FILLER_411_2192 ();
 FILLCELL_X32 FILLER_411_2224 ();
 FILLCELL_X32 FILLER_411_2256 ();
 FILLCELL_X32 FILLER_411_2288 ();
 FILLCELL_X32 FILLER_411_2320 ();
 FILLCELL_X32 FILLER_411_2352 ();
 FILLCELL_X32 FILLER_411_2384 ();
 FILLCELL_X32 FILLER_411_2416 ();
 FILLCELL_X32 FILLER_411_2448 ();
 FILLCELL_X32 FILLER_411_2480 ();
 FILLCELL_X8 FILLER_411_2512 ();
 FILLCELL_X4 FILLER_411_2520 ();
 FILLCELL_X2 FILLER_411_2524 ();
 FILLCELL_X32 FILLER_411_2527 ();
 FILLCELL_X32 FILLER_411_2559 ();
 FILLCELL_X32 FILLER_411_2591 ();
 FILLCELL_X32 FILLER_411_2623 ();
 FILLCELL_X32 FILLER_411_2655 ();
 FILLCELL_X32 FILLER_411_2687 ();
 FILLCELL_X32 FILLER_411_2719 ();
 FILLCELL_X32 FILLER_411_2751 ();
 FILLCELL_X32 FILLER_411_2783 ();
 FILLCELL_X32 FILLER_411_2815 ();
 FILLCELL_X32 FILLER_411_2847 ();
 FILLCELL_X32 FILLER_411_2879 ();
 FILLCELL_X32 FILLER_411_2911 ();
 FILLCELL_X32 FILLER_411_2943 ();
 FILLCELL_X32 FILLER_411_2975 ();
 FILLCELL_X32 FILLER_411_3007 ();
 FILLCELL_X32 FILLER_411_3039 ();
 FILLCELL_X32 FILLER_411_3071 ();
 FILLCELL_X32 FILLER_411_3103 ();
 FILLCELL_X32 FILLER_411_3135 ();
 FILLCELL_X32 FILLER_411_3167 ();
 FILLCELL_X32 FILLER_411_3199 ();
 FILLCELL_X32 FILLER_411_3231 ();
 FILLCELL_X32 FILLER_411_3263 ();
 FILLCELL_X32 FILLER_411_3295 ();
 FILLCELL_X32 FILLER_411_3327 ();
 FILLCELL_X32 FILLER_411_3359 ();
 FILLCELL_X32 FILLER_411_3391 ();
 FILLCELL_X32 FILLER_411_3423 ();
 FILLCELL_X32 FILLER_411_3455 ();
 FILLCELL_X32 FILLER_411_3487 ();
 FILLCELL_X32 FILLER_411_3519 ();
 FILLCELL_X32 FILLER_411_3551 ();
 FILLCELL_X32 FILLER_411_3583 ();
 FILLCELL_X32 FILLER_411_3615 ();
 FILLCELL_X32 FILLER_411_3647 ();
 FILLCELL_X32 FILLER_411_3679 ();
 FILLCELL_X16 FILLER_411_3711 ();
 FILLCELL_X8 FILLER_411_3727 ();
 FILLCELL_X2 FILLER_411_3735 ();
 FILLCELL_X1 FILLER_411_3737 ();
 FILLCELL_X32 FILLER_412_1 ();
 FILLCELL_X32 FILLER_412_33 ();
 FILLCELL_X32 FILLER_412_65 ();
 FILLCELL_X32 FILLER_412_97 ();
 FILLCELL_X32 FILLER_412_129 ();
 FILLCELL_X32 FILLER_412_161 ();
 FILLCELL_X32 FILLER_412_193 ();
 FILLCELL_X32 FILLER_412_225 ();
 FILLCELL_X32 FILLER_412_257 ();
 FILLCELL_X32 FILLER_412_289 ();
 FILLCELL_X32 FILLER_412_321 ();
 FILLCELL_X32 FILLER_412_353 ();
 FILLCELL_X32 FILLER_412_385 ();
 FILLCELL_X32 FILLER_412_417 ();
 FILLCELL_X32 FILLER_412_449 ();
 FILLCELL_X32 FILLER_412_481 ();
 FILLCELL_X32 FILLER_412_513 ();
 FILLCELL_X32 FILLER_412_545 ();
 FILLCELL_X32 FILLER_412_577 ();
 FILLCELL_X16 FILLER_412_609 ();
 FILLCELL_X4 FILLER_412_625 ();
 FILLCELL_X2 FILLER_412_629 ();
 FILLCELL_X32 FILLER_412_632 ();
 FILLCELL_X32 FILLER_412_664 ();
 FILLCELL_X32 FILLER_412_696 ();
 FILLCELL_X32 FILLER_412_728 ();
 FILLCELL_X32 FILLER_412_760 ();
 FILLCELL_X32 FILLER_412_792 ();
 FILLCELL_X32 FILLER_412_824 ();
 FILLCELL_X32 FILLER_412_856 ();
 FILLCELL_X32 FILLER_412_888 ();
 FILLCELL_X32 FILLER_412_920 ();
 FILLCELL_X32 FILLER_412_952 ();
 FILLCELL_X32 FILLER_412_984 ();
 FILLCELL_X32 FILLER_412_1016 ();
 FILLCELL_X32 FILLER_412_1048 ();
 FILLCELL_X32 FILLER_412_1080 ();
 FILLCELL_X32 FILLER_412_1112 ();
 FILLCELL_X32 FILLER_412_1144 ();
 FILLCELL_X32 FILLER_412_1176 ();
 FILLCELL_X32 FILLER_412_1208 ();
 FILLCELL_X32 FILLER_412_1240 ();
 FILLCELL_X32 FILLER_412_1272 ();
 FILLCELL_X32 FILLER_412_1304 ();
 FILLCELL_X32 FILLER_412_1336 ();
 FILLCELL_X32 FILLER_412_1368 ();
 FILLCELL_X32 FILLER_412_1400 ();
 FILLCELL_X32 FILLER_412_1432 ();
 FILLCELL_X32 FILLER_412_1464 ();
 FILLCELL_X32 FILLER_412_1496 ();
 FILLCELL_X32 FILLER_412_1528 ();
 FILLCELL_X32 FILLER_412_1560 ();
 FILLCELL_X32 FILLER_412_1592 ();
 FILLCELL_X32 FILLER_412_1624 ();
 FILLCELL_X32 FILLER_412_1656 ();
 FILLCELL_X32 FILLER_412_1688 ();
 FILLCELL_X32 FILLER_412_1720 ();
 FILLCELL_X32 FILLER_412_1752 ();
 FILLCELL_X32 FILLER_412_1784 ();
 FILLCELL_X32 FILLER_412_1816 ();
 FILLCELL_X32 FILLER_412_1848 ();
 FILLCELL_X8 FILLER_412_1880 ();
 FILLCELL_X4 FILLER_412_1888 ();
 FILLCELL_X2 FILLER_412_1892 ();
 FILLCELL_X32 FILLER_412_1895 ();
 FILLCELL_X32 FILLER_412_1927 ();
 FILLCELL_X32 FILLER_412_1959 ();
 FILLCELL_X32 FILLER_412_1991 ();
 FILLCELL_X32 FILLER_412_2023 ();
 FILLCELL_X32 FILLER_412_2055 ();
 FILLCELL_X32 FILLER_412_2087 ();
 FILLCELL_X32 FILLER_412_2119 ();
 FILLCELL_X32 FILLER_412_2151 ();
 FILLCELL_X32 FILLER_412_2183 ();
 FILLCELL_X32 FILLER_412_2215 ();
 FILLCELL_X32 FILLER_412_2247 ();
 FILLCELL_X32 FILLER_412_2279 ();
 FILLCELL_X32 FILLER_412_2311 ();
 FILLCELL_X32 FILLER_412_2343 ();
 FILLCELL_X32 FILLER_412_2375 ();
 FILLCELL_X32 FILLER_412_2407 ();
 FILLCELL_X32 FILLER_412_2439 ();
 FILLCELL_X32 FILLER_412_2471 ();
 FILLCELL_X32 FILLER_412_2503 ();
 FILLCELL_X32 FILLER_412_2535 ();
 FILLCELL_X32 FILLER_412_2567 ();
 FILLCELL_X32 FILLER_412_2599 ();
 FILLCELL_X32 FILLER_412_2631 ();
 FILLCELL_X32 FILLER_412_2663 ();
 FILLCELL_X32 FILLER_412_2695 ();
 FILLCELL_X32 FILLER_412_2727 ();
 FILLCELL_X32 FILLER_412_2759 ();
 FILLCELL_X32 FILLER_412_2791 ();
 FILLCELL_X32 FILLER_412_2823 ();
 FILLCELL_X32 FILLER_412_2855 ();
 FILLCELL_X32 FILLER_412_2887 ();
 FILLCELL_X32 FILLER_412_2919 ();
 FILLCELL_X32 FILLER_412_2951 ();
 FILLCELL_X32 FILLER_412_2983 ();
 FILLCELL_X32 FILLER_412_3015 ();
 FILLCELL_X32 FILLER_412_3047 ();
 FILLCELL_X32 FILLER_412_3079 ();
 FILLCELL_X32 FILLER_412_3111 ();
 FILLCELL_X8 FILLER_412_3143 ();
 FILLCELL_X4 FILLER_412_3151 ();
 FILLCELL_X2 FILLER_412_3155 ();
 FILLCELL_X32 FILLER_412_3158 ();
 FILLCELL_X32 FILLER_412_3190 ();
 FILLCELL_X32 FILLER_412_3222 ();
 FILLCELL_X32 FILLER_412_3254 ();
 FILLCELL_X32 FILLER_412_3286 ();
 FILLCELL_X32 FILLER_412_3318 ();
 FILLCELL_X32 FILLER_412_3350 ();
 FILLCELL_X32 FILLER_412_3382 ();
 FILLCELL_X32 FILLER_412_3414 ();
 FILLCELL_X32 FILLER_412_3446 ();
 FILLCELL_X32 FILLER_412_3478 ();
 FILLCELL_X32 FILLER_412_3510 ();
 FILLCELL_X32 FILLER_412_3542 ();
 FILLCELL_X32 FILLER_412_3574 ();
 FILLCELL_X32 FILLER_412_3606 ();
 FILLCELL_X32 FILLER_412_3638 ();
 FILLCELL_X32 FILLER_412_3670 ();
 FILLCELL_X32 FILLER_412_3702 ();
 FILLCELL_X4 FILLER_412_3734 ();
 FILLCELL_X32 FILLER_413_1 ();
 FILLCELL_X32 FILLER_413_33 ();
 FILLCELL_X32 FILLER_413_65 ();
 FILLCELL_X32 FILLER_413_97 ();
 FILLCELL_X32 FILLER_413_129 ();
 FILLCELL_X32 FILLER_413_161 ();
 FILLCELL_X32 FILLER_413_193 ();
 FILLCELL_X32 FILLER_413_225 ();
 FILLCELL_X32 FILLER_413_257 ();
 FILLCELL_X32 FILLER_413_289 ();
 FILLCELL_X32 FILLER_413_321 ();
 FILLCELL_X32 FILLER_413_353 ();
 FILLCELL_X32 FILLER_413_385 ();
 FILLCELL_X32 FILLER_413_417 ();
 FILLCELL_X32 FILLER_413_449 ();
 FILLCELL_X32 FILLER_413_481 ();
 FILLCELL_X32 FILLER_413_513 ();
 FILLCELL_X32 FILLER_413_545 ();
 FILLCELL_X32 FILLER_413_577 ();
 FILLCELL_X32 FILLER_413_609 ();
 FILLCELL_X32 FILLER_413_641 ();
 FILLCELL_X32 FILLER_413_673 ();
 FILLCELL_X32 FILLER_413_705 ();
 FILLCELL_X32 FILLER_413_737 ();
 FILLCELL_X32 FILLER_413_769 ();
 FILLCELL_X32 FILLER_413_801 ();
 FILLCELL_X32 FILLER_413_833 ();
 FILLCELL_X32 FILLER_413_865 ();
 FILLCELL_X32 FILLER_413_897 ();
 FILLCELL_X32 FILLER_413_929 ();
 FILLCELL_X32 FILLER_413_961 ();
 FILLCELL_X32 FILLER_413_993 ();
 FILLCELL_X32 FILLER_413_1025 ();
 FILLCELL_X32 FILLER_413_1057 ();
 FILLCELL_X32 FILLER_413_1089 ();
 FILLCELL_X32 FILLER_413_1121 ();
 FILLCELL_X32 FILLER_413_1153 ();
 FILLCELL_X32 FILLER_413_1185 ();
 FILLCELL_X32 FILLER_413_1217 ();
 FILLCELL_X8 FILLER_413_1249 ();
 FILLCELL_X4 FILLER_413_1257 ();
 FILLCELL_X2 FILLER_413_1261 ();
 FILLCELL_X32 FILLER_413_1264 ();
 FILLCELL_X32 FILLER_413_1296 ();
 FILLCELL_X32 FILLER_413_1328 ();
 FILLCELL_X32 FILLER_413_1360 ();
 FILLCELL_X32 FILLER_413_1392 ();
 FILLCELL_X32 FILLER_413_1424 ();
 FILLCELL_X32 FILLER_413_1456 ();
 FILLCELL_X32 FILLER_413_1488 ();
 FILLCELL_X32 FILLER_413_1520 ();
 FILLCELL_X32 FILLER_413_1552 ();
 FILLCELL_X32 FILLER_413_1584 ();
 FILLCELL_X32 FILLER_413_1616 ();
 FILLCELL_X32 FILLER_413_1648 ();
 FILLCELL_X32 FILLER_413_1680 ();
 FILLCELL_X32 FILLER_413_1712 ();
 FILLCELL_X32 FILLER_413_1744 ();
 FILLCELL_X32 FILLER_413_1776 ();
 FILLCELL_X32 FILLER_413_1808 ();
 FILLCELL_X32 FILLER_413_1840 ();
 FILLCELL_X32 FILLER_413_1872 ();
 FILLCELL_X32 FILLER_413_1904 ();
 FILLCELL_X32 FILLER_413_1936 ();
 FILLCELL_X32 FILLER_413_1968 ();
 FILLCELL_X32 FILLER_413_2000 ();
 FILLCELL_X32 FILLER_413_2032 ();
 FILLCELL_X32 FILLER_413_2064 ();
 FILLCELL_X32 FILLER_413_2096 ();
 FILLCELL_X32 FILLER_413_2128 ();
 FILLCELL_X32 FILLER_413_2160 ();
 FILLCELL_X32 FILLER_413_2192 ();
 FILLCELL_X32 FILLER_413_2224 ();
 FILLCELL_X32 FILLER_413_2256 ();
 FILLCELL_X32 FILLER_413_2288 ();
 FILLCELL_X32 FILLER_413_2320 ();
 FILLCELL_X32 FILLER_413_2352 ();
 FILLCELL_X32 FILLER_413_2384 ();
 FILLCELL_X32 FILLER_413_2416 ();
 FILLCELL_X32 FILLER_413_2448 ();
 FILLCELL_X32 FILLER_413_2480 ();
 FILLCELL_X8 FILLER_413_2512 ();
 FILLCELL_X4 FILLER_413_2520 ();
 FILLCELL_X2 FILLER_413_2524 ();
 FILLCELL_X32 FILLER_413_2527 ();
 FILLCELL_X32 FILLER_413_2559 ();
 FILLCELL_X32 FILLER_413_2591 ();
 FILLCELL_X32 FILLER_413_2623 ();
 FILLCELL_X32 FILLER_413_2655 ();
 FILLCELL_X32 FILLER_413_2687 ();
 FILLCELL_X32 FILLER_413_2719 ();
 FILLCELL_X32 FILLER_413_2751 ();
 FILLCELL_X32 FILLER_413_2783 ();
 FILLCELL_X32 FILLER_413_2815 ();
 FILLCELL_X32 FILLER_413_2847 ();
 FILLCELL_X32 FILLER_413_2879 ();
 FILLCELL_X32 FILLER_413_2911 ();
 FILLCELL_X32 FILLER_413_2943 ();
 FILLCELL_X32 FILLER_413_2975 ();
 FILLCELL_X32 FILLER_413_3007 ();
 FILLCELL_X32 FILLER_413_3039 ();
 FILLCELL_X32 FILLER_413_3071 ();
 FILLCELL_X32 FILLER_413_3103 ();
 FILLCELL_X32 FILLER_413_3135 ();
 FILLCELL_X32 FILLER_413_3167 ();
 FILLCELL_X32 FILLER_413_3199 ();
 FILLCELL_X32 FILLER_413_3231 ();
 FILLCELL_X32 FILLER_413_3263 ();
 FILLCELL_X32 FILLER_413_3295 ();
 FILLCELL_X32 FILLER_413_3327 ();
 FILLCELL_X32 FILLER_413_3359 ();
 FILLCELL_X32 FILLER_413_3391 ();
 FILLCELL_X32 FILLER_413_3423 ();
 FILLCELL_X32 FILLER_413_3455 ();
 FILLCELL_X32 FILLER_413_3487 ();
 FILLCELL_X32 FILLER_413_3519 ();
 FILLCELL_X32 FILLER_413_3551 ();
 FILLCELL_X32 FILLER_413_3583 ();
 FILLCELL_X32 FILLER_413_3615 ();
 FILLCELL_X32 FILLER_413_3647 ();
 FILLCELL_X32 FILLER_413_3679 ();
 FILLCELL_X16 FILLER_413_3711 ();
 FILLCELL_X8 FILLER_413_3727 ();
 FILLCELL_X2 FILLER_413_3735 ();
 FILLCELL_X1 FILLER_413_3737 ();
 FILLCELL_X32 FILLER_414_1 ();
 FILLCELL_X32 FILLER_414_33 ();
 FILLCELL_X32 FILLER_414_65 ();
 FILLCELL_X32 FILLER_414_97 ();
 FILLCELL_X32 FILLER_414_129 ();
 FILLCELL_X32 FILLER_414_161 ();
 FILLCELL_X32 FILLER_414_193 ();
 FILLCELL_X32 FILLER_414_225 ();
 FILLCELL_X32 FILLER_414_257 ();
 FILLCELL_X32 FILLER_414_289 ();
 FILLCELL_X32 FILLER_414_321 ();
 FILLCELL_X32 FILLER_414_353 ();
 FILLCELL_X32 FILLER_414_385 ();
 FILLCELL_X32 FILLER_414_417 ();
 FILLCELL_X32 FILLER_414_449 ();
 FILLCELL_X32 FILLER_414_481 ();
 FILLCELL_X32 FILLER_414_513 ();
 FILLCELL_X32 FILLER_414_545 ();
 FILLCELL_X32 FILLER_414_577 ();
 FILLCELL_X16 FILLER_414_609 ();
 FILLCELL_X4 FILLER_414_625 ();
 FILLCELL_X2 FILLER_414_629 ();
 FILLCELL_X32 FILLER_414_632 ();
 FILLCELL_X32 FILLER_414_664 ();
 FILLCELL_X32 FILLER_414_696 ();
 FILLCELL_X32 FILLER_414_728 ();
 FILLCELL_X32 FILLER_414_760 ();
 FILLCELL_X32 FILLER_414_792 ();
 FILLCELL_X32 FILLER_414_824 ();
 FILLCELL_X32 FILLER_414_856 ();
 FILLCELL_X32 FILLER_414_888 ();
 FILLCELL_X32 FILLER_414_920 ();
 FILLCELL_X32 FILLER_414_952 ();
 FILLCELL_X32 FILLER_414_984 ();
 FILLCELL_X32 FILLER_414_1016 ();
 FILLCELL_X32 FILLER_414_1048 ();
 FILLCELL_X32 FILLER_414_1080 ();
 FILLCELL_X32 FILLER_414_1112 ();
 FILLCELL_X32 FILLER_414_1144 ();
 FILLCELL_X32 FILLER_414_1176 ();
 FILLCELL_X32 FILLER_414_1208 ();
 FILLCELL_X32 FILLER_414_1240 ();
 FILLCELL_X32 FILLER_414_1272 ();
 FILLCELL_X32 FILLER_414_1304 ();
 FILLCELL_X32 FILLER_414_1336 ();
 FILLCELL_X32 FILLER_414_1368 ();
 FILLCELL_X32 FILLER_414_1400 ();
 FILLCELL_X32 FILLER_414_1432 ();
 FILLCELL_X32 FILLER_414_1464 ();
 FILLCELL_X32 FILLER_414_1496 ();
 FILLCELL_X32 FILLER_414_1528 ();
 FILLCELL_X32 FILLER_414_1560 ();
 FILLCELL_X32 FILLER_414_1592 ();
 FILLCELL_X32 FILLER_414_1624 ();
 FILLCELL_X32 FILLER_414_1656 ();
 FILLCELL_X32 FILLER_414_1688 ();
 FILLCELL_X32 FILLER_414_1720 ();
 FILLCELL_X32 FILLER_414_1752 ();
 FILLCELL_X32 FILLER_414_1784 ();
 FILLCELL_X32 FILLER_414_1816 ();
 FILLCELL_X32 FILLER_414_1848 ();
 FILLCELL_X8 FILLER_414_1880 ();
 FILLCELL_X4 FILLER_414_1888 ();
 FILLCELL_X2 FILLER_414_1892 ();
 FILLCELL_X32 FILLER_414_1895 ();
 FILLCELL_X32 FILLER_414_1927 ();
 FILLCELL_X32 FILLER_414_1959 ();
 FILLCELL_X32 FILLER_414_1991 ();
 FILLCELL_X32 FILLER_414_2023 ();
 FILLCELL_X32 FILLER_414_2055 ();
 FILLCELL_X32 FILLER_414_2087 ();
 FILLCELL_X32 FILLER_414_2119 ();
 FILLCELL_X32 FILLER_414_2151 ();
 FILLCELL_X32 FILLER_414_2183 ();
 FILLCELL_X32 FILLER_414_2215 ();
 FILLCELL_X32 FILLER_414_2247 ();
 FILLCELL_X32 FILLER_414_2279 ();
 FILLCELL_X32 FILLER_414_2311 ();
 FILLCELL_X32 FILLER_414_2343 ();
 FILLCELL_X32 FILLER_414_2375 ();
 FILLCELL_X32 FILLER_414_2407 ();
 FILLCELL_X32 FILLER_414_2439 ();
 FILLCELL_X32 FILLER_414_2471 ();
 FILLCELL_X32 FILLER_414_2503 ();
 FILLCELL_X32 FILLER_414_2535 ();
 FILLCELL_X32 FILLER_414_2567 ();
 FILLCELL_X32 FILLER_414_2599 ();
 FILLCELL_X32 FILLER_414_2631 ();
 FILLCELL_X32 FILLER_414_2663 ();
 FILLCELL_X32 FILLER_414_2695 ();
 FILLCELL_X32 FILLER_414_2727 ();
 FILLCELL_X32 FILLER_414_2759 ();
 FILLCELL_X32 FILLER_414_2791 ();
 FILLCELL_X32 FILLER_414_2823 ();
 FILLCELL_X32 FILLER_414_2855 ();
 FILLCELL_X32 FILLER_414_2887 ();
 FILLCELL_X32 FILLER_414_2919 ();
 FILLCELL_X32 FILLER_414_2951 ();
 FILLCELL_X32 FILLER_414_2983 ();
 FILLCELL_X32 FILLER_414_3015 ();
 FILLCELL_X32 FILLER_414_3047 ();
 FILLCELL_X32 FILLER_414_3079 ();
 FILLCELL_X32 FILLER_414_3111 ();
 FILLCELL_X8 FILLER_414_3143 ();
 FILLCELL_X4 FILLER_414_3151 ();
 FILLCELL_X2 FILLER_414_3155 ();
 FILLCELL_X32 FILLER_414_3158 ();
 FILLCELL_X32 FILLER_414_3190 ();
 FILLCELL_X32 FILLER_414_3222 ();
 FILLCELL_X32 FILLER_414_3254 ();
 FILLCELL_X32 FILLER_414_3286 ();
 FILLCELL_X32 FILLER_414_3318 ();
 FILLCELL_X32 FILLER_414_3350 ();
 FILLCELL_X32 FILLER_414_3382 ();
 FILLCELL_X32 FILLER_414_3414 ();
 FILLCELL_X32 FILLER_414_3446 ();
 FILLCELL_X32 FILLER_414_3478 ();
 FILLCELL_X32 FILLER_414_3510 ();
 FILLCELL_X32 FILLER_414_3542 ();
 FILLCELL_X32 FILLER_414_3574 ();
 FILLCELL_X32 FILLER_414_3606 ();
 FILLCELL_X32 FILLER_414_3638 ();
 FILLCELL_X32 FILLER_414_3670 ();
 FILLCELL_X32 FILLER_414_3702 ();
 FILLCELL_X4 FILLER_414_3734 ();
 FILLCELL_X32 FILLER_415_1 ();
 FILLCELL_X32 FILLER_415_33 ();
 FILLCELL_X32 FILLER_415_65 ();
 FILLCELL_X32 FILLER_415_97 ();
 FILLCELL_X32 FILLER_415_129 ();
 FILLCELL_X32 FILLER_415_161 ();
 FILLCELL_X32 FILLER_415_193 ();
 FILLCELL_X32 FILLER_415_225 ();
 FILLCELL_X32 FILLER_415_257 ();
 FILLCELL_X32 FILLER_415_289 ();
 FILLCELL_X32 FILLER_415_321 ();
 FILLCELL_X32 FILLER_415_353 ();
 FILLCELL_X32 FILLER_415_385 ();
 FILLCELL_X32 FILLER_415_417 ();
 FILLCELL_X32 FILLER_415_449 ();
 FILLCELL_X32 FILLER_415_481 ();
 FILLCELL_X32 FILLER_415_513 ();
 FILLCELL_X32 FILLER_415_545 ();
 FILLCELL_X32 FILLER_415_577 ();
 FILLCELL_X32 FILLER_415_609 ();
 FILLCELL_X32 FILLER_415_641 ();
 FILLCELL_X32 FILLER_415_673 ();
 FILLCELL_X32 FILLER_415_705 ();
 FILLCELL_X32 FILLER_415_737 ();
 FILLCELL_X32 FILLER_415_769 ();
 FILLCELL_X32 FILLER_415_801 ();
 FILLCELL_X32 FILLER_415_833 ();
 FILLCELL_X32 FILLER_415_865 ();
 FILLCELL_X32 FILLER_415_897 ();
 FILLCELL_X32 FILLER_415_929 ();
 FILLCELL_X32 FILLER_415_961 ();
 FILLCELL_X32 FILLER_415_993 ();
 FILLCELL_X32 FILLER_415_1025 ();
 FILLCELL_X32 FILLER_415_1057 ();
 FILLCELL_X32 FILLER_415_1089 ();
 FILLCELL_X32 FILLER_415_1121 ();
 FILLCELL_X32 FILLER_415_1153 ();
 FILLCELL_X32 FILLER_415_1185 ();
 FILLCELL_X32 FILLER_415_1217 ();
 FILLCELL_X8 FILLER_415_1249 ();
 FILLCELL_X4 FILLER_415_1257 ();
 FILLCELL_X2 FILLER_415_1261 ();
 FILLCELL_X32 FILLER_415_1264 ();
 FILLCELL_X32 FILLER_415_1296 ();
 FILLCELL_X32 FILLER_415_1328 ();
 FILLCELL_X32 FILLER_415_1360 ();
 FILLCELL_X32 FILLER_415_1392 ();
 FILLCELL_X32 FILLER_415_1424 ();
 FILLCELL_X32 FILLER_415_1456 ();
 FILLCELL_X32 FILLER_415_1488 ();
 FILLCELL_X32 FILLER_415_1520 ();
 FILLCELL_X32 FILLER_415_1552 ();
 FILLCELL_X32 FILLER_415_1584 ();
 FILLCELL_X32 FILLER_415_1616 ();
 FILLCELL_X32 FILLER_415_1648 ();
 FILLCELL_X32 FILLER_415_1680 ();
 FILLCELL_X32 FILLER_415_1712 ();
 FILLCELL_X32 FILLER_415_1744 ();
 FILLCELL_X32 FILLER_415_1776 ();
 FILLCELL_X32 FILLER_415_1808 ();
 FILLCELL_X32 FILLER_415_1840 ();
 FILLCELL_X32 FILLER_415_1872 ();
 FILLCELL_X32 FILLER_415_1904 ();
 FILLCELL_X32 FILLER_415_1936 ();
 FILLCELL_X32 FILLER_415_1968 ();
 FILLCELL_X32 FILLER_415_2000 ();
 FILLCELL_X32 FILLER_415_2032 ();
 FILLCELL_X32 FILLER_415_2064 ();
 FILLCELL_X32 FILLER_415_2096 ();
 FILLCELL_X32 FILLER_415_2128 ();
 FILLCELL_X32 FILLER_415_2160 ();
 FILLCELL_X32 FILLER_415_2192 ();
 FILLCELL_X32 FILLER_415_2224 ();
 FILLCELL_X32 FILLER_415_2256 ();
 FILLCELL_X32 FILLER_415_2288 ();
 FILLCELL_X32 FILLER_415_2320 ();
 FILLCELL_X32 FILLER_415_2352 ();
 FILLCELL_X32 FILLER_415_2384 ();
 FILLCELL_X32 FILLER_415_2416 ();
 FILLCELL_X32 FILLER_415_2448 ();
 FILLCELL_X32 FILLER_415_2480 ();
 FILLCELL_X8 FILLER_415_2512 ();
 FILLCELL_X4 FILLER_415_2520 ();
 FILLCELL_X2 FILLER_415_2524 ();
 FILLCELL_X32 FILLER_415_2527 ();
 FILLCELL_X32 FILLER_415_2559 ();
 FILLCELL_X32 FILLER_415_2591 ();
 FILLCELL_X32 FILLER_415_2623 ();
 FILLCELL_X32 FILLER_415_2655 ();
 FILLCELL_X32 FILLER_415_2687 ();
 FILLCELL_X32 FILLER_415_2719 ();
 FILLCELL_X32 FILLER_415_2751 ();
 FILLCELL_X32 FILLER_415_2783 ();
 FILLCELL_X32 FILLER_415_2815 ();
 FILLCELL_X32 FILLER_415_2847 ();
 FILLCELL_X32 FILLER_415_2879 ();
 FILLCELL_X32 FILLER_415_2911 ();
 FILLCELL_X32 FILLER_415_2943 ();
 FILLCELL_X32 FILLER_415_2975 ();
 FILLCELL_X32 FILLER_415_3007 ();
 FILLCELL_X32 FILLER_415_3039 ();
 FILLCELL_X32 FILLER_415_3071 ();
 FILLCELL_X32 FILLER_415_3103 ();
 FILLCELL_X32 FILLER_415_3135 ();
 FILLCELL_X32 FILLER_415_3167 ();
 FILLCELL_X32 FILLER_415_3199 ();
 FILLCELL_X32 FILLER_415_3231 ();
 FILLCELL_X32 FILLER_415_3263 ();
 FILLCELL_X32 FILLER_415_3295 ();
 FILLCELL_X32 FILLER_415_3327 ();
 FILLCELL_X32 FILLER_415_3359 ();
 FILLCELL_X32 FILLER_415_3391 ();
 FILLCELL_X32 FILLER_415_3423 ();
 FILLCELL_X32 FILLER_415_3455 ();
 FILLCELL_X32 FILLER_415_3487 ();
 FILLCELL_X32 FILLER_415_3519 ();
 FILLCELL_X32 FILLER_415_3551 ();
 FILLCELL_X32 FILLER_415_3583 ();
 FILLCELL_X32 FILLER_415_3615 ();
 FILLCELL_X32 FILLER_415_3647 ();
 FILLCELL_X32 FILLER_415_3679 ();
 FILLCELL_X16 FILLER_415_3711 ();
 FILLCELL_X8 FILLER_415_3727 ();
 FILLCELL_X2 FILLER_415_3735 ();
 FILLCELL_X1 FILLER_415_3737 ();
 FILLCELL_X32 FILLER_416_1 ();
 FILLCELL_X32 FILLER_416_33 ();
 FILLCELL_X32 FILLER_416_65 ();
 FILLCELL_X32 FILLER_416_97 ();
 FILLCELL_X32 FILLER_416_129 ();
 FILLCELL_X32 FILLER_416_161 ();
 FILLCELL_X32 FILLER_416_193 ();
 FILLCELL_X32 FILLER_416_225 ();
 FILLCELL_X32 FILLER_416_257 ();
 FILLCELL_X32 FILLER_416_289 ();
 FILLCELL_X32 FILLER_416_321 ();
 FILLCELL_X32 FILLER_416_353 ();
 FILLCELL_X32 FILLER_416_385 ();
 FILLCELL_X32 FILLER_416_417 ();
 FILLCELL_X32 FILLER_416_449 ();
 FILLCELL_X32 FILLER_416_481 ();
 FILLCELL_X32 FILLER_416_513 ();
 FILLCELL_X32 FILLER_416_545 ();
 FILLCELL_X32 FILLER_416_577 ();
 FILLCELL_X16 FILLER_416_609 ();
 FILLCELL_X4 FILLER_416_625 ();
 FILLCELL_X2 FILLER_416_629 ();
 FILLCELL_X32 FILLER_416_632 ();
 FILLCELL_X32 FILLER_416_664 ();
 FILLCELL_X32 FILLER_416_696 ();
 FILLCELL_X32 FILLER_416_728 ();
 FILLCELL_X32 FILLER_416_760 ();
 FILLCELL_X32 FILLER_416_792 ();
 FILLCELL_X32 FILLER_416_824 ();
 FILLCELL_X32 FILLER_416_856 ();
 FILLCELL_X32 FILLER_416_888 ();
 FILLCELL_X32 FILLER_416_920 ();
 FILLCELL_X32 FILLER_416_952 ();
 FILLCELL_X32 FILLER_416_984 ();
 FILLCELL_X32 FILLER_416_1016 ();
 FILLCELL_X32 FILLER_416_1048 ();
 FILLCELL_X32 FILLER_416_1080 ();
 FILLCELL_X32 FILLER_416_1112 ();
 FILLCELL_X32 FILLER_416_1144 ();
 FILLCELL_X32 FILLER_416_1176 ();
 FILLCELL_X32 FILLER_416_1208 ();
 FILLCELL_X32 FILLER_416_1240 ();
 FILLCELL_X32 FILLER_416_1272 ();
 FILLCELL_X32 FILLER_416_1304 ();
 FILLCELL_X32 FILLER_416_1336 ();
 FILLCELL_X32 FILLER_416_1368 ();
 FILLCELL_X32 FILLER_416_1400 ();
 FILLCELL_X32 FILLER_416_1432 ();
 FILLCELL_X32 FILLER_416_1464 ();
 FILLCELL_X32 FILLER_416_1496 ();
 FILLCELL_X32 FILLER_416_1528 ();
 FILLCELL_X32 FILLER_416_1560 ();
 FILLCELL_X32 FILLER_416_1592 ();
 FILLCELL_X32 FILLER_416_1624 ();
 FILLCELL_X32 FILLER_416_1656 ();
 FILLCELL_X32 FILLER_416_1688 ();
 FILLCELL_X32 FILLER_416_1720 ();
 FILLCELL_X32 FILLER_416_1752 ();
 FILLCELL_X32 FILLER_416_1784 ();
 FILLCELL_X32 FILLER_416_1816 ();
 FILLCELL_X32 FILLER_416_1848 ();
 FILLCELL_X8 FILLER_416_1880 ();
 FILLCELL_X4 FILLER_416_1888 ();
 FILLCELL_X2 FILLER_416_1892 ();
 FILLCELL_X32 FILLER_416_1895 ();
 FILLCELL_X32 FILLER_416_1927 ();
 FILLCELL_X32 FILLER_416_1959 ();
 FILLCELL_X32 FILLER_416_1991 ();
 FILLCELL_X32 FILLER_416_2023 ();
 FILLCELL_X32 FILLER_416_2055 ();
 FILLCELL_X32 FILLER_416_2087 ();
 FILLCELL_X32 FILLER_416_2119 ();
 FILLCELL_X32 FILLER_416_2151 ();
 FILLCELL_X32 FILLER_416_2183 ();
 FILLCELL_X32 FILLER_416_2215 ();
 FILLCELL_X32 FILLER_416_2247 ();
 FILLCELL_X32 FILLER_416_2279 ();
 FILLCELL_X32 FILLER_416_2311 ();
 FILLCELL_X32 FILLER_416_2343 ();
 FILLCELL_X32 FILLER_416_2375 ();
 FILLCELL_X32 FILLER_416_2407 ();
 FILLCELL_X32 FILLER_416_2439 ();
 FILLCELL_X32 FILLER_416_2471 ();
 FILLCELL_X32 FILLER_416_2503 ();
 FILLCELL_X32 FILLER_416_2535 ();
 FILLCELL_X32 FILLER_416_2567 ();
 FILLCELL_X32 FILLER_416_2599 ();
 FILLCELL_X32 FILLER_416_2631 ();
 FILLCELL_X32 FILLER_416_2663 ();
 FILLCELL_X32 FILLER_416_2695 ();
 FILLCELL_X32 FILLER_416_2727 ();
 FILLCELL_X32 FILLER_416_2759 ();
 FILLCELL_X32 FILLER_416_2791 ();
 FILLCELL_X32 FILLER_416_2823 ();
 FILLCELL_X32 FILLER_416_2855 ();
 FILLCELL_X32 FILLER_416_2887 ();
 FILLCELL_X32 FILLER_416_2919 ();
 FILLCELL_X32 FILLER_416_2951 ();
 FILLCELL_X32 FILLER_416_2983 ();
 FILLCELL_X32 FILLER_416_3015 ();
 FILLCELL_X32 FILLER_416_3047 ();
 FILLCELL_X32 FILLER_416_3079 ();
 FILLCELL_X32 FILLER_416_3111 ();
 FILLCELL_X8 FILLER_416_3143 ();
 FILLCELL_X4 FILLER_416_3151 ();
 FILLCELL_X2 FILLER_416_3155 ();
 FILLCELL_X32 FILLER_416_3158 ();
 FILLCELL_X32 FILLER_416_3190 ();
 FILLCELL_X32 FILLER_416_3222 ();
 FILLCELL_X32 FILLER_416_3254 ();
 FILLCELL_X32 FILLER_416_3286 ();
 FILLCELL_X32 FILLER_416_3318 ();
 FILLCELL_X32 FILLER_416_3350 ();
 FILLCELL_X32 FILLER_416_3382 ();
 FILLCELL_X32 FILLER_416_3414 ();
 FILLCELL_X32 FILLER_416_3446 ();
 FILLCELL_X32 FILLER_416_3478 ();
 FILLCELL_X32 FILLER_416_3510 ();
 FILLCELL_X32 FILLER_416_3542 ();
 FILLCELL_X32 FILLER_416_3574 ();
 FILLCELL_X32 FILLER_416_3606 ();
 FILLCELL_X32 FILLER_416_3638 ();
 FILLCELL_X32 FILLER_416_3670 ();
 FILLCELL_X32 FILLER_416_3702 ();
 FILLCELL_X4 FILLER_416_3734 ();
 FILLCELL_X32 FILLER_417_1 ();
 FILLCELL_X32 FILLER_417_33 ();
 FILLCELL_X32 FILLER_417_65 ();
 FILLCELL_X32 FILLER_417_97 ();
 FILLCELL_X32 FILLER_417_129 ();
 FILLCELL_X32 FILLER_417_161 ();
 FILLCELL_X32 FILLER_417_193 ();
 FILLCELL_X32 FILLER_417_225 ();
 FILLCELL_X32 FILLER_417_257 ();
 FILLCELL_X32 FILLER_417_289 ();
 FILLCELL_X32 FILLER_417_321 ();
 FILLCELL_X32 FILLER_417_353 ();
 FILLCELL_X32 FILLER_417_385 ();
 FILLCELL_X32 FILLER_417_417 ();
 FILLCELL_X32 FILLER_417_449 ();
 FILLCELL_X32 FILLER_417_481 ();
 FILLCELL_X32 FILLER_417_513 ();
 FILLCELL_X32 FILLER_417_545 ();
 FILLCELL_X32 FILLER_417_577 ();
 FILLCELL_X32 FILLER_417_609 ();
 FILLCELL_X32 FILLER_417_641 ();
 FILLCELL_X32 FILLER_417_673 ();
 FILLCELL_X32 FILLER_417_705 ();
 FILLCELL_X32 FILLER_417_737 ();
 FILLCELL_X32 FILLER_417_769 ();
 FILLCELL_X32 FILLER_417_801 ();
 FILLCELL_X32 FILLER_417_833 ();
 FILLCELL_X32 FILLER_417_865 ();
 FILLCELL_X32 FILLER_417_897 ();
 FILLCELL_X32 FILLER_417_929 ();
 FILLCELL_X32 FILLER_417_961 ();
 FILLCELL_X32 FILLER_417_993 ();
 FILLCELL_X32 FILLER_417_1025 ();
 FILLCELL_X32 FILLER_417_1057 ();
 FILLCELL_X32 FILLER_417_1089 ();
 FILLCELL_X32 FILLER_417_1121 ();
 FILLCELL_X32 FILLER_417_1153 ();
 FILLCELL_X32 FILLER_417_1185 ();
 FILLCELL_X32 FILLER_417_1217 ();
 FILLCELL_X8 FILLER_417_1249 ();
 FILLCELL_X4 FILLER_417_1257 ();
 FILLCELL_X2 FILLER_417_1261 ();
 FILLCELL_X32 FILLER_417_1264 ();
 FILLCELL_X32 FILLER_417_1296 ();
 FILLCELL_X32 FILLER_417_1328 ();
 FILLCELL_X32 FILLER_417_1360 ();
 FILLCELL_X32 FILLER_417_1392 ();
 FILLCELL_X32 FILLER_417_1424 ();
 FILLCELL_X32 FILLER_417_1456 ();
 FILLCELL_X32 FILLER_417_1488 ();
 FILLCELL_X32 FILLER_417_1520 ();
 FILLCELL_X32 FILLER_417_1552 ();
 FILLCELL_X32 FILLER_417_1584 ();
 FILLCELL_X32 FILLER_417_1616 ();
 FILLCELL_X32 FILLER_417_1648 ();
 FILLCELL_X32 FILLER_417_1680 ();
 FILLCELL_X32 FILLER_417_1712 ();
 FILLCELL_X32 FILLER_417_1744 ();
 FILLCELL_X32 FILLER_417_1776 ();
 FILLCELL_X32 FILLER_417_1808 ();
 FILLCELL_X32 FILLER_417_1840 ();
 FILLCELL_X32 FILLER_417_1872 ();
 FILLCELL_X32 FILLER_417_1904 ();
 FILLCELL_X32 FILLER_417_1936 ();
 FILLCELL_X32 FILLER_417_1968 ();
 FILLCELL_X32 FILLER_417_2000 ();
 FILLCELL_X32 FILLER_417_2032 ();
 FILLCELL_X32 FILLER_417_2064 ();
 FILLCELL_X32 FILLER_417_2096 ();
 FILLCELL_X32 FILLER_417_2128 ();
 FILLCELL_X32 FILLER_417_2160 ();
 FILLCELL_X32 FILLER_417_2192 ();
 FILLCELL_X32 FILLER_417_2224 ();
 FILLCELL_X32 FILLER_417_2256 ();
 FILLCELL_X32 FILLER_417_2288 ();
 FILLCELL_X32 FILLER_417_2320 ();
 FILLCELL_X32 FILLER_417_2352 ();
 FILLCELL_X32 FILLER_417_2384 ();
 FILLCELL_X32 FILLER_417_2416 ();
 FILLCELL_X32 FILLER_417_2448 ();
 FILLCELL_X32 FILLER_417_2480 ();
 FILLCELL_X8 FILLER_417_2512 ();
 FILLCELL_X4 FILLER_417_2520 ();
 FILLCELL_X2 FILLER_417_2524 ();
 FILLCELL_X32 FILLER_417_2527 ();
 FILLCELL_X32 FILLER_417_2559 ();
 FILLCELL_X32 FILLER_417_2591 ();
 FILLCELL_X32 FILLER_417_2623 ();
 FILLCELL_X32 FILLER_417_2655 ();
 FILLCELL_X32 FILLER_417_2687 ();
 FILLCELL_X32 FILLER_417_2719 ();
 FILLCELL_X32 FILLER_417_2751 ();
 FILLCELL_X32 FILLER_417_2783 ();
 FILLCELL_X32 FILLER_417_2815 ();
 FILLCELL_X32 FILLER_417_2847 ();
 FILLCELL_X32 FILLER_417_2879 ();
 FILLCELL_X32 FILLER_417_2911 ();
 FILLCELL_X32 FILLER_417_2943 ();
 FILLCELL_X32 FILLER_417_2975 ();
 FILLCELL_X32 FILLER_417_3007 ();
 FILLCELL_X32 FILLER_417_3039 ();
 FILLCELL_X32 FILLER_417_3071 ();
 FILLCELL_X32 FILLER_417_3103 ();
 FILLCELL_X32 FILLER_417_3135 ();
 FILLCELL_X32 FILLER_417_3167 ();
 FILLCELL_X32 FILLER_417_3199 ();
 FILLCELL_X32 FILLER_417_3231 ();
 FILLCELL_X32 FILLER_417_3263 ();
 FILLCELL_X32 FILLER_417_3295 ();
 FILLCELL_X32 FILLER_417_3327 ();
 FILLCELL_X32 FILLER_417_3359 ();
 FILLCELL_X32 FILLER_417_3391 ();
 FILLCELL_X32 FILLER_417_3423 ();
 FILLCELL_X32 FILLER_417_3455 ();
 FILLCELL_X32 FILLER_417_3487 ();
 FILLCELL_X32 FILLER_417_3519 ();
 FILLCELL_X32 FILLER_417_3551 ();
 FILLCELL_X32 FILLER_417_3583 ();
 FILLCELL_X32 FILLER_417_3615 ();
 FILLCELL_X32 FILLER_417_3647 ();
 FILLCELL_X32 FILLER_417_3679 ();
 FILLCELL_X16 FILLER_417_3711 ();
 FILLCELL_X8 FILLER_417_3727 ();
 FILLCELL_X2 FILLER_417_3735 ();
 FILLCELL_X1 FILLER_417_3737 ();
 FILLCELL_X32 FILLER_418_1 ();
 FILLCELL_X32 FILLER_418_33 ();
 FILLCELL_X32 FILLER_418_65 ();
 FILLCELL_X32 FILLER_418_97 ();
 FILLCELL_X32 FILLER_418_129 ();
 FILLCELL_X32 FILLER_418_161 ();
 FILLCELL_X32 FILLER_418_193 ();
 FILLCELL_X32 FILLER_418_225 ();
 FILLCELL_X32 FILLER_418_257 ();
 FILLCELL_X32 FILLER_418_289 ();
 FILLCELL_X32 FILLER_418_321 ();
 FILLCELL_X32 FILLER_418_353 ();
 FILLCELL_X32 FILLER_418_385 ();
 FILLCELL_X32 FILLER_418_417 ();
 FILLCELL_X32 FILLER_418_449 ();
 FILLCELL_X32 FILLER_418_481 ();
 FILLCELL_X32 FILLER_418_513 ();
 FILLCELL_X32 FILLER_418_545 ();
 FILLCELL_X32 FILLER_418_577 ();
 FILLCELL_X16 FILLER_418_609 ();
 FILLCELL_X4 FILLER_418_625 ();
 FILLCELL_X2 FILLER_418_629 ();
 FILLCELL_X32 FILLER_418_632 ();
 FILLCELL_X32 FILLER_418_664 ();
 FILLCELL_X32 FILLER_418_696 ();
 FILLCELL_X32 FILLER_418_728 ();
 FILLCELL_X32 FILLER_418_760 ();
 FILLCELL_X32 FILLER_418_792 ();
 FILLCELL_X32 FILLER_418_824 ();
 FILLCELL_X32 FILLER_418_856 ();
 FILLCELL_X32 FILLER_418_888 ();
 FILLCELL_X32 FILLER_418_920 ();
 FILLCELL_X32 FILLER_418_952 ();
 FILLCELL_X32 FILLER_418_984 ();
 FILLCELL_X32 FILLER_418_1016 ();
 FILLCELL_X32 FILLER_418_1048 ();
 FILLCELL_X32 FILLER_418_1080 ();
 FILLCELL_X32 FILLER_418_1112 ();
 FILLCELL_X32 FILLER_418_1144 ();
 FILLCELL_X32 FILLER_418_1176 ();
 FILLCELL_X32 FILLER_418_1208 ();
 FILLCELL_X32 FILLER_418_1240 ();
 FILLCELL_X32 FILLER_418_1272 ();
 FILLCELL_X32 FILLER_418_1304 ();
 FILLCELL_X32 FILLER_418_1336 ();
 FILLCELL_X32 FILLER_418_1368 ();
 FILLCELL_X32 FILLER_418_1400 ();
 FILLCELL_X32 FILLER_418_1432 ();
 FILLCELL_X32 FILLER_418_1464 ();
 FILLCELL_X32 FILLER_418_1496 ();
 FILLCELL_X32 FILLER_418_1528 ();
 FILLCELL_X32 FILLER_418_1560 ();
 FILLCELL_X32 FILLER_418_1592 ();
 FILLCELL_X32 FILLER_418_1624 ();
 FILLCELL_X32 FILLER_418_1656 ();
 FILLCELL_X32 FILLER_418_1688 ();
 FILLCELL_X32 FILLER_418_1720 ();
 FILLCELL_X32 FILLER_418_1752 ();
 FILLCELL_X32 FILLER_418_1784 ();
 FILLCELL_X32 FILLER_418_1816 ();
 FILLCELL_X32 FILLER_418_1848 ();
 FILLCELL_X8 FILLER_418_1880 ();
 FILLCELL_X4 FILLER_418_1888 ();
 FILLCELL_X2 FILLER_418_1892 ();
 FILLCELL_X32 FILLER_418_1895 ();
 FILLCELL_X32 FILLER_418_1927 ();
 FILLCELL_X32 FILLER_418_1959 ();
 FILLCELL_X32 FILLER_418_1991 ();
 FILLCELL_X32 FILLER_418_2023 ();
 FILLCELL_X32 FILLER_418_2055 ();
 FILLCELL_X32 FILLER_418_2087 ();
 FILLCELL_X32 FILLER_418_2119 ();
 FILLCELL_X32 FILLER_418_2151 ();
 FILLCELL_X32 FILLER_418_2183 ();
 FILLCELL_X32 FILLER_418_2215 ();
 FILLCELL_X32 FILLER_418_2247 ();
 FILLCELL_X32 FILLER_418_2279 ();
 FILLCELL_X32 FILLER_418_2311 ();
 FILLCELL_X32 FILLER_418_2343 ();
 FILLCELL_X32 FILLER_418_2375 ();
 FILLCELL_X32 FILLER_418_2407 ();
 FILLCELL_X32 FILLER_418_2439 ();
 FILLCELL_X32 FILLER_418_2471 ();
 FILLCELL_X32 FILLER_418_2503 ();
 FILLCELL_X32 FILLER_418_2535 ();
 FILLCELL_X32 FILLER_418_2567 ();
 FILLCELL_X32 FILLER_418_2599 ();
 FILLCELL_X32 FILLER_418_2631 ();
 FILLCELL_X32 FILLER_418_2663 ();
 FILLCELL_X32 FILLER_418_2695 ();
 FILLCELL_X32 FILLER_418_2727 ();
 FILLCELL_X32 FILLER_418_2759 ();
 FILLCELL_X32 FILLER_418_2791 ();
 FILLCELL_X32 FILLER_418_2823 ();
 FILLCELL_X32 FILLER_418_2855 ();
 FILLCELL_X32 FILLER_418_2887 ();
 FILLCELL_X32 FILLER_418_2919 ();
 FILLCELL_X32 FILLER_418_2951 ();
 FILLCELL_X32 FILLER_418_2983 ();
 FILLCELL_X32 FILLER_418_3015 ();
 FILLCELL_X32 FILLER_418_3047 ();
 FILLCELL_X32 FILLER_418_3079 ();
 FILLCELL_X32 FILLER_418_3111 ();
 FILLCELL_X8 FILLER_418_3143 ();
 FILLCELL_X4 FILLER_418_3151 ();
 FILLCELL_X2 FILLER_418_3155 ();
 FILLCELL_X32 FILLER_418_3158 ();
 FILLCELL_X32 FILLER_418_3190 ();
 FILLCELL_X32 FILLER_418_3222 ();
 FILLCELL_X32 FILLER_418_3254 ();
 FILLCELL_X32 FILLER_418_3286 ();
 FILLCELL_X32 FILLER_418_3318 ();
 FILLCELL_X32 FILLER_418_3350 ();
 FILLCELL_X32 FILLER_418_3382 ();
 FILLCELL_X32 FILLER_418_3414 ();
 FILLCELL_X32 FILLER_418_3446 ();
 FILLCELL_X32 FILLER_418_3478 ();
 FILLCELL_X32 FILLER_418_3510 ();
 FILLCELL_X32 FILLER_418_3542 ();
 FILLCELL_X32 FILLER_418_3574 ();
 FILLCELL_X32 FILLER_418_3606 ();
 FILLCELL_X32 FILLER_418_3638 ();
 FILLCELL_X32 FILLER_418_3670 ();
 FILLCELL_X32 FILLER_418_3702 ();
 FILLCELL_X4 FILLER_418_3734 ();
 FILLCELL_X32 FILLER_419_1 ();
 FILLCELL_X32 FILLER_419_33 ();
 FILLCELL_X32 FILLER_419_65 ();
 FILLCELL_X32 FILLER_419_97 ();
 FILLCELL_X32 FILLER_419_129 ();
 FILLCELL_X32 FILLER_419_161 ();
 FILLCELL_X32 FILLER_419_193 ();
 FILLCELL_X32 FILLER_419_225 ();
 FILLCELL_X32 FILLER_419_257 ();
 FILLCELL_X32 FILLER_419_289 ();
 FILLCELL_X32 FILLER_419_321 ();
 FILLCELL_X32 FILLER_419_353 ();
 FILLCELL_X32 FILLER_419_385 ();
 FILLCELL_X32 FILLER_419_417 ();
 FILLCELL_X32 FILLER_419_449 ();
 FILLCELL_X32 FILLER_419_481 ();
 FILLCELL_X32 FILLER_419_513 ();
 FILLCELL_X32 FILLER_419_545 ();
 FILLCELL_X32 FILLER_419_577 ();
 FILLCELL_X32 FILLER_419_609 ();
 FILLCELL_X32 FILLER_419_641 ();
 FILLCELL_X32 FILLER_419_673 ();
 FILLCELL_X32 FILLER_419_705 ();
 FILLCELL_X32 FILLER_419_737 ();
 FILLCELL_X32 FILLER_419_769 ();
 FILLCELL_X32 FILLER_419_801 ();
 FILLCELL_X32 FILLER_419_833 ();
 FILLCELL_X32 FILLER_419_865 ();
 FILLCELL_X32 FILLER_419_897 ();
 FILLCELL_X32 FILLER_419_929 ();
 FILLCELL_X32 FILLER_419_961 ();
 FILLCELL_X32 FILLER_419_993 ();
 FILLCELL_X32 FILLER_419_1025 ();
 FILLCELL_X32 FILLER_419_1057 ();
 FILLCELL_X32 FILLER_419_1089 ();
 FILLCELL_X32 FILLER_419_1121 ();
 FILLCELL_X32 FILLER_419_1153 ();
 FILLCELL_X32 FILLER_419_1185 ();
 FILLCELL_X32 FILLER_419_1217 ();
 FILLCELL_X8 FILLER_419_1249 ();
 FILLCELL_X4 FILLER_419_1257 ();
 FILLCELL_X2 FILLER_419_1261 ();
 FILLCELL_X32 FILLER_419_1264 ();
 FILLCELL_X32 FILLER_419_1296 ();
 FILLCELL_X32 FILLER_419_1328 ();
 FILLCELL_X32 FILLER_419_1360 ();
 FILLCELL_X32 FILLER_419_1392 ();
 FILLCELL_X32 FILLER_419_1424 ();
 FILLCELL_X32 FILLER_419_1456 ();
 FILLCELL_X32 FILLER_419_1488 ();
 FILLCELL_X32 FILLER_419_1520 ();
 FILLCELL_X32 FILLER_419_1552 ();
 FILLCELL_X32 FILLER_419_1584 ();
 FILLCELL_X32 FILLER_419_1616 ();
 FILLCELL_X32 FILLER_419_1648 ();
 FILLCELL_X32 FILLER_419_1680 ();
 FILLCELL_X32 FILLER_419_1712 ();
 FILLCELL_X32 FILLER_419_1744 ();
 FILLCELL_X32 FILLER_419_1776 ();
 FILLCELL_X32 FILLER_419_1808 ();
 FILLCELL_X32 FILLER_419_1840 ();
 FILLCELL_X32 FILLER_419_1872 ();
 FILLCELL_X32 FILLER_419_1904 ();
 FILLCELL_X32 FILLER_419_1936 ();
 FILLCELL_X32 FILLER_419_1968 ();
 FILLCELL_X32 FILLER_419_2000 ();
 FILLCELL_X32 FILLER_419_2032 ();
 FILLCELL_X32 FILLER_419_2064 ();
 FILLCELL_X32 FILLER_419_2096 ();
 FILLCELL_X32 FILLER_419_2128 ();
 FILLCELL_X32 FILLER_419_2160 ();
 FILLCELL_X32 FILLER_419_2192 ();
 FILLCELL_X32 FILLER_419_2224 ();
 FILLCELL_X32 FILLER_419_2256 ();
 FILLCELL_X32 FILLER_419_2288 ();
 FILLCELL_X32 FILLER_419_2320 ();
 FILLCELL_X32 FILLER_419_2352 ();
 FILLCELL_X32 FILLER_419_2384 ();
 FILLCELL_X32 FILLER_419_2416 ();
 FILLCELL_X32 FILLER_419_2448 ();
 FILLCELL_X32 FILLER_419_2480 ();
 FILLCELL_X8 FILLER_419_2512 ();
 FILLCELL_X4 FILLER_419_2520 ();
 FILLCELL_X2 FILLER_419_2524 ();
 FILLCELL_X32 FILLER_419_2527 ();
 FILLCELL_X32 FILLER_419_2559 ();
 FILLCELL_X32 FILLER_419_2591 ();
 FILLCELL_X32 FILLER_419_2623 ();
 FILLCELL_X32 FILLER_419_2655 ();
 FILLCELL_X32 FILLER_419_2687 ();
 FILLCELL_X32 FILLER_419_2719 ();
 FILLCELL_X32 FILLER_419_2751 ();
 FILLCELL_X32 FILLER_419_2783 ();
 FILLCELL_X32 FILLER_419_2815 ();
 FILLCELL_X32 FILLER_419_2847 ();
 FILLCELL_X32 FILLER_419_2879 ();
 FILLCELL_X32 FILLER_419_2911 ();
 FILLCELL_X32 FILLER_419_2943 ();
 FILLCELL_X32 FILLER_419_2975 ();
 FILLCELL_X32 FILLER_419_3007 ();
 FILLCELL_X32 FILLER_419_3039 ();
 FILLCELL_X32 FILLER_419_3071 ();
 FILLCELL_X32 FILLER_419_3103 ();
 FILLCELL_X32 FILLER_419_3135 ();
 FILLCELL_X32 FILLER_419_3167 ();
 FILLCELL_X32 FILLER_419_3199 ();
 FILLCELL_X32 FILLER_419_3231 ();
 FILLCELL_X32 FILLER_419_3263 ();
 FILLCELL_X32 FILLER_419_3295 ();
 FILLCELL_X32 FILLER_419_3327 ();
 FILLCELL_X32 FILLER_419_3359 ();
 FILLCELL_X32 FILLER_419_3391 ();
 FILLCELL_X32 FILLER_419_3423 ();
 FILLCELL_X32 FILLER_419_3455 ();
 FILLCELL_X32 FILLER_419_3487 ();
 FILLCELL_X32 FILLER_419_3519 ();
 FILLCELL_X32 FILLER_419_3551 ();
 FILLCELL_X32 FILLER_419_3583 ();
 FILLCELL_X32 FILLER_419_3615 ();
 FILLCELL_X32 FILLER_419_3647 ();
 FILLCELL_X32 FILLER_419_3679 ();
 FILLCELL_X16 FILLER_419_3711 ();
 FILLCELL_X8 FILLER_419_3727 ();
 FILLCELL_X2 FILLER_419_3735 ();
 FILLCELL_X1 FILLER_419_3737 ();
 FILLCELL_X32 FILLER_420_1 ();
 FILLCELL_X32 FILLER_420_33 ();
 FILLCELL_X32 FILLER_420_65 ();
 FILLCELL_X32 FILLER_420_97 ();
 FILLCELL_X32 FILLER_420_129 ();
 FILLCELL_X32 FILLER_420_161 ();
 FILLCELL_X32 FILLER_420_193 ();
 FILLCELL_X32 FILLER_420_225 ();
 FILLCELL_X32 FILLER_420_257 ();
 FILLCELL_X32 FILLER_420_289 ();
 FILLCELL_X32 FILLER_420_321 ();
 FILLCELL_X32 FILLER_420_353 ();
 FILLCELL_X32 FILLER_420_385 ();
 FILLCELL_X32 FILLER_420_417 ();
 FILLCELL_X32 FILLER_420_449 ();
 FILLCELL_X32 FILLER_420_481 ();
 FILLCELL_X32 FILLER_420_513 ();
 FILLCELL_X32 FILLER_420_545 ();
 FILLCELL_X32 FILLER_420_577 ();
 FILLCELL_X16 FILLER_420_609 ();
 FILLCELL_X4 FILLER_420_625 ();
 FILLCELL_X2 FILLER_420_629 ();
 FILLCELL_X32 FILLER_420_632 ();
 FILLCELL_X32 FILLER_420_664 ();
 FILLCELL_X32 FILLER_420_696 ();
 FILLCELL_X32 FILLER_420_728 ();
 FILLCELL_X32 FILLER_420_760 ();
 FILLCELL_X32 FILLER_420_792 ();
 FILLCELL_X32 FILLER_420_824 ();
 FILLCELL_X32 FILLER_420_856 ();
 FILLCELL_X32 FILLER_420_888 ();
 FILLCELL_X32 FILLER_420_920 ();
 FILLCELL_X32 FILLER_420_952 ();
 FILLCELL_X32 FILLER_420_984 ();
 FILLCELL_X32 FILLER_420_1016 ();
 FILLCELL_X32 FILLER_420_1048 ();
 FILLCELL_X32 FILLER_420_1080 ();
 FILLCELL_X32 FILLER_420_1112 ();
 FILLCELL_X32 FILLER_420_1144 ();
 FILLCELL_X32 FILLER_420_1176 ();
 FILLCELL_X32 FILLER_420_1208 ();
 FILLCELL_X32 FILLER_420_1240 ();
 FILLCELL_X32 FILLER_420_1272 ();
 FILLCELL_X32 FILLER_420_1304 ();
 FILLCELL_X32 FILLER_420_1336 ();
 FILLCELL_X32 FILLER_420_1368 ();
 FILLCELL_X32 FILLER_420_1400 ();
 FILLCELL_X32 FILLER_420_1432 ();
 FILLCELL_X32 FILLER_420_1464 ();
 FILLCELL_X32 FILLER_420_1496 ();
 FILLCELL_X32 FILLER_420_1528 ();
 FILLCELL_X32 FILLER_420_1560 ();
 FILLCELL_X32 FILLER_420_1592 ();
 FILLCELL_X32 FILLER_420_1624 ();
 FILLCELL_X32 FILLER_420_1656 ();
 FILLCELL_X32 FILLER_420_1688 ();
 FILLCELL_X32 FILLER_420_1720 ();
 FILLCELL_X32 FILLER_420_1752 ();
 FILLCELL_X32 FILLER_420_1784 ();
 FILLCELL_X32 FILLER_420_1816 ();
 FILLCELL_X32 FILLER_420_1848 ();
 FILLCELL_X8 FILLER_420_1880 ();
 FILLCELL_X4 FILLER_420_1888 ();
 FILLCELL_X2 FILLER_420_1892 ();
 FILLCELL_X32 FILLER_420_1895 ();
 FILLCELL_X32 FILLER_420_1927 ();
 FILLCELL_X32 FILLER_420_1959 ();
 FILLCELL_X32 FILLER_420_1991 ();
 FILLCELL_X32 FILLER_420_2023 ();
 FILLCELL_X32 FILLER_420_2055 ();
 FILLCELL_X32 FILLER_420_2087 ();
 FILLCELL_X32 FILLER_420_2119 ();
 FILLCELL_X32 FILLER_420_2151 ();
 FILLCELL_X32 FILLER_420_2183 ();
 FILLCELL_X32 FILLER_420_2215 ();
 FILLCELL_X32 FILLER_420_2247 ();
 FILLCELL_X32 FILLER_420_2279 ();
 FILLCELL_X32 FILLER_420_2311 ();
 FILLCELL_X32 FILLER_420_2343 ();
 FILLCELL_X32 FILLER_420_2375 ();
 FILLCELL_X32 FILLER_420_2407 ();
 FILLCELL_X32 FILLER_420_2439 ();
 FILLCELL_X32 FILLER_420_2471 ();
 FILLCELL_X32 FILLER_420_2503 ();
 FILLCELL_X32 FILLER_420_2535 ();
 FILLCELL_X32 FILLER_420_2567 ();
 FILLCELL_X32 FILLER_420_2599 ();
 FILLCELL_X32 FILLER_420_2631 ();
 FILLCELL_X32 FILLER_420_2663 ();
 FILLCELL_X32 FILLER_420_2695 ();
 FILLCELL_X32 FILLER_420_2727 ();
 FILLCELL_X32 FILLER_420_2759 ();
 FILLCELL_X32 FILLER_420_2791 ();
 FILLCELL_X32 FILLER_420_2823 ();
 FILLCELL_X32 FILLER_420_2855 ();
 FILLCELL_X32 FILLER_420_2887 ();
 FILLCELL_X32 FILLER_420_2919 ();
 FILLCELL_X32 FILLER_420_2951 ();
 FILLCELL_X32 FILLER_420_2983 ();
 FILLCELL_X32 FILLER_420_3015 ();
 FILLCELL_X32 FILLER_420_3047 ();
 FILLCELL_X32 FILLER_420_3079 ();
 FILLCELL_X32 FILLER_420_3111 ();
 FILLCELL_X8 FILLER_420_3143 ();
 FILLCELL_X4 FILLER_420_3151 ();
 FILLCELL_X2 FILLER_420_3155 ();
 FILLCELL_X32 FILLER_420_3158 ();
 FILLCELL_X32 FILLER_420_3190 ();
 FILLCELL_X32 FILLER_420_3222 ();
 FILLCELL_X32 FILLER_420_3254 ();
 FILLCELL_X32 FILLER_420_3286 ();
 FILLCELL_X32 FILLER_420_3318 ();
 FILLCELL_X32 FILLER_420_3350 ();
 FILLCELL_X32 FILLER_420_3382 ();
 FILLCELL_X32 FILLER_420_3414 ();
 FILLCELL_X32 FILLER_420_3446 ();
 FILLCELL_X32 FILLER_420_3478 ();
 FILLCELL_X32 FILLER_420_3510 ();
 FILLCELL_X32 FILLER_420_3542 ();
 FILLCELL_X32 FILLER_420_3574 ();
 FILLCELL_X32 FILLER_420_3606 ();
 FILLCELL_X32 FILLER_420_3638 ();
 FILLCELL_X32 FILLER_420_3670 ();
 FILLCELL_X32 FILLER_420_3702 ();
 FILLCELL_X4 FILLER_420_3734 ();
 FILLCELL_X32 FILLER_421_1 ();
 FILLCELL_X32 FILLER_421_33 ();
 FILLCELL_X32 FILLER_421_65 ();
 FILLCELL_X32 FILLER_421_97 ();
 FILLCELL_X32 FILLER_421_129 ();
 FILLCELL_X32 FILLER_421_161 ();
 FILLCELL_X32 FILLER_421_193 ();
 FILLCELL_X32 FILLER_421_225 ();
 FILLCELL_X32 FILLER_421_257 ();
 FILLCELL_X32 FILLER_421_289 ();
 FILLCELL_X32 FILLER_421_321 ();
 FILLCELL_X32 FILLER_421_353 ();
 FILLCELL_X32 FILLER_421_385 ();
 FILLCELL_X32 FILLER_421_417 ();
 FILLCELL_X32 FILLER_421_449 ();
 FILLCELL_X32 FILLER_421_481 ();
 FILLCELL_X32 FILLER_421_513 ();
 FILLCELL_X32 FILLER_421_545 ();
 FILLCELL_X32 FILLER_421_577 ();
 FILLCELL_X32 FILLER_421_609 ();
 FILLCELL_X32 FILLER_421_641 ();
 FILLCELL_X32 FILLER_421_673 ();
 FILLCELL_X32 FILLER_421_705 ();
 FILLCELL_X32 FILLER_421_737 ();
 FILLCELL_X32 FILLER_421_769 ();
 FILLCELL_X32 FILLER_421_801 ();
 FILLCELL_X32 FILLER_421_833 ();
 FILLCELL_X32 FILLER_421_865 ();
 FILLCELL_X32 FILLER_421_897 ();
 FILLCELL_X32 FILLER_421_929 ();
 FILLCELL_X32 FILLER_421_961 ();
 FILLCELL_X32 FILLER_421_993 ();
 FILLCELL_X32 FILLER_421_1025 ();
 FILLCELL_X32 FILLER_421_1057 ();
 FILLCELL_X32 FILLER_421_1089 ();
 FILLCELL_X32 FILLER_421_1121 ();
 FILLCELL_X32 FILLER_421_1153 ();
 FILLCELL_X32 FILLER_421_1185 ();
 FILLCELL_X32 FILLER_421_1217 ();
 FILLCELL_X8 FILLER_421_1249 ();
 FILLCELL_X4 FILLER_421_1257 ();
 FILLCELL_X2 FILLER_421_1261 ();
 FILLCELL_X32 FILLER_421_1264 ();
 FILLCELL_X32 FILLER_421_1296 ();
 FILLCELL_X32 FILLER_421_1328 ();
 FILLCELL_X32 FILLER_421_1360 ();
 FILLCELL_X32 FILLER_421_1392 ();
 FILLCELL_X32 FILLER_421_1424 ();
 FILLCELL_X32 FILLER_421_1456 ();
 FILLCELL_X32 FILLER_421_1488 ();
 FILLCELL_X32 FILLER_421_1520 ();
 FILLCELL_X32 FILLER_421_1552 ();
 FILLCELL_X32 FILLER_421_1584 ();
 FILLCELL_X32 FILLER_421_1616 ();
 FILLCELL_X32 FILLER_421_1648 ();
 FILLCELL_X32 FILLER_421_1680 ();
 FILLCELL_X32 FILLER_421_1712 ();
 FILLCELL_X32 FILLER_421_1744 ();
 FILLCELL_X32 FILLER_421_1776 ();
 FILLCELL_X32 FILLER_421_1808 ();
 FILLCELL_X32 FILLER_421_1840 ();
 FILLCELL_X32 FILLER_421_1872 ();
 FILLCELL_X32 FILLER_421_1904 ();
 FILLCELL_X32 FILLER_421_1936 ();
 FILLCELL_X32 FILLER_421_1968 ();
 FILLCELL_X32 FILLER_421_2000 ();
 FILLCELL_X32 FILLER_421_2032 ();
 FILLCELL_X32 FILLER_421_2064 ();
 FILLCELL_X32 FILLER_421_2096 ();
 FILLCELL_X32 FILLER_421_2128 ();
 FILLCELL_X32 FILLER_421_2160 ();
 FILLCELL_X32 FILLER_421_2192 ();
 FILLCELL_X32 FILLER_421_2224 ();
 FILLCELL_X32 FILLER_421_2256 ();
 FILLCELL_X32 FILLER_421_2288 ();
 FILLCELL_X32 FILLER_421_2320 ();
 FILLCELL_X32 FILLER_421_2352 ();
 FILLCELL_X32 FILLER_421_2384 ();
 FILLCELL_X32 FILLER_421_2416 ();
 FILLCELL_X32 FILLER_421_2448 ();
 FILLCELL_X32 FILLER_421_2480 ();
 FILLCELL_X8 FILLER_421_2512 ();
 FILLCELL_X4 FILLER_421_2520 ();
 FILLCELL_X2 FILLER_421_2524 ();
 FILLCELL_X32 FILLER_421_2527 ();
 FILLCELL_X32 FILLER_421_2559 ();
 FILLCELL_X32 FILLER_421_2591 ();
 FILLCELL_X32 FILLER_421_2623 ();
 FILLCELL_X32 FILLER_421_2655 ();
 FILLCELL_X32 FILLER_421_2687 ();
 FILLCELL_X32 FILLER_421_2719 ();
 FILLCELL_X32 FILLER_421_2751 ();
 FILLCELL_X32 FILLER_421_2783 ();
 FILLCELL_X32 FILLER_421_2815 ();
 FILLCELL_X32 FILLER_421_2847 ();
 FILLCELL_X32 FILLER_421_2879 ();
 FILLCELL_X32 FILLER_421_2911 ();
 FILLCELL_X32 FILLER_421_2943 ();
 FILLCELL_X32 FILLER_421_2975 ();
 FILLCELL_X32 FILLER_421_3007 ();
 FILLCELL_X32 FILLER_421_3039 ();
 FILLCELL_X32 FILLER_421_3071 ();
 FILLCELL_X32 FILLER_421_3103 ();
 FILLCELL_X32 FILLER_421_3135 ();
 FILLCELL_X32 FILLER_421_3167 ();
 FILLCELL_X32 FILLER_421_3199 ();
 FILLCELL_X32 FILLER_421_3231 ();
 FILLCELL_X32 FILLER_421_3263 ();
 FILLCELL_X32 FILLER_421_3295 ();
 FILLCELL_X32 FILLER_421_3327 ();
 FILLCELL_X32 FILLER_421_3359 ();
 FILLCELL_X32 FILLER_421_3391 ();
 FILLCELL_X32 FILLER_421_3423 ();
 FILLCELL_X32 FILLER_421_3455 ();
 FILLCELL_X32 FILLER_421_3487 ();
 FILLCELL_X32 FILLER_421_3519 ();
 FILLCELL_X32 FILLER_421_3551 ();
 FILLCELL_X32 FILLER_421_3583 ();
 FILLCELL_X32 FILLER_421_3615 ();
 FILLCELL_X32 FILLER_421_3647 ();
 FILLCELL_X32 FILLER_421_3679 ();
 FILLCELL_X16 FILLER_421_3711 ();
 FILLCELL_X8 FILLER_421_3727 ();
 FILLCELL_X2 FILLER_421_3735 ();
 FILLCELL_X1 FILLER_421_3737 ();
 FILLCELL_X32 FILLER_422_1 ();
 FILLCELL_X32 FILLER_422_33 ();
 FILLCELL_X32 FILLER_422_65 ();
 FILLCELL_X32 FILLER_422_97 ();
 FILLCELL_X32 FILLER_422_129 ();
 FILLCELL_X32 FILLER_422_161 ();
 FILLCELL_X32 FILLER_422_193 ();
 FILLCELL_X32 FILLER_422_225 ();
 FILLCELL_X32 FILLER_422_257 ();
 FILLCELL_X32 FILLER_422_289 ();
 FILLCELL_X32 FILLER_422_321 ();
 FILLCELL_X32 FILLER_422_353 ();
 FILLCELL_X32 FILLER_422_385 ();
 FILLCELL_X32 FILLER_422_417 ();
 FILLCELL_X32 FILLER_422_449 ();
 FILLCELL_X32 FILLER_422_481 ();
 FILLCELL_X32 FILLER_422_513 ();
 FILLCELL_X32 FILLER_422_545 ();
 FILLCELL_X32 FILLER_422_577 ();
 FILLCELL_X16 FILLER_422_609 ();
 FILLCELL_X4 FILLER_422_625 ();
 FILLCELL_X2 FILLER_422_629 ();
 FILLCELL_X32 FILLER_422_632 ();
 FILLCELL_X32 FILLER_422_664 ();
 FILLCELL_X32 FILLER_422_696 ();
 FILLCELL_X32 FILLER_422_728 ();
 FILLCELL_X32 FILLER_422_760 ();
 FILLCELL_X32 FILLER_422_792 ();
 FILLCELL_X32 FILLER_422_824 ();
 FILLCELL_X32 FILLER_422_856 ();
 FILLCELL_X32 FILLER_422_888 ();
 FILLCELL_X32 FILLER_422_920 ();
 FILLCELL_X32 FILLER_422_952 ();
 FILLCELL_X32 FILLER_422_984 ();
 FILLCELL_X32 FILLER_422_1016 ();
 FILLCELL_X32 FILLER_422_1048 ();
 FILLCELL_X32 FILLER_422_1080 ();
 FILLCELL_X32 FILLER_422_1112 ();
 FILLCELL_X32 FILLER_422_1144 ();
 FILLCELL_X32 FILLER_422_1176 ();
 FILLCELL_X32 FILLER_422_1208 ();
 FILLCELL_X32 FILLER_422_1240 ();
 FILLCELL_X32 FILLER_422_1272 ();
 FILLCELL_X32 FILLER_422_1304 ();
 FILLCELL_X32 FILLER_422_1336 ();
 FILLCELL_X32 FILLER_422_1368 ();
 FILLCELL_X32 FILLER_422_1400 ();
 FILLCELL_X32 FILLER_422_1432 ();
 FILLCELL_X32 FILLER_422_1464 ();
 FILLCELL_X32 FILLER_422_1496 ();
 FILLCELL_X32 FILLER_422_1528 ();
 FILLCELL_X32 FILLER_422_1560 ();
 FILLCELL_X32 FILLER_422_1592 ();
 FILLCELL_X32 FILLER_422_1624 ();
 FILLCELL_X32 FILLER_422_1656 ();
 FILLCELL_X32 FILLER_422_1688 ();
 FILLCELL_X32 FILLER_422_1720 ();
 FILLCELL_X32 FILLER_422_1752 ();
 FILLCELL_X32 FILLER_422_1784 ();
 FILLCELL_X32 FILLER_422_1816 ();
 FILLCELL_X32 FILLER_422_1848 ();
 FILLCELL_X8 FILLER_422_1880 ();
 FILLCELL_X4 FILLER_422_1888 ();
 FILLCELL_X2 FILLER_422_1892 ();
 FILLCELL_X32 FILLER_422_1895 ();
 FILLCELL_X32 FILLER_422_1927 ();
 FILLCELL_X32 FILLER_422_1959 ();
 FILLCELL_X32 FILLER_422_1991 ();
 FILLCELL_X32 FILLER_422_2023 ();
 FILLCELL_X32 FILLER_422_2055 ();
 FILLCELL_X32 FILLER_422_2087 ();
 FILLCELL_X32 FILLER_422_2119 ();
 FILLCELL_X32 FILLER_422_2151 ();
 FILLCELL_X32 FILLER_422_2183 ();
 FILLCELL_X32 FILLER_422_2215 ();
 FILLCELL_X32 FILLER_422_2247 ();
 FILLCELL_X32 FILLER_422_2279 ();
 FILLCELL_X32 FILLER_422_2311 ();
 FILLCELL_X32 FILLER_422_2343 ();
 FILLCELL_X32 FILLER_422_2375 ();
 FILLCELL_X32 FILLER_422_2407 ();
 FILLCELL_X32 FILLER_422_2439 ();
 FILLCELL_X32 FILLER_422_2471 ();
 FILLCELL_X32 FILLER_422_2503 ();
 FILLCELL_X32 FILLER_422_2535 ();
 FILLCELL_X32 FILLER_422_2567 ();
 FILLCELL_X32 FILLER_422_2599 ();
 FILLCELL_X32 FILLER_422_2631 ();
 FILLCELL_X32 FILLER_422_2663 ();
 FILLCELL_X32 FILLER_422_2695 ();
 FILLCELL_X32 FILLER_422_2727 ();
 FILLCELL_X32 FILLER_422_2759 ();
 FILLCELL_X32 FILLER_422_2791 ();
 FILLCELL_X32 FILLER_422_2823 ();
 FILLCELL_X32 FILLER_422_2855 ();
 FILLCELL_X32 FILLER_422_2887 ();
 FILLCELL_X32 FILLER_422_2919 ();
 FILLCELL_X32 FILLER_422_2951 ();
 FILLCELL_X32 FILLER_422_2983 ();
 FILLCELL_X32 FILLER_422_3015 ();
 FILLCELL_X32 FILLER_422_3047 ();
 FILLCELL_X32 FILLER_422_3079 ();
 FILLCELL_X32 FILLER_422_3111 ();
 FILLCELL_X8 FILLER_422_3143 ();
 FILLCELL_X4 FILLER_422_3151 ();
 FILLCELL_X2 FILLER_422_3155 ();
 FILLCELL_X32 FILLER_422_3158 ();
 FILLCELL_X32 FILLER_422_3190 ();
 FILLCELL_X32 FILLER_422_3222 ();
 FILLCELL_X32 FILLER_422_3254 ();
 FILLCELL_X32 FILLER_422_3286 ();
 FILLCELL_X32 FILLER_422_3318 ();
 FILLCELL_X32 FILLER_422_3350 ();
 FILLCELL_X32 FILLER_422_3382 ();
 FILLCELL_X32 FILLER_422_3414 ();
 FILLCELL_X32 FILLER_422_3446 ();
 FILLCELL_X32 FILLER_422_3478 ();
 FILLCELL_X32 FILLER_422_3510 ();
 FILLCELL_X32 FILLER_422_3542 ();
 FILLCELL_X32 FILLER_422_3574 ();
 FILLCELL_X32 FILLER_422_3606 ();
 FILLCELL_X32 FILLER_422_3638 ();
 FILLCELL_X32 FILLER_422_3670 ();
 FILLCELL_X32 FILLER_422_3702 ();
 FILLCELL_X4 FILLER_422_3734 ();
 FILLCELL_X32 FILLER_423_1 ();
 FILLCELL_X32 FILLER_423_33 ();
 FILLCELL_X32 FILLER_423_65 ();
 FILLCELL_X32 FILLER_423_97 ();
 FILLCELL_X32 FILLER_423_129 ();
 FILLCELL_X32 FILLER_423_161 ();
 FILLCELL_X32 FILLER_423_193 ();
 FILLCELL_X32 FILLER_423_225 ();
 FILLCELL_X32 FILLER_423_257 ();
 FILLCELL_X32 FILLER_423_289 ();
 FILLCELL_X32 FILLER_423_321 ();
 FILLCELL_X32 FILLER_423_353 ();
 FILLCELL_X32 FILLER_423_385 ();
 FILLCELL_X32 FILLER_423_417 ();
 FILLCELL_X32 FILLER_423_449 ();
 FILLCELL_X32 FILLER_423_481 ();
 FILLCELL_X32 FILLER_423_513 ();
 FILLCELL_X32 FILLER_423_545 ();
 FILLCELL_X32 FILLER_423_577 ();
 FILLCELL_X32 FILLER_423_609 ();
 FILLCELL_X32 FILLER_423_641 ();
 FILLCELL_X32 FILLER_423_673 ();
 FILLCELL_X32 FILLER_423_705 ();
 FILLCELL_X32 FILLER_423_737 ();
 FILLCELL_X32 FILLER_423_769 ();
 FILLCELL_X32 FILLER_423_801 ();
 FILLCELL_X32 FILLER_423_833 ();
 FILLCELL_X32 FILLER_423_865 ();
 FILLCELL_X32 FILLER_423_897 ();
 FILLCELL_X32 FILLER_423_929 ();
 FILLCELL_X32 FILLER_423_961 ();
 FILLCELL_X32 FILLER_423_993 ();
 FILLCELL_X32 FILLER_423_1025 ();
 FILLCELL_X32 FILLER_423_1057 ();
 FILLCELL_X32 FILLER_423_1089 ();
 FILLCELL_X32 FILLER_423_1121 ();
 FILLCELL_X32 FILLER_423_1153 ();
 FILLCELL_X32 FILLER_423_1185 ();
 FILLCELL_X32 FILLER_423_1217 ();
 FILLCELL_X8 FILLER_423_1249 ();
 FILLCELL_X4 FILLER_423_1257 ();
 FILLCELL_X2 FILLER_423_1261 ();
 FILLCELL_X32 FILLER_423_1264 ();
 FILLCELL_X32 FILLER_423_1296 ();
 FILLCELL_X32 FILLER_423_1328 ();
 FILLCELL_X32 FILLER_423_1360 ();
 FILLCELL_X32 FILLER_423_1392 ();
 FILLCELL_X32 FILLER_423_1424 ();
 FILLCELL_X32 FILLER_423_1456 ();
 FILLCELL_X32 FILLER_423_1488 ();
 FILLCELL_X32 FILLER_423_1520 ();
 FILLCELL_X32 FILLER_423_1552 ();
 FILLCELL_X32 FILLER_423_1584 ();
 FILLCELL_X32 FILLER_423_1616 ();
 FILLCELL_X32 FILLER_423_1648 ();
 FILLCELL_X32 FILLER_423_1680 ();
 FILLCELL_X32 FILLER_423_1712 ();
 FILLCELL_X32 FILLER_423_1744 ();
 FILLCELL_X32 FILLER_423_1776 ();
 FILLCELL_X32 FILLER_423_1808 ();
 FILLCELL_X32 FILLER_423_1840 ();
 FILLCELL_X32 FILLER_423_1872 ();
 FILLCELL_X32 FILLER_423_1904 ();
 FILLCELL_X32 FILLER_423_1936 ();
 FILLCELL_X32 FILLER_423_1968 ();
 FILLCELL_X32 FILLER_423_2000 ();
 FILLCELL_X32 FILLER_423_2032 ();
 FILLCELL_X32 FILLER_423_2064 ();
 FILLCELL_X32 FILLER_423_2096 ();
 FILLCELL_X32 FILLER_423_2128 ();
 FILLCELL_X32 FILLER_423_2160 ();
 FILLCELL_X32 FILLER_423_2192 ();
 FILLCELL_X32 FILLER_423_2224 ();
 FILLCELL_X32 FILLER_423_2256 ();
 FILLCELL_X32 FILLER_423_2288 ();
 FILLCELL_X32 FILLER_423_2320 ();
 FILLCELL_X32 FILLER_423_2352 ();
 FILLCELL_X32 FILLER_423_2384 ();
 FILLCELL_X32 FILLER_423_2416 ();
 FILLCELL_X32 FILLER_423_2448 ();
 FILLCELL_X32 FILLER_423_2480 ();
 FILLCELL_X8 FILLER_423_2512 ();
 FILLCELL_X4 FILLER_423_2520 ();
 FILLCELL_X2 FILLER_423_2524 ();
 FILLCELL_X32 FILLER_423_2527 ();
 FILLCELL_X32 FILLER_423_2559 ();
 FILLCELL_X32 FILLER_423_2591 ();
 FILLCELL_X32 FILLER_423_2623 ();
 FILLCELL_X32 FILLER_423_2655 ();
 FILLCELL_X32 FILLER_423_2687 ();
 FILLCELL_X32 FILLER_423_2719 ();
 FILLCELL_X32 FILLER_423_2751 ();
 FILLCELL_X32 FILLER_423_2783 ();
 FILLCELL_X32 FILLER_423_2815 ();
 FILLCELL_X32 FILLER_423_2847 ();
 FILLCELL_X32 FILLER_423_2879 ();
 FILLCELL_X32 FILLER_423_2911 ();
 FILLCELL_X32 FILLER_423_2943 ();
 FILLCELL_X32 FILLER_423_2975 ();
 FILLCELL_X32 FILLER_423_3007 ();
 FILLCELL_X32 FILLER_423_3039 ();
 FILLCELL_X32 FILLER_423_3071 ();
 FILLCELL_X32 FILLER_423_3103 ();
 FILLCELL_X32 FILLER_423_3135 ();
 FILLCELL_X32 FILLER_423_3167 ();
 FILLCELL_X32 FILLER_423_3199 ();
 FILLCELL_X32 FILLER_423_3231 ();
 FILLCELL_X32 FILLER_423_3263 ();
 FILLCELL_X32 FILLER_423_3295 ();
 FILLCELL_X32 FILLER_423_3327 ();
 FILLCELL_X32 FILLER_423_3359 ();
 FILLCELL_X32 FILLER_423_3391 ();
 FILLCELL_X32 FILLER_423_3423 ();
 FILLCELL_X32 FILLER_423_3455 ();
 FILLCELL_X32 FILLER_423_3487 ();
 FILLCELL_X32 FILLER_423_3519 ();
 FILLCELL_X32 FILLER_423_3551 ();
 FILLCELL_X32 FILLER_423_3583 ();
 FILLCELL_X32 FILLER_423_3615 ();
 FILLCELL_X32 FILLER_423_3647 ();
 FILLCELL_X32 FILLER_423_3679 ();
 FILLCELL_X16 FILLER_423_3711 ();
 FILLCELL_X8 FILLER_423_3727 ();
 FILLCELL_X2 FILLER_423_3735 ();
 FILLCELL_X1 FILLER_423_3737 ();
 FILLCELL_X32 FILLER_424_1 ();
 FILLCELL_X32 FILLER_424_33 ();
 FILLCELL_X32 FILLER_424_65 ();
 FILLCELL_X32 FILLER_424_97 ();
 FILLCELL_X32 FILLER_424_129 ();
 FILLCELL_X32 FILLER_424_161 ();
 FILLCELL_X32 FILLER_424_193 ();
 FILLCELL_X32 FILLER_424_225 ();
 FILLCELL_X32 FILLER_424_257 ();
 FILLCELL_X32 FILLER_424_289 ();
 FILLCELL_X32 FILLER_424_321 ();
 FILLCELL_X32 FILLER_424_353 ();
 FILLCELL_X32 FILLER_424_385 ();
 FILLCELL_X32 FILLER_424_417 ();
 FILLCELL_X32 FILLER_424_449 ();
 FILLCELL_X32 FILLER_424_481 ();
 FILLCELL_X32 FILLER_424_513 ();
 FILLCELL_X32 FILLER_424_545 ();
 FILLCELL_X32 FILLER_424_577 ();
 FILLCELL_X16 FILLER_424_609 ();
 FILLCELL_X4 FILLER_424_625 ();
 FILLCELL_X2 FILLER_424_629 ();
 FILLCELL_X32 FILLER_424_632 ();
 FILLCELL_X32 FILLER_424_664 ();
 FILLCELL_X32 FILLER_424_696 ();
 FILLCELL_X32 FILLER_424_728 ();
 FILLCELL_X32 FILLER_424_760 ();
 FILLCELL_X32 FILLER_424_792 ();
 FILLCELL_X32 FILLER_424_824 ();
 FILLCELL_X32 FILLER_424_856 ();
 FILLCELL_X32 FILLER_424_888 ();
 FILLCELL_X32 FILLER_424_920 ();
 FILLCELL_X32 FILLER_424_952 ();
 FILLCELL_X32 FILLER_424_984 ();
 FILLCELL_X32 FILLER_424_1016 ();
 FILLCELL_X32 FILLER_424_1048 ();
 FILLCELL_X32 FILLER_424_1080 ();
 FILLCELL_X32 FILLER_424_1112 ();
 FILLCELL_X32 FILLER_424_1144 ();
 FILLCELL_X32 FILLER_424_1176 ();
 FILLCELL_X32 FILLER_424_1208 ();
 FILLCELL_X32 FILLER_424_1240 ();
 FILLCELL_X32 FILLER_424_1272 ();
 FILLCELL_X32 FILLER_424_1304 ();
 FILLCELL_X32 FILLER_424_1336 ();
 FILLCELL_X32 FILLER_424_1368 ();
 FILLCELL_X32 FILLER_424_1400 ();
 FILLCELL_X32 FILLER_424_1432 ();
 FILLCELL_X32 FILLER_424_1464 ();
 FILLCELL_X32 FILLER_424_1496 ();
 FILLCELL_X32 FILLER_424_1528 ();
 FILLCELL_X32 FILLER_424_1560 ();
 FILLCELL_X32 FILLER_424_1592 ();
 FILLCELL_X32 FILLER_424_1624 ();
 FILLCELL_X32 FILLER_424_1656 ();
 FILLCELL_X32 FILLER_424_1688 ();
 FILLCELL_X32 FILLER_424_1720 ();
 FILLCELL_X32 FILLER_424_1752 ();
 FILLCELL_X32 FILLER_424_1784 ();
 FILLCELL_X32 FILLER_424_1816 ();
 FILLCELL_X32 FILLER_424_1848 ();
 FILLCELL_X8 FILLER_424_1880 ();
 FILLCELL_X4 FILLER_424_1888 ();
 FILLCELL_X2 FILLER_424_1892 ();
 FILLCELL_X32 FILLER_424_1895 ();
 FILLCELL_X32 FILLER_424_1927 ();
 FILLCELL_X32 FILLER_424_1959 ();
 FILLCELL_X32 FILLER_424_1991 ();
 FILLCELL_X32 FILLER_424_2023 ();
 FILLCELL_X32 FILLER_424_2055 ();
 FILLCELL_X32 FILLER_424_2087 ();
 FILLCELL_X32 FILLER_424_2119 ();
 FILLCELL_X32 FILLER_424_2151 ();
 FILLCELL_X32 FILLER_424_2183 ();
 FILLCELL_X32 FILLER_424_2215 ();
 FILLCELL_X32 FILLER_424_2247 ();
 FILLCELL_X32 FILLER_424_2279 ();
 FILLCELL_X32 FILLER_424_2311 ();
 FILLCELL_X32 FILLER_424_2343 ();
 FILLCELL_X32 FILLER_424_2375 ();
 FILLCELL_X32 FILLER_424_2407 ();
 FILLCELL_X32 FILLER_424_2439 ();
 FILLCELL_X32 FILLER_424_2471 ();
 FILLCELL_X32 FILLER_424_2503 ();
 FILLCELL_X32 FILLER_424_2535 ();
 FILLCELL_X32 FILLER_424_2567 ();
 FILLCELL_X32 FILLER_424_2599 ();
 FILLCELL_X32 FILLER_424_2631 ();
 FILLCELL_X32 FILLER_424_2663 ();
 FILLCELL_X32 FILLER_424_2695 ();
 FILLCELL_X32 FILLER_424_2727 ();
 FILLCELL_X32 FILLER_424_2759 ();
 FILLCELL_X32 FILLER_424_2791 ();
 FILLCELL_X32 FILLER_424_2823 ();
 FILLCELL_X32 FILLER_424_2855 ();
 FILLCELL_X32 FILLER_424_2887 ();
 FILLCELL_X32 FILLER_424_2919 ();
 FILLCELL_X32 FILLER_424_2951 ();
 FILLCELL_X32 FILLER_424_2983 ();
 FILLCELL_X32 FILLER_424_3015 ();
 FILLCELL_X32 FILLER_424_3047 ();
 FILLCELL_X32 FILLER_424_3079 ();
 FILLCELL_X32 FILLER_424_3111 ();
 FILLCELL_X8 FILLER_424_3143 ();
 FILLCELL_X4 FILLER_424_3151 ();
 FILLCELL_X2 FILLER_424_3155 ();
 FILLCELL_X32 FILLER_424_3158 ();
 FILLCELL_X32 FILLER_424_3190 ();
 FILLCELL_X32 FILLER_424_3222 ();
 FILLCELL_X32 FILLER_424_3254 ();
 FILLCELL_X32 FILLER_424_3286 ();
 FILLCELL_X32 FILLER_424_3318 ();
 FILLCELL_X32 FILLER_424_3350 ();
 FILLCELL_X32 FILLER_424_3382 ();
 FILLCELL_X32 FILLER_424_3414 ();
 FILLCELL_X32 FILLER_424_3446 ();
 FILLCELL_X32 FILLER_424_3478 ();
 FILLCELL_X32 FILLER_424_3510 ();
 FILLCELL_X32 FILLER_424_3542 ();
 FILLCELL_X32 FILLER_424_3574 ();
 FILLCELL_X32 FILLER_424_3606 ();
 FILLCELL_X32 FILLER_424_3638 ();
 FILLCELL_X32 FILLER_424_3670 ();
 FILLCELL_X32 FILLER_424_3702 ();
 FILLCELL_X4 FILLER_424_3734 ();
 FILLCELL_X32 FILLER_425_1 ();
 FILLCELL_X32 FILLER_425_33 ();
 FILLCELL_X32 FILLER_425_65 ();
 FILLCELL_X32 FILLER_425_97 ();
 FILLCELL_X32 FILLER_425_129 ();
 FILLCELL_X32 FILLER_425_161 ();
 FILLCELL_X32 FILLER_425_193 ();
 FILLCELL_X32 FILLER_425_225 ();
 FILLCELL_X32 FILLER_425_257 ();
 FILLCELL_X32 FILLER_425_289 ();
 FILLCELL_X32 FILLER_425_321 ();
 FILLCELL_X32 FILLER_425_353 ();
 FILLCELL_X32 FILLER_425_385 ();
 FILLCELL_X32 FILLER_425_417 ();
 FILLCELL_X32 FILLER_425_449 ();
 FILLCELL_X32 FILLER_425_481 ();
 FILLCELL_X32 FILLER_425_513 ();
 FILLCELL_X32 FILLER_425_545 ();
 FILLCELL_X32 FILLER_425_577 ();
 FILLCELL_X32 FILLER_425_609 ();
 FILLCELL_X32 FILLER_425_641 ();
 FILLCELL_X32 FILLER_425_673 ();
 FILLCELL_X32 FILLER_425_705 ();
 FILLCELL_X32 FILLER_425_737 ();
 FILLCELL_X32 FILLER_425_769 ();
 FILLCELL_X32 FILLER_425_801 ();
 FILLCELL_X32 FILLER_425_833 ();
 FILLCELL_X32 FILLER_425_865 ();
 FILLCELL_X32 FILLER_425_897 ();
 FILLCELL_X32 FILLER_425_929 ();
 FILLCELL_X32 FILLER_425_961 ();
 FILLCELL_X32 FILLER_425_993 ();
 FILLCELL_X32 FILLER_425_1025 ();
 FILLCELL_X32 FILLER_425_1057 ();
 FILLCELL_X32 FILLER_425_1089 ();
 FILLCELL_X32 FILLER_425_1121 ();
 FILLCELL_X32 FILLER_425_1153 ();
 FILLCELL_X32 FILLER_425_1185 ();
 FILLCELL_X32 FILLER_425_1217 ();
 FILLCELL_X8 FILLER_425_1249 ();
 FILLCELL_X4 FILLER_425_1257 ();
 FILLCELL_X2 FILLER_425_1261 ();
 FILLCELL_X32 FILLER_425_1264 ();
 FILLCELL_X32 FILLER_425_1296 ();
 FILLCELL_X32 FILLER_425_1328 ();
 FILLCELL_X32 FILLER_425_1360 ();
 FILLCELL_X32 FILLER_425_1392 ();
 FILLCELL_X32 FILLER_425_1424 ();
 FILLCELL_X32 FILLER_425_1456 ();
 FILLCELL_X32 FILLER_425_1488 ();
 FILLCELL_X32 FILLER_425_1520 ();
 FILLCELL_X32 FILLER_425_1552 ();
 FILLCELL_X32 FILLER_425_1584 ();
 FILLCELL_X32 FILLER_425_1616 ();
 FILLCELL_X32 FILLER_425_1648 ();
 FILLCELL_X32 FILLER_425_1680 ();
 FILLCELL_X32 FILLER_425_1712 ();
 FILLCELL_X32 FILLER_425_1744 ();
 FILLCELL_X32 FILLER_425_1776 ();
 FILLCELL_X32 FILLER_425_1808 ();
 FILLCELL_X32 FILLER_425_1840 ();
 FILLCELL_X32 FILLER_425_1872 ();
 FILLCELL_X32 FILLER_425_1904 ();
 FILLCELL_X32 FILLER_425_1936 ();
 FILLCELL_X32 FILLER_425_1968 ();
 FILLCELL_X32 FILLER_425_2000 ();
 FILLCELL_X32 FILLER_425_2032 ();
 FILLCELL_X32 FILLER_425_2064 ();
 FILLCELL_X32 FILLER_425_2096 ();
 FILLCELL_X32 FILLER_425_2128 ();
 FILLCELL_X32 FILLER_425_2160 ();
 FILLCELL_X32 FILLER_425_2192 ();
 FILLCELL_X32 FILLER_425_2224 ();
 FILLCELL_X32 FILLER_425_2256 ();
 FILLCELL_X32 FILLER_425_2288 ();
 FILLCELL_X32 FILLER_425_2320 ();
 FILLCELL_X32 FILLER_425_2352 ();
 FILLCELL_X32 FILLER_425_2384 ();
 FILLCELL_X32 FILLER_425_2416 ();
 FILLCELL_X32 FILLER_425_2448 ();
 FILLCELL_X32 FILLER_425_2480 ();
 FILLCELL_X8 FILLER_425_2512 ();
 FILLCELL_X4 FILLER_425_2520 ();
 FILLCELL_X2 FILLER_425_2524 ();
 FILLCELL_X32 FILLER_425_2527 ();
 FILLCELL_X32 FILLER_425_2559 ();
 FILLCELL_X32 FILLER_425_2591 ();
 FILLCELL_X32 FILLER_425_2623 ();
 FILLCELL_X32 FILLER_425_2655 ();
 FILLCELL_X32 FILLER_425_2687 ();
 FILLCELL_X32 FILLER_425_2719 ();
 FILLCELL_X32 FILLER_425_2751 ();
 FILLCELL_X32 FILLER_425_2783 ();
 FILLCELL_X32 FILLER_425_2815 ();
 FILLCELL_X32 FILLER_425_2847 ();
 FILLCELL_X32 FILLER_425_2879 ();
 FILLCELL_X32 FILLER_425_2911 ();
 FILLCELL_X32 FILLER_425_2943 ();
 FILLCELL_X32 FILLER_425_2975 ();
 FILLCELL_X32 FILLER_425_3007 ();
 FILLCELL_X32 FILLER_425_3039 ();
 FILLCELL_X32 FILLER_425_3071 ();
 FILLCELL_X32 FILLER_425_3103 ();
 FILLCELL_X32 FILLER_425_3135 ();
 FILLCELL_X32 FILLER_425_3167 ();
 FILLCELL_X32 FILLER_425_3199 ();
 FILLCELL_X32 FILLER_425_3231 ();
 FILLCELL_X32 FILLER_425_3263 ();
 FILLCELL_X32 FILLER_425_3295 ();
 FILLCELL_X32 FILLER_425_3327 ();
 FILLCELL_X32 FILLER_425_3359 ();
 FILLCELL_X32 FILLER_425_3391 ();
 FILLCELL_X32 FILLER_425_3423 ();
 FILLCELL_X32 FILLER_425_3455 ();
 FILLCELL_X32 FILLER_425_3487 ();
 FILLCELL_X32 FILLER_425_3519 ();
 FILLCELL_X32 FILLER_425_3551 ();
 FILLCELL_X32 FILLER_425_3583 ();
 FILLCELL_X32 FILLER_425_3615 ();
 FILLCELL_X32 FILLER_425_3647 ();
 FILLCELL_X32 FILLER_425_3679 ();
 FILLCELL_X16 FILLER_425_3711 ();
 FILLCELL_X8 FILLER_425_3727 ();
 FILLCELL_X2 FILLER_425_3735 ();
 FILLCELL_X1 FILLER_425_3737 ();
 FILLCELL_X32 FILLER_426_1 ();
 FILLCELL_X32 FILLER_426_33 ();
 FILLCELL_X32 FILLER_426_65 ();
 FILLCELL_X32 FILLER_426_97 ();
 FILLCELL_X32 FILLER_426_129 ();
 FILLCELL_X32 FILLER_426_161 ();
 FILLCELL_X32 FILLER_426_193 ();
 FILLCELL_X32 FILLER_426_225 ();
 FILLCELL_X32 FILLER_426_257 ();
 FILLCELL_X32 FILLER_426_289 ();
 FILLCELL_X32 FILLER_426_321 ();
 FILLCELL_X32 FILLER_426_353 ();
 FILLCELL_X32 FILLER_426_385 ();
 FILLCELL_X32 FILLER_426_417 ();
 FILLCELL_X32 FILLER_426_449 ();
 FILLCELL_X32 FILLER_426_481 ();
 FILLCELL_X32 FILLER_426_513 ();
 FILLCELL_X32 FILLER_426_545 ();
 FILLCELL_X32 FILLER_426_577 ();
 FILLCELL_X16 FILLER_426_609 ();
 FILLCELL_X4 FILLER_426_625 ();
 FILLCELL_X2 FILLER_426_629 ();
 FILLCELL_X32 FILLER_426_632 ();
 FILLCELL_X32 FILLER_426_664 ();
 FILLCELL_X32 FILLER_426_696 ();
 FILLCELL_X32 FILLER_426_728 ();
 FILLCELL_X32 FILLER_426_760 ();
 FILLCELL_X32 FILLER_426_792 ();
 FILLCELL_X32 FILLER_426_824 ();
 FILLCELL_X32 FILLER_426_856 ();
 FILLCELL_X32 FILLER_426_888 ();
 FILLCELL_X32 FILLER_426_920 ();
 FILLCELL_X32 FILLER_426_952 ();
 FILLCELL_X32 FILLER_426_984 ();
 FILLCELL_X32 FILLER_426_1016 ();
 FILLCELL_X32 FILLER_426_1048 ();
 FILLCELL_X32 FILLER_426_1080 ();
 FILLCELL_X32 FILLER_426_1112 ();
 FILLCELL_X32 FILLER_426_1144 ();
 FILLCELL_X32 FILLER_426_1176 ();
 FILLCELL_X32 FILLER_426_1208 ();
 FILLCELL_X32 FILLER_426_1240 ();
 FILLCELL_X32 FILLER_426_1272 ();
 FILLCELL_X32 FILLER_426_1304 ();
 FILLCELL_X32 FILLER_426_1336 ();
 FILLCELL_X32 FILLER_426_1368 ();
 FILLCELL_X32 FILLER_426_1400 ();
 FILLCELL_X32 FILLER_426_1432 ();
 FILLCELL_X32 FILLER_426_1464 ();
 FILLCELL_X32 FILLER_426_1496 ();
 FILLCELL_X32 FILLER_426_1528 ();
 FILLCELL_X32 FILLER_426_1560 ();
 FILLCELL_X32 FILLER_426_1592 ();
 FILLCELL_X32 FILLER_426_1624 ();
 FILLCELL_X32 FILLER_426_1656 ();
 FILLCELL_X32 FILLER_426_1688 ();
 FILLCELL_X32 FILLER_426_1720 ();
 FILLCELL_X32 FILLER_426_1752 ();
 FILLCELL_X32 FILLER_426_1784 ();
 FILLCELL_X32 FILLER_426_1816 ();
 FILLCELL_X32 FILLER_426_1848 ();
 FILLCELL_X8 FILLER_426_1880 ();
 FILLCELL_X4 FILLER_426_1888 ();
 FILLCELL_X2 FILLER_426_1892 ();
 FILLCELL_X32 FILLER_426_1895 ();
 FILLCELL_X32 FILLER_426_1927 ();
 FILLCELL_X32 FILLER_426_1959 ();
 FILLCELL_X32 FILLER_426_1991 ();
 FILLCELL_X32 FILLER_426_2023 ();
 FILLCELL_X32 FILLER_426_2055 ();
 FILLCELL_X32 FILLER_426_2087 ();
 FILLCELL_X32 FILLER_426_2119 ();
 FILLCELL_X32 FILLER_426_2151 ();
 FILLCELL_X32 FILLER_426_2183 ();
 FILLCELL_X32 FILLER_426_2215 ();
 FILLCELL_X32 FILLER_426_2247 ();
 FILLCELL_X32 FILLER_426_2279 ();
 FILLCELL_X32 FILLER_426_2311 ();
 FILLCELL_X32 FILLER_426_2343 ();
 FILLCELL_X32 FILLER_426_2375 ();
 FILLCELL_X32 FILLER_426_2407 ();
 FILLCELL_X32 FILLER_426_2439 ();
 FILLCELL_X32 FILLER_426_2471 ();
 FILLCELL_X32 FILLER_426_2503 ();
 FILLCELL_X32 FILLER_426_2535 ();
 FILLCELL_X32 FILLER_426_2567 ();
 FILLCELL_X32 FILLER_426_2599 ();
 FILLCELL_X32 FILLER_426_2631 ();
 FILLCELL_X32 FILLER_426_2663 ();
 FILLCELL_X32 FILLER_426_2695 ();
 FILLCELL_X32 FILLER_426_2727 ();
 FILLCELL_X32 FILLER_426_2759 ();
 FILLCELL_X32 FILLER_426_2791 ();
 FILLCELL_X32 FILLER_426_2823 ();
 FILLCELL_X32 FILLER_426_2855 ();
 FILLCELL_X32 FILLER_426_2887 ();
 FILLCELL_X32 FILLER_426_2919 ();
 FILLCELL_X32 FILLER_426_2951 ();
 FILLCELL_X32 FILLER_426_2983 ();
 FILLCELL_X32 FILLER_426_3015 ();
 FILLCELL_X32 FILLER_426_3047 ();
 FILLCELL_X32 FILLER_426_3079 ();
 FILLCELL_X32 FILLER_426_3111 ();
 FILLCELL_X8 FILLER_426_3143 ();
 FILLCELL_X4 FILLER_426_3151 ();
 FILLCELL_X2 FILLER_426_3155 ();
 FILLCELL_X32 FILLER_426_3158 ();
 FILLCELL_X32 FILLER_426_3190 ();
 FILLCELL_X32 FILLER_426_3222 ();
 FILLCELL_X32 FILLER_426_3254 ();
 FILLCELL_X32 FILLER_426_3286 ();
 FILLCELL_X32 FILLER_426_3318 ();
 FILLCELL_X32 FILLER_426_3350 ();
 FILLCELL_X32 FILLER_426_3382 ();
 FILLCELL_X32 FILLER_426_3414 ();
 FILLCELL_X32 FILLER_426_3446 ();
 FILLCELL_X32 FILLER_426_3478 ();
 FILLCELL_X32 FILLER_426_3510 ();
 FILLCELL_X32 FILLER_426_3542 ();
 FILLCELL_X32 FILLER_426_3574 ();
 FILLCELL_X32 FILLER_426_3606 ();
 FILLCELL_X32 FILLER_426_3638 ();
 FILLCELL_X32 FILLER_426_3670 ();
 FILLCELL_X32 FILLER_426_3702 ();
 FILLCELL_X4 FILLER_426_3734 ();
 FILLCELL_X32 FILLER_427_1 ();
 FILLCELL_X32 FILLER_427_33 ();
 FILLCELL_X32 FILLER_427_65 ();
 FILLCELL_X32 FILLER_427_97 ();
 FILLCELL_X32 FILLER_427_129 ();
 FILLCELL_X32 FILLER_427_161 ();
 FILLCELL_X32 FILLER_427_193 ();
 FILLCELL_X32 FILLER_427_225 ();
 FILLCELL_X32 FILLER_427_257 ();
 FILLCELL_X32 FILLER_427_289 ();
 FILLCELL_X32 FILLER_427_321 ();
 FILLCELL_X32 FILLER_427_353 ();
 FILLCELL_X32 FILLER_427_385 ();
 FILLCELL_X32 FILLER_427_417 ();
 FILLCELL_X32 FILLER_427_449 ();
 FILLCELL_X32 FILLER_427_481 ();
 FILLCELL_X32 FILLER_427_513 ();
 FILLCELL_X32 FILLER_427_545 ();
 FILLCELL_X32 FILLER_427_577 ();
 FILLCELL_X32 FILLER_427_609 ();
 FILLCELL_X32 FILLER_427_641 ();
 FILLCELL_X32 FILLER_427_673 ();
 FILLCELL_X32 FILLER_427_705 ();
 FILLCELL_X32 FILLER_427_737 ();
 FILLCELL_X32 FILLER_427_769 ();
 FILLCELL_X32 FILLER_427_801 ();
 FILLCELL_X32 FILLER_427_833 ();
 FILLCELL_X32 FILLER_427_865 ();
 FILLCELL_X32 FILLER_427_897 ();
 FILLCELL_X32 FILLER_427_929 ();
 FILLCELL_X32 FILLER_427_961 ();
 FILLCELL_X32 FILLER_427_993 ();
 FILLCELL_X32 FILLER_427_1025 ();
 FILLCELL_X32 FILLER_427_1057 ();
 FILLCELL_X32 FILLER_427_1089 ();
 FILLCELL_X32 FILLER_427_1121 ();
 FILLCELL_X32 FILLER_427_1153 ();
 FILLCELL_X32 FILLER_427_1185 ();
 FILLCELL_X32 FILLER_427_1217 ();
 FILLCELL_X8 FILLER_427_1249 ();
 FILLCELL_X4 FILLER_427_1257 ();
 FILLCELL_X2 FILLER_427_1261 ();
 FILLCELL_X32 FILLER_427_1264 ();
 FILLCELL_X32 FILLER_427_1296 ();
 FILLCELL_X32 FILLER_427_1328 ();
 FILLCELL_X32 FILLER_427_1360 ();
 FILLCELL_X32 FILLER_427_1392 ();
 FILLCELL_X32 FILLER_427_1424 ();
 FILLCELL_X32 FILLER_427_1456 ();
 FILLCELL_X32 FILLER_427_1488 ();
 FILLCELL_X32 FILLER_427_1520 ();
 FILLCELL_X32 FILLER_427_1552 ();
 FILLCELL_X32 FILLER_427_1584 ();
 FILLCELL_X32 FILLER_427_1616 ();
 FILLCELL_X32 FILLER_427_1648 ();
 FILLCELL_X32 FILLER_427_1680 ();
 FILLCELL_X32 FILLER_427_1712 ();
 FILLCELL_X32 FILLER_427_1744 ();
 FILLCELL_X32 FILLER_427_1776 ();
 FILLCELL_X32 FILLER_427_1808 ();
 FILLCELL_X32 FILLER_427_1840 ();
 FILLCELL_X32 FILLER_427_1872 ();
 FILLCELL_X32 FILLER_427_1904 ();
 FILLCELL_X32 FILLER_427_1936 ();
 FILLCELL_X32 FILLER_427_1968 ();
 FILLCELL_X32 FILLER_427_2000 ();
 FILLCELL_X32 FILLER_427_2032 ();
 FILLCELL_X32 FILLER_427_2064 ();
 FILLCELL_X32 FILLER_427_2096 ();
 FILLCELL_X32 FILLER_427_2128 ();
 FILLCELL_X32 FILLER_427_2160 ();
 FILLCELL_X32 FILLER_427_2192 ();
 FILLCELL_X32 FILLER_427_2224 ();
 FILLCELL_X32 FILLER_427_2256 ();
 FILLCELL_X32 FILLER_427_2288 ();
 FILLCELL_X32 FILLER_427_2320 ();
 FILLCELL_X32 FILLER_427_2352 ();
 FILLCELL_X32 FILLER_427_2384 ();
 FILLCELL_X32 FILLER_427_2416 ();
 FILLCELL_X32 FILLER_427_2448 ();
 FILLCELL_X32 FILLER_427_2480 ();
 FILLCELL_X8 FILLER_427_2512 ();
 FILLCELL_X4 FILLER_427_2520 ();
 FILLCELL_X2 FILLER_427_2524 ();
 FILLCELL_X32 FILLER_427_2527 ();
 FILLCELL_X32 FILLER_427_2559 ();
 FILLCELL_X32 FILLER_427_2591 ();
 FILLCELL_X32 FILLER_427_2623 ();
 FILLCELL_X32 FILLER_427_2655 ();
 FILLCELL_X32 FILLER_427_2687 ();
 FILLCELL_X32 FILLER_427_2719 ();
 FILLCELL_X32 FILLER_427_2751 ();
 FILLCELL_X32 FILLER_427_2783 ();
 FILLCELL_X32 FILLER_427_2815 ();
 FILLCELL_X32 FILLER_427_2847 ();
 FILLCELL_X32 FILLER_427_2879 ();
 FILLCELL_X32 FILLER_427_2911 ();
 FILLCELL_X32 FILLER_427_2943 ();
 FILLCELL_X32 FILLER_427_2975 ();
 FILLCELL_X32 FILLER_427_3007 ();
 FILLCELL_X32 FILLER_427_3039 ();
 FILLCELL_X32 FILLER_427_3071 ();
 FILLCELL_X32 FILLER_427_3103 ();
 FILLCELL_X32 FILLER_427_3135 ();
 FILLCELL_X32 FILLER_427_3167 ();
 FILLCELL_X32 FILLER_427_3199 ();
 FILLCELL_X32 FILLER_427_3231 ();
 FILLCELL_X32 FILLER_427_3263 ();
 FILLCELL_X32 FILLER_427_3295 ();
 FILLCELL_X32 FILLER_427_3327 ();
 FILLCELL_X32 FILLER_427_3359 ();
 FILLCELL_X32 FILLER_427_3391 ();
 FILLCELL_X32 FILLER_427_3423 ();
 FILLCELL_X32 FILLER_427_3455 ();
 FILLCELL_X32 FILLER_427_3487 ();
 FILLCELL_X32 FILLER_427_3519 ();
 FILLCELL_X32 FILLER_427_3551 ();
 FILLCELL_X32 FILLER_427_3583 ();
 FILLCELL_X32 FILLER_427_3615 ();
 FILLCELL_X32 FILLER_427_3647 ();
 FILLCELL_X32 FILLER_427_3679 ();
 FILLCELL_X16 FILLER_427_3711 ();
 FILLCELL_X8 FILLER_427_3727 ();
 FILLCELL_X2 FILLER_427_3735 ();
 FILLCELL_X1 FILLER_427_3737 ();
 FILLCELL_X32 FILLER_428_1 ();
 FILLCELL_X32 FILLER_428_33 ();
 FILLCELL_X32 FILLER_428_65 ();
 FILLCELL_X32 FILLER_428_97 ();
 FILLCELL_X32 FILLER_428_129 ();
 FILLCELL_X32 FILLER_428_161 ();
 FILLCELL_X32 FILLER_428_193 ();
 FILLCELL_X32 FILLER_428_225 ();
 FILLCELL_X32 FILLER_428_257 ();
 FILLCELL_X32 FILLER_428_289 ();
 FILLCELL_X32 FILLER_428_321 ();
 FILLCELL_X32 FILLER_428_353 ();
 FILLCELL_X32 FILLER_428_385 ();
 FILLCELL_X32 FILLER_428_417 ();
 FILLCELL_X32 FILLER_428_449 ();
 FILLCELL_X32 FILLER_428_481 ();
 FILLCELL_X32 FILLER_428_513 ();
 FILLCELL_X32 FILLER_428_545 ();
 FILLCELL_X32 FILLER_428_577 ();
 FILLCELL_X16 FILLER_428_609 ();
 FILLCELL_X4 FILLER_428_625 ();
 FILLCELL_X2 FILLER_428_629 ();
 FILLCELL_X32 FILLER_428_632 ();
 FILLCELL_X32 FILLER_428_664 ();
 FILLCELL_X32 FILLER_428_696 ();
 FILLCELL_X32 FILLER_428_728 ();
 FILLCELL_X32 FILLER_428_760 ();
 FILLCELL_X32 FILLER_428_792 ();
 FILLCELL_X32 FILLER_428_824 ();
 FILLCELL_X32 FILLER_428_856 ();
 FILLCELL_X32 FILLER_428_888 ();
 FILLCELL_X32 FILLER_428_920 ();
 FILLCELL_X32 FILLER_428_952 ();
 FILLCELL_X32 FILLER_428_984 ();
 FILLCELL_X32 FILLER_428_1016 ();
 FILLCELL_X32 FILLER_428_1048 ();
 FILLCELL_X32 FILLER_428_1080 ();
 FILLCELL_X32 FILLER_428_1112 ();
 FILLCELL_X32 FILLER_428_1144 ();
 FILLCELL_X32 FILLER_428_1176 ();
 FILLCELL_X32 FILLER_428_1208 ();
 FILLCELL_X32 FILLER_428_1240 ();
 FILLCELL_X32 FILLER_428_1272 ();
 FILLCELL_X32 FILLER_428_1304 ();
 FILLCELL_X32 FILLER_428_1336 ();
 FILLCELL_X32 FILLER_428_1368 ();
 FILLCELL_X32 FILLER_428_1400 ();
 FILLCELL_X32 FILLER_428_1432 ();
 FILLCELL_X32 FILLER_428_1464 ();
 FILLCELL_X32 FILLER_428_1496 ();
 FILLCELL_X32 FILLER_428_1528 ();
 FILLCELL_X32 FILLER_428_1560 ();
 FILLCELL_X32 FILLER_428_1592 ();
 FILLCELL_X32 FILLER_428_1624 ();
 FILLCELL_X32 FILLER_428_1656 ();
 FILLCELL_X32 FILLER_428_1688 ();
 FILLCELL_X32 FILLER_428_1720 ();
 FILLCELL_X32 FILLER_428_1752 ();
 FILLCELL_X32 FILLER_428_1784 ();
 FILLCELL_X32 FILLER_428_1816 ();
 FILLCELL_X32 FILLER_428_1848 ();
 FILLCELL_X8 FILLER_428_1880 ();
 FILLCELL_X4 FILLER_428_1888 ();
 FILLCELL_X2 FILLER_428_1892 ();
 FILLCELL_X32 FILLER_428_1895 ();
 FILLCELL_X32 FILLER_428_1927 ();
 FILLCELL_X32 FILLER_428_1959 ();
 FILLCELL_X32 FILLER_428_1991 ();
 FILLCELL_X32 FILLER_428_2023 ();
 FILLCELL_X32 FILLER_428_2055 ();
 FILLCELL_X32 FILLER_428_2087 ();
 FILLCELL_X32 FILLER_428_2119 ();
 FILLCELL_X32 FILLER_428_2151 ();
 FILLCELL_X32 FILLER_428_2183 ();
 FILLCELL_X32 FILLER_428_2215 ();
 FILLCELL_X32 FILLER_428_2247 ();
 FILLCELL_X32 FILLER_428_2279 ();
 FILLCELL_X32 FILLER_428_2311 ();
 FILLCELL_X32 FILLER_428_2343 ();
 FILLCELL_X32 FILLER_428_2375 ();
 FILLCELL_X32 FILLER_428_2407 ();
 FILLCELL_X32 FILLER_428_2439 ();
 FILLCELL_X32 FILLER_428_2471 ();
 FILLCELL_X32 FILLER_428_2503 ();
 FILLCELL_X32 FILLER_428_2535 ();
 FILLCELL_X32 FILLER_428_2567 ();
 FILLCELL_X32 FILLER_428_2599 ();
 FILLCELL_X32 FILLER_428_2631 ();
 FILLCELL_X32 FILLER_428_2663 ();
 FILLCELL_X32 FILLER_428_2695 ();
 FILLCELL_X32 FILLER_428_2727 ();
 FILLCELL_X32 FILLER_428_2759 ();
 FILLCELL_X32 FILLER_428_2791 ();
 FILLCELL_X32 FILLER_428_2823 ();
 FILLCELL_X32 FILLER_428_2855 ();
 FILLCELL_X32 FILLER_428_2887 ();
 FILLCELL_X32 FILLER_428_2919 ();
 FILLCELL_X32 FILLER_428_2951 ();
 FILLCELL_X32 FILLER_428_2983 ();
 FILLCELL_X32 FILLER_428_3015 ();
 FILLCELL_X32 FILLER_428_3047 ();
 FILLCELL_X32 FILLER_428_3079 ();
 FILLCELL_X32 FILLER_428_3111 ();
 FILLCELL_X8 FILLER_428_3143 ();
 FILLCELL_X4 FILLER_428_3151 ();
 FILLCELL_X2 FILLER_428_3155 ();
 FILLCELL_X32 FILLER_428_3158 ();
 FILLCELL_X32 FILLER_428_3190 ();
 FILLCELL_X32 FILLER_428_3222 ();
 FILLCELL_X32 FILLER_428_3254 ();
 FILLCELL_X32 FILLER_428_3286 ();
 FILLCELL_X32 FILLER_428_3318 ();
 FILLCELL_X32 FILLER_428_3350 ();
 FILLCELL_X32 FILLER_428_3382 ();
 FILLCELL_X32 FILLER_428_3414 ();
 FILLCELL_X32 FILLER_428_3446 ();
 FILLCELL_X32 FILLER_428_3478 ();
 FILLCELL_X32 FILLER_428_3510 ();
 FILLCELL_X32 FILLER_428_3542 ();
 FILLCELL_X32 FILLER_428_3574 ();
 FILLCELL_X32 FILLER_428_3606 ();
 FILLCELL_X32 FILLER_428_3638 ();
 FILLCELL_X32 FILLER_428_3670 ();
 FILLCELL_X32 FILLER_428_3702 ();
 FILLCELL_X4 FILLER_428_3734 ();
 FILLCELL_X32 FILLER_429_1 ();
 FILLCELL_X32 FILLER_429_33 ();
 FILLCELL_X32 FILLER_429_65 ();
 FILLCELL_X32 FILLER_429_97 ();
 FILLCELL_X32 FILLER_429_129 ();
 FILLCELL_X32 FILLER_429_161 ();
 FILLCELL_X32 FILLER_429_193 ();
 FILLCELL_X32 FILLER_429_225 ();
 FILLCELL_X32 FILLER_429_257 ();
 FILLCELL_X32 FILLER_429_289 ();
 FILLCELL_X32 FILLER_429_321 ();
 FILLCELL_X32 FILLER_429_353 ();
 FILLCELL_X32 FILLER_429_385 ();
 FILLCELL_X32 FILLER_429_417 ();
 FILLCELL_X32 FILLER_429_449 ();
 FILLCELL_X32 FILLER_429_481 ();
 FILLCELL_X32 FILLER_429_513 ();
 FILLCELL_X32 FILLER_429_545 ();
 FILLCELL_X32 FILLER_429_577 ();
 FILLCELL_X32 FILLER_429_609 ();
 FILLCELL_X32 FILLER_429_641 ();
 FILLCELL_X32 FILLER_429_673 ();
 FILLCELL_X32 FILLER_429_705 ();
 FILLCELL_X32 FILLER_429_737 ();
 FILLCELL_X32 FILLER_429_769 ();
 FILLCELL_X32 FILLER_429_801 ();
 FILLCELL_X32 FILLER_429_833 ();
 FILLCELL_X32 FILLER_429_865 ();
 FILLCELL_X32 FILLER_429_897 ();
 FILLCELL_X32 FILLER_429_929 ();
 FILLCELL_X32 FILLER_429_961 ();
 FILLCELL_X32 FILLER_429_993 ();
 FILLCELL_X32 FILLER_429_1025 ();
 FILLCELL_X32 FILLER_429_1057 ();
 FILLCELL_X32 FILLER_429_1089 ();
 FILLCELL_X32 FILLER_429_1121 ();
 FILLCELL_X32 FILLER_429_1153 ();
 FILLCELL_X32 FILLER_429_1185 ();
 FILLCELL_X32 FILLER_429_1217 ();
 FILLCELL_X8 FILLER_429_1249 ();
 FILLCELL_X4 FILLER_429_1257 ();
 FILLCELL_X2 FILLER_429_1261 ();
 FILLCELL_X32 FILLER_429_1264 ();
 FILLCELL_X32 FILLER_429_1296 ();
 FILLCELL_X32 FILLER_429_1328 ();
 FILLCELL_X32 FILLER_429_1360 ();
 FILLCELL_X32 FILLER_429_1392 ();
 FILLCELL_X32 FILLER_429_1424 ();
 FILLCELL_X32 FILLER_429_1456 ();
 FILLCELL_X32 FILLER_429_1488 ();
 FILLCELL_X32 FILLER_429_1520 ();
 FILLCELL_X32 FILLER_429_1552 ();
 FILLCELL_X32 FILLER_429_1584 ();
 FILLCELL_X32 FILLER_429_1616 ();
 FILLCELL_X32 FILLER_429_1648 ();
 FILLCELL_X32 FILLER_429_1680 ();
 FILLCELL_X32 FILLER_429_1712 ();
 FILLCELL_X32 FILLER_429_1744 ();
 FILLCELL_X32 FILLER_429_1776 ();
 FILLCELL_X32 FILLER_429_1808 ();
 FILLCELL_X32 FILLER_429_1840 ();
 FILLCELL_X32 FILLER_429_1872 ();
 FILLCELL_X32 FILLER_429_1904 ();
 FILLCELL_X32 FILLER_429_1936 ();
 FILLCELL_X32 FILLER_429_1968 ();
 FILLCELL_X32 FILLER_429_2000 ();
 FILLCELL_X32 FILLER_429_2032 ();
 FILLCELL_X32 FILLER_429_2064 ();
 FILLCELL_X32 FILLER_429_2096 ();
 FILLCELL_X32 FILLER_429_2128 ();
 FILLCELL_X32 FILLER_429_2160 ();
 FILLCELL_X32 FILLER_429_2192 ();
 FILLCELL_X32 FILLER_429_2224 ();
 FILLCELL_X32 FILLER_429_2256 ();
 FILLCELL_X32 FILLER_429_2288 ();
 FILLCELL_X32 FILLER_429_2320 ();
 FILLCELL_X32 FILLER_429_2352 ();
 FILLCELL_X32 FILLER_429_2384 ();
 FILLCELL_X32 FILLER_429_2416 ();
 FILLCELL_X32 FILLER_429_2448 ();
 FILLCELL_X32 FILLER_429_2480 ();
 FILLCELL_X8 FILLER_429_2512 ();
 FILLCELL_X4 FILLER_429_2520 ();
 FILLCELL_X2 FILLER_429_2524 ();
 FILLCELL_X32 FILLER_429_2527 ();
 FILLCELL_X32 FILLER_429_2559 ();
 FILLCELL_X32 FILLER_429_2591 ();
 FILLCELL_X32 FILLER_429_2623 ();
 FILLCELL_X32 FILLER_429_2655 ();
 FILLCELL_X32 FILLER_429_2687 ();
 FILLCELL_X32 FILLER_429_2719 ();
 FILLCELL_X32 FILLER_429_2751 ();
 FILLCELL_X32 FILLER_429_2783 ();
 FILLCELL_X32 FILLER_429_2815 ();
 FILLCELL_X32 FILLER_429_2847 ();
 FILLCELL_X32 FILLER_429_2879 ();
 FILLCELL_X32 FILLER_429_2911 ();
 FILLCELL_X32 FILLER_429_2943 ();
 FILLCELL_X32 FILLER_429_2975 ();
 FILLCELL_X32 FILLER_429_3007 ();
 FILLCELL_X32 FILLER_429_3039 ();
 FILLCELL_X32 FILLER_429_3071 ();
 FILLCELL_X32 FILLER_429_3103 ();
 FILLCELL_X32 FILLER_429_3135 ();
 FILLCELL_X32 FILLER_429_3167 ();
 FILLCELL_X32 FILLER_429_3199 ();
 FILLCELL_X32 FILLER_429_3231 ();
 FILLCELL_X32 FILLER_429_3263 ();
 FILLCELL_X32 FILLER_429_3295 ();
 FILLCELL_X32 FILLER_429_3327 ();
 FILLCELL_X32 FILLER_429_3359 ();
 FILLCELL_X32 FILLER_429_3391 ();
 FILLCELL_X32 FILLER_429_3423 ();
 FILLCELL_X32 FILLER_429_3455 ();
 FILLCELL_X32 FILLER_429_3487 ();
 FILLCELL_X32 FILLER_429_3519 ();
 FILLCELL_X32 FILLER_429_3551 ();
 FILLCELL_X32 FILLER_429_3583 ();
 FILLCELL_X32 FILLER_429_3615 ();
 FILLCELL_X32 FILLER_429_3647 ();
 FILLCELL_X32 FILLER_429_3679 ();
 FILLCELL_X16 FILLER_429_3711 ();
 FILLCELL_X8 FILLER_429_3727 ();
 FILLCELL_X2 FILLER_429_3735 ();
 FILLCELL_X1 FILLER_429_3737 ();
 FILLCELL_X32 FILLER_430_1 ();
 FILLCELL_X32 FILLER_430_33 ();
 FILLCELL_X32 FILLER_430_65 ();
 FILLCELL_X32 FILLER_430_97 ();
 FILLCELL_X32 FILLER_430_129 ();
 FILLCELL_X32 FILLER_430_161 ();
 FILLCELL_X32 FILLER_430_193 ();
 FILLCELL_X32 FILLER_430_225 ();
 FILLCELL_X32 FILLER_430_257 ();
 FILLCELL_X32 FILLER_430_289 ();
 FILLCELL_X32 FILLER_430_321 ();
 FILLCELL_X32 FILLER_430_353 ();
 FILLCELL_X32 FILLER_430_385 ();
 FILLCELL_X32 FILLER_430_417 ();
 FILLCELL_X32 FILLER_430_449 ();
 FILLCELL_X32 FILLER_430_481 ();
 FILLCELL_X32 FILLER_430_513 ();
 FILLCELL_X32 FILLER_430_545 ();
 FILLCELL_X32 FILLER_430_577 ();
 FILLCELL_X16 FILLER_430_609 ();
 FILLCELL_X4 FILLER_430_625 ();
 FILLCELL_X2 FILLER_430_629 ();
 FILLCELL_X32 FILLER_430_632 ();
 FILLCELL_X32 FILLER_430_664 ();
 FILLCELL_X32 FILLER_430_696 ();
 FILLCELL_X32 FILLER_430_728 ();
 FILLCELL_X32 FILLER_430_760 ();
 FILLCELL_X32 FILLER_430_792 ();
 FILLCELL_X32 FILLER_430_824 ();
 FILLCELL_X32 FILLER_430_856 ();
 FILLCELL_X32 FILLER_430_888 ();
 FILLCELL_X32 FILLER_430_920 ();
 FILLCELL_X32 FILLER_430_952 ();
 FILLCELL_X32 FILLER_430_984 ();
 FILLCELL_X32 FILLER_430_1016 ();
 FILLCELL_X32 FILLER_430_1048 ();
 FILLCELL_X32 FILLER_430_1080 ();
 FILLCELL_X32 FILLER_430_1112 ();
 FILLCELL_X32 FILLER_430_1144 ();
 FILLCELL_X32 FILLER_430_1176 ();
 FILLCELL_X32 FILLER_430_1208 ();
 FILLCELL_X32 FILLER_430_1240 ();
 FILLCELL_X32 FILLER_430_1272 ();
 FILLCELL_X32 FILLER_430_1304 ();
 FILLCELL_X32 FILLER_430_1336 ();
 FILLCELL_X32 FILLER_430_1368 ();
 FILLCELL_X32 FILLER_430_1400 ();
 FILLCELL_X32 FILLER_430_1432 ();
 FILLCELL_X32 FILLER_430_1464 ();
 FILLCELL_X32 FILLER_430_1496 ();
 FILLCELL_X32 FILLER_430_1528 ();
 FILLCELL_X32 FILLER_430_1560 ();
 FILLCELL_X32 FILLER_430_1592 ();
 FILLCELL_X32 FILLER_430_1624 ();
 FILLCELL_X32 FILLER_430_1656 ();
 FILLCELL_X32 FILLER_430_1688 ();
 FILLCELL_X32 FILLER_430_1720 ();
 FILLCELL_X32 FILLER_430_1752 ();
 FILLCELL_X32 FILLER_430_1784 ();
 FILLCELL_X32 FILLER_430_1816 ();
 FILLCELL_X32 FILLER_430_1848 ();
 FILLCELL_X8 FILLER_430_1880 ();
 FILLCELL_X4 FILLER_430_1888 ();
 FILLCELL_X2 FILLER_430_1892 ();
 FILLCELL_X32 FILLER_430_1895 ();
 FILLCELL_X32 FILLER_430_1927 ();
 FILLCELL_X32 FILLER_430_1959 ();
 FILLCELL_X32 FILLER_430_1991 ();
 FILLCELL_X32 FILLER_430_2023 ();
 FILLCELL_X32 FILLER_430_2055 ();
 FILLCELL_X32 FILLER_430_2087 ();
 FILLCELL_X32 FILLER_430_2119 ();
 FILLCELL_X32 FILLER_430_2151 ();
 FILLCELL_X32 FILLER_430_2183 ();
 FILLCELL_X32 FILLER_430_2215 ();
 FILLCELL_X32 FILLER_430_2247 ();
 FILLCELL_X32 FILLER_430_2279 ();
 FILLCELL_X32 FILLER_430_2311 ();
 FILLCELL_X32 FILLER_430_2343 ();
 FILLCELL_X32 FILLER_430_2375 ();
 FILLCELL_X32 FILLER_430_2407 ();
 FILLCELL_X32 FILLER_430_2439 ();
 FILLCELL_X32 FILLER_430_2471 ();
 FILLCELL_X32 FILLER_430_2503 ();
 FILLCELL_X32 FILLER_430_2535 ();
 FILLCELL_X32 FILLER_430_2567 ();
 FILLCELL_X32 FILLER_430_2599 ();
 FILLCELL_X32 FILLER_430_2631 ();
 FILLCELL_X32 FILLER_430_2663 ();
 FILLCELL_X32 FILLER_430_2695 ();
 FILLCELL_X32 FILLER_430_2727 ();
 FILLCELL_X32 FILLER_430_2759 ();
 FILLCELL_X32 FILLER_430_2791 ();
 FILLCELL_X32 FILLER_430_2823 ();
 FILLCELL_X32 FILLER_430_2855 ();
 FILLCELL_X32 FILLER_430_2887 ();
 FILLCELL_X32 FILLER_430_2919 ();
 FILLCELL_X32 FILLER_430_2951 ();
 FILLCELL_X32 FILLER_430_2983 ();
 FILLCELL_X32 FILLER_430_3015 ();
 FILLCELL_X32 FILLER_430_3047 ();
 FILLCELL_X32 FILLER_430_3079 ();
 FILLCELL_X32 FILLER_430_3111 ();
 FILLCELL_X8 FILLER_430_3143 ();
 FILLCELL_X4 FILLER_430_3151 ();
 FILLCELL_X2 FILLER_430_3155 ();
 FILLCELL_X32 FILLER_430_3158 ();
 FILLCELL_X32 FILLER_430_3190 ();
 FILLCELL_X32 FILLER_430_3222 ();
 FILLCELL_X32 FILLER_430_3254 ();
 FILLCELL_X32 FILLER_430_3286 ();
 FILLCELL_X32 FILLER_430_3318 ();
 FILLCELL_X32 FILLER_430_3350 ();
 FILLCELL_X32 FILLER_430_3382 ();
 FILLCELL_X32 FILLER_430_3414 ();
 FILLCELL_X32 FILLER_430_3446 ();
 FILLCELL_X32 FILLER_430_3478 ();
 FILLCELL_X32 FILLER_430_3510 ();
 FILLCELL_X32 FILLER_430_3542 ();
 FILLCELL_X32 FILLER_430_3574 ();
 FILLCELL_X32 FILLER_430_3606 ();
 FILLCELL_X32 FILLER_430_3638 ();
 FILLCELL_X32 FILLER_430_3670 ();
 FILLCELL_X32 FILLER_430_3702 ();
 FILLCELL_X4 FILLER_430_3734 ();
 FILLCELL_X32 FILLER_431_1 ();
 FILLCELL_X32 FILLER_431_33 ();
 FILLCELL_X32 FILLER_431_65 ();
 FILLCELL_X32 FILLER_431_97 ();
 FILLCELL_X32 FILLER_431_129 ();
 FILLCELL_X32 FILLER_431_161 ();
 FILLCELL_X32 FILLER_431_193 ();
 FILLCELL_X32 FILLER_431_225 ();
 FILLCELL_X32 FILLER_431_257 ();
 FILLCELL_X32 FILLER_431_289 ();
 FILLCELL_X32 FILLER_431_321 ();
 FILLCELL_X32 FILLER_431_353 ();
 FILLCELL_X32 FILLER_431_385 ();
 FILLCELL_X32 FILLER_431_417 ();
 FILLCELL_X32 FILLER_431_449 ();
 FILLCELL_X32 FILLER_431_481 ();
 FILLCELL_X32 FILLER_431_513 ();
 FILLCELL_X32 FILLER_431_545 ();
 FILLCELL_X32 FILLER_431_577 ();
 FILLCELL_X32 FILLER_431_609 ();
 FILLCELL_X32 FILLER_431_641 ();
 FILLCELL_X32 FILLER_431_673 ();
 FILLCELL_X32 FILLER_431_705 ();
 FILLCELL_X32 FILLER_431_737 ();
 FILLCELL_X32 FILLER_431_769 ();
 FILLCELL_X32 FILLER_431_801 ();
 FILLCELL_X32 FILLER_431_833 ();
 FILLCELL_X32 FILLER_431_865 ();
 FILLCELL_X32 FILLER_431_897 ();
 FILLCELL_X32 FILLER_431_929 ();
 FILLCELL_X32 FILLER_431_961 ();
 FILLCELL_X32 FILLER_431_993 ();
 FILLCELL_X32 FILLER_431_1025 ();
 FILLCELL_X32 FILLER_431_1057 ();
 FILLCELL_X32 FILLER_431_1089 ();
 FILLCELL_X32 FILLER_431_1121 ();
 FILLCELL_X32 FILLER_431_1153 ();
 FILLCELL_X32 FILLER_431_1185 ();
 FILLCELL_X32 FILLER_431_1217 ();
 FILLCELL_X8 FILLER_431_1249 ();
 FILLCELL_X4 FILLER_431_1257 ();
 FILLCELL_X2 FILLER_431_1261 ();
 FILLCELL_X32 FILLER_431_1264 ();
 FILLCELL_X32 FILLER_431_1296 ();
 FILLCELL_X32 FILLER_431_1328 ();
 FILLCELL_X32 FILLER_431_1360 ();
 FILLCELL_X32 FILLER_431_1392 ();
 FILLCELL_X32 FILLER_431_1424 ();
 FILLCELL_X32 FILLER_431_1456 ();
 FILLCELL_X32 FILLER_431_1488 ();
 FILLCELL_X32 FILLER_431_1520 ();
 FILLCELL_X32 FILLER_431_1552 ();
 FILLCELL_X32 FILLER_431_1584 ();
 FILLCELL_X32 FILLER_431_1616 ();
 FILLCELL_X32 FILLER_431_1648 ();
 FILLCELL_X32 FILLER_431_1680 ();
 FILLCELL_X32 FILLER_431_1712 ();
 FILLCELL_X32 FILLER_431_1744 ();
 FILLCELL_X32 FILLER_431_1776 ();
 FILLCELL_X32 FILLER_431_1808 ();
 FILLCELL_X32 FILLER_431_1840 ();
 FILLCELL_X32 FILLER_431_1872 ();
 FILLCELL_X32 FILLER_431_1904 ();
 FILLCELL_X32 FILLER_431_1936 ();
 FILLCELL_X32 FILLER_431_1968 ();
 FILLCELL_X32 FILLER_431_2000 ();
 FILLCELL_X32 FILLER_431_2032 ();
 FILLCELL_X32 FILLER_431_2064 ();
 FILLCELL_X32 FILLER_431_2096 ();
 FILLCELL_X32 FILLER_431_2128 ();
 FILLCELL_X32 FILLER_431_2160 ();
 FILLCELL_X32 FILLER_431_2192 ();
 FILLCELL_X32 FILLER_431_2224 ();
 FILLCELL_X32 FILLER_431_2256 ();
 FILLCELL_X32 FILLER_431_2288 ();
 FILLCELL_X32 FILLER_431_2320 ();
 FILLCELL_X32 FILLER_431_2352 ();
 FILLCELL_X32 FILLER_431_2384 ();
 FILLCELL_X32 FILLER_431_2416 ();
 FILLCELL_X32 FILLER_431_2448 ();
 FILLCELL_X32 FILLER_431_2480 ();
 FILLCELL_X8 FILLER_431_2512 ();
 FILLCELL_X4 FILLER_431_2520 ();
 FILLCELL_X2 FILLER_431_2524 ();
 FILLCELL_X32 FILLER_431_2527 ();
 FILLCELL_X32 FILLER_431_2559 ();
 FILLCELL_X32 FILLER_431_2591 ();
 FILLCELL_X32 FILLER_431_2623 ();
 FILLCELL_X32 FILLER_431_2655 ();
 FILLCELL_X32 FILLER_431_2687 ();
 FILLCELL_X32 FILLER_431_2719 ();
 FILLCELL_X32 FILLER_431_2751 ();
 FILLCELL_X32 FILLER_431_2783 ();
 FILLCELL_X32 FILLER_431_2815 ();
 FILLCELL_X32 FILLER_431_2847 ();
 FILLCELL_X32 FILLER_431_2879 ();
 FILLCELL_X32 FILLER_431_2911 ();
 FILLCELL_X32 FILLER_431_2943 ();
 FILLCELL_X32 FILLER_431_2975 ();
 FILLCELL_X32 FILLER_431_3007 ();
 FILLCELL_X32 FILLER_431_3039 ();
 FILLCELL_X32 FILLER_431_3071 ();
 FILLCELL_X32 FILLER_431_3103 ();
 FILLCELL_X32 FILLER_431_3135 ();
 FILLCELL_X32 FILLER_431_3167 ();
 FILLCELL_X32 FILLER_431_3199 ();
 FILLCELL_X32 FILLER_431_3231 ();
 FILLCELL_X32 FILLER_431_3263 ();
 FILLCELL_X32 FILLER_431_3295 ();
 FILLCELL_X32 FILLER_431_3327 ();
 FILLCELL_X32 FILLER_431_3359 ();
 FILLCELL_X32 FILLER_431_3391 ();
 FILLCELL_X32 FILLER_431_3423 ();
 FILLCELL_X32 FILLER_431_3455 ();
 FILLCELL_X32 FILLER_431_3487 ();
 FILLCELL_X32 FILLER_431_3519 ();
 FILLCELL_X32 FILLER_431_3551 ();
 FILLCELL_X32 FILLER_431_3583 ();
 FILLCELL_X32 FILLER_431_3615 ();
 FILLCELL_X32 FILLER_431_3647 ();
 FILLCELL_X32 FILLER_431_3679 ();
 FILLCELL_X16 FILLER_431_3711 ();
 FILLCELL_X8 FILLER_431_3727 ();
 FILLCELL_X2 FILLER_431_3735 ();
 FILLCELL_X1 FILLER_431_3737 ();
 FILLCELL_X32 FILLER_432_1 ();
 FILLCELL_X32 FILLER_432_33 ();
 FILLCELL_X32 FILLER_432_65 ();
 FILLCELL_X32 FILLER_432_97 ();
 FILLCELL_X32 FILLER_432_129 ();
 FILLCELL_X32 FILLER_432_161 ();
 FILLCELL_X32 FILLER_432_193 ();
 FILLCELL_X32 FILLER_432_225 ();
 FILLCELL_X32 FILLER_432_257 ();
 FILLCELL_X32 FILLER_432_289 ();
 FILLCELL_X32 FILLER_432_321 ();
 FILLCELL_X32 FILLER_432_353 ();
 FILLCELL_X32 FILLER_432_385 ();
 FILLCELL_X32 FILLER_432_417 ();
 FILLCELL_X32 FILLER_432_449 ();
 FILLCELL_X32 FILLER_432_481 ();
 FILLCELL_X32 FILLER_432_513 ();
 FILLCELL_X32 FILLER_432_545 ();
 FILLCELL_X32 FILLER_432_577 ();
 FILLCELL_X16 FILLER_432_609 ();
 FILLCELL_X4 FILLER_432_625 ();
 FILLCELL_X2 FILLER_432_629 ();
 FILLCELL_X32 FILLER_432_632 ();
 FILLCELL_X32 FILLER_432_664 ();
 FILLCELL_X32 FILLER_432_696 ();
 FILLCELL_X32 FILLER_432_728 ();
 FILLCELL_X32 FILLER_432_760 ();
 FILLCELL_X32 FILLER_432_792 ();
 FILLCELL_X32 FILLER_432_824 ();
 FILLCELL_X32 FILLER_432_856 ();
 FILLCELL_X32 FILLER_432_888 ();
 FILLCELL_X32 FILLER_432_920 ();
 FILLCELL_X32 FILLER_432_952 ();
 FILLCELL_X32 FILLER_432_984 ();
 FILLCELL_X32 FILLER_432_1016 ();
 FILLCELL_X32 FILLER_432_1048 ();
 FILLCELL_X32 FILLER_432_1080 ();
 FILLCELL_X32 FILLER_432_1112 ();
 FILLCELL_X32 FILLER_432_1144 ();
 FILLCELL_X32 FILLER_432_1176 ();
 FILLCELL_X32 FILLER_432_1208 ();
 FILLCELL_X32 FILLER_432_1240 ();
 FILLCELL_X32 FILLER_432_1272 ();
 FILLCELL_X32 FILLER_432_1304 ();
 FILLCELL_X32 FILLER_432_1336 ();
 FILLCELL_X32 FILLER_432_1368 ();
 FILLCELL_X32 FILLER_432_1400 ();
 FILLCELL_X32 FILLER_432_1432 ();
 FILLCELL_X32 FILLER_432_1464 ();
 FILLCELL_X32 FILLER_432_1496 ();
 FILLCELL_X32 FILLER_432_1528 ();
 FILLCELL_X32 FILLER_432_1560 ();
 FILLCELL_X32 FILLER_432_1592 ();
 FILLCELL_X32 FILLER_432_1624 ();
 FILLCELL_X32 FILLER_432_1656 ();
 FILLCELL_X32 FILLER_432_1688 ();
 FILLCELL_X32 FILLER_432_1720 ();
 FILLCELL_X32 FILLER_432_1752 ();
 FILLCELL_X32 FILLER_432_1784 ();
 FILLCELL_X32 FILLER_432_1816 ();
 FILLCELL_X32 FILLER_432_1848 ();
 FILLCELL_X8 FILLER_432_1880 ();
 FILLCELL_X4 FILLER_432_1888 ();
 FILLCELL_X2 FILLER_432_1892 ();
 FILLCELL_X32 FILLER_432_1895 ();
 FILLCELL_X32 FILLER_432_1927 ();
 FILLCELL_X32 FILLER_432_1959 ();
 FILLCELL_X32 FILLER_432_1991 ();
 FILLCELL_X32 FILLER_432_2023 ();
 FILLCELL_X32 FILLER_432_2055 ();
 FILLCELL_X32 FILLER_432_2087 ();
 FILLCELL_X32 FILLER_432_2119 ();
 FILLCELL_X32 FILLER_432_2151 ();
 FILLCELL_X32 FILLER_432_2183 ();
 FILLCELL_X32 FILLER_432_2215 ();
 FILLCELL_X32 FILLER_432_2247 ();
 FILLCELL_X32 FILLER_432_2279 ();
 FILLCELL_X32 FILLER_432_2311 ();
 FILLCELL_X32 FILLER_432_2343 ();
 FILLCELL_X32 FILLER_432_2375 ();
 FILLCELL_X32 FILLER_432_2407 ();
 FILLCELL_X32 FILLER_432_2439 ();
 FILLCELL_X32 FILLER_432_2471 ();
 FILLCELL_X32 FILLER_432_2503 ();
 FILLCELL_X32 FILLER_432_2535 ();
 FILLCELL_X32 FILLER_432_2567 ();
 FILLCELL_X32 FILLER_432_2599 ();
 FILLCELL_X32 FILLER_432_2631 ();
 FILLCELL_X32 FILLER_432_2663 ();
 FILLCELL_X32 FILLER_432_2695 ();
 FILLCELL_X32 FILLER_432_2727 ();
 FILLCELL_X32 FILLER_432_2759 ();
 FILLCELL_X32 FILLER_432_2791 ();
 FILLCELL_X32 FILLER_432_2823 ();
 FILLCELL_X32 FILLER_432_2855 ();
 FILLCELL_X32 FILLER_432_2887 ();
 FILLCELL_X32 FILLER_432_2919 ();
 FILLCELL_X32 FILLER_432_2951 ();
 FILLCELL_X32 FILLER_432_2983 ();
 FILLCELL_X32 FILLER_432_3015 ();
 FILLCELL_X32 FILLER_432_3047 ();
 FILLCELL_X32 FILLER_432_3079 ();
 FILLCELL_X32 FILLER_432_3111 ();
 FILLCELL_X8 FILLER_432_3143 ();
 FILLCELL_X4 FILLER_432_3151 ();
 FILLCELL_X2 FILLER_432_3155 ();
 FILLCELL_X32 FILLER_432_3158 ();
 FILLCELL_X32 FILLER_432_3190 ();
 FILLCELL_X32 FILLER_432_3222 ();
 FILLCELL_X32 FILLER_432_3254 ();
 FILLCELL_X32 FILLER_432_3286 ();
 FILLCELL_X32 FILLER_432_3318 ();
 FILLCELL_X32 FILLER_432_3350 ();
 FILLCELL_X32 FILLER_432_3382 ();
 FILLCELL_X32 FILLER_432_3414 ();
 FILLCELL_X32 FILLER_432_3446 ();
 FILLCELL_X32 FILLER_432_3478 ();
 FILLCELL_X32 FILLER_432_3510 ();
 FILLCELL_X32 FILLER_432_3542 ();
 FILLCELL_X32 FILLER_432_3574 ();
 FILLCELL_X32 FILLER_432_3606 ();
 FILLCELL_X32 FILLER_432_3638 ();
 FILLCELL_X32 FILLER_432_3670 ();
 FILLCELL_X32 FILLER_432_3702 ();
 FILLCELL_X4 FILLER_432_3734 ();
 FILLCELL_X32 FILLER_433_1 ();
 FILLCELL_X32 FILLER_433_33 ();
 FILLCELL_X32 FILLER_433_65 ();
 FILLCELL_X32 FILLER_433_97 ();
 FILLCELL_X32 FILLER_433_129 ();
 FILLCELL_X32 FILLER_433_161 ();
 FILLCELL_X32 FILLER_433_193 ();
 FILLCELL_X32 FILLER_433_225 ();
 FILLCELL_X32 FILLER_433_257 ();
 FILLCELL_X32 FILLER_433_289 ();
 FILLCELL_X32 FILLER_433_321 ();
 FILLCELL_X32 FILLER_433_353 ();
 FILLCELL_X32 FILLER_433_385 ();
 FILLCELL_X32 FILLER_433_417 ();
 FILLCELL_X32 FILLER_433_449 ();
 FILLCELL_X32 FILLER_433_481 ();
 FILLCELL_X32 FILLER_433_513 ();
 FILLCELL_X32 FILLER_433_545 ();
 FILLCELL_X32 FILLER_433_577 ();
 FILLCELL_X32 FILLER_433_609 ();
 FILLCELL_X32 FILLER_433_641 ();
 FILLCELL_X32 FILLER_433_673 ();
 FILLCELL_X32 FILLER_433_705 ();
 FILLCELL_X32 FILLER_433_737 ();
 FILLCELL_X32 FILLER_433_769 ();
 FILLCELL_X32 FILLER_433_801 ();
 FILLCELL_X32 FILLER_433_833 ();
 FILLCELL_X32 FILLER_433_865 ();
 FILLCELL_X32 FILLER_433_897 ();
 FILLCELL_X32 FILLER_433_929 ();
 FILLCELL_X32 FILLER_433_961 ();
 FILLCELL_X32 FILLER_433_993 ();
 FILLCELL_X32 FILLER_433_1025 ();
 FILLCELL_X32 FILLER_433_1057 ();
 FILLCELL_X32 FILLER_433_1089 ();
 FILLCELL_X32 FILLER_433_1121 ();
 FILLCELL_X32 FILLER_433_1153 ();
 FILLCELL_X32 FILLER_433_1185 ();
 FILLCELL_X32 FILLER_433_1217 ();
 FILLCELL_X8 FILLER_433_1249 ();
 FILLCELL_X4 FILLER_433_1257 ();
 FILLCELL_X2 FILLER_433_1261 ();
 FILLCELL_X32 FILLER_433_1264 ();
 FILLCELL_X32 FILLER_433_1296 ();
 FILLCELL_X32 FILLER_433_1328 ();
 FILLCELL_X32 FILLER_433_1360 ();
 FILLCELL_X32 FILLER_433_1392 ();
 FILLCELL_X32 FILLER_433_1424 ();
 FILLCELL_X32 FILLER_433_1456 ();
 FILLCELL_X32 FILLER_433_1488 ();
 FILLCELL_X32 FILLER_433_1520 ();
 FILLCELL_X32 FILLER_433_1552 ();
 FILLCELL_X32 FILLER_433_1584 ();
 FILLCELL_X32 FILLER_433_1616 ();
 FILLCELL_X32 FILLER_433_1648 ();
 FILLCELL_X32 FILLER_433_1680 ();
 FILLCELL_X32 FILLER_433_1712 ();
 FILLCELL_X32 FILLER_433_1744 ();
 FILLCELL_X32 FILLER_433_1776 ();
 FILLCELL_X32 FILLER_433_1808 ();
 FILLCELL_X32 FILLER_433_1840 ();
 FILLCELL_X32 FILLER_433_1872 ();
 FILLCELL_X32 FILLER_433_1904 ();
 FILLCELL_X32 FILLER_433_1936 ();
 FILLCELL_X32 FILLER_433_1968 ();
 FILLCELL_X32 FILLER_433_2000 ();
 FILLCELL_X32 FILLER_433_2032 ();
 FILLCELL_X32 FILLER_433_2064 ();
 FILLCELL_X32 FILLER_433_2096 ();
 FILLCELL_X32 FILLER_433_2128 ();
 FILLCELL_X32 FILLER_433_2160 ();
 FILLCELL_X32 FILLER_433_2192 ();
 FILLCELL_X32 FILLER_433_2224 ();
 FILLCELL_X32 FILLER_433_2256 ();
 FILLCELL_X32 FILLER_433_2288 ();
 FILLCELL_X32 FILLER_433_2320 ();
 FILLCELL_X32 FILLER_433_2352 ();
 FILLCELL_X32 FILLER_433_2384 ();
 FILLCELL_X32 FILLER_433_2416 ();
 FILLCELL_X32 FILLER_433_2448 ();
 FILLCELL_X32 FILLER_433_2480 ();
 FILLCELL_X8 FILLER_433_2512 ();
 FILLCELL_X4 FILLER_433_2520 ();
 FILLCELL_X2 FILLER_433_2524 ();
 FILLCELL_X32 FILLER_433_2527 ();
 FILLCELL_X32 FILLER_433_2559 ();
 FILLCELL_X32 FILLER_433_2591 ();
 FILLCELL_X32 FILLER_433_2623 ();
 FILLCELL_X32 FILLER_433_2655 ();
 FILLCELL_X32 FILLER_433_2687 ();
 FILLCELL_X32 FILLER_433_2719 ();
 FILLCELL_X32 FILLER_433_2751 ();
 FILLCELL_X32 FILLER_433_2783 ();
 FILLCELL_X32 FILLER_433_2815 ();
 FILLCELL_X32 FILLER_433_2847 ();
 FILLCELL_X32 FILLER_433_2879 ();
 FILLCELL_X32 FILLER_433_2911 ();
 FILLCELL_X32 FILLER_433_2943 ();
 FILLCELL_X32 FILLER_433_2975 ();
 FILLCELL_X32 FILLER_433_3007 ();
 FILLCELL_X32 FILLER_433_3039 ();
 FILLCELL_X32 FILLER_433_3071 ();
 FILLCELL_X32 FILLER_433_3103 ();
 FILLCELL_X32 FILLER_433_3135 ();
 FILLCELL_X32 FILLER_433_3167 ();
 FILLCELL_X32 FILLER_433_3199 ();
 FILLCELL_X32 FILLER_433_3231 ();
 FILLCELL_X32 FILLER_433_3263 ();
 FILLCELL_X32 FILLER_433_3295 ();
 FILLCELL_X32 FILLER_433_3327 ();
 FILLCELL_X32 FILLER_433_3359 ();
 FILLCELL_X32 FILLER_433_3391 ();
 FILLCELL_X32 FILLER_433_3423 ();
 FILLCELL_X32 FILLER_433_3455 ();
 FILLCELL_X32 FILLER_433_3487 ();
 FILLCELL_X32 FILLER_433_3519 ();
 FILLCELL_X32 FILLER_433_3551 ();
 FILLCELL_X32 FILLER_433_3583 ();
 FILLCELL_X32 FILLER_433_3615 ();
 FILLCELL_X32 FILLER_433_3647 ();
 FILLCELL_X32 FILLER_433_3679 ();
 FILLCELL_X16 FILLER_433_3711 ();
 FILLCELL_X8 FILLER_433_3727 ();
 FILLCELL_X2 FILLER_433_3735 ();
 FILLCELL_X1 FILLER_433_3737 ();
 FILLCELL_X32 FILLER_434_1 ();
 FILLCELL_X32 FILLER_434_33 ();
 FILLCELL_X32 FILLER_434_65 ();
 FILLCELL_X32 FILLER_434_97 ();
 FILLCELL_X32 FILLER_434_129 ();
 FILLCELL_X32 FILLER_434_161 ();
 FILLCELL_X32 FILLER_434_193 ();
 FILLCELL_X32 FILLER_434_225 ();
 FILLCELL_X32 FILLER_434_257 ();
 FILLCELL_X32 FILLER_434_289 ();
 FILLCELL_X32 FILLER_434_321 ();
 FILLCELL_X32 FILLER_434_353 ();
 FILLCELL_X32 FILLER_434_385 ();
 FILLCELL_X32 FILLER_434_417 ();
 FILLCELL_X32 FILLER_434_449 ();
 FILLCELL_X32 FILLER_434_481 ();
 FILLCELL_X32 FILLER_434_513 ();
 FILLCELL_X32 FILLER_434_545 ();
 FILLCELL_X32 FILLER_434_577 ();
 FILLCELL_X16 FILLER_434_609 ();
 FILLCELL_X4 FILLER_434_625 ();
 FILLCELL_X2 FILLER_434_629 ();
 FILLCELL_X32 FILLER_434_632 ();
 FILLCELL_X32 FILLER_434_664 ();
 FILLCELL_X32 FILLER_434_696 ();
 FILLCELL_X32 FILLER_434_728 ();
 FILLCELL_X32 FILLER_434_760 ();
 FILLCELL_X32 FILLER_434_792 ();
 FILLCELL_X32 FILLER_434_824 ();
 FILLCELL_X32 FILLER_434_856 ();
 FILLCELL_X32 FILLER_434_888 ();
 FILLCELL_X32 FILLER_434_920 ();
 FILLCELL_X32 FILLER_434_952 ();
 FILLCELL_X32 FILLER_434_984 ();
 FILLCELL_X32 FILLER_434_1016 ();
 FILLCELL_X32 FILLER_434_1048 ();
 FILLCELL_X32 FILLER_434_1080 ();
 FILLCELL_X32 FILLER_434_1112 ();
 FILLCELL_X32 FILLER_434_1144 ();
 FILLCELL_X32 FILLER_434_1176 ();
 FILLCELL_X32 FILLER_434_1208 ();
 FILLCELL_X32 FILLER_434_1240 ();
 FILLCELL_X32 FILLER_434_1272 ();
 FILLCELL_X32 FILLER_434_1304 ();
 FILLCELL_X32 FILLER_434_1336 ();
 FILLCELL_X32 FILLER_434_1368 ();
 FILLCELL_X32 FILLER_434_1400 ();
 FILLCELL_X32 FILLER_434_1432 ();
 FILLCELL_X32 FILLER_434_1464 ();
 FILLCELL_X32 FILLER_434_1496 ();
 FILLCELL_X32 FILLER_434_1528 ();
 FILLCELL_X32 FILLER_434_1560 ();
 FILLCELL_X32 FILLER_434_1592 ();
 FILLCELL_X32 FILLER_434_1624 ();
 FILLCELL_X32 FILLER_434_1656 ();
 FILLCELL_X32 FILLER_434_1688 ();
 FILLCELL_X32 FILLER_434_1720 ();
 FILLCELL_X32 FILLER_434_1752 ();
 FILLCELL_X32 FILLER_434_1784 ();
 FILLCELL_X32 FILLER_434_1816 ();
 FILLCELL_X32 FILLER_434_1848 ();
 FILLCELL_X8 FILLER_434_1880 ();
 FILLCELL_X4 FILLER_434_1888 ();
 FILLCELL_X2 FILLER_434_1892 ();
 FILLCELL_X32 FILLER_434_1895 ();
 FILLCELL_X32 FILLER_434_1927 ();
 FILLCELL_X32 FILLER_434_1959 ();
 FILLCELL_X32 FILLER_434_1991 ();
 FILLCELL_X32 FILLER_434_2023 ();
 FILLCELL_X32 FILLER_434_2055 ();
 FILLCELL_X32 FILLER_434_2087 ();
 FILLCELL_X32 FILLER_434_2119 ();
 FILLCELL_X32 FILLER_434_2151 ();
 FILLCELL_X32 FILLER_434_2183 ();
 FILLCELL_X32 FILLER_434_2215 ();
 FILLCELL_X32 FILLER_434_2247 ();
 FILLCELL_X32 FILLER_434_2279 ();
 FILLCELL_X32 FILLER_434_2311 ();
 FILLCELL_X32 FILLER_434_2343 ();
 FILLCELL_X32 FILLER_434_2375 ();
 FILLCELL_X32 FILLER_434_2407 ();
 FILLCELL_X32 FILLER_434_2439 ();
 FILLCELL_X32 FILLER_434_2471 ();
 FILLCELL_X32 FILLER_434_2503 ();
 FILLCELL_X32 FILLER_434_2535 ();
 FILLCELL_X32 FILLER_434_2567 ();
 FILLCELL_X32 FILLER_434_2599 ();
 FILLCELL_X32 FILLER_434_2631 ();
 FILLCELL_X32 FILLER_434_2663 ();
 FILLCELL_X32 FILLER_434_2695 ();
 FILLCELL_X32 FILLER_434_2727 ();
 FILLCELL_X32 FILLER_434_2759 ();
 FILLCELL_X32 FILLER_434_2791 ();
 FILLCELL_X32 FILLER_434_2823 ();
 FILLCELL_X32 FILLER_434_2855 ();
 FILLCELL_X32 FILLER_434_2887 ();
 FILLCELL_X32 FILLER_434_2919 ();
 FILLCELL_X32 FILLER_434_2951 ();
 FILLCELL_X32 FILLER_434_2983 ();
 FILLCELL_X32 FILLER_434_3015 ();
 FILLCELL_X32 FILLER_434_3047 ();
 FILLCELL_X32 FILLER_434_3079 ();
 FILLCELL_X32 FILLER_434_3111 ();
 FILLCELL_X8 FILLER_434_3143 ();
 FILLCELL_X4 FILLER_434_3151 ();
 FILLCELL_X2 FILLER_434_3155 ();
 FILLCELL_X32 FILLER_434_3158 ();
 FILLCELL_X32 FILLER_434_3190 ();
 FILLCELL_X32 FILLER_434_3222 ();
 FILLCELL_X32 FILLER_434_3254 ();
 FILLCELL_X32 FILLER_434_3286 ();
 FILLCELL_X32 FILLER_434_3318 ();
 FILLCELL_X32 FILLER_434_3350 ();
 FILLCELL_X32 FILLER_434_3382 ();
 FILLCELL_X32 FILLER_434_3414 ();
 FILLCELL_X32 FILLER_434_3446 ();
 FILLCELL_X32 FILLER_434_3478 ();
 FILLCELL_X32 FILLER_434_3510 ();
 FILLCELL_X32 FILLER_434_3542 ();
 FILLCELL_X32 FILLER_434_3574 ();
 FILLCELL_X32 FILLER_434_3606 ();
 FILLCELL_X32 FILLER_434_3638 ();
 FILLCELL_X32 FILLER_434_3670 ();
 FILLCELL_X32 FILLER_434_3702 ();
 FILLCELL_X4 FILLER_434_3734 ();
 FILLCELL_X32 FILLER_435_1 ();
 FILLCELL_X32 FILLER_435_33 ();
 FILLCELL_X32 FILLER_435_65 ();
 FILLCELL_X32 FILLER_435_97 ();
 FILLCELL_X32 FILLER_435_129 ();
 FILLCELL_X32 FILLER_435_161 ();
 FILLCELL_X32 FILLER_435_193 ();
 FILLCELL_X32 FILLER_435_225 ();
 FILLCELL_X32 FILLER_435_257 ();
 FILLCELL_X32 FILLER_435_289 ();
 FILLCELL_X32 FILLER_435_321 ();
 FILLCELL_X32 FILLER_435_353 ();
 FILLCELL_X32 FILLER_435_385 ();
 FILLCELL_X32 FILLER_435_417 ();
 FILLCELL_X32 FILLER_435_449 ();
 FILLCELL_X32 FILLER_435_481 ();
 FILLCELL_X32 FILLER_435_513 ();
 FILLCELL_X32 FILLER_435_545 ();
 FILLCELL_X32 FILLER_435_577 ();
 FILLCELL_X32 FILLER_435_609 ();
 FILLCELL_X32 FILLER_435_641 ();
 FILLCELL_X32 FILLER_435_673 ();
 FILLCELL_X32 FILLER_435_705 ();
 FILLCELL_X32 FILLER_435_737 ();
 FILLCELL_X32 FILLER_435_769 ();
 FILLCELL_X32 FILLER_435_801 ();
 FILLCELL_X32 FILLER_435_833 ();
 FILLCELL_X32 FILLER_435_865 ();
 FILLCELL_X32 FILLER_435_897 ();
 FILLCELL_X32 FILLER_435_929 ();
 FILLCELL_X32 FILLER_435_961 ();
 FILLCELL_X32 FILLER_435_993 ();
 FILLCELL_X32 FILLER_435_1025 ();
 FILLCELL_X32 FILLER_435_1057 ();
 FILLCELL_X32 FILLER_435_1089 ();
 FILLCELL_X32 FILLER_435_1121 ();
 FILLCELL_X32 FILLER_435_1153 ();
 FILLCELL_X32 FILLER_435_1185 ();
 FILLCELL_X32 FILLER_435_1217 ();
 FILLCELL_X8 FILLER_435_1249 ();
 FILLCELL_X4 FILLER_435_1257 ();
 FILLCELL_X2 FILLER_435_1261 ();
 FILLCELL_X32 FILLER_435_1264 ();
 FILLCELL_X32 FILLER_435_1296 ();
 FILLCELL_X32 FILLER_435_1328 ();
 FILLCELL_X32 FILLER_435_1360 ();
 FILLCELL_X32 FILLER_435_1392 ();
 FILLCELL_X32 FILLER_435_1424 ();
 FILLCELL_X32 FILLER_435_1456 ();
 FILLCELL_X32 FILLER_435_1488 ();
 FILLCELL_X32 FILLER_435_1520 ();
 FILLCELL_X32 FILLER_435_1552 ();
 FILLCELL_X32 FILLER_435_1584 ();
 FILLCELL_X32 FILLER_435_1616 ();
 FILLCELL_X32 FILLER_435_1648 ();
 FILLCELL_X32 FILLER_435_1680 ();
 FILLCELL_X32 FILLER_435_1712 ();
 FILLCELL_X32 FILLER_435_1744 ();
 FILLCELL_X32 FILLER_435_1776 ();
 FILLCELL_X32 FILLER_435_1808 ();
 FILLCELL_X32 FILLER_435_1840 ();
 FILLCELL_X32 FILLER_435_1872 ();
 FILLCELL_X32 FILLER_435_1904 ();
 FILLCELL_X32 FILLER_435_1936 ();
 FILLCELL_X32 FILLER_435_1968 ();
 FILLCELL_X32 FILLER_435_2000 ();
 FILLCELL_X32 FILLER_435_2032 ();
 FILLCELL_X32 FILLER_435_2064 ();
 FILLCELL_X32 FILLER_435_2096 ();
 FILLCELL_X32 FILLER_435_2128 ();
 FILLCELL_X32 FILLER_435_2160 ();
 FILLCELL_X32 FILLER_435_2192 ();
 FILLCELL_X32 FILLER_435_2224 ();
 FILLCELL_X32 FILLER_435_2256 ();
 FILLCELL_X32 FILLER_435_2288 ();
 FILLCELL_X32 FILLER_435_2320 ();
 FILLCELL_X32 FILLER_435_2352 ();
 FILLCELL_X32 FILLER_435_2384 ();
 FILLCELL_X32 FILLER_435_2416 ();
 FILLCELL_X32 FILLER_435_2448 ();
 FILLCELL_X32 FILLER_435_2480 ();
 FILLCELL_X8 FILLER_435_2512 ();
 FILLCELL_X4 FILLER_435_2520 ();
 FILLCELL_X2 FILLER_435_2524 ();
 FILLCELL_X32 FILLER_435_2527 ();
 FILLCELL_X32 FILLER_435_2559 ();
 FILLCELL_X32 FILLER_435_2591 ();
 FILLCELL_X32 FILLER_435_2623 ();
 FILLCELL_X32 FILLER_435_2655 ();
 FILLCELL_X32 FILLER_435_2687 ();
 FILLCELL_X32 FILLER_435_2719 ();
 FILLCELL_X32 FILLER_435_2751 ();
 FILLCELL_X32 FILLER_435_2783 ();
 FILLCELL_X32 FILLER_435_2815 ();
 FILLCELL_X32 FILLER_435_2847 ();
 FILLCELL_X32 FILLER_435_2879 ();
 FILLCELL_X32 FILLER_435_2911 ();
 FILLCELL_X32 FILLER_435_2943 ();
 FILLCELL_X32 FILLER_435_2975 ();
 FILLCELL_X32 FILLER_435_3007 ();
 FILLCELL_X32 FILLER_435_3039 ();
 FILLCELL_X32 FILLER_435_3071 ();
 FILLCELL_X32 FILLER_435_3103 ();
 FILLCELL_X32 FILLER_435_3135 ();
 FILLCELL_X32 FILLER_435_3167 ();
 FILLCELL_X32 FILLER_435_3199 ();
 FILLCELL_X32 FILLER_435_3231 ();
 FILLCELL_X32 FILLER_435_3263 ();
 FILLCELL_X32 FILLER_435_3295 ();
 FILLCELL_X32 FILLER_435_3327 ();
 FILLCELL_X32 FILLER_435_3359 ();
 FILLCELL_X32 FILLER_435_3391 ();
 FILLCELL_X32 FILLER_435_3423 ();
 FILLCELL_X32 FILLER_435_3455 ();
 FILLCELL_X32 FILLER_435_3487 ();
 FILLCELL_X32 FILLER_435_3519 ();
 FILLCELL_X32 FILLER_435_3551 ();
 FILLCELL_X32 FILLER_435_3583 ();
 FILLCELL_X32 FILLER_435_3615 ();
 FILLCELL_X32 FILLER_435_3647 ();
 FILLCELL_X32 FILLER_435_3679 ();
 FILLCELL_X16 FILLER_435_3711 ();
 FILLCELL_X8 FILLER_435_3727 ();
 FILLCELL_X2 FILLER_435_3735 ();
 FILLCELL_X1 FILLER_435_3737 ();
 FILLCELL_X32 FILLER_436_1 ();
 FILLCELL_X32 FILLER_436_33 ();
 FILLCELL_X32 FILLER_436_65 ();
 FILLCELL_X32 FILLER_436_97 ();
 FILLCELL_X32 FILLER_436_129 ();
 FILLCELL_X32 FILLER_436_161 ();
 FILLCELL_X32 FILLER_436_193 ();
 FILLCELL_X32 FILLER_436_225 ();
 FILLCELL_X32 FILLER_436_257 ();
 FILLCELL_X32 FILLER_436_289 ();
 FILLCELL_X32 FILLER_436_321 ();
 FILLCELL_X32 FILLER_436_353 ();
 FILLCELL_X32 FILLER_436_385 ();
 FILLCELL_X32 FILLER_436_417 ();
 FILLCELL_X32 FILLER_436_449 ();
 FILLCELL_X32 FILLER_436_481 ();
 FILLCELL_X32 FILLER_436_513 ();
 FILLCELL_X32 FILLER_436_545 ();
 FILLCELL_X32 FILLER_436_577 ();
 FILLCELL_X16 FILLER_436_609 ();
 FILLCELL_X4 FILLER_436_625 ();
 FILLCELL_X2 FILLER_436_629 ();
 FILLCELL_X32 FILLER_436_632 ();
 FILLCELL_X32 FILLER_436_664 ();
 FILLCELL_X32 FILLER_436_696 ();
 FILLCELL_X32 FILLER_436_728 ();
 FILLCELL_X32 FILLER_436_760 ();
 FILLCELL_X32 FILLER_436_792 ();
 FILLCELL_X32 FILLER_436_824 ();
 FILLCELL_X32 FILLER_436_856 ();
 FILLCELL_X32 FILLER_436_888 ();
 FILLCELL_X32 FILLER_436_920 ();
 FILLCELL_X32 FILLER_436_952 ();
 FILLCELL_X32 FILLER_436_984 ();
 FILLCELL_X32 FILLER_436_1016 ();
 FILLCELL_X32 FILLER_436_1048 ();
 FILLCELL_X32 FILLER_436_1080 ();
 FILLCELL_X32 FILLER_436_1112 ();
 FILLCELL_X32 FILLER_436_1144 ();
 FILLCELL_X32 FILLER_436_1176 ();
 FILLCELL_X32 FILLER_436_1208 ();
 FILLCELL_X32 FILLER_436_1240 ();
 FILLCELL_X32 FILLER_436_1272 ();
 FILLCELL_X32 FILLER_436_1304 ();
 FILLCELL_X32 FILLER_436_1336 ();
 FILLCELL_X32 FILLER_436_1368 ();
 FILLCELL_X32 FILLER_436_1400 ();
 FILLCELL_X32 FILLER_436_1432 ();
 FILLCELL_X32 FILLER_436_1464 ();
 FILLCELL_X32 FILLER_436_1496 ();
 FILLCELL_X32 FILLER_436_1528 ();
 FILLCELL_X32 FILLER_436_1560 ();
 FILLCELL_X32 FILLER_436_1592 ();
 FILLCELL_X32 FILLER_436_1624 ();
 FILLCELL_X32 FILLER_436_1656 ();
 FILLCELL_X32 FILLER_436_1688 ();
 FILLCELL_X32 FILLER_436_1720 ();
 FILLCELL_X32 FILLER_436_1752 ();
 FILLCELL_X32 FILLER_436_1784 ();
 FILLCELL_X32 FILLER_436_1816 ();
 FILLCELL_X32 FILLER_436_1848 ();
 FILLCELL_X8 FILLER_436_1880 ();
 FILLCELL_X4 FILLER_436_1888 ();
 FILLCELL_X2 FILLER_436_1892 ();
 FILLCELL_X32 FILLER_436_1895 ();
 FILLCELL_X32 FILLER_436_1927 ();
 FILLCELL_X32 FILLER_436_1959 ();
 FILLCELL_X32 FILLER_436_1991 ();
 FILLCELL_X32 FILLER_436_2023 ();
 FILLCELL_X32 FILLER_436_2055 ();
 FILLCELL_X32 FILLER_436_2087 ();
 FILLCELL_X32 FILLER_436_2119 ();
 FILLCELL_X32 FILLER_436_2151 ();
 FILLCELL_X32 FILLER_436_2183 ();
 FILLCELL_X32 FILLER_436_2215 ();
 FILLCELL_X32 FILLER_436_2247 ();
 FILLCELL_X32 FILLER_436_2279 ();
 FILLCELL_X32 FILLER_436_2311 ();
 FILLCELL_X32 FILLER_436_2343 ();
 FILLCELL_X32 FILLER_436_2375 ();
 FILLCELL_X32 FILLER_436_2407 ();
 FILLCELL_X32 FILLER_436_2439 ();
 FILLCELL_X32 FILLER_436_2471 ();
 FILLCELL_X32 FILLER_436_2503 ();
 FILLCELL_X32 FILLER_436_2535 ();
 FILLCELL_X32 FILLER_436_2567 ();
 FILLCELL_X32 FILLER_436_2599 ();
 FILLCELL_X32 FILLER_436_2631 ();
 FILLCELL_X32 FILLER_436_2663 ();
 FILLCELL_X32 FILLER_436_2695 ();
 FILLCELL_X32 FILLER_436_2727 ();
 FILLCELL_X32 FILLER_436_2759 ();
 FILLCELL_X32 FILLER_436_2791 ();
 FILLCELL_X32 FILLER_436_2823 ();
 FILLCELL_X32 FILLER_436_2855 ();
 FILLCELL_X32 FILLER_436_2887 ();
 FILLCELL_X32 FILLER_436_2919 ();
 FILLCELL_X32 FILLER_436_2951 ();
 FILLCELL_X32 FILLER_436_2983 ();
 FILLCELL_X32 FILLER_436_3015 ();
 FILLCELL_X32 FILLER_436_3047 ();
 FILLCELL_X32 FILLER_436_3079 ();
 FILLCELL_X32 FILLER_436_3111 ();
 FILLCELL_X8 FILLER_436_3143 ();
 FILLCELL_X4 FILLER_436_3151 ();
 FILLCELL_X2 FILLER_436_3155 ();
 FILLCELL_X32 FILLER_436_3158 ();
 FILLCELL_X32 FILLER_436_3190 ();
 FILLCELL_X32 FILLER_436_3222 ();
 FILLCELL_X32 FILLER_436_3254 ();
 FILLCELL_X32 FILLER_436_3286 ();
 FILLCELL_X32 FILLER_436_3318 ();
 FILLCELL_X32 FILLER_436_3350 ();
 FILLCELL_X32 FILLER_436_3382 ();
 FILLCELL_X32 FILLER_436_3414 ();
 FILLCELL_X32 FILLER_436_3446 ();
 FILLCELL_X32 FILLER_436_3478 ();
 FILLCELL_X32 FILLER_436_3510 ();
 FILLCELL_X32 FILLER_436_3542 ();
 FILLCELL_X32 FILLER_436_3574 ();
 FILLCELL_X32 FILLER_436_3606 ();
 FILLCELL_X32 FILLER_436_3638 ();
 FILLCELL_X32 FILLER_436_3670 ();
 FILLCELL_X32 FILLER_436_3702 ();
 FILLCELL_X4 FILLER_436_3734 ();
 FILLCELL_X32 FILLER_437_1 ();
 FILLCELL_X32 FILLER_437_33 ();
 FILLCELL_X32 FILLER_437_65 ();
 FILLCELL_X32 FILLER_437_97 ();
 FILLCELL_X32 FILLER_437_129 ();
 FILLCELL_X32 FILLER_437_161 ();
 FILLCELL_X32 FILLER_437_193 ();
 FILLCELL_X32 FILLER_437_225 ();
 FILLCELL_X32 FILLER_437_257 ();
 FILLCELL_X32 FILLER_437_289 ();
 FILLCELL_X32 FILLER_437_321 ();
 FILLCELL_X32 FILLER_437_353 ();
 FILLCELL_X32 FILLER_437_385 ();
 FILLCELL_X32 FILLER_437_417 ();
 FILLCELL_X32 FILLER_437_449 ();
 FILLCELL_X32 FILLER_437_481 ();
 FILLCELL_X32 FILLER_437_513 ();
 FILLCELL_X32 FILLER_437_545 ();
 FILLCELL_X32 FILLER_437_577 ();
 FILLCELL_X32 FILLER_437_609 ();
 FILLCELL_X32 FILLER_437_641 ();
 FILLCELL_X32 FILLER_437_673 ();
 FILLCELL_X32 FILLER_437_705 ();
 FILLCELL_X32 FILLER_437_737 ();
 FILLCELL_X32 FILLER_437_769 ();
 FILLCELL_X32 FILLER_437_801 ();
 FILLCELL_X32 FILLER_437_833 ();
 FILLCELL_X32 FILLER_437_865 ();
 FILLCELL_X32 FILLER_437_897 ();
 FILLCELL_X32 FILLER_437_929 ();
 FILLCELL_X32 FILLER_437_961 ();
 FILLCELL_X32 FILLER_437_993 ();
 FILLCELL_X32 FILLER_437_1025 ();
 FILLCELL_X32 FILLER_437_1057 ();
 FILLCELL_X32 FILLER_437_1089 ();
 FILLCELL_X32 FILLER_437_1121 ();
 FILLCELL_X32 FILLER_437_1153 ();
 FILLCELL_X32 FILLER_437_1185 ();
 FILLCELL_X32 FILLER_437_1217 ();
 FILLCELL_X8 FILLER_437_1249 ();
 FILLCELL_X4 FILLER_437_1257 ();
 FILLCELL_X2 FILLER_437_1261 ();
 FILLCELL_X32 FILLER_437_1264 ();
 FILLCELL_X32 FILLER_437_1296 ();
 FILLCELL_X32 FILLER_437_1328 ();
 FILLCELL_X32 FILLER_437_1360 ();
 FILLCELL_X32 FILLER_437_1392 ();
 FILLCELL_X32 FILLER_437_1424 ();
 FILLCELL_X32 FILLER_437_1456 ();
 FILLCELL_X32 FILLER_437_1488 ();
 FILLCELL_X32 FILLER_437_1520 ();
 FILLCELL_X32 FILLER_437_1552 ();
 FILLCELL_X32 FILLER_437_1584 ();
 FILLCELL_X32 FILLER_437_1616 ();
 FILLCELL_X32 FILLER_437_1648 ();
 FILLCELL_X32 FILLER_437_1680 ();
 FILLCELL_X32 FILLER_437_1712 ();
 FILLCELL_X32 FILLER_437_1744 ();
 FILLCELL_X32 FILLER_437_1776 ();
 FILLCELL_X32 FILLER_437_1808 ();
 FILLCELL_X32 FILLER_437_1840 ();
 FILLCELL_X32 FILLER_437_1872 ();
 FILLCELL_X32 FILLER_437_1904 ();
 FILLCELL_X32 FILLER_437_1936 ();
 FILLCELL_X32 FILLER_437_1968 ();
 FILLCELL_X32 FILLER_437_2000 ();
 FILLCELL_X32 FILLER_437_2032 ();
 FILLCELL_X32 FILLER_437_2064 ();
 FILLCELL_X32 FILLER_437_2096 ();
 FILLCELL_X32 FILLER_437_2128 ();
 FILLCELL_X32 FILLER_437_2160 ();
 FILLCELL_X32 FILLER_437_2192 ();
 FILLCELL_X32 FILLER_437_2224 ();
 FILLCELL_X32 FILLER_437_2256 ();
 FILLCELL_X32 FILLER_437_2288 ();
 FILLCELL_X32 FILLER_437_2320 ();
 FILLCELL_X32 FILLER_437_2352 ();
 FILLCELL_X32 FILLER_437_2384 ();
 FILLCELL_X32 FILLER_437_2416 ();
 FILLCELL_X32 FILLER_437_2448 ();
 FILLCELL_X32 FILLER_437_2480 ();
 FILLCELL_X8 FILLER_437_2512 ();
 FILLCELL_X4 FILLER_437_2520 ();
 FILLCELL_X2 FILLER_437_2524 ();
 FILLCELL_X32 FILLER_437_2527 ();
 FILLCELL_X32 FILLER_437_2559 ();
 FILLCELL_X32 FILLER_437_2591 ();
 FILLCELL_X32 FILLER_437_2623 ();
 FILLCELL_X32 FILLER_437_2655 ();
 FILLCELL_X32 FILLER_437_2687 ();
 FILLCELL_X32 FILLER_437_2719 ();
 FILLCELL_X32 FILLER_437_2751 ();
 FILLCELL_X32 FILLER_437_2783 ();
 FILLCELL_X32 FILLER_437_2815 ();
 FILLCELL_X32 FILLER_437_2847 ();
 FILLCELL_X32 FILLER_437_2879 ();
 FILLCELL_X32 FILLER_437_2911 ();
 FILLCELL_X32 FILLER_437_2943 ();
 FILLCELL_X32 FILLER_437_2975 ();
 FILLCELL_X32 FILLER_437_3007 ();
 FILLCELL_X32 FILLER_437_3039 ();
 FILLCELL_X32 FILLER_437_3071 ();
 FILLCELL_X32 FILLER_437_3103 ();
 FILLCELL_X32 FILLER_437_3135 ();
 FILLCELL_X32 FILLER_437_3167 ();
 FILLCELL_X32 FILLER_437_3199 ();
 FILLCELL_X32 FILLER_437_3231 ();
 FILLCELL_X32 FILLER_437_3263 ();
 FILLCELL_X32 FILLER_437_3295 ();
 FILLCELL_X32 FILLER_437_3327 ();
 FILLCELL_X32 FILLER_437_3359 ();
 FILLCELL_X32 FILLER_437_3391 ();
 FILLCELL_X32 FILLER_437_3423 ();
 FILLCELL_X32 FILLER_437_3455 ();
 FILLCELL_X32 FILLER_437_3487 ();
 FILLCELL_X32 FILLER_437_3519 ();
 FILLCELL_X32 FILLER_437_3551 ();
 FILLCELL_X32 FILLER_437_3583 ();
 FILLCELL_X32 FILLER_437_3615 ();
 FILLCELL_X32 FILLER_437_3647 ();
 FILLCELL_X32 FILLER_437_3679 ();
 FILLCELL_X16 FILLER_437_3711 ();
 FILLCELL_X8 FILLER_437_3727 ();
 FILLCELL_X2 FILLER_437_3735 ();
 FILLCELL_X1 FILLER_437_3737 ();
 FILLCELL_X32 FILLER_438_1 ();
 FILLCELL_X32 FILLER_438_33 ();
 FILLCELL_X32 FILLER_438_65 ();
 FILLCELL_X32 FILLER_438_97 ();
 FILLCELL_X32 FILLER_438_129 ();
 FILLCELL_X32 FILLER_438_161 ();
 FILLCELL_X32 FILLER_438_193 ();
 FILLCELL_X32 FILLER_438_225 ();
 FILLCELL_X32 FILLER_438_257 ();
 FILLCELL_X32 FILLER_438_289 ();
 FILLCELL_X32 FILLER_438_321 ();
 FILLCELL_X32 FILLER_438_353 ();
 FILLCELL_X32 FILLER_438_385 ();
 FILLCELL_X32 FILLER_438_417 ();
 FILLCELL_X32 FILLER_438_449 ();
 FILLCELL_X32 FILLER_438_481 ();
 FILLCELL_X32 FILLER_438_513 ();
 FILLCELL_X32 FILLER_438_545 ();
 FILLCELL_X32 FILLER_438_577 ();
 FILLCELL_X16 FILLER_438_609 ();
 FILLCELL_X4 FILLER_438_625 ();
 FILLCELL_X2 FILLER_438_629 ();
 FILLCELL_X32 FILLER_438_632 ();
 FILLCELL_X32 FILLER_438_664 ();
 FILLCELL_X32 FILLER_438_696 ();
 FILLCELL_X32 FILLER_438_728 ();
 FILLCELL_X32 FILLER_438_760 ();
 FILLCELL_X32 FILLER_438_792 ();
 FILLCELL_X32 FILLER_438_824 ();
 FILLCELL_X32 FILLER_438_856 ();
 FILLCELL_X32 FILLER_438_888 ();
 FILLCELL_X32 FILLER_438_920 ();
 FILLCELL_X32 FILLER_438_952 ();
 FILLCELL_X32 FILLER_438_984 ();
 FILLCELL_X32 FILLER_438_1016 ();
 FILLCELL_X32 FILLER_438_1048 ();
 FILLCELL_X32 FILLER_438_1080 ();
 FILLCELL_X32 FILLER_438_1112 ();
 FILLCELL_X32 FILLER_438_1144 ();
 FILLCELL_X32 FILLER_438_1176 ();
 FILLCELL_X32 FILLER_438_1208 ();
 FILLCELL_X32 FILLER_438_1240 ();
 FILLCELL_X32 FILLER_438_1272 ();
 FILLCELL_X32 FILLER_438_1304 ();
 FILLCELL_X32 FILLER_438_1336 ();
 FILLCELL_X32 FILLER_438_1368 ();
 FILLCELL_X32 FILLER_438_1400 ();
 FILLCELL_X32 FILLER_438_1432 ();
 FILLCELL_X32 FILLER_438_1464 ();
 FILLCELL_X32 FILLER_438_1496 ();
 FILLCELL_X32 FILLER_438_1528 ();
 FILLCELL_X32 FILLER_438_1560 ();
 FILLCELL_X32 FILLER_438_1592 ();
 FILLCELL_X32 FILLER_438_1624 ();
 FILLCELL_X32 FILLER_438_1656 ();
 FILLCELL_X32 FILLER_438_1688 ();
 FILLCELL_X32 FILLER_438_1720 ();
 FILLCELL_X32 FILLER_438_1752 ();
 FILLCELL_X32 FILLER_438_1784 ();
 FILLCELL_X32 FILLER_438_1816 ();
 FILLCELL_X32 FILLER_438_1848 ();
 FILLCELL_X8 FILLER_438_1880 ();
 FILLCELL_X4 FILLER_438_1888 ();
 FILLCELL_X2 FILLER_438_1892 ();
 FILLCELL_X32 FILLER_438_1895 ();
 FILLCELL_X32 FILLER_438_1927 ();
 FILLCELL_X32 FILLER_438_1959 ();
 FILLCELL_X32 FILLER_438_1991 ();
 FILLCELL_X32 FILLER_438_2023 ();
 FILLCELL_X32 FILLER_438_2055 ();
 FILLCELL_X32 FILLER_438_2087 ();
 FILLCELL_X32 FILLER_438_2119 ();
 FILLCELL_X32 FILLER_438_2151 ();
 FILLCELL_X32 FILLER_438_2183 ();
 FILLCELL_X32 FILLER_438_2215 ();
 FILLCELL_X32 FILLER_438_2247 ();
 FILLCELL_X32 FILLER_438_2279 ();
 FILLCELL_X32 FILLER_438_2311 ();
 FILLCELL_X32 FILLER_438_2343 ();
 FILLCELL_X32 FILLER_438_2375 ();
 FILLCELL_X32 FILLER_438_2407 ();
 FILLCELL_X32 FILLER_438_2439 ();
 FILLCELL_X32 FILLER_438_2471 ();
 FILLCELL_X32 FILLER_438_2503 ();
 FILLCELL_X32 FILLER_438_2535 ();
 FILLCELL_X32 FILLER_438_2567 ();
 FILLCELL_X32 FILLER_438_2599 ();
 FILLCELL_X32 FILLER_438_2631 ();
 FILLCELL_X32 FILLER_438_2663 ();
 FILLCELL_X32 FILLER_438_2695 ();
 FILLCELL_X32 FILLER_438_2727 ();
 FILLCELL_X32 FILLER_438_2759 ();
 FILLCELL_X32 FILLER_438_2791 ();
 FILLCELL_X32 FILLER_438_2823 ();
 FILLCELL_X32 FILLER_438_2855 ();
 FILLCELL_X32 FILLER_438_2887 ();
 FILLCELL_X32 FILLER_438_2919 ();
 FILLCELL_X32 FILLER_438_2951 ();
 FILLCELL_X32 FILLER_438_2983 ();
 FILLCELL_X32 FILLER_438_3015 ();
 FILLCELL_X32 FILLER_438_3047 ();
 FILLCELL_X32 FILLER_438_3079 ();
 FILLCELL_X32 FILLER_438_3111 ();
 FILLCELL_X8 FILLER_438_3143 ();
 FILLCELL_X4 FILLER_438_3151 ();
 FILLCELL_X2 FILLER_438_3155 ();
 FILLCELL_X32 FILLER_438_3158 ();
 FILLCELL_X32 FILLER_438_3190 ();
 FILLCELL_X32 FILLER_438_3222 ();
 FILLCELL_X32 FILLER_438_3254 ();
 FILLCELL_X32 FILLER_438_3286 ();
 FILLCELL_X32 FILLER_438_3318 ();
 FILLCELL_X32 FILLER_438_3350 ();
 FILLCELL_X32 FILLER_438_3382 ();
 FILLCELL_X32 FILLER_438_3414 ();
 FILLCELL_X32 FILLER_438_3446 ();
 FILLCELL_X32 FILLER_438_3478 ();
 FILLCELL_X32 FILLER_438_3510 ();
 FILLCELL_X32 FILLER_438_3542 ();
 FILLCELL_X32 FILLER_438_3574 ();
 FILLCELL_X32 FILLER_438_3606 ();
 FILLCELL_X32 FILLER_438_3638 ();
 FILLCELL_X32 FILLER_438_3670 ();
 FILLCELL_X32 FILLER_438_3702 ();
 FILLCELL_X4 FILLER_438_3734 ();
 FILLCELL_X32 FILLER_439_1 ();
 FILLCELL_X32 FILLER_439_33 ();
 FILLCELL_X32 FILLER_439_65 ();
 FILLCELL_X32 FILLER_439_97 ();
 FILLCELL_X32 FILLER_439_129 ();
 FILLCELL_X32 FILLER_439_161 ();
 FILLCELL_X32 FILLER_439_193 ();
 FILLCELL_X32 FILLER_439_225 ();
 FILLCELL_X32 FILLER_439_257 ();
 FILLCELL_X32 FILLER_439_289 ();
 FILLCELL_X32 FILLER_439_321 ();
 FILLCELL_X32 FILLER_439_353 ();
 FILLCELL_X32 FILLER_439_385 ();
 FILLCELL_X32 FILLER_439_417 ();
 FILLCELL_X32 FILLER_439_449 ();
 FILLCELL_X32 FILLER_439_481 ();
 FILLCELL_X32 FILLER_439_513 ();
 FILLCELL_X32 FILLER_439_545 ();
 FILLCELL_X32 FILLER_439_577 ();
 FILLCELL_X32 FILLER_439_609 ();
 FILLCELL_X32 FILLER_439_641 ();
 FILLCELL_X32 FILLER_439_673 ();
 FILLCELL_X32 FILLER_439_705 ();
 FILLCELL_X32 FILLER_439_737 ();
 FILLCELL_X32 FILLER_439_769 ();
 FILLCELL_X32 FILLER_439_801 ();
 FILLCELL_X32 FILLER_439_833 ();
 FILLCELL_X32 FILLER_439_865 ();
 FILLCELL_X32 FILLER_439_897 ();
 FILLCELL_X32 FILLER_439_929 ();
 FILLCELL_X32 FILLER_439_961 ();
 FILLCELL_X32 FILLER_439_993 ();
 FILLCELL_X32 FILLER_439_1025 ();
 FILLCELL_X32 FILLER_439_1057 ();
 FILLCELL_X32 FILLER_439_1089 ();
 FILLCELL_X32 FILLER_439_1121 ();
 FILLCELL_X32 FILLER_439_1153 ();
 FILLCELL_X32 FILLER_439_1185 ();
 FILLCELL_X32 FILLER_439_1217 ();
 FILLCELL_X8 FILLER_439_1249 ();
 FILLCELL_X4 FILLER_439_1257 ();
 FILLCELL_X2 FILLER_439_1261 ();
 FILLCELL_X32 FILLER_439_1264 ();
 FILLCELL_X32 FILLER_439_1296 ();
 FILLCELL_X32 FILLER_439_1328 ();
 FILLCELL_X32 FILLER_439_1360 ();
 FILLCELL_X32 FILLER_439_1392 ();
 FILLCELL_X32 FILLER_439_1424 ();
 FILLCELL_X32 FILLER_439_1456 ();
 FILLCELL_X32 FILLER_439_1488 ();
 FILLCELL_X32 FILLER_439_1520 ();
 FILLCELL_X32 FILLER_439_1552 ();
 FILLCELL_X32 FILLER_439_1584 ();
 FILLCELL_X32 FILLER_439_1616 ();
 FILLCELL_X32 FILLER_439_1648 ();
 FILLCELL_X32 FILLER_439_1680 ();
 FILLCELL_X32 FILLER_439_1712 ();
 FILLCELL_X32 FILLER_439_1744 ();
 FILLCELL_X32 FILLER_439_1776 ();
 FILLCELL_X32 FILLER_439_1808 ();
 FILLCELL_X32 FILLER_439_1840 ();
 FILLCELL_X32 FILLER_439_1872 ();
 FILLCELL_X32 FILLER_439_1904 ();
 FILLCELL_X32 FILLER_439_1936 ();
 FILLCELL_X32 FILLER_439_1968 ();
 FILLCELL_X32 FILLER_439_2000 ();
 FILLCELL_X32 FILLER_439_2032 ();
 FILLCELL_X32 FILLER_439_2064 ();
 FILLCELL_X32 FILLER_439_2096 ();
 FILLCELL_X32 FILLER_439_2128 ();
 FILLCELL_X32 FILLER_439_2160 ();
 FILLCELL_X32 FILLER_439_2192 ();
 FILLCELL_X32 FILLER_439_2224 ();
 FILLCELL_X32 FILLER_439_2256 ();
 FILLCELL_X32 FILLER_439_2288 ();
 FILLCELL_X32 FILLER_439_2320 ();
 FILLCELL_X32 FILLER_439_2352 ();
 FILLCELL_X32 FILLER_439_2384 ();
 FILLCELL_X32 FILLER_439_2416 ();
 FILLCELL_X32 FILLER_439_2448 ();
 FILLCELL_X32 FILLER_439_2480 ();
 FILLCELL_X8 FILLER_439_2512 ();
 FILLCELL_X4 FILLER_439_2520 ();
 FILLCELL_X2 FILLER_439_2524 ();
 FILLCELL_X32 FILLER_439_2527 ();
 FILLCELL_X32 FILLER_439_2559 ();
 FILLCELL_X32 FILLER_439_2591 ();
 FILLCELL_X32 FILLER_439_2623 ();
 FILLCELL_X32 FILLER_439_2655 ();
 FILLCELL_X32 FILLER_439_2687 ();
 FILLCELL_X32 FILLER_439_2719 ();
 FILLCELL_X32 FILLER_439_2751 ();
 FILLCELL_X32 FILLER_439_2783 ();
 FILLCELL_X32 FILLER_439_2815 ();
 FILLCELL_X32 FILLER_439_2847 ();
 FILLCELL_X32 FILLER_439_2879 ();
 FILLCELL_X32 FILLER_439_2911 ();
 FILLCELL_X32 FILLER_439_2943 ();
 FILLCELL_X32 FILLER_439_2975 ();
 FILLCELL_X32 FILLER_439_3007 ();
 FILLCELL_X32 FILLER_439_3039 ();
 FILLCELL_X32 FILLER_439_3071 ();
 FILLCELL_X32 FILLER_439_3103 ();
 FILLCELL_X32 FILLER_439_3135 ();
 FILLCELL_X32 FILLER_439_3167 ();
 FILLCELL_X32 FILLER_439_3199 ();
 FILLCELL_X32 FILLER_439_3231 ();
 FILLCELL_X32 FILLER_439_3263 ();
 FILLCELL_X32 FILLER_439_3295 ();
 FILLCELL_X32 FILLER_439_3327 ();
 FILLCELL_X32 FILLER_439_3359 ();
 FILLCELL_X32 FILLER_439_3391 ();
 FILLCELL_X32 FILLER_439_3423 ();
 FILLCELL_X32 FILLER_439_3455 ();
 FILLCELL_X32 FILLER_439_3487 ();
 FILLCELL_X32 FILLER_439_3519 ();
 FILLCELL_X32 FILLER_439_3551 ();
 FILLCELL_X32 FILLER_439_3583 ();
 FILLCELL_X32 FILLER_439_3615 ();
 FILLCELL_X32 FILLER_439_3647 ();
 FILLCELL_X32 FILLER_439_3679 ();
 FILLCELL_X16 FILLER_439_3711 ();
 FILLCELL_X8 FILLER_439_3727 ();
 FILLCELL_X2 FILLER_439_3735 ();
 FILLCELL_X1 FILLER_439_3737 ();
 FILLCELL_X32 FILLER_440_1 ();
 FILLCELL_X32 FILLER_440_33 ();
 FILLCELL_X32 FILLER_440_65 ();
 FILLCELL_X32 FILLER_440_97 ();
 FILLCELL_X32 FILLER_440_129 ();
 FILLCELL_X32 FILLER_440_161 ();
 FILLCELL_X32 FILLER_440_193 ();
 FILLCELL_X32 FILLER_440_225 ();
 FILLCELL_X32 FILLER_440_257 ();
 FILLCELL_X32 FILLER_440_289 ();
 FILLCELL_X32 FILLER_440_321 ();
 FILLCELL_X32 FILLER_440_353 ();
 FILLCELL_X32 FILLER_440_385 ();
 FILLCELL_X32 FILLER_440_417 ();
 FILLCELL_X32 FILLER_440_449 ();
 FILLCELL_X32 FILLER_440_481 ();
 FILLCELL_X32 FILLER_440_513 ();
 FILLCELL_X32 FILLER_440_545 ();
 FILLCELL_X32 FILLER_440_577 ();
 FILLCELL_X16 FILLER_440_609 ();
 FILLCELL_X4 FILLER_440_625 ();
 FILLCELL_X2 FILLER_440_629 ();
 FILLCELL_X32 FILLER_440_632 ();
 FILLCELL_X32 FILLER_440_664 ();
 FILLCELL_X32 FILLER_440_696 ();
 FILLCELL_X32 FILLER_440_728 ();
 FILLCELL_X32 FILLER_440_760 ();
 FILLCELL_X32 FILLER_440_792 ();
 FILLCELL_X32 FILLER_440_824 ();
 FILLCELL_X32 FILLER_440_856 ();
 FILLCELL_X32 FILLER_440_888 ();
 FILLCELL_X32 FILLER_440_920 ();
 FILLCELL_X32 FILLER_440_952 ();
 FILLCELL_X32 FILLER_440_984 ();
 FILLCELL_X32 FILLER_440_1016 ();
 FILLCELL_X32 FILLER_440_1048 ();
 FILLCELL_X32 FILLER_440_1080 ();
 FILLCELL_X32 FILLER_440_1112 ();
 FILLCELL_X32 FILLER_440_1144 ();
 FILLCELL_X32 FILLER_440_1176 ();
 FILLCELL_X32 FILLER_440_1208 ();
 FILLCELL_X32 FILLER_440_1240 ();
 FILLCELL_X32 FILLER_440_1272 ();
 FILLCELL_X32 FILLER_440_1304 ();
 FILLCELL_X32 FILLER_440_1336 ();
 FILLCELL_X32 FILLER_440_1368 ();
 FILLCELL_X32 FILLER_440_1400 ();
 FILLCELL_X32 FILLER_440_1432 ();
 FILLCELL_X32 FILLER_440_1464 ();
 FILLCELL_X32 FILLER_440_1496 ();
 FILLCELL_X32 FILLER_440_1528 ();
 FILLCELL_X32 FILLER_440_1560 ();
 FILLCELL_X32 FILLER_440_1592 ();
 FILLCELL_X32 FILLER_440_1624 ();
 FILLCELL_X32 FILLER_440_1656 ();
 FILLCELL_X32 FILLER_440_1688 ();
 FILLCELL_X32 FILLER_440_1720 ();
 FILLCELL_X32 FILLER_440_1752 ();
 FILLCELL_X32 FILLER_440_1784 ();
 FILLCELL_X32 FILLER_440_1816 ();
 FILLCELL_X32 FILLER_440_1848 ();
 FILLCELL_X8 FILLER_440_1880 ();
 FILLCELL_X4 FILLER_440_1888 ();
 FILLCELL_X2 FILLER_440_1892 ();
 FILLCELL_X32 FILLER_440_1895 ();
 FILLCELL_X32 FILLER_440_1927 ();
 FILLCELL_X32 FILLER_440_1959 ();
 FILLCELL_X32 FILLER_440_1991 ();
 FILLCELL_X32 FILLER_440_2023 ();
 FILLCELL_X32 FILLER_440_2055 ();
 FILLCELL_X32 FILLER_440_2087 ();
 FILLCELL_X32 FILLER_440_2119 ();
 FILLCELL_X32 FILLER_440_2151 ();
 FILLCELL_X32 FILLER_440_2183 ();
 FILLCELL_X32 FILLER_440_2215 ();
 FILLCELL_X32 FILLER_440_2247 ();
 FILLCELL_X32 FILLER_440_2279 ();
 FILLCELL_X32 FILLER_440_2311 ();
 FILLCELL_X32 FILLER_440_2343 ();
 FILLCELL_X32 FILLER_440_2375 ();
 FILLCELL_X32 FILLER_440_2407 ();
 FILLCELL_X32 FILLER_440_2439 ();
 FILLCELL_X32 FILLER_440_2471 ();
 FILLCELL_X32 FILLER_440_2503 ();
 FILLCELL_X32 FILLER_440_2535 ();
 FILLCELL_X32 FILLER_440_2567 ();
 FILLCELL_X32 FILLER_440_2599 ();
 FILLCELL_X32 FILLER_440_2631 ();
 FILLCELL_X32 FILLER_440_2663 ();
 FILLCELL_X32 FILLER_440_2695 ();
 FILLCELL_X32 FILLER_440_2727 ();
 FILLCELL_X32 FILLER_440_2759 ();
 FILLCELL_X32 FILLER_440_2791 ();
 FILLCELL_X32 FILLER_440_2823 ();
 FILLCELL_X32 FILLER_440_2855 ();
 FILLCELL_X32 FILLER_440_2887 ();
 FILLCELL_X32 FILLER_440_2919 ();
 FILLCELL_X32 FILLER_440_2951 ();
 FILLCELL_X32 FILLER_440_2983 ();
 FILLCELL_X32 FILLER_440_3015 ();
 FILLCELL_X32 FILLER_440_3047 ();
 FILLCELL_X32 FILLER_440_3079 ();
 FILLCELL_X32 FILLER_440_3111 ();
 FILLCELL_X8 FILLER_440_3143 ();
 FILLCELL_X4 FILLER_440_3151 ();
 FILLCELL_X2 FILLER_440_3155 ();
 FILLCELL_X32 FILLER_440_3158 ();
 FILLCELL_X32 FILLER_440_3190 ();
 FILLCELL_X32 FILLER_440_3222 ();
 FILLCELL_X32 FILLER_440_3254 ();
 FILLCELL_X32 FILLER_440_3286 ();
 FILLCELL_X32 FILLER_440_3318 ();
 FILLCELL_X32 FILLER_440_3350 ();
 FILLCELL_X32 FILLER_440_3382 ();
 FILLCELL_X32 FILLER_440_3414 ();
 FILLCELL_X32 FILLER_440_3446 ();
 FILLCELL_X32 FILLER_440_3478 ();
 FILLCELL_X32 FILLER_440_3510 ();
 FILLCELL_X32 FILLER_440_3542 ();
 FILLCELL_X32 FILLER_440_3574 ();
 FILLCELL_X32 FILLER_440_3606 ();
 FILLCELL_X32 FILLER_440_3638 ();
 FILLCELL_X32 FILLER_440_3670 ();
 FILLCELL_X32 FILLER_440_3702 ();
 FILLCELL_X4 FILLER_440_3734 ();
 FILLCELL_X32 FILLER_441_1 ();
 FILLCELL_X32 FILLER_441_33 ();
 FILLCELL_X32 FILLER_441_65 ();
 FILLCELL_X32 FILLER_441_97 ();
 FILLCELL_X32 FILLER_441_129 ();
 FILLCELL_X32 FILLER_441_161 ();
 FILLCELL_X32 FILLER_441_193 ();
 FILLCELL_X32 FILLER_441_225 ();
 FILLCELL_X32 FILLER_441_257 ();
 FILLCELL_X32 FILLER_441_289 ();
 FILLCELL_X32 FILLER_441_321 ();
 FILLCELL_X32 FILLER_441_353 ();
 FILLCELL_X32 FILLER_441_385 ();
 FILLCELL_X32 FILLER_441_417 ();
 FILLCELL_X32 FILLER_441_449 ();
 FILLCELL_X32 FILLER_441_481 ();
 FILLCELL_X32 FILLER_441_513 ();
 FILLCELL_X32 FILLER_441_545 ();
 FILLCELL_X32 FILLER_441_577 ();
 FILLCELL_X32 FILLER_441_609 ();
 FILLCELL_X32 FILLER_441_641 ();
 FILLCELL_X32 FILLER_441_673 ();
 FILLCELL_X32 FILLER_441_705 ();
 FILLCELL_X32 FILLER_441_737 ();
 FILLCELL_X32 FILLER_441_769 ();
 FILLCELL_X32 FILLER_441_801 ();
 FILLCELL_X32 FILLER_441_833 ();
 FILLCELL_X32 FILLER_441_865 ();
 FILLCELL_X32 FILLER_441_897 ();
 FILLCELL_X32 FILLER_441_929 ();
 FILLCELL_X32 FILLER_441_961 ();
 FILLCELL_X32 FILLER_441_993 ();
 FILLCELL_X32 FILLER_441_1025 ();
 FILLCELL_X32 FILLER_441_1057 ();
 FILLCELL_X32 FILLER_441_1089 ();
 FILLCELL_X32 FILLER_441_1121 ();
 FILLCELL_X32 FILLER_441_1153 ();
 FILLCELL_X32 FILLER_441_1185 ();
 FILLCELL_X32 FILLER_441_1217 ();
 FILLCELL_X8 FILLER_441_1249 ();
 FILLCELL_X4 FILLER_441_1257 ();
 FILLCELL_X2 FILLER_441_1261 ();
 FILLCELL_X32 FILLER_441_1264 ();
 FILLCELL_X32 FILLER_441_1296 ();
 FILLCELL_X32 FILLER_441_1328 ();
 FILLCELL_X32 FILLER_441_1360 ();
 FILLCELL_X32 FILLER_441_1392 ();
 FILLCELL_X32 FILLER_441_1424 ();
 FILLCELL_X32 FILLER_441_1456 ();
 FILLCELL_X32 FILLER_441_1488 ();
 FILLCELL_X32 FILLER_441_1520 ();
 FILLCELL_X32 FILLER_441_1552 ();
 FILLCELL_X32 FILLER_441_1584 ();
 FILLCELL_X32 FILLER_441_1616 ();
 FILLCELL_X32 FILLER_441_1648 ();
 FILLCELL_X32 FILLER_441_1680 ();
 FILLCELL_X32 FILLER_441_1712 ();
 FILLCELL_X32 FILLER_441_1744 ();
 FILLCELL_X32 FILLER_441_1776 ();
 FILLCELL_X32 FILLER_441_1808 ();
 FILLCELL_X32 FILLER_441_1840 ();
 FILLCELL_X32 FILLER_441_1872 ();
 FILLCELL_X32 FILLER_441_1904 ();
 FILLCELL_X32 FILLER_441_1936 ();
 FILLCELL_X32 FILLER_441_1968 ();
 FILLCELL_X32 FILLER_441_2000 ();
 FILLCELL_X32 FILLER_441_2032 ();
 FILLCELL_X32 FILLER_441_2064 ();
 FILLCELL_X32 FILLER_441_2096 ();
 FILLCELL_X32 FILLER_441_2128 ();
 FILLCELL_X32 FILLER_441_2160 ();
 FILLCELL_X32 FILLER_441_2192 ();
 FILLCELL_X32 FILLER_441_2224 ();
 FILLCELL_X32 FILLER_441_2256 ();
 FILLCELL_X32 FILLER_441_2288 ();
 FILLCELL_X32 FILLER_441_2320 ();
 FILLCELL_X32 FILLER_441_2352 ();
 FILLCELL_X32 FILLER_441_2384 ();
 FILLCELL_X32 FILLER_441_2416 ();
 FILLCELL_X32 FILLER_441_2448 ();
 FILLCELL_X32 FILLER_441_2480 ();
 FILLCELL_X8 FILLER_441_2512 ();
 FILLCELL_X4 FILLER_441_2520 ();
 FILLCELL_X2 FILLER_441_2524 ();
 FILLCELL_X32 FILLER_441_2527 ();
 FILLCELL_X32 FILLER_441_2559 ();
 FILLCELL_X32 FILLER_441_2591 ();
 FILLCELL_X32 FILLER_441_2623 ();
 FILLCELL_X32 FILLER_441_2655 ();
 FILLCELL_X32 FILLER_441_2687 ();
 FILLCELL_X32 FILLER_441_2719 ();
 FILLCELL_X32 FILLER_441_2751 ();
 FILLCELL_X32 FILLER_441_2783 ();
 FILLCELL_X32 FILLER_441_2815 ();
 FILLCELL_X32 FILLER_441_2847 ();
 FILLCELL_X32 FILLER_441_2879 ();
 FILLCELL_X32 FILLER_441_2911 ();
 FILLCELL_X32 FILLER_441_2943 ();
 FILLCELL_X32 FILLER_441_2975 ();
 FILLCELL_X32 FILLER_441_3007 ();
 FILLCELL_X32 FILLER_441_3039 ();
 FILLCELL_X32 FILLER_441_3071 ();
 FILLCELL_X32 FILLER_441_3103 ();
 FILLCELL_X32 FILLER_441_3135 ();
 FILLCELL_X32 FILLER_441_3167 ();
 FILLCELL_X32 FILLER_441_3199 ();
 FILLCELL_X32 FILLER_441_3231 ();
 FILLCELL_X32 FILLER_441_3263 ();
 FILLCELL_X32 FILLER_441_3295 ();
 FILLCELL_X32 FILLER_441_3327 ();
 FILLCELL_X32 FILLER_441_3359 ();
 FILLCELL_X32 FILLER_441_3391 ();
 FILLCELL_X32 FILLER_441_3423 ();
 FILLCELL_X32 FILLER_441_3455 ();
 FILLCELL_X32 FILLER_441_3487 ();
 FILLCELL_X32 FILLER_441_3519 ();
 FILLCELL_X32 FILLER_441_3551 ();
 FILLCELL_X32 FILLER_441_3583 ();
 FILLCELL_X32 FILLER_441_3615 ();
 FILLCELL_X32 FILLER_441_3647 ();
 FILLCELL_X32 FILLER_441_3679 ();
 FILLCELL_X16 FILLER_441_3711 ();
 FILLCELL_X8 FILLER_441_3727 ();
 FILLCELL_X2 FILLER_441_3735 ();
 FILLCELL_X1 FILLER_441_3737 ();
 FILLCELL_X32 FILLER_442_1 ();
 FILLCELL_X32 FILLER_442_33 ();
 FILLCELL_X32 FILLER_442_65 ();
 FILLCELL_X32 FILLER_442_97 ();
 FILLCELL_X32 FILLER_442_129 ();
 FILLCELL_X32 FILLER_442_161 ();
 FILLCELL_X32 FILLER_442_193 ();
 FILLCELL_X32 FILLER_442_225 ();
 FILLCELL_X32 FILLER_442_257 ();
 FILLCELL_X32 FILLER_442_289 ();
 FILLCELL_X32 FILLER_442_321 ();
 FILLCELL_X32 FILLER_442_353 ();
 FILLCELL_X32 FILLER_442_385 ();
 FILLCELL_X32 FILLER_442_417 ();
 FILLCELL_X32 FILLER_442_449 ();
 FILLCELL_X32 FILLER_442_481 ();
 FILLCELL_X32 FILLER_442_513 ();
 FILLCELL_X32 FILLER_442_545 ();
 FILLCELL_X32 FILLER_442_577 ();
 FILLCELL_X16 FILLER_442_609 ();
 FILLCELL_X4 FILLER_442_625 ();
 FILLCELL_X2 FILLER_442_629 ();
 FILLCELL_X32 FILLER_442_632 ();
 FILLCELL_X32 FILLER_442_664 ();
 FILLCELL_X32 FILLER_442_696 ();
 FILLCELL_X32 FILLER_442_728 ();
 FILLCELL_X32 FILLER_442_760 ();
 FILLCELL_X32 FILLER_442_792 ();
 FILLCELL_X32 FILLER_442_824 ();
 FILLCELL_X32 FILLER_442_856 ();
 FILLCELL_X32 FILLER_442_888 ();
 FILLCELL_X32 FILLER_442_920 ();
 FILLCELL_X32 FILLER_442_952 ();
 FILLCELL_X32 FILLER_442_984 ();
 FILLCELL_X32 FILLER_442_1016 ();
 FILLCELL_X32 FILLER_442_1048 ();
 FILLCELL_X32 FILLER_442_1080 ();
 FILLCELL_X32 FILLER_442_1112 ();
 FILLCELL_X32 FILLER_442_1144 ();
 FILLCELL_X32 FILLER_442_1176 ();
 FILLCELL_X32 FILLER_442_1208 ();
 FILLCELL_X32 FILLER_442_1240 ();
 FILLCELL_X32 FILLER_442_1272 ();
 FILLCELL_X32 FILLER_442_1304 ();
 FILLCELL_X32 FILLER_442_1336 ();
 FILLCELL_X32 FILLER_442_1368 ();
 FILLCELL_X32 FILLER_442_1400 ();
 FILLCELL_X32 FILLER_442_1432 ();
 FILLCELL_X32 FILLER_442_1464 ();
 FILLCELL_X32 FILLER_442_1496 ();
 FILLCELL_X32 FILLER_442_1528 ();
 FILLCELL_X32 FILLER_442_1560 ();
 FILLCELL_X32 FILLER_442_1592 ();
 FILLCELL_X32 FILLER_442_1624 ();
 FILLCELL_X32 FILLER_442_1656 ();
 FILLCELL_X32 FILLER_442_1688 ();
 FILLCELL_X32 FILLER_442_1720 ();
 FILLCELL_X32 FILLER_442_1752 ();
 FILLCELL_X32 FILLER_442_1784 ();
 FILLCELL_X32 FILLER_442_1816 ();
 FILLCELL_X32 FILLER_442_1848 ();
 FILLCELL_X8 FILLER_442_1880 ();
 FILLCELL_X4 FILLER_442_1888 ();
 FILLCELL_X2 FILLER_442_1892 ();
 FILLCELL_X32 FILLER_442_1895 ();
 FILLCELL_X32 FILLER_442_1927 ();
 FILLCELL_X32 FILLER_442_1959 ();
 FILLCELL_X32 FILLER_442_1991 ();
 FILLCELL_X32 FILLER_442_2023 ();
 FILLCELL_X32 FILLER_442_2055 ();
 FILLCELL_X32 FILLER_442_2087 ();
 FILLCELL_X32 FILLER_442_2119 ();
 FILLCELL_X32 FILLER_442_2151 ();
 FILLCELL_X32 FILLER_442_2183 ();
 FILLCELL_X32 FILLER_442_2215 ();
 FILLCELL_X32 FILLER_442_2247 ();
 FILLCELL_X32 FILLER_442_2279 ();
 FILLCELL_X32 FILLER_442_2311 ();
 FILLCELL_X32 FILLER_442_2343 ();
 FILLCELL_X32 FILLER_442_2375 ();
 FILLCELL_X32 FILLER_442_2407 ();
 FILLCELL_X32 FILLER_442_2439 ();
 FILLCELL_X32 FILLER_442_2471 ();
 FILLCELL_X32 FILLER_442_2503 ();
 FILLCELL_X32 FILLER_442_2535 ();
 FILLCELL_X32 FILLER_442_2567 ();
 FILLCELL_X32 FILLER_442_2599 ();
 FILLCELL_X32 FILLER_442_2631 ();
 FILLCELL_X32 FILLER_442_2663 ();
 FILLCELL_X32 FILLER_442_2695 ();
 FILLCELL_X32 FILLER_442_2727 ();
 FILLCELL_X32 FILLER_442_2759 ();
 FILLCELL_X32 FILLER_442_2791 ();
 FILLCELL_X32 FILLER_442_2823 ();
 FILLCELL_X32 FILLER_442_2855 ();
 FILLCELL_X32 FILLER_442_2887 ();
 FILLCELL_X32 FILLER_442_2919 ();
 FILLCELL_X32 FILLER_442_2951 ();
 FILLCELL_X32 FILLER_442_2983 ();
 FILLCELL_X32 FILLER_442_3015 ();
 FILLCELL_X32 FILLER_442_3047 ();
 FILLCELL_X32 FILLER_442_3079 ();
 FILLCELL_X32 FILLER_442_3111 ();
 FILLCELL_X8 FILLER_442_3143 ();
 FILLCELL_X4 FILLER_442_3151 ();
 FILLCELL_X2 FILLER_442_3155 ();
 FILLCELL_X32 FILLER_442_3158 ();
 FILLCELL_X32 FILLER_442_3190 ();
 FILLCELL_X32 FILLER_442_3222 ();
 FILLCELL_X32 FILLER_442_3254 ();
 FILLCELL_X32 FILLER_442_3286 ();
 FILLCELL_X32 FILLER_442_3318 ();
 FILLCELL_X32 FILLER_442_3350 ();
 FILLCELL_X32 FILLER_442_3382 ();
 FILLCELL_X32 FILLER_442_3414 ();
 FILLCELL_X32 FILLER_442_3446 ();
 FILLCELL_X32 FILLER_442_3478 ();
 FILLCELL_X32 FILLER_442_3510 ();
 FILLCELL_X32 FILLER_442_3542 ();
 FILLCELL_X32 FILLER_442_3574 ();
 FILLCELL_X32 FILLER_442_3606 ();
 FILLCELL_X32 FILLER_442_3638 ();
 FILLCELL_X32 FILLER_442_3670 ();
 FILLCELL_X32 FILLER_442_3702 ();
 FILLCELL_X4 FILLER_442_3734 ();
 FILLCELL_X32 FILLER_443_1 ();
 FILLCELL_X32 FILLER_443_33 ();
 FILLCELL_X32 FILLER_443_65 ();
 FILLCELL_X32 FILLER_443_97 ();
 FILLCELL_X32 FILLER_443_129 ();
 FILLCELL_X32 FILLER_443_161 ();
 FILLCELL_X32 FILLER_443_193 ();
 FILLCELL_X32 FILLER_443_225 ();
 FILLCELL_X32 FILLER_443_257 ();
 FILLCELL_X32 FILLER_443_289 ();
 FILLCELL_X32 FILLER_443_321 ();
 FILLCELL_X32 FILLER_443_353 ();
 FILLCELL_X32 FILLER_443_385 ();
 FILLCELL_X32 FILLER_443_417 ();
 FILLCELL_X32 FILLER_443_449 ();
 FILLCELL_X32 FILLER_443_481 ();
 FILLCELL_X32 FILLER_443_513 ();
 FILLCELL_X32 FILLER_443_545 ();
 FILLCELL_X32 FILLER_443_577 ();
 FILLCELL_X32 FILLER_443_609 ();
 FILLCELL_X32 FILLER_443_641 ();
 FILLCELL_X32 FILLER_443_673 ();
 FILLCELL_X32 FILLER_443_705 ();
 FILLCELL_X32 FILLER_443_737 ();
 FILLCELL_X32 FILLER_443_769 ();
 FILLCELL_X32 FILLER_443_801 ();
 FILLCELL_X32 FILLER_443_833 ();
 FILLCELL_X32 FILLER_443_865 ();
 FILLCELL_X32 FILLER_443_897 ();
 FILLCELL_X32 FILLER_443_929 ();
 FILLCELL_X32 FILLER_443_961 ();
 FILLCELL_X32 FILLER_443_993 ();
 FILLCELL_X32 FILLER_443_1025 ();
 FILLCELL_X32 FILLER_443_1057 ();
 FILLCELL_X32 FILLER_443_1089 ();
 FILLCELL_X32 FILLER_443_1121 ();
 FILLCELL_X32 FILLER_443_1153 ();
 FILLCELL_X32 FILLER_443_1185 ();
 FILLCELL_X32 FILLER_443_1217 ();
 FILLCELL_X8 FILLER_443_1249 ();
 FILLCELL_X4 FILLER_443_1257 ();
 FILLCELL_X2 FILLER_443_1261 ();
 FILLCELL_X32 FILLER_443_1264 ();
 FILLCELL_X32 FILLER_443_1296 ();
 FILLCELL_X32 FILLER_443_1328 ();
 FILLCELL_X32 FILLER_443_1360 ();
 FILLCELL_X32 FILLER_443_1392 ();
 FILLCELL_X32 FILLER_443_1424 ();
 FILLCELL_X32 FILLER_443_1456 ();
 FILLCELL_X32 FILLER_443_1488 ();
 FILLCELL_X32 FILLER_443_1520 ();
 FILLCELL_X32 FILLER_443_1552 ();
 FILLCELL_X32 FILLER_443_1584 ();
 FILLCELL_X32 FILLER_443_1616 ();
 FILLCELL_X32 FILLER_443_1648 ();
 FILLCELL_X32 FILLER_443_1680 ();
 FILLCELL_X32 FILLER_443_1712 ();
 FILLCELL_X32 FILLER_443_1744 ();
 FILLCELL_X32 FILLER_443_1776 ();
 FILLCELL_X32 FILLER_443_1808 ();
 FILLCELL_X32 FILLER_443_1840 ();
 FILLCELL_X32 FILLER_443_1872 ();
 FILLCELL_X32 FILLER_443_1904 ();
 FILLCELL_X32 FILLER_443_1936 ();
 FILLCELL_X32 FILLER_443_1968 ();
 FILLCELL_X32 FILLER_443_2000 ();
 FILLCELL_X32 FILLER_443_2032 ();
 FILLCELL_X32 FILLER_443_2064 ();
 FILLCELL_X32 FILLER_443_2096 ();
 FILLCELL_X32 FILLER_443_2128 ();
 FILLCELL_X32 FILLER_443_2160 ();
 FILLCELL_X32 FILLER_443_2192 ();
 FILLCELL_X32 FILLER_443_2224 ();
 FILLCELL_X32 FILLER_443_2256 ();
 FILLCELL_X32 FILLER_443_2288 ();
 FILLCELL_X32 FILLER_443_2320 ();
 FILLCELL_X32 FILLER_443_2352 ();
 FILLCELL_X32 FILLER_443_2384 ();
 FILLCELL_X32 FILLER_443_2416 ();
 FILLCELL_X32 FILLER_443_2448 ();
 FILLCELL_X32 FILLER_443_2480 ();
 FILLCELL_X8 FILLER_443_2512 ();
 FILLCELL_X4 FILLER_443_2520 ();
 FILLCELL_X2 FILLER_443_2524 ();
 FILLCELL_X32 FILLER_443_2527 ();
 FILLCELL_X32 FILLER_443_2559 ();
 FILLCELL_X32 FILLER_443_2591 ();
 FILLCELL_X32 FILLER_443_2623 ();
 FILLCELL_X32 FILLER_443_2655 ();
 FILLCELL_X32 FILLER_443_2687 ();
 FILLCELL_X32 FILLER_443_2719 ();
 FILLCELL_X32 FILLER_443_2751 ();
 FILLCELL_X32 FILLER_443_2783 ();
 FILLCELL_X32 FILLER_443_2815 ();
 FILLCELL_X32 FILLER_443_2847 ();
 FILLCELL_X32 FILLER_443_2879 ();
 FILLCELL_X32 FILLER_443_2911 ();
 FILLCELL_X32 FILLER_443_2943 ();
 FILLCELL_X32 FILLER_443_2975 ();
 FILLCELL_X32 FILLER_443_3007 ();
 FILLCELL_X32 FILLER_443_3039 ();
 FILLCELL_X32 FILLER_443_3071 ();
 FILLCELL_X32 FILLER_443_3103 ();
 FILLCELL_X32 FILLER_443_3135 ();
 FILLCELL_X32 FILLER_443_3167 ();
 FILLCELL_X32 FILLER_443_3199 ();
 FILLCELL_X32 FILLER_443_3231 ();
 FILLCELL_X32 FILLER_443_3263 ();
 FILLCELL_X32 FILLER_443_3295 ();
 FILLCELL_X32 FILLER_443_3327 ();
 FILLCELL_X32 FILLER_443_3359 ();
 FILLCELL_X32 FILLER_443_3391 ();
 FILLCELL_X32 FILLER_443_3423 ();
 FILLCELL_X32 FILLER_443_3455 ();
 FILLCELL_X32 FILLER_443_3487 ();
 FILLCELL_X32 FILLER_443_3519 ();
 FILLCELL_X32 FILLER_443_3551 ();
 FILLCELL_X32 FILLER_443_3583 ();
 FILLCELL_X32 FILLER_443_3615 ();
 FILLCELL_X32 FILLER_443_3647 ();
 FILLCELL_X32 FILLER_443_3679 ();
 FILLCELL_X16 FILLER_443_3711 ();
 FILLCELL_X8 FILLER_443_3727 ();
 FILLCELL_X2 FILLER_443_3735 ();
 FILLCELL_X1 FILLER_443_3737 ();
 FILLCELL_X32 FILLER_444_1 ();
 FILLCELL_X32 FILLER_444_33 ();
 FILLCELL_X32 FILLER_444_65 ();
 FILLCELL_X32 FILLER_444_97 ();
 FILLCELL_X32 FILLER_444_129 ();
 FILLCELL_X32 FILLER_444_161 ();
 FILLCELL_X32 FILLER_444_193 ();
 FILLCELL_X32 FILLER_444_225 ();
 FILLCELL_X32 FILLER_444_257 ();
 FILLCELL_X32 FILLER_444_289 ();
 FILLCELL_X32 FILLER_444_321 ();
 FILLCELL_X32 FILLER_444_353 ();
 FILLCELL_X32 FILLER_444_385 ();
 FILLCELL_X32 FILLER_444_417 ();
 FILLCELL_X32 FILLER_444_449 ();
 FILLCELL_X32 FILLER_444_481 ();
 FILLCELL_X32 FILLER_444_513 ();
 FILLCELL_X32 FILLER_444_545 ();
 FILLCELL_X32 FILLER_444_577 ();
 FILLCELL_X16 FILLER_444_609 ();
 FILLCELL_X4 FILLER_444_625 ();
 FILLCELL_X2 FILLER_444_629 ();
 FILLCELL_X32 FILLER_444_632 ();
 FILLCELL_X32 FILLER_444_664 ();
 FILLCELL_X32 FILLER_444_696 ();
 FILLCELL_X32 FILLER_444_728 ();
 FILLCELL_X32 FILLER_444_760 ();
 FILLCELL_X32 FILLER_444_792 ();
 FILLCELL_X32 FILLER_444_824 ();
 FILLCELL_X32 FILLER_444_856 ();
 FILLCELL_X32 FILLER_444_888 ();
 FILLCELL_X32 FILLER_444_920 ();
 FILLCELL_X32 FILLER_444_952 ();
 FILLCELL_X32 FILLER_444_984 ();
 FILLCELL_X32 FILLER_444_1016 ();
 FILLCELL_X32 FILLER_444_1048 ();
 FILLCELL_X32 FILLER_444_1080 ();
 FILLCELL_X32 FILLER_444_1112 ();
 FILLCELL_X32 FILLER_444_1144 ();
 FILLCELL_X32 FILLER_444_1176 ();
 FILLCELL_X32 FILLER_444_1208 ();
 FILLCELL_X32 FILLER_444_1240 ();
 FILLCELL_X32 FILLER_444_1272 ();
 FILLCELL_X32 FILLER_444_1304 ();
 FILLCELL_X32 FILLER_444_1336 ();
 FILLCELL_X32 FILLER_444_1368 ();
 FILLCELL_X32 FILLER_444_1400 ();
 FILLCELL_X32 FILLER_444_1432 ();
 FILLCELL_X32 FILLER_444_1464 ();
 FILLCELL_X32 FILLER_444_1496 ();
 FILLCELL_X32 FILLER_444_1528 ();
 FILLCELL_X32 FILLER_444_1560 ();
 FILLCELL_X32 FILLER_444_1592 ();
 FILLCELL_X32 FILLER_444_1624 ();
 FILLCELL_X32 FILLER_444_1656 ();
 FILLCELL_X32 FILLER_444_1688 ();
 FILLCELL_X32 FILLER_444_1720 ();
 FILLCELL_X32 FILLER_444_1752 ();
 FILLCELL_X32 FILLER_444_1784 ();
 FILLCELL_X32 FILLER_444_1816 ();
 FILLCELL_X32 FILLER_444_1848 ();
 FILLCELL_X8 FILLER_444_1880 ();
 FILLCELL_X4 FILLER_444_1888 ();
 FILLCELL_X2 FILLER_444_1892 ();
 FILLCELL_X32 FILLER_444_1895 ();
 FILLCELL_X32 FILLER_444_1927 ();
 FILLCELL_X32 FILLER_444_1959 ();
 FILLCELL_X32 FILLER_444_1991 ();
 FILLCELL_X32 FILLER_444_2023 ();
 FILLCELL_X32 FILLER_444_2055 ();
 FILLCELL_X32 FILLER_444_2087 ();
 FILLCELL_X32 FILLER_444_2119 ();
 FILLCELL_X32 FILLER_444_2151 ();
 FILLCELL_X32 FILLER_444_2183 ();
 FILLCELL_X32 FILLER_444_2215 ();
 FILLCELL_X32 FILLER_444_2247 ();
 FILLCELL_X32 FILLER_444_2279 ();
 FILLCELL_X32 FILLER_444_2311 ();
 FILLCELL_X32 FILLER_444_2343 ();
 FILLCELL_X32 FILLER_444_2375 ();
 FILLCELL_X32 FILLER_444_2407 ();
 FILLCELL_X32 FILLER_444_2439 ();
 FILLCELL_X32 FILLER_444_2471 ();
 FILLCELL_X32 FILLER_444_2503 ();
 FILLCELL_X32 FILLER_444_2535 ();
 FILLCELL_X32 FILLER_444_2567 ();
 FILLCELL_X32 FILLER_444_2599 ();
 FILLCELL_X32 FILLER_444_2631 ();
 FILLCELL_X32 FILLER_444_2663 ();
 FILLCELL_X32 FILLER_444_2695 ();
 FILLCELL_X32 FILLER_444_2727 ();
 FILLCELL_X32 FILLER_444_2759 ();
 FILLCELL_X32 FILLER_444_2791 ();
 FILLCELL_X32 FILLER_444_2823 ();
 FILLCELL_X32 FILLER_444_2855 ();
 FILLCELL_X32 FILLER_444_2887 ();
 FILLCELL_X32 FILLER_444_2919 ();
 FILLCELL_X32 FILLER_444_2951 ();
 FILLCELL_X32 FILLER_444_2983 ();
 FILLCELL_X32 FILLER_444_3015 ();
 FILLCELL_X32 FILLER_444_3047 ();
 FILLCELL_X32 FILLER_444_3079 ();
 FILLCELL_X32 FILLER_444_3111 ();
 FILLCELL_X8 FILLER_444_3143 ();
 FILLCELL_X4 FILLER_444_3151 ();
 FILLCELL_X2 FILLER_444_3155 ();
 FILLCELL_X32 FILLER_444_3158 ();
 FILLCELL_X32 FILLER_444_3190 ();
 FILLCELL_X32 FILLER_444_3222 ();
 FILLCELL_X32 FILLER_444_3254 ();
 FILLCELL_X32 FILLER_444_3286 ();
 FILLCELL_X32 FILLER_444_3318 ();
 FILLCELL_X32 FILLER_444_3350 ();
 FILLCELL_X32 FILLER_444_3382 ();
 FILLCELL_X32 FILLER_444_3414 ();
 FILLCELL_X32 FILLER_444_3446 ();
 FILLCELL_X32 FILLER_444_3478 ();
 FILLCELL_X32 FILLER_444_3510 ();
 FILLCELL_X32 FILLER_444_3542 ();
 FILLCELL_X32 FILLER_444_3574 ();
 FILLCELL_X32 FILLER_444_3606 ();
 FILLCELL_X32 FILLER_444_3638 ();
 FILLCELL_X32 FILLER_444_3670 ();
 FILLCELL_X32 FILLER_444_3702 ();
 FILLCELL_X4 FILLER_444_3734 ();
 FILLCELL_X32 FILLER_445_1 ();
 FILLCELL_X32 FILLER_445_33 ();
 FILLCELL_X32 FILLER_445_65 ();
 FILLCELL_X32 FILLER_445_97 ();
 FILLCELL_X32 FILLER_445_129 ();
 FILLCELL_X32 FILLER_445_161 ();
 FILLCELL_X32 FILLER_445_193 ();
 FILLCELL_X32 FILLER_445_225 ();
 FILLCELL_X32 FILLER_445_257 ();
 FILLCELL_X32 FILLER_445_289 ();
 FILLCELL_X32 FILLER_445_321 ();
 FILLCELL_X32 FILLER_445_353 ();
 FILLCELL_X32 FILLER_445_385 ();
 FILLCELL_X32 FILLER_445_417 ();
 FILLCELL_X32 FILLER_445_449 ();
 FILLCELL_X32 FILLER_445_481 ();
 FILLCELL_X32 FILLER_445_513 ();
 FILLCELL_X32 FILLER_445_545 ();
 FILLCELL_X32 FILLER_445_577 ();
 FILLCELL_X32 FILLER_445_609 ();
 FILLCELL_X32 FILLER_445_641 ();
 FILLCELL_X32 FILLER_445_673 ();
 FILLCELL_X32 FILLER_445_705 ();
 FILLCELL_X32 FILLER_445_737 ();
 FILLCELL_X32 FILLER_445_769 ();
 FILLCELL_X32 FILLER_445_801 ();
 FILLCELL_X32 FILLER_445_833 ();
 FILLCELL_X32 FILLER_445_865 ();
 FILLCELL_X32 FILLER_445_897 ();
 FILLCELL_X32 FILLER_445_929 ();
 FILLCELL_X32 FILLER_445_961 ();
 FILLCELL_X32 FILLER_445_993 ();
 FILLCELL_X32 FILLER_445_1025 ();
 FILLCELL_X32 FILLER_445_1057 ();
 FILLCELL_X32 FILLER_445_1089 ();
 FILLCELL_X32 FILLER_445_1121 ();
 FILLCELL_X32 FILLER_445_1153 ();
 FILLCELL_X32 FILLER_445_1185 ();
 FILLCELL_X32 FILLER_445_1217 ();
 FILLCELL_X8 FILLER_445_1249 ();
 FILLCELL_X4 FILLER_445_1257 ();
 FILLCELL_X2 FILLER_445_1261 ();
 FILLCELL_X32 FILLER_445_1264 ();
 FILLCELL_X32 FILLER_445_1296 ();
 FILLCELL_X32 FILLER_445_1328 ();
 FILLCELL_X32 FILLER_445_1360 ();
 FILLCELL_X32 FILLER_445_1392 ();
 FILLCELL_X32 FILLER_445_1424 ();
 FILLCELL_X32 FILLER_445_1456 ();
 FILLCELL_X32 FILLER_445_1488 ();
 FILLCELL_X32 FILLER_445_1520 ();
 FILLCELL_X32 FILLER_445_1552 ();
 FILLCELL_X32 FILLER_445_1584 ();
 FILLCELL_X32 FILLER_445_1616 ();
 FILLCELL_X32 FILLER_445_1648 ();
 FILLCELL_X32 FILLER_445_1680 ();
 FILLCELL_X32 FILLER_445_1712 ();
 FILLCELL_X32 FILLER_445_1744 ();
 FILLCELL_X32 FILLER_445_1776 ();
 FILLCELL_X32 FILLER_445_1808 ();
 FILLCELL_X32 FILLER_445_1840 ();
 FILLCELL_X32 FILLER_445_1872 ();
 FILLCELL_X32 FILLER_445_1904 ();
 FILLCELL_X32 FILLER_445_1936 ();
 FILLCELL_X32 FILLER_445_1968 ();
 FILLCELL_X32 FILLER_445_2000 ();
 FILLCELL_X32 FILLER_445_2032 ();
 FILLCELL_X32 FILLER_445_2064 ();
 FILLCELL_X32 FILLER_445_2096 ();
 FILLCELL_X32 FILLER_445_2128 ();
 FILLCELL_X32 FILLER_445_2160 ();
 FILLCELL_X32 FILLER_445_2192 ();
 FILLCELL_X32 FILLER_445_2224 ();
 FILLCELL_X32 FILLER_445_2256 ();
 FILLCELL_X32 FILLER_445_2288 ();
 FILLCELL_X32 FILLER_445_2320 ();
 FILLCELL_X32 FILLER_445_2352 ();
 FILLCELL_X32 FILLER_445_2384 ();
 FILLCELL_X32 FILLER_445_2416 ();
 FILLCELL_X32 FILLER_445_2448 ();
 FILLCELL_X32 FILLER_445_2480 ();
 FILLCELL_X8 FILLER_445_2512 ();
 FILLCELL_X4 FILLER_445_2520 ();
 FILLCELL_X2 FILLER_445_2524 ();
 FILLCELL_X32 FILLER_445_2527 ();
 FILLCELL_X32 FILLER_445_2559 ();
 FILLCELL_X32 FILLER_445_2591 ();
 FILLCELL_X32 FILLER_445_2623 ();
 FILLCELL_X32 FILLER_445_2655 ();
 FILLCELL_X32 FILLER_445_2687 ();
 FILLCELL_X32 FILLER_445_2719 ();
 FILLCELL_X32 FILLER_445_2751 ();
 FILLCELL_X32 FILLER_445_2783 ();
 FILLCELL_X32 FILLER_445_2815 ();
 FILLCELL_X32 FILLER_445_2847 ();
 FILLCELL_X32 FILLER_445_2879 ();
 FILLCELL_X32 FILLER_445_2911 ();
 FILLCELL_X32 FILLER_445_2943 ();
 FILLCELL_X32 FILLER_445_2975 ();
 FILLCELL_X32 FILLER_445_3007 ();
 FILLCELL_X32 FILLER_445_3039 ();
 FILLCELL_X32 FILLER_445_3071 ();
 FILLCELL_X32 FILLER_445_3103 ();
 FILLCELL_X32 FILLER_445_3135 ();
 FILLCELL_X32 FILLER_445_3167 ();
 FILLCELL_X32 FILLER_445_3199 ();
 FILLCELL_X32 FILLER_445_3231 ();
 FILLCELL_X32 FILLER_445_3263 ();
 FILLCELL_X32 FILLER_445_3295 ();
 FILLCELL_X32 FILLER_445_3327 ();
 FILLCELL_X32 FILLER_445_3359 ();
 FILLCELL_X32 FILLER_445_3391 ();
 FILLCELL_X32 FILLER_445_3423 ();
 FILLCELL_X32 FILLER_445_3455 ();
 FILLCELL_X32 FILLER_445_3487 ();
 FILLCELL_X32 FILLER_445_3519 ();
 FILLCELL_X32 FILLER_445_3551 ();
 FILLCELL_X32 FILLER_445_3583 ();
 FILLCELL_X32 FILLER_445_3615 ();
 FILLCELL_X32 FILLER_445_3647 ();
 FILLCELL_X32 FILLER_445_3679 ();
 FILLCELL_X16 FILLER_445_3711 ();
 FILLCELL_X8 FILLER_445_3727 ();
 FILLCELL_X2 FILLER_445_3735 ();
 FILLCELL_X1 FILLER_445_3737 ();
 FILLCELL_X32 FILLER_446_1 ();
 FILLCELL_X32 FILLER_446_33 ();
 FILLCELL_X32 FILLER_446_65 ();
 FILLCELL_X32 FILLER_446_97 ();
 FILLCELL_X32 FILLER_446_129 ();
 FILLCELL_X32 FILLER_446_161 ();
 FILLCELL_X32 FILLER_446_193 ();
 FILLCELL_X32 FILLER_446_225 ();
 FILLCELL_X32 FILLER_446_257 ();
 FILLCELL_X32 FILLER_446_289 ();
 FILLCELL_X32 FILLER_446_321 ();
 FILLCELL_X32 FILLER_446_353 ();
 FILLCELL_X32 FILLER_446_385 ();
 FILLCELL_X32 FILLER_446_417 ();
 FILLCELL_X32 FILLER_446_449 ();
 FILLCELL_X32 FILLER_446_481 ();
 FILLCELL_X32 FILLER_446_513 ();
 FILLCELL_X32 FILLER_446_545 ();
 FILLCELL_X32 FILLER_446_577 ();
 FILLCELL_X16 FILLER_446_609 ();
 FILLCELL_X4 FILLER_446_625 ();
 FILLCELL_X2 FILLER_446_629 ();
 FILLCELL_X32 FILLER_446_632 ();
 FILLCELL_X32 FILLER_446_664 ();
 FILLCELL_X32 FILLER_446_696 ();
 FILLCELL_X32 FILLER_446_728 ();
 FILLCELL_X32 FILLER_446_760 ();
 FILLCELL_X32 FILLER_446_792 ();
 FILLCELL_X32 FILLER_446_824 ();
 FILLCELL_X32 FILLER_446_856 ();
 FILLCELL_X32 FILLER_446_888 ();
 FILLCELL_X32 FILLER_446_920 ();
 FILLCELL_X32 FILLER_446_952 ();
 FILLCELL_X32 FILLER_446_984 ();
 FILLCELL_X32 FILLER_446_1016 ();
 FILLCELL_X32 FILLER_446_1048 ();
 FILLCELL_X32 FILLER_446_1080 ();
 FILLCELL_X32 FILLER_446_1112 ();
 FILLCELL_X32 FILLER_446_1144 ();
 FILLCELL_X32 FILLER_446_1176 ();
 FILLCELL_X32 FILLER_446_1208 ();
 FILLCELL_X32 FILLER_446_1240 ();
 FILLCELL_X32 FILLER_446_1272 ();
 FILLCELL_X32 FILLER_446_1304 ();
 FILLCELL_X32 FILLER_446_1336 ();
 FILLCELL_X32 FILLER_446_1368 ();
 FILLCELL_X32 FILLER_446_1400 ();
 FILLCELL_X32 FILLER_446_1432 ();
 FILLCELL_X32 FILLER_446_1464 ();
 FILLCELL_X32 FILLER_446_1496 ();
 FILLCELL_X32 FILLER_446_1528 ();
 FILLCELL_X32 FILLER_446_1560 ();
 FILLCELL_X32 FILLER_446_1592 ();
 FILLCELL_X32 FILLER_446_1624 ();
 FILLCELL_X32 FILLER_446_1656 ();
 FILLCELL_X32 FILLER_446_1688 ();
 FILLCELL_X32 FILLER_446_1720 ();
 FILLCELL_X32 FILLER_446_1752 ();
 FILLCELL_X32 FILLER_446_1784 ();
 FILLCELL_X32 FILLER_446_1816 ();
 FILLCELL_X32 FILLER_446_1848 ();
 FILLCELL_X8 FILLER_446_1880 ();
 FILLCELL_X4 FILLER_446_1888 ();
 FILLCELL_X2 FILLER_446_1892 ();
 FILLCELL_X32 FILLER_446_1895 ();
 FILLCELL_X32 FILLER_446_1927 ();
 FILLCELL_X32 FILLER_446_1959 ();
 FILLCELL_X32 FILLER_446_1991 ();
 FILLCELL_X32 FILLER_446_2023 ();
 FILLCELL_X32 FILLER_446_2055 ();
 FILLCELL_X32 FILLER_446_2087 ();
 FILLCELL_X32 FILLER_446_2119 ();
 FILLCELL_X32 FILLER_446_2151 ();
 FILLCELL_X32 FILLER_446_2183 ();
 FILLCELL_X32 FILLER_446_2215 ();
 FILLCELL_X32 FILLER_446_2247 ();
 FILLCELL_X32 FILLER_446_2279 ();
 FILLCELL_X32 FILLER_446_2311 ();
 FILLCELL_X32 FILLER_446_2343 ();
 FILLCELL_X32 FILLER_446_2375 ();
 FILLCELL_X32 FILLER_446_2407 ();
 FILLCELL_X32 FILLER_446_2439 ();
 FILLCELL_X32 FILLER_446_2471 ();
 FILLCELL_X32 FILLER_446_2503 ();
 FILLCELL_X32 FILLER_446_2535 ();
 FILLCELL_X32 FILLER_446_2567 ();
 FILLCELL_X32 FILLER_446_2599 ();
 FILLCELL_X32 FILLER_446_2631 ();
 FILLCELL_X32 FILLER_446_2663 ();
 FILLCELL_X32 FILLER_446_2695 ();
 FILLCELL_X32 FILLER_446_2727 ();
 FILLCELL_X32 FILLER_446_2759 ();
 FILLCELL_X32 FILLER_446_2791 ();
 FILLCELL_X32 FILLER_446_2823 ();
 FILLCELL_X32 FILLER_446_2855 ();
 FILLCELL_X32 FILLER_446_2887 ();
 FILLCELL_X32 FILLER_446_2919 ();
 FILLCELL_X32 FILLER_446_2951 ();
 FILLCELL_X32 FILLER_446_2983 ();
 FILLCELL_X32 FILLER_446_3015 ();
 FILLCELL_X32 FILLER_446_3047 ();
 FILLCELL_X32 FILLER_446_3079 ();
 FILLCELL_X32 FILLER_446_3111 ();
 FILLCELL_X8 FILLER_446_3143 ();
 FILLCELL_X4 FILLER_446_3151 ();
 FILLCELL_X2 FILLER_446_3155 ();
 FILLCELL_X32 FILLER_446_3158 ();
 FILLCELL_X32 FILLER_446_3190 ();
 FILLCELL_X32 FILLER_446_3222 ();
 FILLCELL_X32 FILLER_446_3254 ();
 FILLCELL_X32 FILLER_446_3286 ();
 FILLCELL_X32 FILLER_446_3318 ();
 FILLCELL_X32 FILLER_446_3350 ();
 FILLCELL_X32 FILLER_446_3382 ();
 FILLCELL_X32 FILLER_446_3414 ();
 FILLCELL_X32 FILLER_446_3446 ();
 FILLCELL_X32 FILLER_446_3478 ();
 FILLCELL_X32 FILLER_446_3510 ();
 FILLCELL_X32 FILLER_446_3542 ();
 FILLCELL_X32 FILLER_446_3574 ();
 FILLCELL_X32 FILLER_446_3606 ();
 FILLCELL_X32 FILLER_446_3638 ();
 FILLCELL_X32 FILLER_446_3670 ();
 FILLCELL_X32 FILLER_446_3702 ();
 FILLCELL_X4 FILLER_446_3734 ();
 FILLCELL_X32 FILLER_447_1 ();
 FILLCELL_X32 FILLER_447_33 ();
 FILLCELL_X32 FILLER_447_65 ();
 FILLCELL_X32 FILLER_447_97 ();
 FILLCELL_X32 FILLER_447_129 ();
 FILLCELL_X32 FILLER_447_161 ();
 FILLCELL_X32 FILLER_447_193 ();
 FILLCELL_X32 FILLER_447_225 ();
 FILLCELL_X32 FILLER_447_257 ();
 FILLCELL_X32 FILLER_447_289 ();
 FILLCELL_X32 FILLER_447_321 ();
 FILLCELL_X32 FILLER_447_353 ();
 FILLCELL_X32 FILLER_447_385 ();
 FILLCELL_X32 FILLER_447_417 ();
 FILLCELL_X32 FILLER_447_449 ();
 FILLCELL_X32 FILLER_447_481 ();
 FILLCELL_X32 FILLER_447_513 ();
 FILLCELL_X32 FILLER_447_545 ();
 FILLCELL_X32 FILLER_447_577 ();
 FILLCELL_X32 FILLER_447_609 ();
 FILLCELL_X32 FILLER_447_641 ();
 FILLCELL_X32 FILLER_447_673 ();
 FILLCELL_X32 FILLER_447_705 ();
 FILLCELL_X32 FILLER_447_737 ();
 FILLCELL_X32 FILLER_447_769 ();
 FILLCELL_X32 FILLER_447_801 ();
 FILLCELL_X32 FILLER_447_833 ();
 FILLCELL_X32 FILLER_447_865 ();
 FILLCELL_X32 FILLER_447_897 ();
 FILLCELL_X32 FILLER_447_929 ();
 FILLCELL_X32 FILLER_447_961 ();
 FILLCELL_X32 FILLER_447_993 ();
 FILLCELL_X32 FILLER_447_1025 ();
 FILLCELL_X32 FILLER_447_1057 ();
 FILLCELL_X32 FILLER_447_1089 ();
 FILLCELL_X32 FILLER_447_1121 ();
 FILLCELL_X32 FILLER_447_1153 ();
 FILLCELL_X32 FILLER_447_1185 ();
 FILLCELL_X32 FILLER_447_1217 ();
 FILLCELL_X8 FILLER_447_1249 ();
 FILLCELL_X4 FILLER_447_1257 ();
 FILLCELL_X2 FILLER_447_1261 ();
 FILLCELL_X32 FILLER_447_1264 ();
 FILLCELL_X32 FILLER_447_1296 ();
 FILLCELL_X32 FILLER_447_1328 ();
 FILLCELL_X32 FILLER_447_1360 ();
 FILLCELL_X32 FILLER_447_1392 ();
 FILLCELL_X32 FILLER_447_1424 ();
 FILLCELL_X32 FILLER_447_1456 ();
 FILLCELL_X32 FILLER_447_1488 ();
 FILLCELL_X32 FILLER_447_1520 ();
 FILLCELL_X32 FILLER_447_1552 ();
 FILLCELL_X32 FILLER_447_1584 ();
 FILLCELL_X32 FILLER_447_1616 ();
 FILLCELL_X32 FILLER_447_1648 ();
 FILLCELL_X32 FILLER_447_1680 ();
 FILLCELL_X32 FILLER_447_1712 ();
 FILLCELL_X32 FILLER_447_1744 ();
 FILLCELL_X32 FILLER_447_1776 ();
 FILLCELL_X32 FILLER_447_1808 ();
 FILLCELL_X32 FILLER_447_1840 ();
 FILLCELL_X32 FILLER_447_1872 ();
 FILLCELL_X32 FILLER_447_1904 ();
 FILLCELL_X32 FILLER_447_1936 ();
 FILLCELL_X32 FILLER_447_1968 ();
 FILLCELL_X32 FILLER_447_2000 ();
 FILLCELL_X32 FILLER_447_2032 ();
 FILLCELL_X32 FILLER_447_2064 ();
 FILLCELL_X32 FILLER_447_2096 ();
 FILLCELL_X32 FILLER_447_2128 ();
 FILLCELL_X32 FILLER_447_2160 ();
 FILLCELL_X32 FILLER_447_2192 ();
 FILLCELL_X32 FILLER_447_2224 ();
 FILLCELL_X32 FILLER_447_2256 ();
 FILLCELL_X32 FILLER_447_2288 ();
 FILLCELL_X32 FILLER_447_2320 ();
 FILLCELL_X32 FILLER_447_2352 ();
 FILLCELL_X32 FILLER_447_2384 ();
 FILLCELL_X32 FILLER_447_2416 ();
 FILLCELL_X32 FILLER_447_2448 ();
 FILLCELL_X32 FILLER_447_2480 ();
 FILLCELL_X8 FILLER_447_2512 ();
 FILLCELL_X4 FILLER_447_2520 ();
 FILLCELL_X2 FILLER_447_2524 ();
 FILLCELL_X32 FILLER_447_2527 ();
 FILLCELL_X32 FILLER_447_2559 ();
 FILLCELL_X32 FILLER_447_2591 ();
 FILLCELL_X32 FILLER_447_2623 ();
 FILLCELL_X32 FILLER_447_2655 ();
 FILLCELL_X32 FILLER_447_2687 ();
 FILLCELL_X32 FILLER_447_2719 ();
 FILLCELL_X32 FILLER_447_2751 ();
 FILLCELL_X32 FILLER_447_2783 ();
 FILLCELL_X32 FILLER_447_2815 ();
 FILLCELL_X32 FILLER_447_2847 ();
 FILLCELL_X32 FILLER_447_2879 ();
 FILLCELL_X32 FILLER_447_2911 ();
 FILLCELL_X32 FILLER_447_2943 ();
 FILLCELL_X32 FILLER_447_2975 ();
 FILLCELL_X32 FILLER_447_3007 ();
 FILLCELL_X32 FILLER_447_3039 ();
 FILLCELL_X32 FILLER_447_3071 ();
 FILLCELL_X32 FILLER_447_3103 ();
 FILLCELL_X32 FILLER_447_3135 ();
 FILLCELL_X32 FILLER_447_3167 ();
 FILLCELL_X32 FILLER_447_3199 ();
 FILLCELL_X32 FILLER_447_3231 ();
 FILLCELL_X32 FILLER_447_3263 ();
 FILLCELL_X32 FILLER_447_3295 ();
 FILLCELL_X32 FILLER_447_3327 ();
 FILLCELL_X32 FILLER_447_3359 ();
 FILLCELL_X32 FILLER_447_3391 ();
 FILLCELL_X32 FILLER_447_3423 ();
 FILLCELL_X32 FILLER_447_3455 ();
 FILLCELL_X32 FILLER_447_3487 ();
 FILLCELL_X32 FILLER_447_3519 ();
 FILLCELL_X32 FILLER_447_3551 ();
 FILLCELL_X32 FILLER_447_3583 ();
 FILLCELL_X32 FILLER_447_3615 ();
 FILLCELL_X32 FILLER_447_3647 ();
 FILLCELL_X32 FILLER_447_3679 ();
 FILLCELL_X16 FILLER_447_3711 ();
 FILLCELL_X8 FILLER_447_3727 ();
 FILLCELL_X2 FILLER_447_3735 ();
 FILLCELL_X1 FILLER_447_3737 ();
 FILLCELL_X32 FILLER_448_1 ();
 FILLCELL_X32 FILLER_448_33 ();
 FILLCELL_X32 FILLER_448_65 ();
 FILLCELL_X32 FILLER_448_97 ();
 FILLCELL_X32 FILLER_448_129 ();
 FILLCELL_X32 FILLER_448_161 ();
 FILLCELL_X32 FILLER_448_193 ();
 FILLCELL_X32 FILLER_448_225 ();
 FILLCELL_X32 FILLER_448_257 ();
 FILLCELL_X32 FILLER_448_289 ();
 FILLCELL_X32 FILLER_448_321 ();
 FILLCELL_X32 FILLER_448_353 ();
 FILLCELL_X32 FILLER_448_385 ();
 FILLCELL_X32 FILLER_448_417 ();
 FILLCELL_X32 FILLER_448_449 ();
 FILLCELL_X32 FILLER_448_481 ();
 FILLCELL_X32 FILLER_448_513 ();
 FILLCELL_X32 FILLER_448_545 ();
 FILLCELL_X32 FILLER_448_577 ();
 FILLCELL_X16 FILLER_448_609 ();
 FILLCELL_X4 FILLER_448_625 ();
 FILLCELL_X2 FILLER_448_629 ();
 FILLCELL_X32 FILLER_448_632 ();
 FILLCELL_X32 FILLER_448_664 ();
 FILLCELL_X32 FILLER_448_696 ();
 FILLCELL_X32 FILLER_448_728 ();
 FILLCELL_X32 FILLER_448_760 ();
 FILLCELL_X32 FILLER_448_792 ();
 FILLCELL_X32 FILLER_448_824 ();
 FILLCELL_X32 FILLER_448_856 ();
 FILLCELL_X32 FILLER_448_888 ();
 FILLCELL_X32 FILLER_448_920 ();
 FILLCELL_X32 FILLER_448_952 ();
 FILLCELL_X32 FILLER_448_984 ();
 FILLCELL_X32 FILLER_448_1016 ();
 FILLCELL_X32 FILLER_448_1048 ();
 FILLCELL_X32 FILLER_448_1080 ();
 FILLCELL_X32 FILLER_448_1112 ();
 FILLCELL_X32 FILLER_448_1144 ();
 FILLCELL_X32 FILLER_448_1176 ();
 FILLCELL_X32 FILLER_448_1208 ();
 FILLCELL_X32 FILLER_448_1240 ();
 FILLCELL_X32 FILLER_448_1272 ();
 FILLCELL_X32 FILLER_448_1304 ();
 FILLCELL_X32 FILLER_448_1336 ();
 FILLCELL_X32 FILLER_448_1368 ();
 FILLCELL_X32 FILLER_448_1400 ();
 FILLCELL_X32 FILLER_448_1432 ();
 FILLCELL_X32 FILLER_448_1464 ();
 FILLCELL_X32 FILLER_448_1496 ();
 FILLCELL_X32 FILLER_448_1528 ();
 FILLCELL_X32 FILLER_448_1560 ();
 FILLCELL_X32 FILLER_448_1592 ();
 FILLCELL_X32 FILLER_448_1624 ();
 FILLCELL_X32 FILLER_448_1656 ();
 FILLCELL_X32 FILLER_448_1688 ();
 FILLCELL_X32 FILLER_448_1720 ();
 FILLCELL_X32 FILLER_448_1752 ();
 FILLCELL_X32 FILLER_448_1784 ();
 FILLCELL_X32 FILLER_448_1816 ();
 FILLCELL_X32 FILLER_448_1848 ();
 FILLCELL_X8 FILLER_448_1880 ();
 FILLCELL_X4 FILLER_448_1888 ();
 FILLCELL_X2 FILLER_448_1892 ();
 FILLCELL_X32 FILLER_448_1895 ();
 FILLCELL_X32 FILLER_448_1927 ();
 FILLCELL_X32 FILLER_448_1959 ();
 FILLCELL_X32 FILLER_448_1991 ();
 FILLCELL_X32 FILLER_448_2023 ();
 FILLCELL_X32 FILLER_448_2055 ();
 FILLCELL_X32 FILLER_448_2087 ();
 FILLCELL_X32 FILLER_448_2119 ();
 FILLCELL_X32 FILLER_448_2151 ();
 FILLCELL_X32 FILLER_448_2183 ();
 FILLCELL_X32 FILLER_448_2215 ();
 FILLCELL_X32 FILLER_448_2247 ();
 FILLCELL_X32 FILLER_448_2279 ();
 FILLCELL_X32 FILLER_448_2311 ();
 FILLCELL_X32 FILLER_448_2343 ();
 FILLCELL_X32 FILLER_448_2375 ();
 FILLCELL_X32 FILLER_448_2407 ();
 FILLCELL_X32 FILLER_448_2439 ();
 FILLCELL_X32 FILLER_448_2471 ();
 FILLCELL_X32 FILLER_448_2503 ();
 FILLCELL_X32 FILLER_448_2535 ();
 FILLCELL_X32 FILLER_448_2567 ();
 FILLCELL_X32 FILLER_448_2599 ();
 FILLCELL_X32 FILLER_448_2631 ();
 FILLCELL_X32 FILLER_448_2663 ();
 FILLCELL_X32 FILLER_448_2695 ();
 FILLCELL_X32 FILLER_448_2727 ();
 FILLCELL_X32 FILLER_448_2759 ();
 FILLCELL_X32 FILLER_448_2791 ();
 FILLCELL_X32 FILLER_448_2823 ();
 FILLCELL_X32 FILLER_448_2855 ();
 FILLCELL_X32 FILLER_448_2887 ();
 FILLCELL_X32 FILLER_448_2919 ();
 FILLCELL_X32 FILLER_448_2951 ();
 FILLCELL_X32 FILLER_448_2983 ();
 FILLCELL_X32 FILLER_448_3015 ();
 FILLCELL_X32 FILLER_448_3047 ();
 FILLCELL_X32 FILLER_448_3079 ();
 FILLCELL_X32 FILLER_448_3111 ();
 FILLCELL_X8 FILLER_448_3143 ();
 FILLCELL_X4 FILLER_448_3151 ();
 FILLCELL_X2 FILLER_448_3155 ();
 FILLCELL_X32 FILLER_448_3158 ();
 FILLCELL_X32 FILLER_448_3190 ();
 FILLCELL_X32 FILLER_448_3222 ();
 FILLCELL_X32 FILLER_448_3254 ();
 FILLCELL_X32 FILLER_448_3286 ();
 FILLCELL_X32 FILLER_448_3318 ();
 FILLCELL_X32 FILLER_448_3350 ();
 FILLCELL_X32 FILLER_448_3382 ();
 FILLCELL_X32 FILLER_448_3414 ();
 FILLCELL_X32 FILLER_448_3446 ();
 FILLCELL_X32 FILLER_448_3478 ();
 FILLCELL_X32 FILLER_448_3510 ();
 FILLCELL_X32 FILLER_448_3542 ();
 FILLCELL_X32 FILLER_448_3574 ();
 FILLCELL_X32 FILLER_448_3606 ();
 FILLCELL_X32 FILLER_448_3638 ();
 FILLCELL_X32 FILLER_448_3670 ();
 FILLCELL_X32 FILLER_448_3702 ();
 FILLCELL_X4 FILLER_448_3734 ();
 FILLCELL_X32 FILLER_449_1 ();
 FILLCELL_X32 FILLER_449_33 ();
 FILLCELL_X32 FILLER_449_65 ();
 FILLCELL_X32 FILLER_449_97 ();
 FILLCELL_X32 FILLER_449_129 ();
 FILLCELL_X32 FILLER_449_161 ();
 FILLCELL_X32 FILLER_449_193 ();
 FILLCELL_X32 FILLER_449_225 ();
 FILLCELL_X32 FILLER_449_257 ();
 FILLCELL_X32 FILLER_449_289 ();
 FILLCELL_X32 FILLER_449_321 ();
 FILLCELL_X32 FILLER_449_353 ();
 FILLCELL_X32 FILLER_449_385 ();
 FILLCELL_X32 FILLER_449_417 ();
 FILLCELL_X32 FILLER_449_449 ();
 FILLCELL_X32 FILLER_449_481 ();
 FILLCELL_X32 FILLER_449_513 ();
 FILLCELL_X32 FILLER_449_545 ();
 FILLCELL_X32 FILLER_449_577 ();
 FILLCELL_X32 FILLER_449_609 ();
 FILLCELL_X32 FILLER_449_641 ();
 FILLCELL_X32 FILLER_449_673 ();
 FILLCELL_X32 FILLER_449_705 ();
 FILLCELL_X32 FILLER_449_737 ();
 FILLCELL_X32 FILLER_449_769 ();
 FILLCELL_X32 FILLER_449_801 ();
 FILLCELL_X32 FILLER_449_833 ();
 FILLCELL_X32 FILLER_449_865 ();
 FILLCELL_X32 FILLER_449_897 ();
 FILLCELL_X32 FILLER_449_929 ();
 FILLCELL_X32 FILLER_449_961 ();
 FILLCELL_X32 FILLER_449_993 ();
 FILLCELL_X32 FILLER_449_1025 ();
 FILLCELL_X32 FILLER_449_1057 ();
 FILLCELL_X32 FILLER_449_1089 ();
 FILLCELL_X32 FILLER_449_1121 ();
 FILLCELL_X32 FILLER_449_1153 ();
 FILLCELL_X32 FILLER_449_1185 ();
 FILLCELL_X32 FILLER_449_1217 ();
 FILLCELL_X8 FILLER_449_1249 ();
 FILLCELL_X4 FILLER_449_1257 ();
 FILLCELL_X2 FILLER_449_1261 ();
 FILLCELL_X32 FILLER_449_1264 ();
 FILLCELL_X32 FILLER_449_1296 ();
 FILLCELL_X32 FILLER_449_1328 ();
 FILLCELL_X32 FILLER_449_1360 ();
 FILLCELL_X32 FILLER_449_1392 ();
 FILLCELL_X32 FILLER_449_1424 ();
 FILLCELL_X32 FILLER_449_1456 ();
 FILLCELL_X32 FILLER_449_1488 ();
 FILLCELL_X32 FILLER_449_1520 ();
 FILLCELL_X32 FILLER_449_1552 ();
 FILLCELL_X32 FILLER_449_1584 ();
 FILLCELL_X32 FILLER_449_1616 ();
 FILLCELL_X32 FILLER_449_1648 ();
 FILLCELL_X32 FILLER_449_1680 ();
 FILLCELL_X32 FILLER_449_1712 ();
 FILLCELL_X32 FILLER_449_1744 ();
 FILLCELL_X32 FILLER_449_1776 ();
 FILLCELL_X32 FILLER_449_1808 ();
 FILLCELL_X32 FILLER_449_1840 ();
 FILLCELL_X32 FILLER_449_1872 ();
 FILLCELL_X32 FILLER_449_1904 ();
 FILLCELL_X32 FILLER_449_1936 ();
 FILLCELL_X32 FILLER_449_1968 ();
 FILLCELL_X32 FILLER_449_2000 ();
 FILLCELL_X32 FILLER_449_2032 ();
 FILLCELL_X32 FILLER_449_2064 ();
 FILLCELL_X32 FILLER_449_2096 ();
 FILLCELL_X32 FILLER_449_2128 ();
 FILLCELL_X32 FILLER_449_2160 ();
 FILLCELL_X32 FILLER_449_2192 ();
 FILLCELL_X32 FILLER_449_2224 ();
 FILLCELL_X32 FILLER_449_2256 ();
 FILLCELL_X32 FILLER_449_2288 ();
 FILLCELL_X32 FILLER_449_2320 ();
 FILLCELL_X32 FILLER_449_2352 ();
 FILLCELL_X32 FILLER_449_2384 ();
 FILLCELL_X32 FILLER_449_2416 ();
 FILLCELL_X32 FILLER_449_2448 ();
 FILLCELL_X32 FILLER_449_2480 ();
 FILLCELL_X8 FILLER_449_2512 ();
 FILLCELL_X4 FILLER_449_2520 ();
 FILLCELL_X2 FILLER_449_2524 ();
 FILLCELL_X32 FILLER_449_2527 ();
 FILLCELL_X32 FILLER_449_2559 ();
 FILLCELL_X32 FILLER_449_2591 ();
 FILLCELL_X32 FILLER_449_2623 ();
 FILLCELL_X32 FILLER_449_2655 ();
 FILLCELL_X32 FILLER_449_2687 ();
 FILLCELL_X32 FILLER_449_2719 ();
 FILLCELL_X32 FILLER_449_2751 ();
 FILLCELL_X32 FILLER_449_2783 ();
 FILLCELL_X32 FILLER_449_2815 ();
 FILLCELL_X32 FILLER_449_2847 ();
 FILLCELL_X32 FILLER_449_2879 ();
 FILLCELL_X32 FILLER_449_2911 ();
 FILLCELL_X32 FILLER_449_2943 ();
 FILLCELL_X32 FILLER_449_2975 ();
 FILLCELL_X32 FILLER_449_3007 ();
 FILLCELL_X32 FILLER_449_3039 ();
 FILLCELL_X32 FILLER_449_3071 ();
 FILLCELL_X32 FILLER_449_3103 ();
 FILLCELL_X32 FILLER_449_3135 ();
 FILLCELL_X32 FILLER_449_3167 ();
 FILLCELL_X32 FILLER_449_3199 ();
 FILLCELL_X32 FILLER_449_3231 ();
 FILLCELL_X32 FILLER_449_3263 ();
 FILLCELL_X32 FILLER_449_3295 ();
 FILLCELL_X32 FILLER_449_3327 ();
 FILLCELL_X32 FILLER_449_3359 ();
 FILLCELL_X32 FILLER_449_3391 ();
 FILLCELL_X32 FILLER_449_3423 ();
 FILLCELL_X32 FILLER_449_3455 ();
 FILLCELL_X32 FILLER_449_3487 ();
 FILLCELL_X32 FILLER_449_3519 ();
 FILLCELL_X32 FILLER_449_3551 ();
 FILLCELL_X32 FILLER_449_3583 ();
 FILLCELL_X32 FILLER_449_3615 ();
 FILLCELL_X32 FILLER_449_3647 ();
 FILLCELL_X32 FILLER_449_3679 ();
 FILLCELL_X16 FILLER_449_3711 ();
 FILLCELL_X8 FILLER_449_3727 ();
 FILLCELL_X2 FILLER_449_3735 ();
 FILLCELL_X1 FILLER_449_3737 ();
 FILLCELL_X32 FILLER_450_1 ();
 FILLCELL_X32 FILLER_450_33 ();
 FILLCELL_X32 FILLER_450_65 ();
 FILLCELL_X32 FILLER_450_97 ();
 FILLCELL_X32 FILLER_450_129 ();
 FILLCELL_X32 FILLER_450_161 ();
 FILLCELL_X32 FILLER_450_193 ();
 FILLCELL_X32 FILLER_450_225 ();
 FILLCELL_X32 FILLER_450_257 ();
 FILLCELL_X32 FILLER_450_289 ();
 FILLCELL_X32 FILLER_450_321 ();
 FILLCELL_X32 FILLER_450_353 ();
 FILLCELL_X32 FILLER_450_385 ();
 FILLCELL_X32 FILLER_450_417 ();
 FILLCELL_X32 FILLER_450_449 ();
 FILLCELL_X32 FILLER_450_481 ();
 FILLCELL_X32 FILLER_450_513 ();
 FILLCELL_X32 FILLER_450_545 ();
 FILLCELL_X32 FILLER_450_577 ();
 FILLCELL_X16 FILLER_450_609 ();
 FILLCELL_X4 FILLER_450_625 ();
 FILLCELL_X2 FILLER_450_629 ();
 FILLCELL_X32 FILLER_450_632 ();
 FILLCELL_X32 FILLER_450_664 ();
 FILLCELL_X32 FILLER_450_696 ();
 FILLCELL_X32 FILLER_450_728 ();
 FILLCELL_X32 FILLER_450_760 ();
 FILLCELL_X32 FILLER_450_792 ();
 FILLCELL_X32 FILLER_450_824 ();
 FILLCELL_X32 FILLER_450_856 ();
 FILLCELL_X32 FILLER_450_888 ();
 FILLCELL_X32 FILLER_450_920 ();
 FILLCELL_X32 FILLER_450_952 ();
 FILLCELL_X32 FILLER_450_984 ();
 FILLCELL_X32 FILLER_450_1016 ();
 FILLCELL_X32 FILLER_450_1048 ();
 FILLCELL_X32 FILLER_450_1080 ();
 FILLCELL_X32 FILLER_450_1112 ();
 FILLCELL_X32 FILLER_450_1144 ();
 FILLCELL_X32 FILLER_450_1176 ();
 FILLCELL_X32 FILLER_450_1208 ();
 FILLCELL_X32 FILLER_450_1240 ();
 FILLCELL_X32 FILLER_450_1272 ();
 FILLCELL_X32 FILLER_450_1304 ();
 FILLCELL_X32 FILLER_450_1336 ();
 FILLCELL_X32 FILLER_450_1368 ();
 FILLCELL_X32 FILLER_450_1400 ();
 FILLCELL_X32 FILLER_450_1432 ();
 FILLCELL_X32 FILLER_450_1464 ();
 FILLCELL_X32 FILLER_450_1496 ();
 FILLCELL_X32 FILLER_450_1528 ();
 FILLCELL_X32 FILLER_450_1560 ();
 FILLCELL_X32 FILLER_450_1592 ();
 FILLCELL_X32 FILLER_450_1624 ();
 FILLCELL_X32 FILLER_450_1656 ();
 FILLCELL_X32 FILLER_450_1688 ();
 FILLCELL_X32 FILLER_450_1720 ();
 FILLCELL_X32 FILLER_450_1752 ();
 FILLCELL_X32 FILLER_450_1784 ();
 FILLCELL_X32 FILLER_450_1816 ();
 FILLCELL_X32 FILLER_450_1848 ();
 FILLCELL_X8 FILLER_450_1880 ();
 FILLCELL_X4 FILLER_450_1888 ();
 FILLCELL_X2 FILLER_450_1892 ();
 FILLCELL_X32 FILLER_450_1895 ();
 FILLCELL_X32 FILLER_450_1927 ();
 FILLCELL_X32 FILLER_450_1959 ();
 FILLCELL_X32 FILLER_450_1991 ();
 FILLCELL_X32 FILLER_450_2023 ();
 FILLCELL_X32 FILLER_450_2055 ();
 FILLCELL_X32 FILLER_450_2087 ();
 FILLCELL_X32 FILLER_450_2119 ();
 FILLCELL_X32 FILLER_450_2151 ();
 FILLCELL_X32 FILLER_450_2183 ();
 FILLCELL_X32 FILLER_450_2215 ();
 FILLCELL_X32 FILLER_450_2247 ();
 FILLCELL_X32 FILLER_450_2279 ();
 FILLCELL_X32 FILLER_450_2311 ();
 FILLCELL_X32 FILLER_450_2343 ();
 FILLCELL_X32 FILLER_450_2375 ();
 FILLCELL_X32 FILLER_450_2407 ();
 FILLCELL_X32 FILLER_450_2439 ();
 FILLCELL_X32 FILLER_450_2471 ();
 FILLCELL_X32 FILLER_450_2503 ();
 FILLCELL_X32 FILLER_450_2535 ();
 FILLCELL_X32 FILLER_450_2567 ();
 FILLCELL_X32 FILLER_450_2599 ();
 FILLCELL_X32 FILLER_450_2631 ();
 FILLCELL_X32 FILLER_450_2663 ();
 FILLCELL_X32 FILLER_450_2695 ();
 FILLCELL_X32 FILLER_450_2727 ();
 FILLCELL_X32 FILLER_450_2759 ();
 FILLCELL_X32 FILLER_450_2791 ();
 FILLCELL_X32 FILLER_450_2823 ();
 FILLCELL_X32 FILLER_450_2855 ();
 FILLCELL_X32 FILLER_450_2887 ();
 FILLCELL_X32 FILLER_450_2919 ();
 FILLCELL_X32 FILLER_450_2951 ();
 FILLCELL_X32 FILLER_450_2983 ();
 FILLCELL_X32 FILLER_450_3015 ();
 FILLCELL_X32 FILLER_450_3047 ();
 FILLCELL_X32 FILLER_450_3079 ();
 FILLCELL_X32 FILLER_450_3111 ();
 FILLCELL_X8 FILLER_450_3143 ();
 FILLCELL_X4 FILLER_450_3151 ();
 FILLCELL_X2 FILLER_450_3155 ();
 FILLCELL_X32 FILLER_450_3158 ();
 FILLCELL_X32 FILLER_450_3190 ();
 FILLCELL_X32 FILLER_450_3222 ();
 FILLCELL_X32 FILLER_450_3254 ();
 FILLCELL_X32 FILLER_450_3286 ();
 FILLCELL_X32 FILLER_450_3318 ();
 FILLCELL_X32 FILLER_450_3350 ();
 FILLCELL_X32 FILLER_450_3382 ();
 FILLCELL_X32 FILLER_450_3414 ();
 FILLCELL_X32 FILLER_450_3446 ();
 FILLCELL_X32 FILLER_450_3478 ();
 FILLCELL_X32 FILLER_450_3510 ();
 FILLCELL_X32 FILLER_450_3542 ();
 FILLCELL_X32 FILLER_450_3574 ();
 FILLCELL_X32 FILLER_450_3606 ();
 FILLCELL_X32 FILLER_450_3638 ();
 FILLCELL_X32 FILLER_450_3670 ();
 FILLCELL_X32 FILLER_450_3702 ();
 FILLCELL_X4 FILLER_450_3734 ();
 FILLCELL_X32 FILLER_451_1 ();
 FILLCELL_X32 FILLER_451_33 ();
 FILLCELL_X32 FILLER_451_65 ();
 FILLCELL_X32 FILLER_451_97 ();
 FILLCELL_X32 FILLER_451_129 ();
 FILLCELL_X32 FILLER_451_161 ();
 FILLCELL_X32 FILLER_451_193 ();
 FILLCELL_X32 FILLER_451_225 ();
 FILLCELL_X32 FILLER_451_257 ();
 FILLCELL_X32 FILLER_451_289 ();
 FILLCELL_X32 FILLER_451_321 ();
 FILLCELL_X32 FILLER_451_353 ();
 FILLCELL_X32 FILLER_451_385 ();
 FILLCELL_X32 FILLER_451_417 ();
 FILLCELL_X32 FILLER_451_449 ();
 FILLCELL_X32 FILLER_451_481 ();
 FILLCELL_X32 FILLER_451_513 ();
 FILLCELL_X32 FILLER_451_545 ();
 FILLCELL_X32 FILLER_451_577 ();
 FILLCELL_X32 FILLER_451_609 ();
 FILLCELL_X32 FILLER_451_641 ();
 FILLCELL_X32 FILLER_451_673 ();
 FILLCELL_X32 FILLER_451_705 ();
 FILLCELL_X32 FILLER_451_737 ();
 FILLCELL_X32 FILLER_451_769 ();
 FILLCELL_X32 FILLER_451_801 ();
 FILLCELL_X32 FILLER_451_833 ();
 FILLCELL_X32 FILLER_451_865 ();
 FILLCELL_X32 FILLER_451_897 ();
 FILLCELL_X32 FILLER_451_929 ();
 FILLCELL_X32 FILLER_451_961 ();
 FILLCELL_X32 FILLER_451_993 ();
 FILLCELL_X32 FILLER_451_1025 ();
 FILLCELL_X32 FILLER_451_1057 ();
 FILLCELL_X32 FILLER_451_1089 ();
 FILLCELL_X32 FILLER_451_1121 ();
 FILLCELL_X32 FILLER_451_1153 ();
 FILLCELL_X32 FILLER_451_1185 ();
 FILLCELL_X32 FILLER_451_1217 ();
 FILLCELL_X8 FILLER_451_1249 ();
 FILLCELL_X4 FILLER_451_1257 ();
 FILLCELL_X2 FILLER_451_1261 ();
 FILLCELL_X32 FILLER_451_1264 ();
 FILLCELL_X32 FILLER_451_1296 ();
 FILLCELL_X32 FILLER_451_1328 ();
 FILLCELL_X32 FILLER_451_1360 ();
 FILLCELL_X32 FILLER_451_1392 ();
 FILLCELL_X32 FILLER_451_1424 ();
 FILLCELL_X32 FILLER_451_1456 ();
 FILLCELL_X32 FILLER_451_1488 ();
 FILLCELL_X32 FILLER_451_1520 ();
 FILLCELL_X32 FILLER_451_1552 ();
 FILLCELL_X32 FILLER_451_1584 ();
 FILLCELL_X32 FILLER_451_1616 ();
 FILLCELL_X32 FILLER_451_1648 ();
 FILLCELL_X32 FILLER_451_1680 ();
 FILLCELL_X32 FILLER_451_1712 ();
 FILLCELL_X32 FILLER_451_1744 ();
 FILLCELL_X32 FILLER_451_1776 ();
 FILLCELL_X32 FILLER_451_1808 ();
 FILLCELL_X32 FILLER_451_1840 ();
 FILLCELL_X32 FILLER_451_1872 ();
 FILLCELL_X32 FILLER_451_1904 ();
 FILLCELL_X32 FILLER_451_1936 ();
 FILLCELL_X32 FILLER_451_1968 ();
 FILLCELL_X32 FILLER_451_2000 ();
 FILLCELL_X32 FILLER_451_2032 ();
 FILLCELL_X32 FILLER_451_2064 ();
 FILLCELL_X32 FILLER_451_2096 ();
 FILLCELL_X32 FILLER_451_2128 ();
 FILLCELL_X32 FILLER_451_2160 ();
 FILLCELL_X32 FILLER_451_2192 ();
 FILLCELL_X32 FILLER_451_2224 ();
 FILLCELL_X32 FILLER_451_2256 ();
 FILLCELL_X32 FILLER_451_2288 ();
 FILLCELL_X32 FILLER_451_2320 ();
 FILLCELL_X32 FILLER_451_2352 ();
 FILLCELL_X32 FILLER_451_2384 ();
 FILLCELL_X32 FILLER_451_2416 ();
 FILLCELL_X32 FILLER_451_2448 ();
 FILLCELL_X32 FILLER_451_2480 ();
 FILLCELL_X8 FILLER_451_2512 ();
 FILLCELL_X4 FILLER_451_2520 ();
 FILLCELL_X2 FILLER_451_2524 ();
 FILLCELL_X32 FILLER_451_2527 ();
 FILLCELL_X32 FILLER_451_2559 ();
 FILLCELL_X32 FILLER_451_2591 ();
 FILLCELL_X32 FILLER_451_2623 ();
 FILLCELL_X32 FILLER_451_2655 ();
 FILLCELL_X32 FILLER_451_2687 ();
 FILLCELL_X32 FILLER_451_2719 ();
 FILLCELL_X32 FILLER_451_2751 ();
 FILLCELL_X32 FILLER_451_2783 ();
 FILLCELL_X32 FILLER_451_2815 ();
 FILLCELL_X32 FILLER_451_2847 ();
 FILLCELL_X32 FILLER_451_2879 ();
 FILLCELL_X32 FILLER_451_2911 ();
 FILLCELL_X32 FILLER_451_2943 ();
 FILLCELL_X32 FILLER_451_2975 ();
 FILLCELL_X32 FILLER_451_3007 ();
 FILLCELL_X32 FILLER_451_3039 ();
 FILLCELL_X32 FILLER_451_3071 ();
 FILLCELL_X32 FILLER_451_3103 ();
 FILLCELL_X32 FILLER_451_3135 ();
 FILLCELL_X32 FILLER_451_3167 ();
 FILLCELL_X32 FILLER_451_3199 ();
 FILLCELL_X32 FILLER_451_3231 ();
 FILLCELL_X32 FILLER_451_3263 ();
 FILLCELL_X32 FILLER_451_3295 ();
 FILLCELL_X32 FILLER_451_3327 ();
 FILLCELL_X32 FILLER_451_3359 ();
 FILLCELL_X32 FILLER_451_3391 ();
 FILLCELL_X32 FILLER_451_3423 ();
 FILLCELL_X32 FILLER_451_3455 ();
 FILLCELL_X32 FILLER_451_3487 ();
 FILLCELL_X32 FILLER_451_3519 ();
 FILLCELL_X32 FILLER_451_3551 ();
 FILLCELL_X32 FILLER_451_3583 ();
 FILLCELL_X32 FILLER_451_3615 ();
 FILLCELL_X32 FILLER_451_3647 ();
 FILLCELL_X32 FILLER_451_3679 ();
 FILLCELL_X16 FILLER_451_3711 ();
 FILLCELL_X8 FILLER_451_3727 ();
 FILLCELL_X2 FILLER_451_3735 ();
 FILLCELL_X1 FILLER_451_3737 ();
 FILLCELL_X32 FILLER_452_1 ();
 FILLCELL_X32 FILLER_452_33 ();
 FILLCELL_X32 FILLER_452_65 ();
 FILLCELL_X32 FILLER_452_97 ();
 FILLCELL_X32 FILLER_452_129 ();
 FILLCELL_X32 FILLER_452_161 ();
 FILLCELL_X32 FILLER_452_193 ();
 FILLCELL_X32 FILLER_452_225 ();
 FILLCELL_X32 FILLER_452_257 ();
 FILLCELL_X32 FILLER_452_289 ();
 FILLCELL_X32 FILLER_452_321 ();
 FILLCELL_X32 FILLER_452_353 ();
 FILLCELL_X32 FILLER_452_385 ();
 FILLCELL_X32 FILLER_452_417 ();
 FILLCELL_X32 FILLER_452_449 ();
 FILLCELL_X32 FILLER_452_481 ();
 FILLCELL_X32 FILLER_452_513 ();
 FILLCELL_X32 FILLER_452_545 ();
 FILLCELL_X32 FILLER_452_577 ();
 FILLCELL_X16 FILLER_452_609 ();
 FILLCELL_X4 FILLER_452_625 ();
 FILLCELL_X2 FILLER_452_629 ();
 FILLCELL_X32 FILLER_452_632 ();
 FILLCELL_X32 FILLER_452_664 ();
 FILLCELL_X32 FILLER_452_696 ();
 FILLCELL_X32 FILLER_452_728 ();
 FILLCELL_X32 FILLER_452_760 ();
 FILLCELL_X32 FILLER_452_792 ();
 FILLCELL_X32 FILLER_452_824 ();
 FILLCELL_X32 FILLER_452_856 ();
 FILLCELL_X32 FILLER_452_888 ();
 FILLCELL_X32 FILLER_452_920 ();
 FILLCELL_X32 FILLER_452_952 ();
 FILLCELL_X32 FILLER_452_984 ();
 FILLCELL_X32 FILLER_452_1016 ();
 FILLCELL_X32 FILLER_452_1048 ();
 FILLCELL_X32 FILLER_452_1080 ();
 FILLCELL_X32 FILLER_452_1112 ();
 FILLCELL_X32 FILLER_452_1144 ();
 FILLCELL_X32 FILLER_452_1176 ();
 FILLCELL_X32 FILLER_452_1208 ();
 FILLCELL_X32 FILLER_452_1240 ();
 FILLCELL_X32 FILLER_452_1272 ();
 FILLCELL_X32 FILLER_452_1304 ();
 FILLCELL_X32 FILLER_452_1336 ();
 FILLCELL_X32 FILLER_452_1368 ();
 FILLCELL_X32 FILLER_452_1400 ();
 FILLCELL_X32 FILLER_452_1432 ();
 FILLCELL_X32 FILLER_452_1464 ();
 FILLCELL_X32 FILLER_452_1496 ();
 FILLCELL_X32 FILLER_452_1528 ();
 FILLCELL_X32 FILLER_452_1560 ();
 FILLCELL_X32 FILLER_452_1592 ();
 FILLCELL_X32 FILLER_452_1624 ();
 FILLCELL_X32 FILLER_452_1656 ();
 FILLCELL_X32 FILLER_452_1688 ();
 FILLCELL_X32 FILLER_452_1720 ();
 FILLCELL_X32 FILLER_452_1752 ();
 FILLCELL_X32 FILLER_452_1784 ();
 FILLCELL_X32 FILLER_452_1816 ();
 FILLCELL_X32 FILLER_452_1848 ();
 FILLCELL_X8 FILLER_452_1880 ();
 FILLCELL_X4 FILLER_452_1888 ();
 FILLCELL_X2 FILLER_452_1892 ();
 FILLCELL_X32 FILLER_452_1895 ();
 FILLCELL_X32 FILLER_452_1927 ();
 FILLCELL_X32 FILLER_452_1959 ();
 FILLCELL_X32 FILLER_452_1991 ();
 FILLCELL_X32 FILLER_452_2023 ();
 FILLCELL_X32 FILLER_452_2055 ();
 FILLCELL_X32 FILLER_452_2087 ();
 FILLCELL_X32 FILLER_452_2119 ();
 FILLCELL_X32 FILLER_452_2151 ();
 FILLCELL_X32 FILLER_452_2183 ();
 FILLCELL_X32 FILLER_452_2215 ();
 FILLCELL_X32 FILLER_452_2247 ();
 FILLCELL_X32 FILLER_452_2279 ();
 FILLCELL_X32 FILLER_452_2311 ();
 FILLCELL_X32 FILLER_452_2343 ();
 FILLCELL_X32 FILLER_452_2375 ();
 FILLCELL_X32 FILLER_452_2407 ();
 FILLCELL_X32 FILLER_452_2439 ();
 FILLCELL_X32 FILLER_452_2471 ();
 FILLCELL_X32 FILLER_452_2503 ();
 FILLCELL_X32 FILLER_452_2535 ();
 FILLCELL_X32 FILLER_452_2567 ();
 FILLCELL_X32 FILLER_452_2599 ();
 FILLCELL_X32 FILLER_452_2631 ();
 FILLCELL_X32 FILLER_452_2663 ();
 FILLCELL_X32 FILLER_452_2695 ();
 FILLCELL_X32 FILLER_452_2727 ();
 FILLCELL_X32 FILLER_452_2759 ();
 FILLCELL_X32 FILLER_452_2791 ();
 FILLCELL_X32 FILLER_452_2823 ();
 FILLCELL_X32 FILLER_452_2855 ();
 FILLCELL_X32 FILLER_452_2887 ();
 FILLCELL_X32 FILLER_452_2919 ();
 FILLCELL_X32 FILLER_452_2951 ();
 FILLCELL_X32 FILLER_452_2983 ();
 FILLCELL_X32 FILLER_452_3015 ();
 FILLCELL_X32 FILLER_452_3047 ();
 FILLCELL_X32 FILLER_452_3079 ();
 FILLCELL_X32 FILLER_452_3111 ();
 FILLCELL_X8 FILLER_452_3143 ();
 FILLCELL_X4 FILLER_452_3151 ();
 FILLCELL_X2 FILLER_452_3155 ();
 FILLCELL_X32 FILLER_452_3158 ();
 FILLCELL_X32 FILLER_452_3190 ();
 FILLCELL_X32 FILLER_452_3222 ();
 FILLCELL_X32 FILLER_452_3254 ();
 FILLCELL_X32 FILLER_452_3286 ();
 FILLCELL_X32 FILLER_452_3318 ();
 FILLCELL_X32 FILLER_452_3350 ();
 FILLCELL_X32 FILLER_452_3382 ();
 FILLCELL_X32 FILLER_452_3414 ();
 FILLCELL_X32 FILLER_452_3446 ();
 FILLCELL_X32 FILLER_452_3478 ();
 FILLCELL_X32 FILLER_452_3510 ();
 FILLCELL_X32 FILLER_452_3542 ();
 FILLCELL_X32 FILLER_452_3574 ();
 FILLCELL_X32 FILLER_452_3606 ();
 FILLCELL_X32 FILLER_452_3638 ();
 FILLCELL_X32 FILLER_452_3670 ();
 FILLCELL_X32 FILLER_452_3702 ();
 FILLCELL_X4 FILLER_452_3734 ();
 FILLCELL_X32 FILLER_453_1 ();
 FILLCELL_X32 FILLER_453_33 ();
 FILLCELL_X32 FILLER_453_65 ();
 FILLCELL_X32 FILLER_453_97 ();
 FILLCELL_X32 FILLER_453_129 ();
 FILLCELL_X32 FILLER_453_161 ();
 FILLCELL_X32 FILLER_453_193 ();
 FILLCELL_X32 FILLER_453_225 ();
 FILLCELL_X32 FILLER_453_257 ();
 FILLCELL_X32 FILLER_453_289 ();
 FILLCELL_X32 FILLER_453_321 ();
 FILLCELL_X32 FILLER_453_353 ();
 FILLCELL_X32 FILLER_453_385 ();
 FILLCELL_X32 FILLER_453_417 ();
 FILLCELL_X32 FILLER_453_449 ();
 FILLCELL_X32 FILLER_453_481 ();
 FILLCELL_X32 FILLER_453_513 ();
 FILLCELL_X32 FILLER_453_545 ();
 FILLCELL_X32 FILLER_453_577 ();
 FILLCELL_X32 FILLER_453_609 ();
 FILLCELL_X32 FILLER_453_641 ();
 FILLCELL_X32 FILLER_453_673 ();
 FILLCELL_X32 FILLER_453_705 ();
 FILLCELL_X32 FILLER_453_737 ();
 FILLCELL_X32 FILLER_453_769 ();
 FILLCELL_X32 FILLER_453_801 ();
 FILLCELL_X32 FILLER_453_833 ();
 FILLCELL_X32 FILLER_453_865 ();
 FILLCELL_X32 FILLER_453_897 ();
 FILLCELL_X32 FILLER_453_929 ();
 FILLCELL_X32 FILLER_453_961 ();
 FILLCELL_X32 FILLER_453_993 ();
 FILLCELL_X32 FILLER_453_1025 ();
 FILLCELL_X32 FILLER_453_1057 ();
 FILLCELL_X32 FILLER_453_1089 ();
 FILLCELL_X32 FILLER_453_1121 ();
 FILLCELL_X32 FILLER_453_1153 ();
 FILLCELL_X32 FILLER_453_1185 ();
 FILLCELL_X32 FILLER_453_1217 ();
 FILLCELL_X8 FILLER_453_1249 ();
 FILLCELL_X4 FILLER_453_1257 ();
 FILLCELL_X2 FILLER_453_1261 ();
 FILLCELL_X32 FILLER_453_1264 ();
 FILLCELL_X32 FILLER_453_1296 ();
 FILLCELL_X32 FILLER_453_1328 ();
 FILLCELL_X32 FILLER_453_1360 ();
 FILLCELL_X32 FILLER_453_1392 ();
 FILLCELL_X32 FILLER_453_1424 ();
 FILLCELL_X32 FILLER_453_1456 ();
 FILLCELL_X32 FILLER_453_1488 ();
 FILLCELL_X32 FILLER_453_1520 ();
 FILLCELL_X32 FILLER_453_1552 ();
 FILLCELL_X32 FILLER_453_1584 ();
 FILLCELL_X32 FILLER_453_1616 ();
 FILLCELL_X32 FILLER_453_1648 ();
 FILLCELL_X32 FILLER_453_1680 ();
 FILLCELL_X32 FILLER_453_1712 ();
 FILLCELL_X32 FILLER_453_1744 ();
 FILLCELL_X32 FILLER_453_1776 ();
 FILLCELL_X32 FILLER_453_1808 ();
 FILLCELL_X32 FILLER_453_1840 ();
 FILLCELL_X32 FILLER_453_1872 ();
 FILLCELL_X32 FILLER_453_1904 ();
 FILLCELL_X32 FILLER_453_1936 ();
 FILLCELL_X32 FILLER_453_1968 ();
 FILLCELL_X32 FILLER_453_2000 ();
 FILLCELL_X32 FILLER_453_2032 ();
 FILLCELL_X32 FILLER_453_2064 ();
 FILLCELL_X32 FILLER_453_2096 ();
 FILLCELL_X32 FILLER_453_2128 ();
 FILLCELL_X32 FILLER_453_2160 ();
 FILLCELL_X32 FILLER_453_2192 ();
 FILLCELL_X32 FILLER_453_2224 ();
 FILLCELL_X32 FILLER_453_2256 ();
 FILLCELL_X32 FILLER_453_2288 ();
 FILLCELL_X32 FILLER_453_2320 ();
 FILLCELL_X32 FILLER_453_2352 ();
 FILLCELL_X32 FILLER_453_2384 ();
 FILLCELL_X32 FILLER_453_2416 ();
 FILLCELL_X32 FILLER_453_2448 ();
 FILLCELL_X32 FILLER_453_2480 ();
 FILLCELL_X8 FILLER_453_2512 ();
 FILLCELL_X4 FILLER_453_2520 ();
 FILLCELL_X2 FILLER_453_2524 ();
 FILLCELL_X32 FILLER_453_2527 ();
 FILLCELL_X32 FILLER_453_2559 ();
 FILLCELL_X32 FILLER_453_2591 ();
 FILLCELL_X32 FILLER_453_2623 ();
 FILLCELL_X32 FILLER_453_2655 ();
 FILLCELL_X32 FILLER_453_2687 ();
 FILLCELL_X32 FILLER_453_2719 ();
 FILLCELL_X32 FILLER_453_2751 ();
 FILLCELL_X32 FILLER_453_2783 ();
 FILLCELL_X32 FILLER_453_2815 ();
 FILLCELL_X32 FILLER_453_2847 ();
 FILLCELL_X32 FILLER_453_2879 ();
 FILLCELL_X32 FILLER_453_2911 ();
 FILLCELL_X32 FILLER_453_2943 ();
 FILLCELL_X32 FILLER_453_2975 ();
 FILLCELL_X32 FILLER_453_3007 ();
 FILLCELL_X32 FILLER_453_3039 ();
 FILLCELL_X32 FILLER_453_3071 ();
 FILLCELL_X32 FILLER_453_3103 ();
 FILLCELL_X32 FILLER_453_3135 ();
 FILLCELL_X32 FILLER_453_3167 ();
 FILLCELL_X32 FILLER_453_3199 ();
 FILLCELL_X32 FILLER_453_3231 ();
 FILLCELL_X32 FILLER_453_3263 ();
 FILLCELL_X32 FILLER_453_3295 ();
 FILLCELL_X32 FILLER_453_3327 ();
 FILLCELL_X32 FILLER_453_3359 ();
 FILLCELL_X32 FILLER_453_3391 ();
 FILLCELL_X32 FILLER_453_3423 ();
 FILLCELL_X32 FILLER_453_3455 ();
 FILLCELL_X32 FILLER_453_3487 ();
 FILLCELL_X32 FILLER_453_3519 ();
 FILLCELL_X32 FILLER_453_3551 ();
 FILLCELL_X32 FILLER_453_3583 ();
 FILLCELL_X32 FILLER_453_3615 ();
 FILLCELL_X32 FILLER_453_3647 ();
 FILLCELL_X32 FILLER_453_3679 ();
 FILLCELL_X16 FILLER_453_3711 ();
 FILLCELL_X8 FILLER_453_3727 ();
 FILLCELL_X2 FILLER_453_3735 ();
 FILLCELL_X1 FILLER_453_3737 ();
 FILLCELL_X32 FILLER_454_1 ();
 FILLCELL_X32 FILLER_454_33 ();
 FILLCELL_X32 FILLER_454_65 ();
 FILLCELL_X32 FILLER_454_97 ();
 FILLCELL_X32 FILLER_454_129 ();
 FILLCELL_X32 FILLER_454_161 ();
 FILLCELL_X32 FILLER_454_193 ();
 FILLCELL_X32 FILLER_454_225 ();
 FILLCELL_X32 FILLER_454_257 ();
 FILLCELL_X32 FILLER_454_289 ();
 FILLCELL_X32 FILLER_454_321 ();
 FILLCELL_X32 FILLER_454_353 ();
 FILLCELL_X32 FILLER_454_385 ();
 FILLCELL_X32 FILLER_454_417 ();
 FILLCELL_X32 FILLER_454_449 ();
 FILLCELL_X32 FILLER_454_481 ();
 FILLCELL_X32 FILLER_454_513 ();
 FILLCELL_X32 FILLER_454_545 ();
 FILLCELL_X32 FILLER_454_577 ();
 FILLCELL_X16 FILLER_454_609 ();
 FILLCELL_X4 FILLER_454_625 ();
 FILLCELL_X2 FILLER_454_629 ();
 FILLCELL_X32 FILLER_454_632 ();
 FILLCELL_X32 FILLER_454_664 ();
 FILLCELL_X32 FILLER_454_696 ();
 FILLCELL_X32 FILLER_454_728 ();
 FILLCELL_X32 FILLER_454_760 ();
 FILLCELL_X32 FILLER_454_792 ();
 FILLCELL_X32 FILLER_454_824 ();
 FILLCELL_X32 FILLER_454_856 ();
 FILLCELL_X32 FILLER_454_888 ();
 FILLCELL_X32 FILLER_454_920 ();
 FILLCELL_X32 FILLER_454_952 ();
 FILLCELL_X32 FILLER_454_984 ();
 FILLCELL_X32 FILLER_454_1016 ();
 FILLCELL_X32 FILLER_454_1048 ();
 FILLCELL_X32 FILLER_454_1080 ();
 FILLCELL_X32 FILLER_454_1112 ();
 FILLCELL_X32 FILLER_454_1144 ();
 FILLCELL_X32 FILLER_454_1176 ();
 FILLCELL_X32 FILLER_454_1208 ();
 FILLCELL_X32 FILLER_454_1240 ();
 FILLCELL_X32 FILLER_454_1272 ();
 FILLCELL_X32 FILLER_454_1304 ();
 FILLCELL_X32 FILLER_454_1336 ();
 FILLCELL_X32 FILLER_454_1368 ();
 FILLCELL_X32 FILLER_454_1400 ();
 FILLCELL_X32 FILLER_454_1432 ();
 FILLCELL_X32 FILLER_454_1464 ();
 FILLCELL_X32 FILLER_454_1496 ();
 FILLCELL_X32 FILLER_454_1528 ();
 FILLCELL_X32 FILLER_454_1560 ();
 FILLCELL_X32 FILLER_454_1592 ();
 FILLCELL_X32 FILLER_454_1624 ();
 FILLCELL_X32 FILLER_454_1656 ();
 FILLCELL_X32 FILLER_454_1688 ();
 FILLCELL_X32 FILLER_454_1720 ();
 FILLCELL_X32 FILLER_454_1752 ();
 FILLCELL_X32 FILLER_454_1784 ();
 FILLCELL_X32 FILLER_454_1816 ();
 FILLCELL_X32 FILLER_454_1848 ();
 FILLCELL_X8 FILLER_454_1880 ();
 FILLCELL_X4 FILLER_454_1888 ();
 FILLCELL_X2 FILLER_454_1892 ();
 FILLCELL_X32 FILLER_454_1895 ();
 FILLCELL_X32 FILLER_454_1927 ();
 FILLCELL_X32 FILLER_454_1959 ();
 FILLCELL_X32 FILLER_454_1991 ();
 FILLCELL_X32 FILLER_454_2023 ();
 FILLCELL_X32 FILLER_454_2055 ();
 FILLCELL_X32 FILLER_454_2087 ();
 FILLCELL_X32 FILLER_454_2119 ();
 FILLCELL_X32 FILLER_454_2151 ();
 FILLCELL_X32 FILLER_454_2183 ();
 FILLCELL_X32 FILLER_454_2215 ();
 FILLCELL_X32 FILLER_454_2247 ();
 FILLCELL_X32 FILLER_454_2279 ();
 FILLCELL_X32 FILLER_454_2311 ();
 FILLCELL_X32 FILLER_454_2343 ();
 FILLCELL_X32 FILLER_454_2375 ();
 FILLCELL_X32 FILLER_454_2407 ();
 FILLCELL_X32 FILLER_454_2439 ();
 FILLCELL_X32 FILLER_454_2471 ();
 FILLCELL_X32 FILLER_454_2503 ();
 FILLCELL_X32 FILLER_454_2535 ();
 FILLCELL_X32 FILLER_454_2567 ();
 FILLCELL_X32 FILLER_454_2599 ();
 FILLCELL_X32 FILLER_454_2631 ();
 FILLCELL_X32 FILLER_454_2663 ();
 FILLCELL_X32 FILLER_454_2695 ();
 FILLCELL_X32 FILLER_454_2727 ();
 FILLCELL_X32 FILLER_454_2759 ();
 FILLCELL_X32 FILLER_454_2791 ();
 FILLCELL_X32 FILLER_454_2823 ();
 FILLCELL_X32 FILLER_454_2855 ();
 FILLCELL_X32 FILLER_454_2887 ();
 FILLCELL_X32 FILLER_454_2919 ();
 FILLCELL_X32 FILLER_454_2951 ();
 FILLCELL_X32 FILLER_454_2983 ();
 FILLCELL_X32 FILLER_454_3015 ();
 FILLCELL_X32 FILLER_454_3047 ();
 FILLCELL_X32 FILLER_454_3079 ();
 FILLCELL_X32 FILLER_454_3111 ();
 FILLCELL_X8 FILLER_454_3143 ();
 FILLCELL_X4 FILLER_454_3151 ();
 FILLCELL_X2 FILLER_454_3155 ();
 FILLCELL_X32 FILLER_454_3158 ();
 FILLCELL_X32 FILLER_454_3190 ();
 FILLCELL_X32 FILLER_454_3222 ();
 FILLCELL_X32 FILLER_454_3254 ();
 FILLCELL_X32 FILLER_454_3286 ();
 FILLCELL_X32 FILLER_454_3318 ();
 FILLCELL_X32 FILLER_454_3350 ();
 FILLCELL_X32 FILLER_454_3382 ();
 FILLCELL_X32 FILLER_454_3414 ();
 FILLCELL_X32 FILLER_454_3446 ();
 FILLCELL_X32 FILLER_454_3478 ();
 FILLCELL_X32 FILLER_454_3510 ();
 FILLCELL_X32 FILLER_454_3542 ();
 FILLCELL_X32 FILLER_454_3574 ();
 FILLCELL_X32 FILLER_454_3606 ();
 FILLCELL_X32 FILLER_454_3638 ();
 FILLCELL_X32 FILLER_454_3670 ();
 FILLCELL_X32 FILLER_454_3702 ();
 FILLCELL_X4 FILLER_454_3734 ();
 FILLCELL_X32 FILLER_455_1 ();
 FILLCELL_X32 FILLER_455_33 ();
 FILLCELL_X32 FILLER_455_65 ();
 FILLCELL_X32 FILLER_455_97 ();
 FILLCELL_X32 FILLER_455_129 ();
 FILLCELL_X32 FILLER_455_161 ();
 FILLCELL_X32 FILLER_455_193 ();
 FILLCELL_X32 FILLER_455_225 ();
 FILLCELL_X32 FILLER_455_257 ();
 FILLCELL_X32 FILLER_455_289 ();
 FILLCELL_X32 FILLER_455_321 ();
 FILLCELL_X32 FILLER_455_353 ();
 FILLCELL_X32 FILLER_455_385 ();
 FILLCELL_X32 FILLER_455_417 ();
 FILLCELL_X32 FILLER_455_449 ();
 FILLCELL_X32 FILLER_455_481 ();
 FILLCELL_X32 FILLER_455_513 ();
 FILLCELL_X32 FILLER_455_545 ();
 FILLCELL_X32 FILLER_455_577 ();
 FILLCELL_X32 FILLER_455_609 ();
 FILLCELL_X32 FILLER_455_641 ();
 FILLCELL_X32 FILLER_455_673 ();
 FILLCELL_X32 FILLER_455_705 ();
 FILLCELL_X32 FILLER_455_737 ();
 FILLCELL_X32 FILLER_455_769 ();
 FILLCELL_X32 FILLER_455_801 ();
 FILLCELL_X32 FILLER_455_833 ();
 FILLCELL_X32 FILLER_455_865 ();
 FILLCELL_X32 FILLER_455_897 ();
 FILLCELL_X32 FILLER_455_929 ();
 FILLCELL_X32 FILLER_455_961 ();
 FILLCELL_X32 FILLER_455_993 ();
 FILLCELL_X32 FILLER_455_1025 ();
 FILLCELL_X32 FILLER_455_1057 ();
 FILLCELL_X32 FILLER_455_1089 ();
 FILLCELL_X32 FILLER_455_1121 ();
 FILLCELL_X32 FILLER_455_1153 ();
 FILLCELL_X32 FILLER_455_1185 ();
 FILLCELL_X32 FILLER_455_1217 ();
 FILLCELL_X8 FILLER_455_1249 ();
 FILLCELL_X4 FILLER_455_1257 ();
 FILLCELL_X2 FILLER_455_1261 ();
 FILLCELL_X32 FILLER_455_1264 ();
 FILLCELL_X32 FILLER_455_1296 ();
 FILLCELL_X32 FILLER_455_1328 ();
 FILLCELL_X32 FILLER_455_1360 ();
 FILLCELL_X32 FILLER_455_1392 ();
 FILLCELL_X32 FILLER_455_1424 ();
 FILLCELL_X32 FILLER_455_1456 ();
 FILLCELL_X32 FILLER_455_1488 ();
 FILLCELL_X32 FILLER_455_1520 ();
 FILLCELL_X32 FILLER_455_1552 ();
 FILLCELL_X32 FILLER_455_1584 ();
 FILLCELL_X32 FILLER_455_1616 ();
 FILLCELL_X32 FILLER_455_1648 ();
 FILLCELL_X32 FILLER_455_1680 ();
 FILLCELL_X32 FILLER_455_1712 ();
 FILLCELL_X32 FILLER_455_1744 ();
 FILLCELL_X32 FILLER_455_1776 ();
 FILLCELL_X32 FILLER_455_1808 ();
 FILLCELL_X32 FILLER_455_1840 ();
 FILLCELL_X32 FILLER_455_1872 ();
 FILLCELL_X32 FILLER_455_1904 ();
 FILLCELL_X32 FILLER_455_1936 ();
 FILLCELL_X32 FILLER_455_1968 ();
 FILLCELL_X32 FILLER_455_2000 ();
 FILLCELL_X32 FILLER_455_2032 ();
 FILLCELL_X32 FILLER_455_2064 ();
 FILLCELL_X32 FILLER_455_2096 ();
 FILLCELL_X32 FILLER_455_2128 ();
 FILLCELL_X32 FILLER_455_2160 ();
 FILLCELL_X32 FILLER_455_2192 ();
 FILLCELL_X32 FILLER_455_2224 ();
 FILLCELL_X32 FILLER_455_2256 ();
 FILLCELL_X32 FILLER_455_2288 ();
 FILLCELL_X32 FILLER_455_2320 ();
 FILLCELL_X32 FILLER_455_2352 ();
 FILLCELL_X32 FILLER_455_2384 ();
 FILLCELL_X32 FILLER_455_2416 ();
 FILLCELL_X32 FILLER_455_2448 ();
 FILLCELL_X32 FILLER_455_2480 ();
 FILLCELL_X8 FILLER_455_2512 ();
 FILLCELL_X4 FILLER_455_2520 ();
 FILLCELL_X2 FILLER_455_2524 ();
 FILLCELL_X32 FILLER_455_2527 ();
 FILLCELL_X32 FILLER_455_2559 ();
 FILLCELL_X32 FILLER_455_2591 ();
 FILLCELL_X32 FILLER_455_2623 ();
 FILLCELL_X32 FILLER_455_2655 ();
 FILLCELL_X32 FILLER_455_2687 ();
 FILLCELL_X32 FILLER_455_2719 ();
 FILLCELL_X32 FILLER_455_2751 ();
 FILLCELL_X32 FILLER_455_2783 ();
 FILLCELL_X32 FILLER_455_2815 ();
 FILLCELL_X32 FILLER_455_2847 ();
 FILLCELL_X32 FILLER_455_2879 ();
 FILLCELL_X32 FILLER_455_2911 ();
 FILLCELL_X32 FILLER_455_2943 ();
 FILLCELL_X32 FILLER_455_2975 ();
 FILLCELL_X32 FILLER_455_3007 ();
 FILLCELL_X32 FILLER_455_3039 ();
 FILLCELL_X32 FILLER_455_3071 ();
 FILLCELL_X32 FILLER_455_3103 ();
 FILLCELL_X32 FILLER_455_3135 ();
 FILLCELL_X32 FILLER_455_3167 ();
 FILLCELL_X32 FILLER_455_3199 ();
 FILLCELL_X32 FILLER_455_3231 ();
 FILLCELL_X32 FILLER_455_3263 ();
 FILLCELL_X32 FILLER_455_3295 ();
 FILLCELL_X32 FILLER_455_3327 ();
 FILLCELL_X32 FILLER_455_3359 ();
 FILLCELL_X32 FILLER_455_3391 ();
 FILLCELL_X32 FILLER_455_3423 ();
 FILLCELL_X32 FILLER_455_3455 ();
 FILLCELL_X32 FILLER_455_3487 ();
 FILLCELL_X32 FILLER_455_3519 ();
 FILLCELL_X32 FILLER_455_3551 ();
 FILLCELL_X32 FILLER_455_3583 ();
 FILLCELL_X32 FILLER_455_3615 ();
 FILLCELL_X32 FILLER_455_3647 ();
 FILLCELL_X32 FILLER_455_3679 ();
 FILLCELL_X16 FILLER_455_3711 ();
 FILLCELL_X8 FILLER_455_3727 ();
 FILLCELL_X2 FILLER_455_3735 ();
 FILLCELL_X1 FILLER_455_3737 ();
 FILLCELL_X32 FILLER_456_1 ();
 FILLCELL_X32 FILLER_456_33 ();
 FILLCELL_X32 FILLER_456_65 ();
 FILLCELL_X32 FILLER_456_97 ();
 FILLCELL_X32 FILLER_456_129 ();
 FILLCELL_X32 FILLER_456_161 ();
 FILLCELL_X32 FILLER_456_193 ();
 FILLCELL_X32 FILLER_456_225 ();
 FILLCELL_X32 FILLER_456_257 ();
 FILLCELL_X32 FILLER_456_289 ();
 FILLCELL_X32 FILLER_456_321 ();
 FILLCELL_X32 FILLER_456_353 ();
 FILLCELL_X32 FILLER_456_385 ();
 FILLCELL_X32 FILLER_456_417 ();
 FILLCELL_X32 FILLER_456_449 ();
 FILLCELL_X32 FILLER_456_481 ();
 FILLCELL_X32 FILLER_456_513 ();
 FILLCELL_X32 FILLER_456_545 ();
 FILLCELL_X32 FILLER_456_577 ();
 FILLCELL_X16 FILLER_456_609 ();
 FILLCELL_X4 FILLER_456_625 ();
 FILLCELL_X2 FILLER_456_629 ();
 FILLCELL_X32 FILLER_456_632 ();
 FILLCELL_X32 FILLER_456_664 ();
 FILLCELL_X32 FILLER_456_696 ();
 FILLCELL_X32 FILLER_456_728 ();
 FILLCELL_X32 FILLER_456_760 ();
 FILLCELL_X32 FILLER_456_792 ();
 FILLCELL_X32 FILLER_456_824 ();
 FILLCELL_X32 FILLER_456_856 ();
 FILLCELL_X32 FILLER_456_888 ();
 FILLCELL_X32 FILLER_456_920 ();
 FILLCELL_X32 FILLER_456_952 ();
 FILLCELL_X32 FILLER_456_984 ();
 FILLCELL_X32 FILLER_456_1016 ();
 FILLCELL_X32 FILLER_456_1048 ();
 FILLCELL_X32 FILLER_456_1080 ();
 FILLCELL_X32 FILLER_456_1112 ();
 FILLCELL_X32 FILLER_456_1144 ();
 FILLCELL_X32 FILLER_456_1176 ();
 FILLCELL_X32 FILLER_456_1208 ();
 FILLCELL_X32 FILLER_456_1240 ();
 FILLCELL_X32 FILLER_456_1272 ();
 FILLCELL_X32 FILLER_456_1304 ();
 FILLCELL_X32 FILLER_456_1336 ();
 FILLCELL_X32 FILLER_456_1368 ();
 FILLCELL_X32 FILLER_456_1400 ();
 FILLCELL_X32 FILLER_456_1432 ();
 FILLCELL_X32 FILLER_456_1464 ();
 FILLCELL_X32 FILLER_456_1496 ();
 FILLCELL_X32 FILLER_456_1528 ();
 FILLCELL_X32 FILLER_456_1560 ();
 FILLCELL_X32 FILLER_456_1592 ();
 FILLCELL_X32 FILLER_456_1624 ();
 FILLCELL_X32 FILLER_456_1656 ();
 FILLCELL_X32 FILLER_456_1688 ();
 FILLCELL_X32 FILLER_456_1720 ();
 FILLCELL_X32 FILLER_456_1752 ();
 FILLCELL_X32 FILLER_456_1784 ();
 FILLCELL_X32 FILLER_456_1816 ();
 FILLCELL_X32 FILLER_456_1848 ();
 FILLCELL_X8 FILLER_456_1880 ();
 FILLCELL_X4 FILLER_456_1888 ();
 FILLCELL_X2 FILLER_456_1892 ();
 FILLCELL_X32 FILLER_456_1895 ();
 FILLCELL_X32 FILLER_456_1927 ();
 FILLCELL_X32 FILLER_456_1959 ();
 FILLCELL_X32 FILLER_456_1991 ();
 FILLCELL_X32 FILLER_456_2023 ();
 FILLCELL_X32 FILLER_456_2055 ();
 FILLCELL_X32 FILLER_456_2087 ();
 FILLCELL_X32 FILLER_456_2119 ();
 FILLCELL_X32 FILLER_456_2151 ();
 FILLCELL_X32 FILLER_456_2183 ();
 FILLCELL_X32 FILLER_456_2215 ();
 FILLCELL_X32 FILLER_456_2247 ();
 FILLCELL_X32 FILLER_456_2279 ();
 FILLCELL_X32 FILLER_456_2311 ();
 FILLCELL_X32 FILLER_456_2343 ();
 FILLCELL_X32 FILLER_456_2375 ();
 FILLCELL_X32 FILLER_456_2407 ();
 FILLCELL_X32 FILLER_456_2439 ();
 FILLCELL_X32 FILLER_456_2471 ();
 FILLCELL_X32 FILLER_456_2503 ();
 FILLCELL_X32 FILLER_456_2535 ();
 FILLCELL_X32 FILLER_456_2567 ();
 FILLCELL_X32 FILLER_456_2599 ();
 FILLCELL_X32 FILLER_456_2631 ();
 FILLCELL_X32 FILLER_456_2663 ();
 FILLCELL_X32 FILLER_456_2695 ();
 FILLCELL_X32 FILLER_456_2727 ();
 FILLCELL_X32 FILLER_456_2759 ();
 FILLCELL_X32 FILLER_456_2791 ();
 FILLCELL_X32 FILLER_456_2823 ();
 FILLCELL_X32 FILLER_456_2855 ();
 FILLCELL_X32 FILLER_456_2887 ();
 FILLCELL_X32 FILLER_456_2919 ();
 FILLCELL_X32 FILLER_456_2951 ();
 FILLCELL_X32 FILLER_456_2983 ();
 FILLCELL_X32 FILLER_456_3015 ();
 FILLCELL_X32 FILLER_456_3047 ();
 FILLCELL_X32 FILLER_456_3079 ();
 FILLCELL_X32 FILLER_456_3111 ();
 FILLCELL_X8 FILLER_456_3143 ();
 FILLCELL_X4 FILLER_456_3151 ();
 FILLCELL_X2 FILLER_456_3155 ();
 FILLCELL_X32 FILLER_456_3158 ();
 FILLCELL_X32 FILLER_456_3190 ();
 FILLCELL_X32 FILLER_456_3222 ();
 FILLCELL_X32 FILLER_456_3254 ();
 FILLCELL_X32 FILLER_456_3286 ();
 FILLCELL_X32 FILLER_456_3318 ();
 FILLCELL_X32 FILLER_456_3350 ();
 FILLCELL_X32 FILLER_456_3382 ();
 FILLCELL_X32 FILLER_456_3414 ();
 FILLCELL_X32 FILLER_456_3446 ();
 FILLCELL_X32 FILLER_456_3478 ();
 FILLCELL_X32 FILLER_456_3510 ();
 FILLCELL_X32 FILLER_456_3542 ();
 FILLCELL_X32 FILLER_456_3574 ();
 FILLCELL_X32 FILLER_456_3606 ();
 FILLCELL_X32 FILLER_456_3638 ();
 FILLCELL_X32 FILLER_456_3670 ();
 FILLCELL_X32 FILLER_456_3702 ();
 FILLCELL_X4 FILLER_456_3734 ();
 FILLCELL_X32 FILLER_457_1 ();
 FILLCELL_X32 FILLER_457_33 ();
 FILLCELL_X32 FILLER_457_65 ();
 FILLCELL_X32 FILLER_457_97 ();
 FILLCELL_X32 FILLER_457_129 ();
 FILLCELL_X32 FILLER_457_161 ();
 FILLCELL_X32 FILLER_457_193 ();
 FILLCELL_X32 FILLER_457_225 ();
 FILLCELL_X32 FILLER_457_257 ();
 FILLCELL_X32 FILLER_457_289 ();
 FILLCELL_X32 FILLER_457_321 ();
 FILLCELL_X32 FILLER_457_353 ();
 FILLCELL_X32 FILLER_457_385 ();
 FILLCELL_X32 FILLER_457_417 ();
 FILLCELL_X32 FILLER_457_449 ();
 FILLCELL_X32 FILLER_457_481 ();
 FILLCELL_X32 FILLER_457_513 ();
 FILLCELL_X32 FILLER_457_545 ();
 FILLCELL_X32 FILLER_457_577 ();
 FILLCELL_X32 FILLER_457_609 ();
 FILLCELL_X32 FILLER_457_641 ();
 FILLCELL_X32 FILLER_457_673 ();
 FILLCELL_X32 FILLER_457_705 ();
 FILLCELL_X32 FILLER_457_737 ();
 FILLCELL_X32 FILLER_457_769 ();
 FILLCELL_X32 FILLER_457_801 ();
 FILLCELL_X32 FILLER_457_833 ();
 FILLCELL_X32 FILLER_457_865 ();
 FILLCELL_X32 FILLER_457_897 ();
 FILLCELL_X32 FILLER_457_929 ();
 FILLCELL_X32 FILLER_457_961 ();
 FILLCELL_X32 FILLER_457_993 ();
 FILLCELL_X32 FILLER_457_1025 ();
 FILLCELL_X32 FILLER_457_1057 ();
 FILLCELL_X32 FILLER_457_1089 ();
 FILLCELL_X32 FILLER_457_1121 ();
 FILLCELL_X32 FILLER_457_1153 ();
 FILLCELL_X32 FILLER_457_1185 ();
 FILLCELL_X32 FILLER_457_1217 ();
 FILLCELL_X8 FILLER_457_1249 ();
 FILLCELL_X4 FILLER_457_1257 ();
 FILLCELL_X2 FILLER_457_1261 ();
 FILLCELL_X32 FILLER_457_1264 ();
 FILLCELL_X32 FILLER_457_1296 ();
 FILLCELL_X32 FILLER_457_1328 ();
 FILLCELL_X32 FILLER_457_1360 ();
 FILLCELL_X32 FILLER_457_1392 ();
 FILLCELL_X32 FILLER_457_1424 ();
 FILLCELL_X32 FILLER_457_1456 ();
 FILLCELL_X32 FILLER_457_1488 ();
 FILLCELL_X32 FILLER_457_1520 ();
 FILLCELL_X32 FILLER_457_1552 ();
 FILLCELL_X32 FILLER_457_1584 ();
 FILLCELL_X32 FILLER_457_1616 ();
 FILLCELL_X32 FILLER_457_1648 ();
 FILLCELL_X32 FILLER_457_1680 ();
 FILLCELL_X32 FILLER_457_1712 ();
 FILLCELL_X32 FILLER_457_1744 ();
 FILLCELL_X32 FILLER_457_1776 ();
 FILLCELL_X32 FILLER_457_1808 ();
 FILLCELL_X32 FILLER_457_1840 ();
 FILLCELL_X32 FILLER_457_1872 ();
 FILLCELL_X32 FILLER_457_1904 ();
 FILLCELL_X32 FILLER_457_1936 ();
 FILLCELL_X32 FILLER_457_1968 ();
 FILLCELL_X32 FILLER_457_2000 ();
 FILLCELL_X32 FILLER_457_2032 ();
 FILLCELL_X32 FILLER_457_2064 ();
 FILLCELL_X32 FILLER_457_2096 ();
 FILLCELL_X32 FILLER_457_2128 ();
 FILLCELL_X32 FILLER_457_2160 ();
 FILLCELL_X32 FILLER_457_2192 ();
 FILLCELL_X32 FILLER_457_2224 ();
 FILLCELL_X32 FILLER_457_2256 ();
 FILLCELL_X32 FILLER_457_2288 ();
 FILLCELL_X32 FILLER_457_2320 ();
 FILLCELL_X32 FILLER_457_2352 ();
 FILLCELL_X32 FILLER_457_2384 ();
 FILLCELL_X32 FILLER_457_2416 ();
 FILLCELL_X32 FILLER_457_2448 ();
 FILLCELL_X32 FILLER_457_2480 ();
 FILLCELL_X8 FILLER_457_2512 ();
 FILLCELL_X4 FILLER_457_2520 ();
 FILLCELL_X2 FILLER_457_2524 ();
 FILLCELL_X32 FILLER_457_2527 ();
 FILLCELL_X32 FILLER_457_2559 ();
 FILLCELL_X32 FILLER_457_2591 ();
 FILLCELL_X32 FILLER_457_2623 ();
 FILLCELL_X32 FILLER_457_2655 ();
 FILLCELL_X32 FILLER_457_2687 ();
 FILLCELL_X32 FILLER_457_2719 ();
 FILLCELL_X32 FILLER_457_2751 ();
 FILLCELL_X32 FILLER_457_2783 ();
 FILLCELL_X32 FILLER_457_2815 ();
 FILLCELL_X32 FILLER_457_2847 ();
 FILLCELL_X32 FILLER_457_2879 ();
 FILLCELL_X32 FILLER_457_2911 ();
 FILLCELL_X32 FILLER_457_2943 ();
 FILLCELL_X32 FILLER_457_2975 ();
 FILLCELL_X32 FILLER_457_3007 ();
 FILLCELL_X32 FILLER_457_3039 ();
 FILLCELL_X32 FILLER_457_3071 ();
 FILLCELL_X32 FILLER_457_3103 ();
 FILLCELL_X32 FILLER_457_3135 ();
 FILLCELL_X32 FILLER_457_3167 ();
 FILLCELL_X32 FILLER_457_3199 ();
 FILLCELL_X32 FILLER_457_3231 ();
 FILLCELL_X32 FILLER_457_3263 ();
 FILLCELL_X32 FILLER_457_3295 ();
 FILLCELL_X32 FILLER_457_3327 ();
 FILLCELL_X32 FILLER_457_3359 ();
 FILLCELL_X32 FILLER_457_3391 ();
 FILLCELL_X32 FILLER_457_3423 ();
 FILLCELL_X32 FILLER_457_3455 ();
 FILLCELL_X32 FILLER_457_3487 ();
 FILLCELL_X32 FILLER_457_3519 ();
 FILLCELL_X32 FILLER_457_3551 ();
 FILLCELL_X32 FILLER_457_3583 ();
 FILLCELL_X32 FILLER_457_3615 ();
 FILLCELL_X32 FILLER_457_3647 ();
 FILLCELL_X32 FILLER_457_3679 ();
 FILLCELL_X16 FILLER_457_3711 ();
 FILLCELL_X8 FILLER_457_3727 ();
 FILLCELL_X2 FILLER_457_3735 ();
 FILLCELL_X1 FILLER_457_3737 ();
 FILLCELL_X32 FILLER_458_1 ();
 FILLCELL_X32 FILLER_458_33 ();
 FILLCELL_X32 FILLER_458_65 ();
 FILLCELL_X32 FILLER_458_97 ();
 FILLCELL_X32 FILLER_458_129 ();
 FILLCELL_X32 FILLER_458_161 ();
 FILLCELL_X32 FILLER_458_193 ();
 FILLCELL_X32 FILLER_458_225 ();
 FILLCELL_X32 FILLER_458_257 ();
 FILLCELL_X32 FILLER_458_289 ();
 FILLCELL_X32 FILLER_458_321 ();
 FILLCELL_X32 FILLER_458_353 ();
 FILLCELL_X32 FILLER_458_385 ();
 FILLCELL_X32 FILLER_458_417 ();
 FILLCELL_X32 FILLER_458_449 ();
 FILLCELL_X32 FILLER_458_481 ();
 FILLCELL_X32 FILLER_458_513 ();
 FILLCELL_X32 FILLER_458_545 ();
 FILLCELL_X32 FILLER_458_577 ();
 FILLCELL_X16 FILLER_458_609 ();
 FILLCELL_X4 FILLER_458_625 ();
 FILLCELL_X2 FILLER_458_629 ();
 FILLCELL_X32 FILLER_458_632 ();
 FILLCELL_X32 FILLER_458_664 ();
 FILLCELL_X32 FILLER_458_696 ();
 FILLCELL_X32 FILLER_458_728 ();
 FILLCELL_X32 FILLER_458_760 ();
 FILLCELL_X32 FILLER_458_792 ();
 FILLCELL_X32 FILLER_458_824 ();
 FILLCELL_X32 FILLER_458_856 ();
 FILLCELL_X32 FILLER_458_888 ();
 FILLCELL_X32 FILLER_458_920 ();
 FILLCELL_X32 FILLER_458_952 ();
 FILLCELL_X32 FILLER_458_984 ();
 FILLCELL_X32 FILLER_458_1016 ();
 FILLCELL_X32 FILLER_458_1048 ();
 FILLCELL_X32 FILLER_458_1080 ();
 FILLCELL_X32 FILLER_458_1112 ();
 FILLCELL_X32 FILLER_458_1144 ();
 FILLCELL_X32 FILLER_458_1176 ();
 FILLCELL_X32 FILLER_458_1208 ();
 FILLCELL_X32 FILLER_458_1240 ();
 FILLCELL_X32 FILLER_458_1272 ();
 FILLCELL_X32 FILLER_458_1304 ();
 FILLCELL_X32 FILLER_458_1336 ();
 FILLCELL_X32 FILLER_458_1368 ();
 FILLCELL_X32 FILLER_458_1400 ();
 FILLCELL_X32 FILLER_458_1432 ();
 FILLCELL_X32 FILLER_458_1464 ();
 FILLCELL_X32 FILLER_458_1496 ();
 FILLCELL_X32 FILLER_458_1528 ();
 FILLCELL_X32 FILLER_458_1560 ();
 FILLCELL_X32 FILLER_458_1592 ();
 FILLCELL_X32 FILLER_458_1624 ();
 FILLCELL_X32 FILLER_458_1656 ();
 FILLCELL_X32 FILLER_458_1688 ();
 FILLCELL_X32 FILLER_458_1720 ();
 FILLCELL_X32 FILLER_458_1752 ();
 FILLCELL_X32 FILLER_458_1784 ();
 FILLCELL_X32 FILLER_458_1816 ();
 FILLCELL_X32 FILLER_458_1848 ();
 FILLCELL_X8 FILLER_458_1880 ();
 FILLCELL_X4 FILLER_458_1888 ();
 FILLCELL_X2 FILLER_458_1892 ();
 FILLCELL_X32 FILLER_458_1895 ();
 FILLCELL_X32 FILLER_458_1927 ();
 FILLCELL_X32 FILLER_458_1959 ();
 FILLCELL_X32 FILLER_458_1991 ();
 FILLCELL_X32 FILLER_458_2023 ();
 FILLCELL_X32 FILLER_458_2055 ();
 FILLCELL_X32 FILLER_458_2087 ();
 FILLCELL_X32 FILLER_458_2119 ();
 FILLCELL_X32 FILLER_458_2151 ();
 FILLCELL_X32 FILLER_458_2183 ();
 FILLCELL_X32 FILLER_458_2215 ();
 FILLCELL_X32 FILLER_458_2247 ();
 FILLCELL_X32 FILLER_458_2279 ();
 FILLCELL_X32 FILLER_458_2311 ();
 FILLCELL_X32 FILLER_458_2343 ();
 FILLCELL_X32 FILLER_458_2375 ();
 FILLCELL_X32 FILLER_458_2407 ();
 FILLCELL_X32 FILLER_458_2439 ();
 FILLCELL_X32 FILLER_458_2471 ();
 FILLCELL_X32 FILLER_458_2503 ();
 FILLCELL_X32 FILLER_458_2535 ();
 FILLCELL_X32 FILLER_458_2567 ();
 FILLCELL_X32 FILLER_458_2599 ();
 FILLCELL_X32 FILLER_458_2631 ();
 FILLCELL_X32 FILLER_458_2663 ();
 FILLCELL_X32 FILLER_458_2695 ();
 FILLCELL_X32 FILLER_458_2727 ();
 FILLCELL_X32 FILLER_458_2759 ();
 FILLCELL_X32 FILLER_458_2791 ();
 FILLCELL_X32 FILLER_458_2823 ();
 FILLCELL_X32 FILLER_458_2855 ();
 FILLCELL_X32 FILLER_458_2887 ();
 FILLCELL_X32 FILLER_458_2919 ();
 FILLCELL_X32 FILLER_458_2951 ();
 FILLCELL_X32 FILLER_458_2983 ();
 FILLCELL_X32 FILLER_458_3015 ();
 FILLCELL_X32 FILLER_458_3047 ();
 FILLCELL_X32 FILLER_458_3079 ();
 FILLCELL_X32 FILLER_458_3111 ();
 FILLCELL_X8 FILLER_458_3143 ();
 FILLCELL_X4 FILLER_458_3151 ();
 FILLCELL_X2 FILLER_458_3155 ();
 FILLCELL_X32 FILLER_458_3158 ();
 FILLCELL_X32 FILLER_458_3190 ();
 FILLCELL_X32 FILLER_458_3222 ();
 FILLCELL_X32 FILLER_458_3254 ();
 FILLCELL_X32 FILLER_458_3286 ();
 FILLCELL_X32 FILLER_458_3318 ();
 FILLCELL_X32 FILLER_458_3350 ();
 FILLCELL_X32 FILLER_458_3382 ();
 FILLCELL_X32 FILLER_458_3414 ();
 FILLCELL_X32 FILLER_458_3446 ();
 FILLCELL_X32 FILLER_458_3478 ();
 FILLCELL_X32 FILLER_458_3510 ();
 FILLCELL_X32 FILLER_458_3542 ();
 FILLCELL_X32 FILLER_458_3574 ();
 FILLCELL_X32 FILLER_458_3606 ();
 FILLCELL_X32 FILLER_458_3638 ();
 FILLCELL_X32 FILLER_458_3670 ();
 FILLCELL_X32 FILLER_458_3702 ();
 FILLCELL_X4 FILLER_458_3734 ();
 FILLCELL_X32 FILLER_459_1 ();
 FILLCELL_X32 FILLER_459_33 ();
 FILLCELL_X32 FILLER_459_65 ();
 FILLCELL_X32 FILLER_459_97 ();
 FILLCELL_X32 FILLER_459_129 ();
 FILLCELL_X32 FILLER_459_161 ();
 FILLCELL_X32 FILLER_459_193 ();
 FILLCELL_X32 FILLER_459_225 ();
 FILLCELL_X32 FILLER_459_257 ();
 FILLCELL_X32 FILLER_459_289 ();
 FILLCELL_X32 FILLER_459_321 ();
 FILLCELL_X32 FILLER_459_353 ();
 FILLCELL_X32 FILLER_459_385 ();
 FILLCELL_X32 FILLER_459_417 ();
 FILLCELL_X32 FILLER_459_449 ();
 FILLCELL_X32 FILLER_459_481 ();
 FILLCELL_X32 FILLER_459_513 ();
 FILLCELL_X32 FILLER_459_545 ();
 FILLCELL_X32 FILLER_459_577 ();
 FILLCELL_X32 FILLER_459_609 ();
 FILLCELL_X32 FILLER_459_641 ();
 FILLCELL_X32 FILLER_459_673 ();
 FILLCELL_X32 FILLER_459_705 ();
 FILLCELL_X32 FILLER_459_737 ();
 FILLCELL_X32 FILLER_459_769 ();
 FILLCELL_X32 FILLER_459_801 ();
 FILLCELL_X32 FILLER_459_833 ();
 FILLCELL_X32 FILLER_459_865 ();
 FILLCELL_X32 FILLER_459_897 ();
 FILLCELL_X32 FILLER_459_929 ();
 FILLCELL_X32 FILLER_459_961 ();
 FILLCELL_X32 FILLER_459_993 ();
 FILLCELL_X32 FILLER_459_1025 ();
 FILLCELL_X32 FILLER_459_1057 ();
 FILLCELL_X32 FILLER_459_1089 ();
 FILLCELL_X32 FILLER_459_1121 ();
 FILLCELL_X32 FILLER_459_1153 ();
 FILLCELL_X32 FILLER_459_1185 ();
 FILLCELL_X32 FILLER_459_1217 ();
 FILLCELL_X8 FILLER_459_1249 ();
 FILLCELL_X4 FILLER_459_1257 ();
 FILLCELL_X2 FILLER_459_1261 ();
 FILLCELL_X32 FILLER_459_1264 ();
 FILLCELL_X32 FILLER_459_1296 ();
 FILLCELL_X32 FILLER_459_1328 ();
 FILLCELL_X32 FILLER_459_1360 ();
 FILLCELL_X32 FILLER_459_1392 ();
 FILLCELL_X32 FILLER_459_1424 ();
 FILLCELL_X32 FILLER_459_1456 ();
 FILLCELL_X32 FILLER_459_1488 ();
 FILLCELL_X32 FILLER_459_1520 ();
 FILLCELL_X32 FILLER_459_1552 ();
 FILLCELL_X32 FILLER_459_1584 ();
 FILLCELL_X32 FILLER_459_1616 ();
 FILLCELL_X32 FILLER_459_1648 ();
 FILLCELL_X32 FILLER_459_1680 ();
 FILLCELL_X32 FILLER_459_1712 ();
 FILLCELL_X32 FILLER_459_1744 ();
 FILLCELL_X32 FILLER_459_1776 ();
 FILLCELL_X32 FILLER_459_1808 ();
 FILLCELL_X32 FILLER_459_1840 ();
 FILLCELL_X32 FILLER_459_1872 ();
 FILLCELL_X32 FILLER_459_1904 ();
 FILLCELL_X32 FILLER_459_1936 ();
 FILLCELL_X32 FILLER_459_1968 ();
 FILLCELL_X32 FILLER_459_2000 ();
 FILLCELL_X32 FILLER_459_2032 ();
 FILLCELL_X32 FILLER_459_2064 ();
 FILLCELL_X32 FILLER_459_2096 ();
 FILLCELL_X32 FILLER_459_2128 ();
 FILLCELL_X32 FILLER_459_2160 ();
 FILLCELL_X32 FILLER_459_2192 ();
 FILLCELL_X32 FILLER_459_2224 ();
 FILLCELL_X32 FILLER_459_2256 ();
 FILLCELL_X32 FILLER_459_2288 ();
 FILLCELL_X32 FILLER_459_2320 ();
 FILLCELL_X32 FILLER_459_2352 ();
 FILLCELL_X32 FILLER_459_2384 ();
 FILLCELL_X32 FILLER_459_2416 ();
 FILLCELL_X32 FILLER_459_2448 ();
 FILLCELL_X32 FILLER_459_2480 ();
 FILLCELL_X8 FILLER_459_2512 ();
 FILLCELL_X4 FILLER_459_2520 ();
 FILLCELL_X2 FILLER_459_2524 ();
 FILLCELL_X32 FILLER_459_2527 ();
 FILLCELL_X32 FILLER_459_2559 ();
 FILLCELL_X32 FILLER_459_2591 ();
 FILLCELL_X32 FILLER_459_2623 ();
 FILLCELL_X32 FILLER_459_2655 ();
 FILLCELL_X32 FILLER_459_2687 ();
 FILLCELL_X32 FILLER_459_2719 ();
 FILLCELL_X32 FILLER_459_2751 ();
 FILLCELL_X32 FILLER_459_2783 ();
 FILLCELL_X32 FILLER_459_2815 ();
 FILLCELL_X32 FILLER_459_2847 ();
 FILLCELL_X32 FILLER_459_2879 ();
 FILLCELL_X32 FILLER_459_2911 ();
 FILLCELL_X32 FILLER_459_2943 ();
 FILLCELL_X32 FILLER_459_2975 ();
 FILLCELL_X32 FILLER_459_3007 ();
 FILLCELL_X32 FILLER_459_3039 ();
 FILLCELL_X32 FILLER_459_3071 ();
 FILLCELL_X32 FILLER_459_3103 ();
 FILLCELL_X32 FILLER_459_3135 ();
 FILLCELL_X32 FILLER_459_3167 ();
 FILLCELL_X32 FILLER_459_3199 ();
 FILLCELL_X32 FILLER_459_3231 ();
 FILLCELL_X32 FILLER_459_3263 ();
 FILLCELL_X32 FILLER_459_3295 ();
 FILLCELL_X32 FILLER_459_3327 ();
 FILLCELL_X32 FILLER_459_3359 ();
 FILLCELL_X32 FILLER_459_3391 ();
 FILLCELL_X32 FILLER_459_3423 ();
 FILLCELL_X32 FILLER_459_3455 ();
 FILLCELL_X32 FILLER_459_3487 ();
 FILLCELL_X32 FILLER_459_3519 ();
 FILLCELL_X32 FILLER_459_3551 ();
 FILLCELL_X32 FILLER_459_3583 ();
 FILLCELL_X32 FILLER_459_3615 ();
 FILLCELL_X32 FILLER_459_3647 ();
 FILLCELL_X32 FILLER_459_3679 ();
 FILLCELL_X16 FILLER_459_3711 ();
 FILLCELL_X8 FILLER_459_3727 ();
 FILLCELL_X2 FILLER_459_3735 ();
 FILLCELL_X1 FILLER_459_3737 ();
 FILLCELL_X32 FILLER_460_1 ();
 FILLCELL_X32 FILLER_460_33 ();
 FILLCELL_X32 FILLER_460_65 ();
 FILLCELL_X32 FILLER_460_97 ();
 FILLCELL_X32 FILLER_460_129 ();
 FILLCELL_X32 FILLER_460_161 ();
 FILLCELL_X32 FILLER_460_193 ();
 FILLCELL_X32 FILLER_460_225 ();
 FILLCELL_X32 FILLER_460_257 ();
 FILLCELL_X32 FILLER_460_289 ();
 FILLCELL_X32 FILLER_460_321 ();
 FILLCELL_X32 FILLER_460_353 ();
 FILLCELL_X32 FILLER_460_385 ();
 FILLCELL_X32 FILLER_460_417 ();
 FILLCELL_X32 FILLER_460_449 ();
 FILLCELL_X32 FILLER_460_481 ();
 FILLCELL_X32 FILLER_460_513 ();
 FILLCELL_X32 FILLER_460_545 ();
 FILLCELL_X32 FILLER_460_577 ();
 FILLCELL_X16 FILLER_460_609 ();
 FILLCELL_X4 FILLER_460_625 ();
 FILLCELL_X2 FILLER_460_629 ();
 FILLCELL_X32 FILLER_460_632 ();
 FILLCELL_X32 FILLER_460_664 ();
 FILLCELL_X32 FILLER_460_696 ();
 FILLCELL_X32 FILLER_460_728 ();
 FILLCELL_X32 FILLER_460_760 ();
 FILLCELL_X32 FILLER_460_792 ();
 FILLCELL_X32 FILLER_460_824 ();
 FILLCELL_X32 FILLER_460_856 ();
 FILLCELL_X32 FILLER_460_888 ();
 FILLCELL_X32 FILLER_460_920 ();
 FILLCELL_X32 FILLER_460_952 ();
 FILLCELL_X32 FILLER_460_984 ();
 FILLCELL_X32 FILLER_460_1016 ();
 FILLCELL_X32 FILLER_460_1048 ();
 FILLCELL_X32 FILLER_460_1080 ();
 FILLCELL_X32 FILLER_460_1112 ();
 FILLCELL_X32 FILLER_460_1144 ();
 FILLCELL_X32 FILLER_460_1176 ();
 FILLCELL_X32 FILLER_460_1208 ();
 FILLCELL_X32 FILLER_460_1240 ();
 FILLCELL_X32 FILLER_460_1272 ();
 FILLCELL_X32 FILLER_460_1304 ();
 FILLCELL_X32 FILLER_460_1336 ();
 FILLCELL_X32 FILLER_460_1368 ();
 FILLCELL_X32 FILLER_460_1400 ();
 FILLCELL_X32 FILLER_460_1432 ();
 FILLCELL_X32 FILLER_460_1464 ();
 FILLCELL_X32 FILLER_460_1496 ();
 FILLCELL_X32 FILLER_460_1528 ();
 FILLCELL_X32 FILLER_460_1560 ();
 FILLCELL_X32 FILLER_460_1592 ();
 FILLCELL_X32 FILLER_460_1624 ();
 FILLCELL_X32 FILLER_460_1656 ();
 FILLCELL_X32 FILLER_460_1688 ();
 FILLCELL_X32 FILLER_460_1720 ();
 FILLCELL_X32 FILLER_460_1752 ();
 FILLCELL_X32 FILLER_460_1784 ();
 FILLCELL_X32 FILLER_460_1816 ();
 FILLCELL_X32 FILLER_460_1848 ();
 FILLCELL_X8 FILLER_460_1880 ();
 FILLCELL_X4 FILLER_460_1888 ();
 FILLCELL_X2 FILLER_460_1892 ();
 FILLCELL_X32 FILLER_460_1895 ();
 FILLCELL_X32 FILLER_460_1927 ();
 FILLCELL_X32 FILLER_460_1959 ();
 FILLCELL_X32 FILLER_460_1991 ();
 FILLCELL_X32 FILLER_460_2023 ();
 FILLCELL_X32 FILLER_460_2055 ();
 FILLCELL_X32 FILLER_460_2087 ();
 FILLCELL_X32 FILLER_460_2119 ();
 FILLCELL_X32 FILLER_460_2151 ();
 FILLCELL_X32 FILLER_460_2183 ();
 FILLCELL_X32 FILLER_460_2215 ();
 FILLCELL_X32 FILLER_460_2247 ();
 FILLCELL_X32 FILLER_460_2279 ();
 FILLCELL_X32 FILLER_460_2311 ();
 FILLCELL_X32 FILLER_460_2343 ();
 FILLCELL_X32 FILLER_460_2375 ();
 FILLCELL_X32 FILLER_460_2407 ();
 FILLCELL_X32 FILLER_460_2439 ();
 FILLCELL_X32 FILLER_460_2471 ();
 FILLCELL_X32 FILLER_460_2503 ();
 FILLCELL_X32 FILLER_460_2535 ();
 FILLCELL_X32 FILLER_460_2567 ();
 FILLCELL_X32 FILLER_460_2599 ();
 FILLCELL_X32 FILLER_460_2631 ();
 FILLCELL_X32 FILLER_460_2663 ();
 FILLCELL_X32 FILLER_460_2695 ();
 FILLCELL_X32 FILLER_460_2727 ();
 FILLCELL_X32 FILLER_460_2759 ();
 FILLCELL_X32 FILLER_460_2791 ();
 FILLCELL_X32 FILLER_460_2823 ();
 FILLCELL_X32 FILLER_460_2855 ();
 FILLCELL_X32 FILLER_460_2887 ();
 FILLCELL_X32 FILLER_460_2919 ();
 FILLCELL_X32 FILLER_460_2951 ();
 FILLCELL_X32 FILLER_460_2983 ();
 FILLCELL_X32 FILLER_460_3015 ();
 FILLCELL_X32 FILLER_460_3047 ();
 FILLCELL_X32 FILLER_460_3079 ();
 FILLCELL_X32 FILLER_460_3111 ();
 FILLCELL_X8 FILLER_460_3143 ();
 FILLCELL_X4 FILLER_460_3151 ();
 FILLCELL_X2 FILLER_460_3155 ();
 FILLCELL_X32 FILLER_460_3158 ();
 FILLCELL_X32 FILLER_460_3190 ();
 FILLCELL_X32 FILLER_460_3222 ();
 FILLCELL_X32 FILLER_460_3254 ();
 FILLCELL_X32 FILLER_460_3286 ();
 FILLCELL_X32 FILLER_460_3318 ();
 FILLCELL_X32 FILLER_460_3350 ();
 FILLCELL_X32 FILLER_460_3382 ();
 FILLCELL_X32 FILLER_460_3414 ();
 FILLCELL_X32 FILLER_460_3446 ();
 FILLCELL_X32 FILLER_460_3478 ();
 FILLCELL_X32 FILLER_460_3510 ();
 FILLCELL_X32 FILLER_460_3542 ();
 FILLCELL_X32 FILLER_460_3574 ();
 FILLCELL_X32 FILLER_460_3606 ();
 FILLCELL_X32 FILLER_460_3638 ();
 FILLCELL_X32 FILLER_460_3670 ();
 FILLCELL_X32 FILLER_460_3702 ();
 FILLCELL_X4 FILLER_460_3734 ();
 FILLCELL_X32 FILLER_461_1 ();
 FILLCELL_X32 FILLER_461_33 ();
 FILLCELL_X32 FILLER_461_65 ();
 FILLCELL_X32 FILLER_461_97 ();
 FILLCELL_X32 FILLER_461_129 ();
 FILLCELL_X32 FILLER_461_161 ();
 FILLCELL_X32 FILLER_461_193 ();
 FILLCELL_X32 FILLER_461_225 ();
 FILLCELL_X32 FILLER_461_257 ();
 FILLCELL_X32 FILLER_461_289 ();
 FILLCELL_X32 FILLER_461_321 ();
 FILLCELL_X32 FILLER_461_353 ();
 FILLCELL_X32 FILLER_461_385 ();
 FILLCELL_X32 FILLER_461_417 ();
 FILLCELL_X32 FILLER_461_449 ();
 FILLCELL_X32 FILLER_461_481 ();
 FILLCELL_X32 FILLER_461_513 ();
 FILLCELL_X32 FILLER_461_545 ();
 FILLCELL_X32 FILLER_461_577 ();
 FILLCELL_X32 FILLER_461_609 ();
 FILLCELL_X32 FILLER_461_641 ();
 FILLCELL_X32 FILLER_461_673 ();
 FILLCELL_X32 FILLER_461_705 ();
 FILLCELL_X32 FILLER_461_737 ();
 FILLCELL_X32 FILLER_461_769 ();
 FILLCELL_X32 FILLER_461_801 ();
 FILLCELL_X32 FILLER_461_833 ();
 FILLCELL_X32 FILLER_461_865 ();
 FILLCELL_X32 FILLER_461_897 ();
 FILLCELL_X32 FILLER_461_929 ();
 FILLCELL_X32 FILLER_461_961 ();
 FILLCELL_X32 FILLER_461_993 ();
 FILLCELL_X32 FILLER_461_1025 ();
 FILLCELL_X32 FILLER_461_1057 ();
 FILLCELL_X32 FILLER_461_1089 ();
 FILLCELL_X32 FILLER_461_1121 ();
 FILLCELL_X32 FILLER_461_1153 ();
 FILLCELL_X32 FILLER_461_1185 ();
 FILLCELL_X32 FILLER_461_1217 ();
 FILLCELL_X8 FILLER_461_1249 ();
 FILLCELL_X4 FILLER_461_1257 ();
 FILLCELL_X2 FILLER_461_1261 ();
 FILLCELL_X32 FILLER_461_1264 ();
 FILLCELL_X32 FILLER_461_1296 ();
 FILLCELL_X32 FILLER_461_1328 ();
 FILLCELL_X32 FILLER_461_1360 ();
 FILLCELL_X32 FILLER_461_1392 ();
 FILLCELL_X32 FILLER_461_1424 ();
 FILLCELL_X32 FILLER_461_1456 ();
 FILLCELL_X32 FILLER_461_1488 ();
 FILLCELL_X32 FILLER_461_1520 ();
 FILLCELL_X32 FILLER_461_1552 ();
 FILLCELL_X32 FILLER_461_1584 ();
 FILLCELL_X32 FILLER_461_1616 ();
 FILLCELL_X32 FILLER_461_1648 ();
 FILLCELL_X32 FILLER_461_1680 ();
 FILLCELL_X32 FILLER_461_1712 ();
 FILLCELL_X32 FILLER_461_1744 ();
 FILLCELL_X32 FILLER_461_1776 ();
 FILLCELL_X32 FILLER_461_1808 ();
 FILLCELL_X32 FILLER_461_1840 ();
 FILLCELL_X32 FILLER_461_1872 ();
 FILLCELL_X32 FILLER_461_1904 ();
 FILLCELL_X32 FILLER_461_1936 ();
 FILLCELL_X32 FILLER_461_1968 ();
 FILLCELL_X32 FILLER_461_2000 ();
 FILLCELL_X32 FILLER_461_2032 ();
 FILLCELL_X32 FILLER_461_2064 ();
 FILLCELL_X32 FILLER_461_2096 ();
 FILLCELL_X32 FILLER_461_2128 ();
 FILLCELL_X32 FILLER_461_2160 ();
 FILLCELL_X32 FILLER_461_2192 ();
 FILLCELL_X32 FILLER_461_2224 ();
 FILLCELL_X32 FILLER_461_2256 ();
 FILLCELL_X32 FILLER_461_2288 ();
 FILLCELL_X32 FILLER_461_2320 ();
 FILLCELL_X32 FILLER_461_2352 ();
 FILLCELL_X32 FILLER_461_2384 ();
 FILLCELL_X32 FILLER_461_2416 ();
 FILLCELL_X32 FILLER_461_2448 ();
 FILLCELL_X32 FILLER_461_2480 ();
 FILLCELL_X8 FILLER_461_2512 ();
 FILLCELL_X4 FILLER_461_2520 ();
 FILLCELL_X2 FILLER_461_2524 ();
 FILLCELL_X32 FILLER_461_2527 ();
 FILLCELL_X32 FILLER_461_2559 ();
 FILLCELL_X32 FILLER_461_2591 ();
 FILLCELL_X32 FILLER_461_2623 ();
 FILLCELL_X32 FILLER_461_2655 ();
 FILLCELL_X32 FILLER_461_2687 ();
 FILLCELL_X32 FILLER_461_2719 ();
 FILLCELL_X32 FILLER_461_2751 ();
 FILLCELL_X32 FILLER_461_2783 ();
 FILLCELL_X32 FILLER_461_2815 ();
 FILLCELL_X32 FILLER_461_2847 ();
 FILLCELL_X32 FILLER_461_2879 ();
 FILLCELL_X32 FILLER_461_2911 ();
 FILLCELL_X32 FILLER_461_2943 ();
 FILLCELL_X32 FILLER_461_2975 ();
 FILLCELL_X32 FILLER_461_3007 ();
 FILLCELL_X32 FILLER_461_3039 ();
 FILLCELL_X32 FILLER_461_3071 ();
 FILLCELL_X32 FILLER_461_3103 ();
 FILLCELL_X32 FILLER_461_3135 ();
 FILLCELL_X32 FILLER_461_3167 ();
 FILLCELL_X32 FILLER_461_3199 ();
 FILLCELL_X32 FILLER_461_3231 ();
 FILLCELL_X32 FILLER_461_3263 ();
 FILLCELL_X32 FILLER_461_3295 ();
 FILLCELL_X32 FILLER_461_3327 ();
 FILLCELL_X32 FILLER_461_3359 ();
 FILLCELL_X32 FILLER_461_3391 ();
 FILLCELL_X32 FILLER_461_3423 ();
 FILLCELL_X32 FILLER_461_3455 ();
 FILLCELL_X32 FILLER_461_3487 ();
 FILLCELL_X32 FILLER_461_3519 ();
 FILLCELL_X32 FILLER_461_3551 ();
 FILLCELL_X32 FILLER_461_3583 ();
 FILLCELL_X32 FILLER_461_3615 ();
 FILLCELL_X32 FILLER_461_3647 ();
 FILLCELL_X32 FILLER_461_3679 ();
 FILLCELL_X16 FILLER_461_3711 ();
 FILLCELL_X8 FILLER_461_3727 ();
 FILLCELL_X2 FILLER_461_3735 ();
 FILLCELL_X1 FILLER_461_3737 ();
 FILLCELL_X32 FILLER_462_1 ();
 FILLCELL_X32 FILLER_462_33 ();
 FILLCELL_X32 FILLER_462_65 ();
 FILLCELL_X32 FILLER_462_97 ();
 FILLCELL_X32 FILLER_462_129 ();
 FILLCELL_X32 FILLER_462_161 ();
 FILLCELL_X32 FILLER_462_193 ();
 FILLCELL_X32 FILLER_462_225 ();
 FILLCELL_X32 FILLER_462_257 ();
 FILLCELL_X32 FILLER_462_289 ();
 FILLCELL_X32 FILLER_462_321 ();
 FILLCELL_X32 FILLER_462_353 ();
 FILLCELL_X32 FILLER_462_385 ();
 FILLCELL_X32 FILLER_462_417 ();
 FILLCELL_X32 FILLER_462_449 ();
 FILLCELL_X32 FILLER_462_481 ();
 FILLCELL_X32 FILLER_462_513 ();
 FILLCELL_X32 FILLER_462_545 ();
 FILLCELL_X32 FILLER_462_577 ();
 FILLCELL_X16 FILLER_462_609 ();
 FILLCELL_X4 FILLER_462_625 ();
 FILLCELL_X2 FILLER_462_629 ();
 FILLCELL_X32 FILLER_462_632 ();
 FILLCELL_X32 FILLER_462_664 ();
 FILLCELL_X32 FILLER_462_696 ();
 FILLCELL_X32 FILLER_462_728 ();
 FILLCELL_X32 FILLER_462_760 ();
 FILLCELL_X32 FILLER_462_792 ();
 FILLCELL_X32 FILLER_462_824 ();
 FILLCELL_X32 FILLER_462_856 ();
 FILLCELL_X32 FILLER_462_888 ();
 FILLCELL_X32 FILLER_462_920 ();
 FILLCELL_X32 FILLER_462_952 ();
 FILLCELL_X32 FILLER_462_984 ();
 FILLCELL_X32 FILLER_462_1016 ();
 FILLCELL_X32 FILLER_462_1048 ();
 FILLCELL_X32 FILLER_462_1080 ();
 FILLCELL_X32 FILLER_462_1112 ();
 FILLCELL_X32 FILLER_462_1144 ();
 FILLCELL_X32 FILLER_462_1176 ();
 FILLCELL_X32 FILLER_462_1208 ();
 FILLCELL_X32 FILLER_462_1240 ();
 FILLCELL_X32 FILLER_462_1272 ();
 FILLCELL_X32 FILLER_462_1304 ();
 FILLCELL_X32 FILLER_462_1336 ();
 FILLCELL_X32 FILLER_462_1368 ();
 FILLCELL_X32 FILLER_462_1400 ();
 FILLCELL_X32 FILLER_462_1432 ();
 FILLCELL_X32 FILLER_462_1464 ();
 FILLCELL_X32 FILLER_462_1496 ();
 FILLCELL_X32 FILLER_462_1528 ();
 FILLCELL_X32 FILLER_462_1560 ();
 FILLCELL_X32 FILLER_462_1592 ();
 FILLCELL_X32 FILLER_462_1624 ();
 FILLCELL_X32 FILLER_462_1656 ();
 FILLCELL_X32 FILLER_462_1688 ();
 FILLCELL_X32 FILLER_462_1720 ();
 FILLCELL_X32 FILLER_462_1752 ();
 FILLCELL_X32 FILLER_462_1784 ();
 FILLCELL_X32 FILLER_462_1816 ();
 FILLCELL_X32 FILLER_462_1848 ();
 FILLCELL_X8 FILLER_462_1880 ();
 FILLCELL_X4 FILLER_462_1888 ();
 FILLCELL_X2 FILLER_462_1892 ();
 FILLCELL_X32 FILLER_462_1895 ();
 FILLCELL_X32 FILLER_462_1927 ();
 FILLCELL_X32 FILLER_462_1959 ();
 FILLCELL_X32 FILLER_462_1991 ();
 FILLCELL_X32 FILLER_462_2023 ();
 FILLCELL_X32 FILLER_462_2055 ();
 FILLCELL_X32 FILLER_462_2087 ();
 FILLCELL_X32 FILLER_462_2119 ();
 FILLCELL_X32 FILLER_462_2151 ();
 FILLCELL_X32 FILLER_462_2183 ();
 FILLCELL_X32 FILLER_462_2215 ();
 FILLCELL_X32 FILLER_462_2247 ();
 FILLCELL_X32 FILLER_462_2279 ();
 FILLCELL_X32 FILLER_462_2311 ();
 FILLCELL_X32 FILLER_462_2343 ();
 FILLCELL_X32 FILLER_462_2375 ();
 FILLCELL_X32 FILLER_462_2407 ();
 FILLCELL_X32 FILLER_462_2439 ();
 FILLCELL_X32 FILLER_462_2471 ();
 FILLCELL_X32 FILLER_462_2503 ();
 FILLCELL_X32 FILLER_462_2535 ();
 FILLCELL_X32 FILLER_462_2567 ();
 FILLCELL_X32 FILLER_462_2599 ();
 FILLCELL_X32 FILLER_462_2631 ();
 FILLCELL_X32 FILLER_462_2663 ();
 FILLCELL_X32 FILLER_462_2695 ();
 FILLCELL_X32 FILLER_462_2727 ();
 FILLCELL_X32 FILLER_462_2759 ();
 FILLCELL_X32 FILLER_462_2791 ();
 FILLCELL_X32 FILLER_462_2823 ();
 FILLCELL_X32 FILLER_462_2855 ();
 FILLCELL_X32 FILLER_462_2887 ();
 FILLCELL_X32 FILLER_462_2919 ();
 FILLCELL_X32 FILLER_462_2951 ();
 FILLCELL_X32 FILLER_462_2983 ();
 FILLCELL_X32 FILLER_462_3015 ();
 FILLCELL_X32 FILLER_462_3047 ();
 FILLCELL_X32 FILLER_462_3079 ();
 FILLCELL_X32 FILLER_462_3111 ();
 FILLCELL_X8 FILLER_462_3143 ();
 FILLCELL_X4 FILLER_462_3151 ();
 FILLCELL_X2 FILLER_462_3155 ();
 FILLCELL_X32 FILLER_462_3158 ();
 FILLCELL_X32 FILLER_462_3190 ();
 FILLCELL_X32 FILLER_462_3222 ();
 FILLCELL_X32 FILLER_462_3254 ();
 FILLCELL_X32 FILLER_462_3286 ();
 FILLCELL_X32 FILLER_462_3318 ();
 FILLCELL_X32 FILLER_462_3350 ();
 FILLCELL_X32 FILLER_462_3382 ();
 FILLCELL_X32 FILLER_462_3414 ();
 FILLCELL_X32 FILLER_462_3446 ();
 FILLCELL_X32 FILLER_462_3478 ();
 FILLCELL_X32 FILLER_462_3510 ();
 FILLCELL_X32 FILLER_462_3542 ();
 FILLCELL_X32 FILLER_462_3574 ();
 FILLCELL_X32 FILLER_462_3606 ();
 FILLCELL_X32 FILLER_462_3638 ();
 FILLCELL_X32 FILLER_462_3670 ();
 FILLCELL_X32 FILLER_462_3702 ();
 FILLCELL_X4 FILLER_462_3734 ();
 FILLCELL_X32 FILLER_463_1 ();
 FILLCELL_X32 FILLER_463_33 ();
 FILLCELL_X32 FILLER_463_65 ();
 FILLCELL_X32 FILLER_463_97 ();
 FILLCELL_X32 FILLER_463_129 ();
 FILLCELL_X32 FILLER_463_161 ();
 FILLCELL_X32 FILLER_463_193 ();
 FILLCELL_X32 FILLER_463_225 ();
 FILLCELL_X32 FILLER_463_257 ();
 FILLCELL_X32 FILLER_463_289 ();
 FILLCELL_X32 FILLER_463_321 ();
 FILLCELL_X32 FILLER_463_353 ();
 FILLCELL_X32 FILLER_463_385 ();
 FILLCELL_X32 FILLER_463_417 ();
 FILLCELL_X32 FILLER_463_449 ();
 FILLCELL_X32 FILLER_463_481 ();
 FILLCELL_X32 FILLER_463_513 ();
 FILLCELL_X32 FILLER_463_545 ();
 FILLCELL_X32 FILLER_463_577 ();
 FILLCELL_X32 FILLER_463_609 ();
 FILLCELL_X32 FILLER_463_641 ();
 FILLCELL_X32 FILLER_463_673 ();
 FILLCELL_X32 FILLER_463_705 ();
 FILLCELL_X32 FILLER_463_737 ();
 FILLCELL_X32 FILLER_463_769 ();
 FILLCELL_X32 FILLER_463_801 ();
 FILLCELL_X32 FILLER_463_833 ();
 FILLCELL_X32 FILLER_463_865 ();
 FILLCELL_X32 FILLER_463_897 ();
 FILLCELL_X32 FILLER_463_929 ();
 FILLCELL_X32 FILLER_463_961 ();
 FILLCELL_X32 FILLER_463_993 ();
 FILLCELL_X32 FILLER_463_1025 ();
 FILLCELL_X32 FILLER_463_1057 ();
 FILLCELL_X32 FILLER_463_1089 ();
 FILLCELL_X32 FILLER_463_1121 ();
 FILLCELL_X32 FILLER_463_1153 ();
 FILLCELL_X32 FILLER_463_1185 ();
 FILLCELL_X32 FILLER_463_1217 ();
 FILLCELL_X8 FILLER_463_1249 ();
 FILLCELL_X4 FILLER_463_1257 ();
 FILLCELL_X2 FILLER_463_1261 ();
 FILLCELL_X32 FILLER_463_1264 ();
 FILLCELL_X32 FILLER_463_1296 ();
 FILLCELL_X32 FILLER_463_1328 ();
 FILLCELL_X32 FILLER_463_1360 ();
 FILLCELL_X32 FILLER_463_1392 ();
 FILLCELL_X32 FILLER_463_1424 ();
 FILLCELL_X32 FILLER_463_1456 ();
 FILLCELL_X32 FILLER_463_1488 ();
 FILLCELL_X32 FILLER_463_1520 ();
 FILLCELL_X32 FILLER_463_1552 ();
 FILLCELL_X32 FILLER_463_1584 ();
 FILLCELL_X32 FILLER_463_1616 ();
 FILLCELL_X32 FILLER_463_1648 ();
 FILLCELL_X32 FILLER_463_1680 ();
 FILLCELL_X32 FILLER_463_1712 ();
 FILLCELL_X32 FILLER_463_1744 ();
 FILLCELL_X32 FILLER_463_1776 ();
 FILLCELL_X32 FILLER_463_1808 ();
 FILLCELL_X32 FILLER_463_1840 ();
 FILLCELL_X32 FILLER_463_1872 ();
 FILLCELL_X32 FILLER_463_1904 ();
 FILLCELL_X32 FILLER_463_1936 ();
 FILLCELL_X32 FILLER_463_1968 ();
 FILLCELL_X32 FILLER_463_2000 ();
 FILLCELL_X32 FILLER_463_2032 ();
 FILLCELL_X32 FILLER_463_2064 ();
 FILLCELL_X32 FILLER_463_2096 ();
 FILLCELL_X32 FILLER_463_2128 ();
 FILLCELL_X32 FILLER_463_2160 ();
 FILLCELL_X32 FILLER_463_2192 ();
 FILLCELL_X32 FILLER_463_2224 ();
 FILLCELL_X32 FILLER_463_2256 ();
 FILLCELL_X32 FILLER_463_2288 ();
 FILLCELL_X32 FILLER_463_2320 ();
 FILLCELL_X32 FILLER_463_2352 ();
 FILLCELL_X32 FILLER_463_2384 ();
 FILLCELL_X32 FILLER_463_2416 ();
 FILLCELL_X32 FILLER_463_2448 ();
 FILLCELL_X32 FILLER_463_2480 ();
 FILLCELL_X8 FILLER_463_2512 ();
 FILLCELL_X4 FILLER_463_2520 ();
 FILLCELL_X2 FILLER_463_2524 ();
 FILLCELL_X32 FILLER_463_2527 ();
 FILLCELL_X32 FILLER_463_2559 ();
 FILLCELL_X32 FILLER_463_2591 ();
 FILLCELL_X32 FILLER_463_2623 ();
 FILLCELL_X32 FILLER_463_2655 ();
 FILLCELL_X32 FILLER_463_2687 ();
 FILLCELL_X32 FILLER_463_2719 ();
 FILLCELL_X32 FILLER_463_2751 ();
 FILLCELL_X32 FILLER_463_2783 ();
 FILLCELL_X32 FILLER_463_2815 ();
 FILLCELL_X32 FILLER_463_2847 ();
 FILLCELL_X32 FILLER_463_2879 ();
 FILLCELL_X32 FILLER_463_2911 ();
 FILLCELL_X32 FILLER_463_2943 ();
 FILLCELL_X32 FILLER_463_2975 ();
 FILLCELL_X32 FILLER_463_3007 ();
 FILLCELL_X32 FILLER_463_3039 ();
 FILLCELL_X32 FILLER_463_3071 ();
 FILLCELL_X32 FILLER_463_3103 ();
 FILLCELL_X32 FILLER_463_3135 ();
 FILLCELL_X32 FILLER_463_3167 ();
 FILLCELL_X32 FILLER_463_3199 ();
 FILLCELL_X32 FILLER_463_3231 ();
 FILLCELL_X32 FILLER_463_3263 ();
 FILLCELL_X32 FILLER_463_3295 ();
 FILLCELL_X32 FILLER_463_3327 ();
 FILLCELL_X32 FILLER_463_3359 ();
 FILLCELL_X32 FILLER_463_3391 ();
 FILLCELL_X32 FILLER_463_3423 ();
 FILLCELL_X32 FILLER_463_3455 ();
 FILLCELL_X32 FILLER_463_3487 ();
 FILLCELL_X32 FILLER_463_3519 ();
 FILLCELL_X32 FILLER_463_3551 ();
 FILLCELL_X32 FILLER_463_3583 ();
 FILLCELL_X32 FILLER_463_3615 ();
 FILLCELL_X32 FILLER_463_3647 ();
 FILLCELL_X32 FILLER_463_3679 ();
 FILLCELL_X16 FILLER_463_3711 ();
 FILLCELL_X8 FILLER_463_3727 ();
 FILLCELL_X2 FILLER_463_3735 ();
 FILLCELL_X1 FILLER_463_3737 ();
 FILLCELL_X32 FILLER_464_1 ();
 FILLCELL_X32 FILLER_464_33 ();
 FILLCELL_X32 FILLER_464_65 ();
 FILLCELL_X32 FILLER_464_97 ();
 FILLCELL_X32 FILLER_464_129 ();
 FILLCELL_X32 FILLER_464_161 ();
 FILLCELL_X32 FILLER_464_193 ();
 FILLCELL_X32 FILLER_464_225 ();
 FILLCELL_X32 FILLER_464_257 ();
 FILLCELL_X32 FILLER_464_289 ();
 FILLCELL_X32 FILLER_464_321 ();
 FILLCELL_X32 FILLER_464_353 ();
 FILLCELL_X32 FILLER_464_385 ();
 FILLCELL_X32 FILLER_464_417 ();
 FILLCELL_X32 FILLER_464_449 ();
 FILLCELL_X32 FILLER_464_481 ();
 FILLCELL_X32 FILLER_464_513 ();
 FILLCELL_X32 FILLER_464_545 ();
 FILLCELL_X32 FILLER_464_577 ();
 FILLCELL_X16 FILLER_464_609 ();
 FILLCELL_X4 FILLER_464_625 ();
 FILLCELL_X2 FILLER_464_629 ();
 FILLCELL_X32 FILLER_464_632 ();
 FILLCELL_X32 FILLER_464_664 ();
 FILLCELL_X32 FILLER_464_696 ();
 FILLCELL_X32 FILLER_464_728 ();
 FILLCELL_X32 FILLER_464_760 ();
 FILLCELL_X32 FILLER_464_792 ();
 FILLCELL_X32 FILLER_464_824 ();
 FILLCELL_X32 FILLER_464_856 ();
 FILLCELL_X32 FILLER_464_888 ();
 FILLCELL_X32 FILLER_464_920 ();
 FILLCELL_X32 FILLER_464_952 ();
 FILLCELL_X32 FILLER_464_984 ();
 FILLCELL_X32 FILLER_464_1016 ();
 FILLCELL_X32 FILLER_464_1048 ();
 FILLCELL_X32 FILLER_464_1080 ();
 FILLCELL_X32 FILLER_464_1112 ();
 FILLCELL_X32 FILLER_464_1144 ();
 FILLCELL_X32 FILLER_464_1176 ();
 FILLCELL_X32 FILLER_464_1208 ();
 FILLCELL_X32 FILLER_464_1240 ();
 FILLCELL_X32 FILLER_464_1272 ();
 FILLCELL_X32 FILLER_464_1304 ();
 FILLCELL_X32 FILLER_464_1336 ();
 FILLCELL_X32 FILLER_464_1368 ();
 FILLCELL_X32 FILLER_464_1400 ();
 FILLCELL_X32 FILLER_464_1432 ();
 FILLCELL_X32 FILLER_464_1464 ();
 FILLCELL_X32 FILLER_464_1496 ();
 FILLCELL_X32 FILLER_464_1528 ();
 FILLCELL_X32 FILLER_464_1560 ();
 FILLCELL_X32 FILLER_464_1592 ();
 FILLCELL_X32 FILLER_464_1624 ();
 FILLCELL_X32 FILLER_464_1656 ();
 FILLCELL_X32 FILLER_464_1688 ();
 FILLCELL_X32 FILLER_464_1720 ();
 FILLCELL_X32 FILLER_464_1752 ();
 FILLCELL_X32 FILLER_464_1784 ();
 FILLCELL_X32 FILLER_464_1816 ();
 FILLCELL_X32 FILLER_464_1848 ();
 FILLCELL_X8 FILLER_464_1880 ();
 FILLCELL_X4 FILLER_464_1888 ();
 FILLCELL_X2 FILLER_464_1892 ();
 FILLCELL_X32 FILLER_464_1895 ();
 FILLCELL_X32 FILLER_464_1927 ();
 FILLCELL_X32 FILLER_464_1959 ();
 FILLCELL_X32 FILLER_464_1991 ();
 FILLCELL_X32 FILLER_464_2023 ();
 FILLCELL_X32 FILLER_464_2055 ();
 FILLCELL_X32 FILLER_464_2087 ();
 FILLCELL_X32 FILLER_464_2119 ();
 FILLCELL_X32 FILLER_464_2151 ();
 FILLCELL_X32 FILLER_464_2183 ();
 FILLCELL_X32 FILLER_464_2215 ();
 FILLCELL_X32 FILLER_464_2247 ();
 FILLCELL_X32 FILLER_464_2279 ();
 FILLCELL_X32 FILLER_464_2311 ();
 FILLCELL_X32 FILLER_464_2343 ();
 FILLCELL_X32 FILLER_464_2375 ();
 FILLCELL_X32 FILLER_464_2407 ();
 FILLCELL_X32 FILLER_464_2439 ();
 FILLCELL_X32 FILLER_464_2471 ();
 FILLCELL_X32 FILLER_464_2503 ();
 FILLCELL_X32 FILLER_464_2535 ();
 FILLCELL_X32 FILLER_464_2567 ();
 FILLCELL_X32 FILLER_464_2599 ();
 FILLCELL_X32 FILLER_464_2631 ();
 FILLCELL_X32 FILLER_464_2663 ();
 FILLCELL_X32 FILLER_464_2695 ();
 FILLCELL_X32 FILLER_464_2727 ();
 FILLCELL_X32 FILLER_464_2759 ();
 FILLCELL_X32 FILLER_464_2791 ();
 FILLCELL_X32 FILLER_464_2823 ();
 FILLCELL_X32 FILLER_464_2855 ();
 FILLCELL_X32 FILLER_464_2887 ();
 FILLCELL_X32 FILLER_464_2919 ();
 FILLCELL_X32 FILLER_464_2951 ();
 FILLCELL_X32 FILLER_464_2983 ();
 FILLCELL_X32 FILLER_464_3015 ();
 FILLCELL_X32 FILLER_464_3047 ();
 FILLCELL_X32 FILLER_464_3079 ();
 FILLCELL_X32 FILLER_464_3111 ();
 FILLCELL_X8 FILLER_464_3143 ();
 FILLCELL_X4 FILLER_464_3151 ();
 FILLCELL_X2 FILLER_464_3155 ();
 FILLCELL_X32 FILLER_464_3158 ();
 FILLCELL_X32 FILLER_464_3190 ();
 FILLCELL_X32 FILLER_464_3222 ();
 FILLCELL_X32 FILLER_464_3254 ();
 FILLCELL_X32 FILLER_464_3286 ();
 FILLCELL_X32 FILLER_464_3318 ();
 FILLCELL_X32 FILLER_464_3350 ();
 FILLCELL_X32 FILLER_464_3382 ();
 FILLCELL_X32 FILLER_464_3414 ();
 FILLCELL_X32 FILLER_464_3446 ();
 FILLCELL_X32 FILLER_464_3478 ();
 FILLCELL_X32 FILLER_464_3510 ();
 FILLCELL_X32 FILLER_464_3542 ();
 FILLCELL_X32 FILLER_464_3574 ();
 FILLCELL_X32 FILLER_464_3606 ();
 FILLCELL_X32 FILLER_464_3638 ();
 FILLCELL_X32 FILLER_464_3670 ();
 FILLCELL_X32 FILLER_464_3702 ();
 FILLCELL_X4 FILLER_464_3734 ();
 FILLCELL_X32 FILLER_465_1 ();
 FILLCELL_X32 FILLER_465_33 ();
 FILLCELL_X32 FILLER_465_65 ();
 FILLCELL_X32 FILLER_465_97 ();
 FILLCELL_X32 FILLER_465_129 ();
 FILLCELL_X32 FILLER_465_161 ();
 FILLCELL_X32 FILLER_465_193 ();
 FILLCELL_X32 FILLER_465_225 ();
 FILLCELL_X32 FILLER_465_257 ();
 FILLCELL_X32 FILLER_465_289 ();
 FILLCELL_X32 FILLER_465_321 ();
 FILLCELL_X32 FILLER_465_353 ();
 FILLCELL_X32 FILLER_465_385 ();
 FILLCELL_X32 FILLER_465_417 ();
 FILLCELL_X32 FILLER_465_449 ();
 FILLCELL_X32 FILLER_465_481 ();
 FILLCELL_X32 FILLER_465_513 ();
 FILLCELL_X32 FILLER_465_545 ();
 FILLCELL_X32 FILLER_465_577 ();
 FILLCELL_X32 FILLER_465_609 ();
 FILLCELL_X32 FILLER_465_641 ();
 FILLCELL_X32 FILLER_465_673 ();
 FILLCELL_X32 FILLER_465_705 ();
 FILLCELL_X32 FILLER_465_737 ();
 FILLCELL_X32 FILLER_465_769 ();
 FILLCELL_X32 FILLER_465_801 ();
 FILLCELL_X32 FILLER_465_833 ();
 FILLCELL_X32 FILLER_465_865 ();
 FILLCELL_X32 FILLER_465_897 ();
 FILLCELL_X32 FILLER_465_929 ();
 FILLCELL_X32 FILLER_465_961 ();
 FILLCELL_X32 FILLER_465_993 ();
 FILLCELL_X32 FILLER_465_1025 ();
 FILLCELL_X32 FILLER_465_1057 ();
 FILLCELL_X32 FILLER_465_1089 ();
 FILLCELL_X32 FILLER_465_1121 ();
 FILLCELL_X32 FILLER_465_1153 ();
 FILLCELL_X32 FILLER_465_1185 ();
 FILLCELL_X32 FILLER_465_1217 ();
 FILLCELL_X8 FILLER_465_1249 ();
 FILLCELL_X4 FILLER_465_1257 ();
 FILLCELL_X2 FILLER_465_1261 ();
 FILLCELL_X32 FILLER_465_1264 ();
 FILLCELL_X32 FILLER_465_1296 ();
 FILLCELL_X32 FILLER_465_1328 ();
 FILLCELL_X32 FILLER_465_1360 ();
 FILLCELL_X32 FILLER_465_1392 ();
 FILLCELL_X32 FILLER_465_1424 ();
 FILLCELL_X32 FILLER_465_1456 ();
 FILLCELL_X32 FILLER_465_1488 ();
 FILLCELL_X32 FILLER_465_1520 ();
 FILLCELL_X32 FILLER_465_1552 ();
 FILLCELL_X32 FILLER_465_1584 ();
 FILLCELL_X32 FILLER_465_1616 ();
 FILLCELL_X32 FILLER_465_1648 ();
 FILLCELL_X32 FILLER_465_1680 ();
 FILLCELL_X32 FILLER_465_1712 ();
 FILLCELL_X32 FILLER_465_1744 ();
 FILLCELL_X32 FILLER_465_1776 ();
 FILLCELL_X32 FILLER_465_1808 ();
 FILLCELL_X32 FILLER_465_1840 ();
 FILLCELL_X32 FILLER_465_1872 ();
 FILLCELL_X32 FILLER_465_1904 ();
 FILLCELL_X32 FILLER_465_1936 ();
 FILLCELL_X32 FILLER_465_1968 ();
 FILLCELL_X32 FILLER_465_2000 ();
 FILLCELL_X32 FILLER_465_2032 ();
 FILLCELL_X32 FILLER_465_2064 ();
 FILLCELL_X32 FILLER_465_2096 ();
 FILLCELL_X32 FILLER_465_2128 ();
 FILLCELL_X32 FILLER_465_2160 ();
 FILLCELL_X32 FILLER_465_2192 ();
 FILLCELL_X32 FILLER_465_2224 ();
 FILLCELL_X32 FILLER_465_2256 ();
 FILLCELL_X32 FILLER_465_2288 ();
 FILLCELL_X32 FILLER_465_2320 ();
 FILLCELL_X32 FILLER_465_2352 ();
 FILLCELL_X32 FILLER_465_2384 ();
 FILLCELL_X32 FILLER_465_2416 ();
 FILLCELL_X32 FILLER_465_2448 ();
 FILLCELL_X32 FILLER_465_2480 ();
 FILLCELL_X8 FILLER_465_2512 ();
 FILLCELL_X4 FILLER_465_2520 ();
 FILLCELL_X2 FILLER_465_2524 ();
 FILLCELL_X32 FILLER_465_2527 ();
 FILLCELL_X32 FILLER_465_2559 ();
 FILLCELL_X32 FILLER_465_2591 ();
 FILLCELL_X32 FILLER_465_2623 ();
 FILLCELL_X32 FILLER_465_2655 ();
 FILLCELL_X32 FILLER_465_2687 ();
 FILLCELL_X32 FILLER_465_2719 ();
 FILLCELL_X32 FILLER_465_2751 ();
 FILLCELL_X32 FILLER_465_2783 ();
 FILLCELL_X32 FILLER_465_2815 ();
 FILLCELL_X32 FILLER_465_2847 ();
 FILLCELL_X32 FILLER_465_2879 ();
 FILLCELL_X32 FILLER_465_2911 ();
 FILLCELL_X32 FILLER_465_2943 ();
 FILLCELL_X32 FILLER_465_2975 ();
 FILLCELL_X32 FILLER_465_3007 ();
 FILLCELL_X32 FILLER_465_3039 ();
 FILLCELL_X32 FILLER_465_3071 ();
 FILLCELL_X32 FILLER_465_3103 ();
 FILLCELL_X32 FILLER_465_3135 ();
 FILLCELL_X32 FILLER_465_3167 ();
 FILLCELL_X32 FILLER_465_3199 ();
 FILLCELL_X32 FILLER_465_3231 ();
 FILLCELL_X32 FILLER_465_3263 ();
 FILLCELL_X32 FILLER_465_3295 ();
 FILLCELL_X32 FILLER_465_3327 ();
 FILLCELL_X32 FILLER_465_3359 ();
 FILLCELL_X32 FILLER_465_3391 ();
 FILLCELL_X32 FILLER_465_3423 ();
 FILLCELL_X32 FILLER_465_3455 ();
 FILLCELL_X32 FILLER_465_3487 ();
 FILLCELL_X32 FILLER_465_3519 ();
 FILLCELL_X32 FILLER_465_3551 ();
 FILLCELL_X32 FILLER_465_3583 ();
 FILLCELL_X32 FILLER_465_3615 ();
 FILLCELL_X32 FILLER_465_3647 ();
 FILLCELL_X32 FILLER_465_3679 ();
 FILLCELL_X16 FILLER_465_3711 ();
 FILLCELL_X8 FILLER_465_3727 ();
 FILLCELL_X2 FILLER_465_3735 ();
 FILLCELL_X1 FILLER_465_3737 ();
 FILLCELL_X32 FILLER_466_1 ();
 FILLCELL_X32 FILLER_466_33 ();
 FILLCELL_X32 FILLER_466_65 ();
 FILLCELL_X32 FILLER_466_97 ();
 FILLCELL_X32 FILLER_466_129 ();
 FILLCELL_X32 FILLER_466_161 ();
 FILLCELL_X32 FILLER_466_193 ();
 FILLCELL_X32 FILLER_466_225 ();
 FILLCELL_X32 FILLER_466_257 ();
 FILLCELL_X32 FILLER_466_289 ();
 FILLCELL_X32 FILLER_466_321 ();
 FILLCELL_X32 FILLER_466_353 ();
 FILLCELL_X32 FILLER_466_385 ();
 FILLCELL_X32 FILLER_466_417 ();
 FILLCELL_X32 FILLER_466_449 ();
 FILLCELL_X32 FILLER_466_481 ();
 FILLCELL_X32 FILLER_466_513 ();
 FILLCELL_X32 FILLER_466_545 ();
 FILLCELL_X32 FILLER_466_577 ();
 FILLCELL_X16 FILLER_466_609 ();
 FILLCELL_X4 FILLER_466_625 ();
 FILLCELL_X2 FILLER_466_629 ();
 FILLCELL_X32 FILLER_466_632 ();
 FILLCELL_X32 FILLER_466_664 ();
 FILLCELL_X32 FILLER_466_696 ();
 FILLCELL_X32 FILLER_466_728 ();
 FILLCELL_X32 FILLER_466_760 ();
 FILLCELL_X32 FILLER_466_792 ();
 FILLCELL_X32 FILLER_466_824 ();
 FILLCELL_X32 FILLER_466_856 ();
 FILLCELL_X32 FILLER_466_888 ();
 FILLCELL_X32 FILLER_466_920 ();
 FILLCELL_X32 FILLER_466_952 ();
 FILLCELL_X32 FILLER_466_984 ();
 FILLCELL_X32 FILLER_466_1016 ();
 FILLCELL_X32 FILLER_466_1048 ();
 FILLCELL_X32 FILLER_466_1080 ();
 FILLCELL_X32 FILLER_466_1112 ();
 FILLCELL_X32 FILLER_466_1144 ();
 FILLCELL_X32 FILLER_466_1176 ();
 FILLCELL_X32 FILLER_466_1208 ();
 FILLCELL_X32 FILLER_466_1240 ();
 FILLCELL_X32 FILLER_466_1272 ();
 FILLCELL_X32 FILLER_466_1304 ();
 FILLCELL_X32 FILLER_466_1336 ();
 FILLCELL_X32 FILLER_466_1368 ();
 FILLCELL_X32 FILLER_466_1400 ();
 FILLCELL_X32 FILLER_466_1432 ();
 FILLCELL_X32 FILLER_466_1464 ();
 FILLCELL_X32 FILLER_466_1496 ();
 FILLCELL_X32 FILLER_466_1528 ();
 FILLCELL_X32 FILLER_466_1560 ();
 FILLCELL_X32 FILLER_466_1592 ();
 FILLCELL_X32 FILLER_466_1624 ();
 FILLCELL_X32 FILLER_466_1656 ();
 FILLCELL_X32 FILLER_466_1688 ();
 FILLCELL_X32 FILLER_466_1720 ();
 FILLCELL_X32 FILLER_466_1752 ();
 FILLCELL_X32 FILLER_466_1784 ();
 FILLCELL_X32 FILLER_466_1816 ();
 FILLCELL_X32 FILLER_466_1848 ();
 FILLCELL_X8 FILLER_466_1880 ();
 FILLCELL_X4 FILLER_466_1888 ();
 FILLCELL_X2 FILLER_466_1892 ();
 FILLCELL_X32 FILLER_466_1895 ();
 FILLCELL_X32 FILLER_466_1927 ();
 FILLCELL_X32 FILLER_466_1959 ();
 FILLCELL_X32 FILLER_466_1991 ();
 FILLCELL_X32 FILLER_466_2023 ();
 FILLCELL_X32 FILLER_466_2055 ();
 FILLCELL_X32 FILLER_466_2087 ();
 FILLCELL_X32 FILLER_466_2119 ();
 FILLCELL_X32 FILLER_466_2151 ();
 FILLCELL_X32 FILLER_466_2183 ();
 FILLCELL_X32 FILLER_466_2215 ();
 FILLCELL_X32 FILLER_466_2247 ();
 FILLCELL_X32 FILLER_466_2279 ();
 FILLCELL_X32 FILLER_466_2311 ();
 FILLCELL_X32 FILLER_466_2343 ();
 FILLCELL_X32 FILLER_466_2375 ();
 FILLCELL_X32 FILLER_466_2407 ();
 FILLCELL_X32 FILLER_466_2439 ();
 FILLCELL_X32 FILLER_466_2471 ();
 FILLCELL_X32 FILLER_466_2503 ();
 FILLCELL_X32 FILLER_466_2535 ();
 FILLCELL_X32 FILLER_466_2567 ();
 FILLCELL_X32 FILLER_466_2599 ();
 FILLCELL_X32 FILLER_466_2631 ();
 FILLCELL_X32 FILLER_466_2663 ();
 FILLCELL_X32 FILLER_466_2695 ();
 FILLCELL_X32 FILLER_466_2727 ();
 FILLCELL_X32 FILLER_466_2759 ();
 FILLCELL_X32 FILLER_466_2791 ();
 FILLCELL_X32 FILLER_466_2823 ();
 FILLCELL_X32 FILLER_466_2855 ();
 FILLCELL_X32 FILLER_466_2887 ();
 FILLCELL_X32 FILLER_466_2919 ();
 FILLCELL_X32 FILLER_466_2951 ();
 FILLCELL_X32 FILLER_466_2983 ();
 FILLCELL_X32 FILLER_466_3015 ();
 FILLCELL_X32 FILLER_466_3047 ();
 FILLCELL_X32 FILLER_466_3079 ();
 FILLCELL_X32 FILLER_466_3111 ();
 FILLCELL_X8 FILLER_466_3143 ();
 FILLCELL_X4 FILLER_466_3151 ();
 FILLCELL_X2 FILLER_466_3155 ();
 FILLCELL_X32 FILLER_466_3158 ();
 FILLCELL_X32 FILLER_466_3190 ();
 FILLCELL_X32 FILLER_466_3222 ();
 FILLCELL_X32 FILLER_466_3254 ();
 FILLCELL_X32 FILLER_466_3286 ();
 FILLCELL_X32 FILLER_466_3318 ();
 FILLCELL_X32 FILLER_466_3350 ();
 FILLCELL_X32 FILLER_466_3382 ();
 FILLCELL_X32 FILLER_466_3414 ();
 FILLCELL_X32 FILLER_466_3446 ();
 FILLCELL_X32 FILLER_466_3478 ();
 FILLCELL_X32 FILLER_466_3510 ();
 FILLCELL_X32 FILLER_466_3542 ();
 FILLCELL_X32 FILLER_466_3574 ();
 FILLCELL_X32 FILLER_466_3606 ();
 FILLCELL_X32 FILLER_466_3638 ();
 FILLCELL_X32 FILLER_466_3670 ();
 FILLCELL_X32 FILLER_466_3702 ();
 FILLCELL_X4 FILLER_466_3734 ();
 FILLCELL_X32 FILLER_467_1 ();
 FILLCELL_X32 FILLER_467_33 ();
 FILLCELL_X32 FILLER_467_65 ();
 FILLCELL_X32 FILLER_467_97 ();
 FILLCELL_X32 FILLER_467_129 ();
 FILLCELL_X32 FILLER_467_161 ();
 FILLCELL_X32 FILLER_467_193 ();
 FILLCELL_X32 FILLER_467_225 ();
 FILLCELL_X32 FILLER_467_257 ();
 FILLCELL_X32 FILLER_467_289 ();
 FILLCELL_X32 FILLER_467_321 ();
 FILLCELL_X32 FILLER_467_353 ();
 FILLCELL_X32 FILLER_467_385 ();
 FILLCELL_X32 FILLER_467_417 ();
 FILLCELL_X32 FILLER_467_449 ();
 FILLCELL_X32 FILLER_467_481 ();
 FILLCELL_X32 FILLER_467_513 ();
 FILLCELL_X32 FILLER_467_545 ();
 FILLCELL_X32 FILLER_467_577 ();
 FILLCELL_X32 FILLER_467_609 ();
 FILLCELL_X32 FILLER_467_641 ();
 FILLCELL_X32 FILLER_467_673 ();
 FILLCELL_X32 FILLER_467_705 ();
 FILLCELL_X32 FILLER_467_737 ();
 FILLCELL_X32 FILLER_467_769 ();
 FILLCELL_X32 FILLER_467_801 ();
 FILLCELL_X32 FILLER_467_833 ();
 FILLCELL_X32 FILLER_467_865 ();
 FILLCELL_X32 FILLER_467_897 ();
 FILLCELL_X32 FILLER_467_929 ();
 FILLCELL_X32 FILLER_467_961 ();
 FILLCELL_X32 FILLER_467_993 ();
 FILLCELL_X32 FILLER_467_1025 ();
 FILLCELL_X32 FILLER_467_1057 ();
 FILLCELL_X32 FILLER_467_1089 ();
 FILLCELL_X32 FILLER_467_1121 ();
 FILLCELL_X32 FILLER_467_1153 ();
 FILLCELL_X32 FILLER_467_1185 ();
 FILLCELL_X32 FILLER_467_1217 ();
 FILLCELL_X8 FILLER_467_1249 ();
 FILLCELL_X4 FILLER_467_1257 ();
 FILLCELL_X2 FILLER_467_1261 ();
 FILLCELL_X32 FILLER_467_1264 ();
 FILLCELL_X32 FILLER_467_1296 ();
 FILLCELL_X32 FILLER_467_1328 ();
 FILLCELL_X32 FILLER_467_1360 ();
 FILLCELL_X32 FILLER_467_1392 ();
 FILLCELL_X32 FILLER_467_1424 ();
 FILLCELL_X32 FILLER_467_1456 ();
 FILLCELL_X32 FILLER_467_1488 ();
 FILLCELL_X32 FILLER_467_1520 ();
 FILLCELL_X32 FILLER_467_1552 ();
 FILLCELL_X32 FILLER_467_1584 ();
 FILLCELL_X32 FILLER_467_1616 ();
 FILLCELL_X32 FILLER_467_1648 ();
 FILLCELL_X32 FILLER_467_1680 ();
 FILLCELL_X32 FILLER_467_1712 ();
 FILLCELL_X32 FILLER_467_1744 ();
 FILLCELL_X32 FILLER_467_1776 ();
 FILLCELL_X32 FILLER_467_1808 ();
 FILLCELL_X32 FILLER_467_1840 ();
 FILLCELL_X32 FILLER_467_1872 ();
 FILLCELL_X32 FILLER_467_1904 ();
 FILLCELL_X32 FILLER_467_1936 ();
 FILLCELL_X32 FILLER_467_1968 ();
 FILLCELL_X32 FILLER_467_2000 ();
 FILLCELL_X32 FILLER_467_2032 ();
 FILLCELL_X32 FILLER_467_2064 ();
 FILLCELL_X32 FILLER_467_2096 ();
 FILLCELL_X32 FILLER_467_2128 ();
 FILLCELL_X32 FILLER_467_2160 ();
 FILLCELL_X32 FILLER_467_2192 ();
 FILLCELL_X32 FILLER_467_2224 ();
 FILLCELL_X32 FILLER_467_2256 ();
 FILLCELL_X32 FILLER_467_2288 ();
 FILLCELL_X32 FILLER_467_2320 ();
 FILLCELL_X32 FILLER_467_2352 ();
 FILLCELL_X32 FILLER_467_2384 ();
 FILLCELL_X32 FILLER_467_2416 ();
 FILLCELL_X32 FILLER_467_2448 ();
 FILLCELL_X32 FILLER_467_2480 ();
 FILLCELL_X8 FILLER_467_2512 ();
 FILLCELL_X4 FILLER_467_2520 ();
 FILLCELL_X2 FILLER_467_2524 ();
 FILLCELL_X32 FILLER_467_2527 ();
 FILLCELL_X32 FILLER_467_2559 ();
 FILLCELL_X32 FILLER_467_2591 ();
 FILLCELL_X32 FILLER_467_2623 ();
 FILLCELL_X32 FILLER_467_2655 ();
 FILLCELL_X32 FILLER_467_2687 ();
 FILLCELL_X32 FILLER_467_2719 ();
 FILLCELL_X32 FILLER_467_2751 ();
 FILLCELL_X32 FILLER_467_2783 ();
 FILLCELL_X32 FILLER_467_2815 ();
 FILLCELL_X32 FILLER_467_2847 ();
 FILLCELL_X32 FILLER_467_2879 ();
 FILLCELL_X32 FILLER_467_2911 ();
 FILLCELL_X32 FILLER_467_2943 ();
 FILLCELL_X32 FILLER_467_2975 ();
 FILLCELL_X32 FILLER_467_3007 ();
 FILLCELL_X32 FILLER_467_3039 ();
 FILLCELL_X32 FILLER_467_3071 ();
 FILLCELL_X32 FILLER_467_3103 ();
 FILLCELL_X32 FILLER_467_3135 ();
 FILLCELL_X32 FILLER_467_3167 ();
 FILLCELL_X32 FILLER_467_3199 ();
 FILLCELL_X32 FILLER_467_3231 ();
 FILLCELL_X32 FILLER_467_3263 ();
 FILLCELL_X32 FILLER_467_3295 ();
 FILLCELL_X32 FILLER_467_3327 ();
 FILLCELL_X32 FILLER_467_3359 ();
 FILLCELL_X32 FILLER_467_3391 ();
 FILLCELL_X32 FILLER_467_3423 ();
 FILLCELL_X32 FILLER_467_3455 ();
 FILLCELL_X32 FILLER_467_3487 ();
 FILLCELL_X32 FILLER_467_3519 ();
 FILLCELL_X32 FILLER_467_3551 ();
 FILLCELL_X32 FILLER_467_3583 ();
 FILLCELL_X32 FILLER_467_3615 ();
 FILLCELL_X32 FILLER_467_3647 ();
 FILLCELL_X32 FILLER_467_3679 ();
 FILLCELL_X16 FILLER_467_3711 ();
 FILLCELL_X8 FILLER_467_3727 ();
 FILLCELL_X2 FILLER_467_3735 ();
 FILLCELL_X1 FILLER_467_3737 ();
 FILLCELL_X32 FILLER_468_1 ();
 FILLCELL_X32 FILLER_468_33 ();
 FILLCELL_X32 FILLER_468_65 ();
 FILLCELL_X32 FILLER_468_97 ();
 FILLCELL_X32 FILLER_468_129 ();
 FILLCELL_X32 FILLER_468_161 ();
 FILLCELL_X32 FILLER_468_193 ();
 FILLCELL_X32 FILLER_468_225 ();
 FILLCELL_X32 FILLER_468_257 ();
 FILLCELL_X32 FILLER_468_289 ();
 FILLCELL_X32 FILLER_468_321 ();
 FILLCELL_X32 FILLER_468_353 ();
 FILLCELL_X32 FILLER_468_385 ();
 FILLCELL_X32 FILLER_468_417 ();
 FILLCELL_X32 FILLER_468_449 ();
 FILLCELL_X32 FILLER_468_481 ();
 FILLCELL_X32 FILLER_468_513 ();
 FILLCELL_X32 FILLER_468_545 ();
 FILLCELL_X32 FILLER_468_577 ();
 FILLCELL_X16 FILLER_468_609 ();
 FILLCELL_X4 FILLER_468_625 ();
 FILLCELL_X2 FILLER_468_629 ();
 FILLCELL_X32 FILLER_468_632 ();
 FILLCELL_X32 FILLER_468_664 ();
 FILLCELL_X32 FILLER_468_696 ();
 FILLCELL_X32 FILLER_468_728 ();
 FILLCELL_X32 FILLER_468_760 ();
 FILLCELL_X32 FILLER_468_792 ();
 FILLCELL_X32 FILLER_468_824 ();
 FILLCELL_X32 FILLER_468_856 ();
 FILLCELL_X32 FILLER_468_888 ();
 FILLCELL_X32 FILLER_468_920 ();
 FILLCELL_X32 FILLER_468_952 ();
 FILLCELL_X32 FILLER_468_984 ();
 FILLCELL_X32 FILLER_468_1016 ();
 FILLCELL_X32 FILLER_468_1048 ();
 FILLCELL_X32 FILLER_468_1080 ();
 FILLCELL_X32 FILLER_468_1112 ();
 FILLCELL_X32 FILLER_468_1144 ();
 FILLCELL_X32 FILLER_468_1176 ();
 FILLCELL_X32 FILLER_468_1208 ();
 FILLCELL_X32 FILLER_468_1240 ();
 FILLCELL_X32 FILLER_468_1272 ();
 FILLCELL_X32 FILLER_468_1304 ();
 FILLCELL_X32 FILLER_468_1336 ();
 FILLCELL_X32 FILLER_468_1368 ();
 FILLCELL_X32 FILLER_468_1400 ();
 FILLCELL_X32 FILLER_468_1432 ();
 FILLCELL_X32 FILLER_468_1464 ();
 FILLCELL_X32 FILLER_468_1496 ();
 FILLCELL_X32 FILLER_468_1528 ();
 FILLCELL_X32 FILLER_468_1560 ();
 FILLCELL_X32 FILLER_468_1592 ();
 FILLCELL_X32 FILLER_468_1624 ();
 FILLCELL_X32 FILLER_468_1656 ();
 FILLCELL_X32 FILLER_468_1688 ();
 FILLCELL_X32 FILLER_468_1720 ();
 FILLCELL_X32 FILLER_468_1752 ();
 FILLCELL_X32 FILLER_468_1784 ();
 FILLCELL_X32 FILLER_468_1816 ();
 FILLCELL_X32 FILLER_468_1848 ();
 FILLCELL_X8 FILLER_468_1880 ();
 FILLCELL_X4 FILLER_468_1888 ();
 FILLCELL_X2 FILLER_468_1892 ();
 FILLCELL_X32 FILLER_468_1895 ();
 FILLCELL_X32 FILLER_468_1927 ();
 FILLCELL_X32 FILLER_468_1959 ();
 FILLCELL_X32 FILLER_468_1991 ();
 FILLCELL_X32 FILLER_468_2023 ();
 FILLCELL_X32 FILLER_468_2055 ();
 FILLCELL_X32 FILLER_468_2087 ();
 FILLCELL_X32 FILLER_468_2119 ();
 FILLCELL_X32 FILLER_468_2151 ();
 FILLCELL_X32 FILLER_468_2183 ();
 FILLCELL_X32 FILLER_468_2215 ();
 FILLCELL_X32 FILLER_468_2247 ();
 FILLCELL_X32 FILLER_468_2279 ();
 FILLCELL_X32 FILLER_468_2311 ();
 FILLCELL_X32 FILLER_468_2343 ();
 FILLCELL_X32 FILLER_468_2375 ();
 FILLCELL_X32 FILLER_468_2407 ();
 FILLCELL_X32 FILLER_468_2439 ();
 FILLCELL_X32 FILLER_468_2471 ();
 FILLCELL_X32 FILLER_468_2503 ();
 FILLCELL_X32 FILLER_468_2535 ();
 FILLCELL_X32 FILLER_468_2567 ();
 FILLCELL_X32 FILLER_468_2599 ();
 FILLCELL_X32 FILLER_468_2631 ();
 FILLCELL_X32 FILLER_468_2663 ();
 FILLCELL_X32 FILLER_468_2695 ();
 FILLCELL_X32 FILLER_468_2727 ();
 FILLCELL_X32 FILLER_468_2759 ();
 FILLCELL_X32 FILLER_468_2791 ();
 FILLCELL_X32 FILLER_468_2823 ();
 FILLCELL_X32 FILLER_468_2855 ();
 FILLCELL_X32 FILLER_468_2887 ();
 FILLCELL_X32 FILLER_468_2919 ();
 FILLCELL_X32 FILLER_468_2951 ();
 FILLCELL_X32 FILLER_468_2983 ();
 FILLCELL_X32 FILLER_468_3015 ();
 FILLCELL_X32 FILLER_468_3047 ();
 FILLCELL_X32 FILLER_468_3079 ();
 FILLCELL_X32 FILLER_468_3111 ();
 FILLCELL_X8 FILLER_468_3143 ();
 FILLCELL_X4 FILLER_468_3151 ();
 FILLCELL_X2 FILLER_468_3155 ();
 FILLCELL_X32 FILLER_468_3158 ();
 FILLCELL_X32 FILLER_468_3190 ();
 FILLCELL_X32 FILLER_468_3222 ();
 FILLCELL_X32 FILLER_468_3254 ();
 FILLCELL_X32 FILLER_468_3286 ();
 FILLCELL_X32 FILLER_468_3318 ();
 FILLCELL_X32 FILLER_468_3350 ();
 FILLCELL_X32 FILLER_468_3382 ();
 FILLCELL_X32 FILLER_468_3414 ();
 FILLCELL_X32 FILLER_468_3446 ();
 FILLCELL_X32 FILLER_468_3478 ();
 FILLCELL_X32 FILLER_468_3510 ();
 FILLCELL_X32 FILLER_468_3542 ();
 FILLCELL_X32 FILLER_468_3574 ();
 FILLCELL_X32 FILLER_468_3606 ();
 FILLCELL_X32 FILLER_468_3638 ();
 FILLCELL_X32 FILLER_468_3670 ();
 FILLCELL_X32 FILLER_468_3702 ();
 FILLCELL_X4 FILLER_468_3734 ();
 FILLCELL_X32 FILLER_469_1 ();
 FILLCELL_X32 FILLER_469_33 ();
 FILLCELL_X32 FILLER_469_65 ();
 FILLCELL_X32 FILLER_469_97 ();
 FILLCELL_X32 FILLER_469_129 ();
 FILLCELL_X32 FILLER_469_161 ();
 FILLCELL_X32 FILLER_469_193 ();
 FILLCELL_X32 FILLER_469_225 ();
 FILLCELL_X32 FILLER_469_257 ();
 FILLCELL_X32 FILLER_469_289 ();
 FILLCELL_X32 FILLER_469_321 ();
 FILLCELL_X32 FILLER_469_353 ();
 FILLCELL_X32 FILLER_469_385 ();
 FILLCELL_X32 FILLER_469_417 ();
 FILLCELL_X32 FILLER_469_449 ();
 FILLCELL_X32 FILLER_469_481 ();
 FILLCELL_X32 FILLER_469_513 ();
 FILLCELL_X32 FILLER_469_545 ();
 FILLCELL_X32 FILLER_469_577 ();
 FILLCELL_X32 FILLER_469_609 ();
 FILLCELL_X32 FILLER_469_641 ();
 FILLCELL_X32 FILLER_469_673 ();
 FILLCELL_X32 FILLER_469_705 ();
 FILLCELL_X32 FILLER_469_737 ();
 FILLCELL_X32 FILLER_469_769 ();
 FILLCELL_X32 FILLER_469_801 ();
 FILLCELL_X32 FILLER_469_833 ();
 FILLCELL_X32 FILLER_469_865 ();
 FILLCELL_X32 FILLER_469_897 ();
 FILLCELL_X32 FILLER_469_929 ();
 FILLCELL_X32 FILLER_469_961 ();
 FILLCELL_X32 FILLER_469_993 ();
 FILLCELL_X32 FILLER_469_1025 ();
 FILLCELL_X32 FILLER_469_1057 ();
 FILLCELL_X32 FILLER_469_1089 ();
 FILLCELL_X32 FILLER_469_1121 ();
 FILLCELL_X32 FILLER_469_1153 ();
 FILLCELL_X32 FILLER_469_1185 ();
 FILLCELL_X32 FILLER_469_1217 ();
 FILLCELL_X8 FILLER_469_1249 ();
 FILLCELL_X4 FILLER_469_1257 ();
 FILLCELL_X2 FILLER_469_1261 ();
 FILLCELL_X32 FILLER_469_1264 ();
 FILLCELL_X32 FILLER_469_1296 ();
 FILLCELL_X32 FILLER_469_1328 ();
 FILLCELL_X32 FILLER_469_1360 ();
 FILLCELL_X32 FILLER_469_1392 ();
 FILLCELL_X32 FILLER_469_1424 ();
 FILLCELL_X32 FILLER_469_1456 ();
 FILLCELL_X32 FILLER_469_1488 ();
 FILLCELL_X32 FILLER_469_1520 ();
 FILLCELL_X32 FILLER_469_1552 ();
 FILLCELL_X32 FILLER_469_1584 ();
 FILLCELL_X32 FILLER_469_1616 ();
 FILLCELL_X32 FILLER_469_1648 ();
 FILLCELL_X32 FILLER_469_1680 ();
 FILLCELL_X32 FILLER_469_1712 ();
 FILLCELL_X32 FILLER_469_1744 ();
 FILLCELL_X32 FILLER_469_1776 ();
 FILLCELL_X32 FILLER_469_1808 ();
 FILLCELL_X32 FILLER_469_1840 ();
 FILLCELL_X32 FILLER_469_1872 ();
 FILLCELL_X32 FILLER_469_1904 ();
 FILLCELL_X32 FILLER_469_1936 ();
 FILLCELL_X32 FILLER_469_1968 ();
 FILLCELL_X32 FILLER_469_2000 ();
 FILLCELL_X32 FILLER_469_2032 ();
 FILLCELL_X32 FILLER_469_2064 ();
 FILLCELL_X32 FILLER_469_2096 ();
 FILLCELL_X32 FILLER_469_2128 ();
 FILLCELL_X32 FILLER_469_2160 ();
 FILLCELL_X32 FILLER_469_2192 ();
 FILLCELL_X32 FILLER_469_2224 ();
 FILLCELL_X32 FILLER_469_2256 ();
 FILLCELL_X32 FILLER_469_2288 ();
 FILLCELL_X32 FILLER_469_2320 ();
 FILLCELL_X32 FILLER_469_2352 ();
 FILLCELL_X32 FILLER_469_2384 ();
 FILLCELL_X32 FILLER_469_2416 ();
 FILLCELL_X32 FILLER_469_2448 ();
 FILLCELL_X32 FILLER_469_2480 ();
 FILLCELL_X8 FILLER_469_2512 ();
 FILLCELL_X4 FILLER_469_2520 ();
 FILLCELL_X2 FILLER_469_2524 ();
 FILLCELL_X32 FILLER_469_2527 ();
 FILLCELL_X32 FILLER_469_2559 ();
 FILLCELL_X32 FILLER_469_2591 ();
 FILLCELL_X32 FILLER_469_2623 ();
 FILLCELL_X32 FILLER_469_2655 ();
 FILLCELL_X32 FILLER_469_2687 ();
 FILLCELL_X32 FILLER_469_2719 ();
 FILLCELL_X32 FILLER_469_2751 ();
 FILLCELL_X32 FILLER_469_2783 ();
 FILLCELL_X32 FILLER_469_2815 ();
 FILLCELL_X32 FILLER_469_2847 ();
 FILLCELL_X32 FILLER_469_2879 ();
 FILLCELL_X32 FILLER_469_2911 ();
 FILLCELL_X32 FILLER_469_2943 ();
 FILLCELL_X32 FILLER_469_2975 ();
 FILLCELL_X32 FILLER_469_3007 ();
 FILLCELL_X32 FILLER_469_3039 ();
 FILLCELL_X32 FILLER_469_3071 ();
 FILLCELL_X32 FILLER_469_3103 ();
 FILLCELL_X32 FILLER_469_3135 ();
 FILLCELL_X32 FILLER_469_3167 ();
 FILLCELL_X32 FILLER_469_3199 ();
 FILLCELL_X32 FILLER_469_3231 ();
 FILLCELL_X32 FILLER_469_3263 ();
 FILLCELL_X32 FILLER_469_3295 ();
 FILLCELL_X32 FILLER_469_3327 ();
 FILLCELL_X32 FILLER_469_3359 ();
 FILLCELL_X32 FILLER_469_3391 ();
 FILLCELL_X32 FILLER_469_3423 ();
 FILLCELL_X32 FILLER_469_3455 ();
 FILLCELL_X32 FILLER_469_3487 ();
 FILLCELL_X32 FILLER_469_3519 ();
 FILLCELL_X32 FILLER_469_3551 ();
 FILLCELL_X32 FILLER_469_3583 ();
 FILLCELL_X32 FILLER_469_3615 ();
 FILLCELL_X32 FILLER_469_3647 ();
 FILLCELL_X32 FILLER_469_3679 ();
 FILLCELL_X16 FILLER_469_3711 ();
 FILLCELL_X8 FILLER_469_3727 ();
 FILLCELL_X2 FILLER_469_3735 ();
 FILLCELL_X1 FILLER_469_3737 ();
 FILLCELL_X32 FILLER_470_1 ();
 FILLCELL_X32 FILLER_470_33 ();
 FILLCELL_X32 FILLER_470_65 ();
 FILLCELL_X32 FILLER_470_97 ();
 FILLCELL_X32 FILLER_470_129 ();
 FILLCELL_X32 FILLER_470_161 ();
 FILLCELL_X32 FILLER_470_193 ();
 FILLCELL_X32 FILLER_470_225 ();
 FILLCELL_X32 FILLER_470_257 ();
 FILLCELL_X32 FILLER_470_289 ();
 FILLCELL_X32 FILLER_470_321 ();
 FILLCELL_X32 FILLER_470_353 ();
 FILLCELL_X32 FILLER_470_385 ();
 FILLCELL_X32 FILLER_470_417 ();
 FILLCELL_X32 FILLER_470_449 ();
 FILLCELL_X32 FILLER_470_481 ();
 FILLCELL_X32 FILLER_470_513 ();
 FILLCELL_X32 FILLER_470_545 ();
 FILLCELL_X32 FILLER_470_577 ();
 FILLCELL_X16 FILLER_470_609 ();
 FILLCELL_X4 FILLER_470_625 ();
 FILLCELL_X2 FILLER_470_629 ();
 FILLCELL_X32 FILLER_470_632 ();
 FILLCELL_X32 FILLER_470_664 ();
 FILLCELL_X32 FILLER_470_696 ();
 FILLCELL_X32 FILLER_470_728 ();
 FILLCELL_X32 FILLER_470_760 ();
 FILLCELL_X32 FILLER_470_792 ();
 FILLCELL_X32 FILLER_470_824 ();
 FILLCELL_X32 FILLER_470_856 ();
 FILLCELL_X32 FILLER_470_888 ();
 FILLCELL_X32 FILLER_470_920 ();
 FILLCELL_X32 FILLER_470_952 ();
 FILLCELL_X32 FILLER_470_984 ();
 FILLCELL_X32 FILLER_470_1016 ();
 FILLCELL_X32 FILLER_470_1048 ();
 FILLCELL_X32 FILLER_470_1080 ();
 FILLCELL_X32 FILLER_470_1112 ();
 FILLCELL_X32 FILLER_470_1144 ();
 FILLCELL_X32 FILLER_470_1176 ();
 FILLCELL_X32 FILLER_470_1208 ();
 FILLCELL_X32 FILLER_470_1240 ();
 FILLCELL_X32 FILLER_470_1272 ();
 FILLCELL_X32 FILLER_470_1304 ();
 FILLCELL_X32 FILLER_470_1336 ();
 FILLCELL_X32 FILLER_470_1368 ();
 FILLCELL_X32 FILLER_470_1400 ();
 FILLCELL_X32 FILLER_470_1432 ();
 FILLCELL_X32 FILLER_470_1464 ();
 FILLCELL_X32 FILLER_470_1496 ();
 FILLCELL_X32 FILLER_470_1528 ();
 FILLCELL_X32 FILLER_470_1560 ();
 FILLCELL_X32 FILLER_470_1592 ();
 FILLCELL_X32 FILLER_470_1624 ();
 FILLCELL_X32 FILLER_470_1656 ();
 FILLCELL_X32 FILLER_470_1688 ();
 FILLCELL_X32 FILLER_470_1720 ();
 FILLCELL_X32 FILLER_470_1752 ();
 FILLCELL_X32 FILLER_470_1784 ();
 FILLCELL_X32 FILLER_470_1816 ();
 FILLCELL_X32 FILLER_470_1848 ();
 FILLCELL_X8 FILLER_470_1880 ();
 FILLCELL_X4 FILLER_470_1888 ();
 FILLCELL_X2 FILLER_470_1892 ();
 FILLCELL_X32 FILLER_470_1895 ();
 FILLCELL_X32 FILLER_470_1927 ();
 FILLCELL_X32 FILLER_470_1959 ();
 FILLCELL_X32 FILLER_470_1991 ();
 FILLCELL_X32 FILLER_470_2023 ();
 FILLCELL_X32 FILLER_470_2055 ();
 FILLCELL_X32 FILLER_470_2087 ();
 FILLCELL_X32 FILLER_470_2119 ();
 FILLCELL_X32 FILLER_470_2151 ();
 FILLCELL_X32 FILLER_470_2183 ();
 FILLCELL_X32 FILLER_470_2215 ();
 FILLCELL_X32 FILLER_470_2247 ();
 FILLCELL_X32 FILLER_470_2279 ();
 FILLCELL_X32 FILLER_470_2311 ();
 FILLCELL_X32 FILLER_470_2343 ();
 FILLCELL_X32 FILLER_470_2375 ();
 FILLCELL_X32 FILLER_470_2407 ();
 FILLCELL_X32 FILLER_470_2439 ();
 FILLCELL_X32 FILLER_470_2471 ();
 FILLCELL_X32 FILLER_470_2503 ();
 FILLCELL_X32 FILLER_470_2535 ();
 FILLCELL_X32 FILLER_470_2567 ();
 FILLCELL_X32 FILLER_470_2599 ();
 FILLCELL_X32 FILLER_470_2631 ();
 FILLCELL_X32 FILLER_470_2663 ();
 FILLCELL_X32 FILLER_470_2695 ();
 FILLCELL_X32 FILLER_470_2727 ();
 FILLCELL_X32 FILLER_470_2759 ();
 FILLCELL_X32 FILLER_470_2791 ();
 FILLCELL_X32 FILLER_470_2823 ();
 FILLCELL_X32 FILLER_470_2855 ();
 FILLCELL_X32 FILLER_470_2887 ();
 FILLCELL_X32 FILLER_470_2919 ();
 FILLCELL_X32 FILLER_470_2951 ();
 FILLCELL_X32 FILLER_470_2983 ();
 FILLCELL_X32 FILLER_470_3015 ();
 FILLCELL_X32 FILLER_470_3047 ();
 FILLCELL_X32 FILLER_470_3079 ();
 FILLCELL_X32 FILLER_470_3111 ();
 FILLCELL_X8 FILLER_470_3143 ();
 FILLCELL_X4 FILLER_470_3151 ();
 FILLCELL_X2 FILLER_470_3155 ();
 FILLCELL_X32 FILLER_470_3158 ();
 FILLCELL_X32 FILLER_470_3190 ();
 FILLCELL_X32 FILLER_470_3222 ();
 FILLCELL_X32 FILLER_470_3254 ();
 FILLCELL_X32 FILLER_470_3286 ();
 FILLCELL_X32 FILLER_470_3318 ();
 FILLCELL_X32 FILLER_470_3350 ();
 FILLCELL_X32 FILLER_470_3382 ();
 FILLCELL_X32 FILLER_470_3414 ();
 FILLCELL_X32 FILLER_470_3446 ();
 FILLCELL_X32 FILLER_470_3478 ();
 FILLCELL_X32 FILLER_470_3510 ();
 FILLCELL_X32 FILLER_470_3542 ();
 FILLCELL_X32 FILLER_470_3574 ();
 FILLCELL_X32 FILLER_470_3606 ();
 FILLCELL_X32 FILLER_470_3638 ();
 FILLCELL_X32 FILLER_470_3670 ();
 FILLCELL_X32 FILLER_470_3702 ();
 FILLCELL_X4 FILLER_470_3734 ();
 FILLCELL_X32 FILLER_471_1 ();
 FILLCELL_X32 FILLER_471_33 ();
 FILLCELL_X32 FILLER_471_65 ();
 FILLCELL_X32 FILLER_471_97 ();
 FILLCELL_X32 FILLER_471_129 ();
 FILLCELL_X32 FILLER_471_161 ();
 FILLCELL_X32 FILLER_471_193 ();
 FILLCELL_X32 FILLER_471_225 ();
 FILLCELL_X32 FILLER_471_257 ();
 FILLCELL_X32 FILLER_471_289 ();
 FILLCELL_X32 FILLER_471_321 ();
 FILLCELL_X32 FILLER_471_353 ();
 FILLCELL_X32 FILLER_471_385 ();
 FILLCELL_X32 FILLER_471_417 ();
 FILLCELL_X32 FILLER_471_449 ();
 FILLCELL_X32 FILLER_471_481 ();
 FILLCELL_X32 FILLER_471_513 ();
 FILLCELL_X32 FILLER_471_545 ();
 FILLCELL_X32 FILLER_471_577 ();
 FILLCELL_X32 FILLER_471_609 ();
 FILLCELL_X32 FILLER_471_641 ();
 FILLCELL_X32 FILLER_471_673 ();
 FILLCELL_X32 FILLER_471_705 ();
 FILLCELL_X32 FILLER_471_737 ();
 FILLCELL_X32 FILLER_471_769 ();
 FILLCELL_X32 FILLER_471_801 ();
 FILLCELL_X32 FILLER_471_833 ();
 FILLCELL_X32 FILLER_471_865 ();
 FILLCELL_X32 FILLER_471_897 ();
 FILLCELL_X32 FILLER_471_929 ();
 FILLCELL_X32 FILLER_471_961 ();
 FILLCELL_X32 FILLER_471_993 ();
 FILLCELL_X32 FILLER_471_1025 ();
 FILLCELL_X32 FILLER_471_1057 ();
 FILLCELL_X32 FILLER_471_1089 ();
 FILLCELL_X32 FILLER_471_1121 ();
 FILLCELL_X32 FILLER_471_1153 ();
 FILLCELL_X32 FILLER_471_1185 ();
 FILLCELL_X32 FILLER_471_1217 ();
 FILLCELL_X8 FILLER_471_1249 ();
 FILLCELL_X4 FILLER_471_1257 ();
 FILLCELL_X2 FILLER_471_1261 ();
 FILLCELL_X32 FILLER_471_1264 ();
 FILLCELL_X32 FILLER_471_1296 ();
 FILLCELL_X32 FILLER_471_1328 ();
 FILLCELL_X32 FILLER_471_1360 ();
 FILLCELL_X32 FILLER_471_1392 ();
 FILLCELL_X32 FILLER_471_1424 ();
 FILLCELL_X32 FILLER_471_1456 ();
 FILLCELL_X32 FILLER_471_1488 ();
 FILLCELL_X32 FILLER_471_1520 ();
 FILLCELL_X32 FILLER_471_1552 ();
 FILLCELL_X32 FILLER_471_1584 ();
 FILLCELL_X32 FILLER_471_1616 ();
 FILLCELL_X32 FILLER_471_1648 ();
 FILLCELL_X32 FILLER_471_1680 ();
 FILLCELL_X32 FILLER_471_1712 ();
 FILLCELL_X32 FILLER_471_1744 ();
 FILLCELL_X32 FILLER_471_1776 ();
 FILLCELL_X32 FILLER_471_1808 ();
 FILLCELL_X32 FILLER_471_1840 ();
 FILLCELL_X32 FILLER_471_1872 ();
 FILLCELL_X32 FILLER_471_1904 ();
 FILLCELL_X32 FILLER_471_1936 ();
 FILLCELL_X32 FILLER_471_1968 ();
 FILLCELL_X32 FILLER_471_2000 ();
 FILLCELL_X32 FILLER_471_2032 ();
 FILLCELL_X32 FILLER_471_2064 ();
 FILLCELL_X32 FILLER_471_2096 ();
 FILLCELL_X32 FILLER_471_2128 ();
 FILLCELL_X32 FILLER_471_2160 ();
 FILLCELL_X32 FILLER_471_2192 ();
 FILLCELL_X32 FILLER_471_2224 ();
 FILLCELL_X32 FILLER_471_2256 ();
 FILLCELL_X32 FILLER_471_2288 ();
 FILLCELL_X32 FILLER_471_2320 ();
 FILLCELL_X32 FILLER_471_2352 ();
 FILLCELL_X32 FILLER_471_2384 ();
 FILLCELL_X32 FILLER_471_2416 ();
 FILLCELL_X32 FILLER_471_2448 ();
 FILLCELL_X32 FILLER_471_2480 ();
 FILLCELL_X8 FILLER_471_2512 ();
 FILLCELL_X4 FILLER_471_2520 ();
 FILLCELL_X2 FILLER_471_2524 ();
 FILLCELL_X32 FILLER_471_2527 ();
 FILLCELL_X32 FILLER_471_2559 ();
 FILLCELL_X32 FILLER_471_2591 ();
 FILLCELL_X32 FILLER_471_2623 ();
 FILLCELL_X32 FILLER_471_2655 ();
 FILLCELL_X32 FILLER_471_2687 ();
 FILLCELL_X32 FILLER_471_2719 ();
 FILLCELL_X32 FILLER_471_2751 ();
 FILLCELL_X32 FILLER_471_2783 ();
 FILLCELL_X32 FILLER_471_2815 ();
 FILLCELL_X32 FILLER_471_2847 ();
 FILLCELL_X32 FILLER_471_2879 ();
 FILLCELL_X32 FILLER_471_2911 ();
 FILLCELL_X32 FILLER_471_2943 ();
 FILLCELL_X32 FILLER_471_2975 ();
 FILLCELL_X32 FILLER_471_3007 ();
 FILLCELL_X32 FILLER_471_3039 ();
 FILLCELL_X32 FILLER_471_3071 ();
 FILLCELL_X32 FILLER_471_3103 ();
 FILLCELL_X32 FILLER_471_3135 ();
 FILLCELL_X32 FILLER_471_3167 ();
 FILLCELL_X32 FILLER_471_3199 ();
 FILLCELL_X32 FILLER_471_3231 ();
 FILLCELL_X32 FILLER_471_3263 ();
 FILLCELL_X32 FILLER_471_3295 ();
 FILLCELL_X32 FILLER_471_3327 ();
 FILLCELL_X32 FILLER_471_3359 ();
 FILLCELL_X32 FILLER_471_3391 ();
 FILLCELL_X32 FILLER_471_3423 ();
 FILLCELL_X32 FILLER_471_3455 ();
 FILLCELL_X32 FILLER_471_3487 ();
 FILLCELL_X32 FILLER_471_3519 ();
 FILLCELL_X32 FILLER_471_3551 ();
 FILLCELL_X32 FILLER_471_3583 ();
 FILLCELL_X32 FILLER_471_3615 ();
 FILLCELL_X32 FILLER_471_3647 ();
 FILLCELL_X32 FILLER_471_3679 ();
 FILLCELL_X16 FILLER_471_3711 ();
 FILLCELL_X8 FILLER_471_3727 ();
 FILLCELL_X2 FILLER_471_3735 ();
 FILLCELL_X1 FILLER_471_3737 ();
 FILLCELL_X32 FILLER_472_1 ();
 FILLCELL_X32 FILLER_472_33 ();
 FILLCELL_X32 FILLER_472_65 ();
 FILLCELL_X32 FILLER_472_97 ();
 FILLCELL_X32 FILLER_472_129 ();
 FILLCELL_X32 FILLER_472_161 ();
 FILLCELL_X32 FILLER_472_193 ();
 FILLCELL_X32 FILLER_472_225 ();
 FILLCELL_X32 FILLER_472_257 ();
 FILLCELL_X32 FILLER_472_289 ();
 FILLCELL_X32 FILLER_472_321 ();
 FILLCELL_X32 FILLER_472_353 ();
 FILLCELL_X32 FILLER_472_385 ();
 FILLCELL_X32 FILLER_472_417 ();
 FILLCELL_X32 FILLER_472_449 ();
 FILLCELL_X32 FILLER_472_481 ();
 FILLCELL_X32 FILLER_472_513 ();
 FILLCELL_X32 FILLER_472_545 ();
 FILLCELL_X32 FILLER_472_577 ();
 FILLCELL_X16 FILLER_472_609 ();
 FILLCELL_X4 FILLER_472_625 ();
 FILLCELL_X2 FILLER_472_629 ();
 FILLCELL_X32 FILLER_472_632 ();
 FILLCELL_X32 FILLER_472_664 ();
 FILLCELL_X32 FILLER_472_696 ();
 FILLCELL_X32 FILLER_472_728 ();
 FILLCELL_X32 FILLER_472_760 ();
 FILLCELL_X32 FILLER_472_792 ();
 FILLCELL_X32 FILLER_472_824 ();
 FILLCELL_X32 FILLER_472_856 ();
 FILLCELL_X32 FILLER_472_888 ();
 FILLCELL_X32 FILLER_472_920 ();
 FILLCELL_X32 FILLER_472_952 ();
 FILLCELL_X32 FILLER_472_984 ();
 FILLCELL_X32 FILLER_472_1016 ();
 FILLCELL_X32 FILLER_472_1048 ();
 FILLCELL_X32 FILLER_472_1080 ();
 FILLCELL_X32 FILLER_472_1112 ();
 FILLCELL_X32 FILLER_472_1144 ();
 FILLCELL_X32 FILLER_472_1176 ();
 FILLCELL_X32 FILLER_472_1208 ();
 FILLCELL_X32 FILLER_472_1240 ();
 FILLCELL_X32 FILLER_472_1272 ();
 FILLCELL_X32 FILLER_472_1304 ();
 FILLCELL_X32 FILLER_472_1336 ();
 FILLCELL_X32 FILLER_472_1368 ();
 FILLCELL_X32 FILLER_472_1400 ();
 FILLCELL_X32 FILLER_472_1432 ();
 FILLCELL_X32 FILLER_472_1464 ();
 FILLCELL_X32 FILLER_472_1496 ();
 FILLCELL_X32 FILLER_472_1528 ();
 FILLCELL_X32 FILLER_472_1560 ();
 FILLCELL_X32 FILLER_472_1592 ();
 FILLCELL_X32 FILLER_472_1624 ();
 FILLCELL_X32 FILLER_472_1656 ();
 FILLCELL_X32 FILLER_472_1688 ();
 FILLCELL_X32 FILLER_472_1720 ();
 FILLCELL_X32 FILLER_472_1752 ();
 FILLCELL_X32 FILLER_472_1784 ();
 FILLCELL_X32 FILLER_472_1816 ();
 FILLCELL_X32 FILLER_472_1848 ();
 FILLCELL_X8 FILLER_472_1880 ();
 FILLCELL_X4 FILLER_472_1888 ();
 FILLCELL_X2 FILLER_472_1892 ();
 FILLCELL_X32 FILLER_472_1895 ();
 FILLCELL_X32 FILLER_472_1927 ();
 FILLCELL_X32 FILLER_472_1959 ();
 FILLCELL_X32 FILLER_472_1991 ();
 FILLCELL_X32 FILLER_472_2023 ();
 FILLCELL_X32 FILLER_472_2055 ();
 FILLCELL_X32 FILLER_472_2087 ();
 FILLCELL_X32 FILLER_472_2119 ();
 FILLCELL_X32 FILLER_472_2151 ();
 FILLCELL_X32 FILLER_472_2183 ();
 FILLCELL_X32 FILLER_472_2215 ();
 FILLCELL_X32 FILLER_472_2247 ();
 FILLCELL_X32 FILLER_472_2279 ();
 FILLCELL_X32 FILLER_472_2311 ();
 FILLCELL_X32 FILLER_472_2343 ();
 FILLCELL_X32 FILLER_472_2375 ();
 FILLCELL_X32 FILLER_472_2407 ();
 FILLCELL_X32 FILLER_472_2439 ();
 FILLCELL_X32 FILLER_472_2471 ();
 FILLCELL_X32 FILLER_472_2503 ();
 FILLCELL_X32 FILLER_472_2535 ();
 FILLCELL_X32 FILLER_472_2567 ();
 FILLCELL_X32 FILLER_472_2599 ();
 FILLCELL_X32 FILLER_472_2631 ();
 FILLCELL_X32 FILLER_472_2663 ();
 FILLCELL_X32 FILLER_472_2695 ();
 FILLCELL_X32 FILLER_472_2727 ();
 FILLCELL_X32 FILLER_472_2759 ();
 FILLCELL_X32 FILLER_472_2791 ();
 FILLCELL_X32 FILLER_472_2823 ();
 FILLCELL_X32 FILLER_472_2855 ();
 FILLCELL_X32 FILLER_472_2887 ();
 FILLCELL_X32 FILLER_472_2919 ();
 FILLCELL_X32 FILLER_472_2951 ();
 FILLCELL_X32 FILLER_472_2983 ();
 FILLCELL_X32 FILLER_472_3015 ();
 FILLCELL_X32 FILLER_472_3047 ();
 FILLCELL_X32 FILLER_472_3079 ();
 FILLCELL_X32 FILLER_472_3111 ();
 FILLCELL_X8 FILLER_472_3143 ();
 FILLCELL_X4 FILLER_472_3151 ();
 FILLCELL_X2 FILLER_472_3155 ();
 FILLCELL_X32 FILLER_472_3158 ();
 FILLCELL_X32 FILLER_472_3190 ();
 FILLCELL_X32 FILLER_472_3222 ();
 FILLCELL_X32 FILLER_472_3254 ();
 FILLCELL_X32 FILLER_472_3286 ();
 FILLCELL_X32 FILLER_472_3318 ();
 FILLCELL_X32 FILLER_472_3350 ();
 FILLCELL_X32 FILLER_472_3382 ();
 FILLCELL_X32 FILLER_472_3414 ();
 FILLCELL_X32 FILLER_472_3446 ();
 FILLCELL_X32 FILLER_472_3478 ();
 FILLCELL_X32 FILLER_472_3510 ();
 FILLCELL_X32 FILLER_472_3542 ();
 FILLCELL_X32 FILLER_472_3574 ();
 FILLCELL_X32 FILLER_472_3606 ();
 FILLCELL_X32 FILLER_472_3638 ();
 FILLCELL_X32 FILLER_472_3670 ();
 FILLCELL_X32 FILLER_472_3702 ();
 FILLCELL_X4 FILLER_472_3734 ();
 FILLCELL_X32 FILLER_473_1 ();
 FILLCELL_X32 FILLER_473_33 ();
 FILLCELL_X32 FILLER_473_65 ();
 FILLCELL_X32 FILLER_473_97 ();
 FILLCELL_X32 FILLER_473_129 ();
 FILLCELL_X32 FILLER_473_161 ();
 FILLCELL_X32 FILLER_473_193 ();
 FILLCELL_X32 FILLER_473_225 ();
 FILLCELL_X32 FILLER_473_257 ();
 FILLCELL_X32 FILLER_473_289 ();
 FILLCELL_X32 FILLER_473_321 ();
 FILLCELL_X32 FILLER_473_353 ();
 FILLCELL_X32 FILLER_473_385 ();
 FILLCELL_X32 FILLER_473_417 ();
 FILLCELL_X32 FILLER_473_449 ();
 FILLCELL_X32 FILLER_473_481 ();
 FILLCELL_X32 FILLER_473_513 ();
 FILLCELL_X32 FILLER_473_545 ();
 FILLCELL_X32 FILLER_473_577 ();
 FILLCELL_X32 FILLER_473_609 ();
 FILLCELL_X32 FILLER_473_641 ();
 FILLCELL_X32 FILLER_473_673 ();
 FILLCELL_X32 FILLER_473_705 ();
 FILLCELL_X32 FILLER_473_737 ();
 FILLCELL_X32 FILLER_473_769 ();
 FILLCELL_X32 FILLER_473_801 ();
 FILLCELL_X32 FILLER_473_833 ();
 FILLCELL_X32 FILLER_473_865 ();
 FILLCELL_X32 FILLER_473_897 ();
 FILLCELL_X32 FILLER_473_929 ();
 FILLCELL_X32 FILLER_473_961 ();
 FILLCELL_X32 FILLER_473_993 ();
 FILLCELL_X32 FILLER_473_1025 ();
 FILLCELL_X32 FILLER_473_1057 ();
 FILLCELL_X32 FILLER_473_1089 ();
 FILLCELL_X32 FILLER_473_1121 ();
 FILLCELL_X32 FILLER_473_1153 ();
 FILLCELL_X32 FILLER_473_1185 ();
 FILLCELL_X32 FILLER_473_1217 ();
 FILLCELL_X8 FILLER_473_1249 ();
 FILLCELL_X4 FILLER_473_1257 ();
 FILLCELL_X2 FILLER_473_1261 ();
 FILLCELL_X32 FILLER_473_1264 ();
 FILLCELL_X32 FILLER_473_1296 ();
 FILLCELL_X32 FILLER_473_1328 ();
 FILLCELL_X32 FILLER_473_1360 ();
 FILLCELL_X32 FILLER_473_1392 ();
 FILLCELL_X32 FILLER_473_1424 ();
 FILLCELL_X32 FILLER_473_1456 ();
 FILLCELL_X32 FILLER_473_1488 ();
 FILLCELL_X32 FILLER_473_1520 ();
 FILLCELL_X32 FILLER_473_1552 ();
 FILLCELL_X32 FILLER_473_1584 ();
 FILLCELL_X32 FILLER_473_1616 ();
 FILLCELL_X32 FILLER_473_1648 ();
 FILLCELL_X32 FILLER_473_1680 ();
 FILLCELL_X32 FILLER_473_1712 ();
 FILLCELL_X32 FILLER_473_1744 ();
 FILLCELL_X32 FILLER_473_1776 ();
 FILLCELL_X32 FILLER_473_1808 ();
 FILLCELL_X32 FILLER_473_1840 ();
 FILLCELL_X32 FILLER_473_1872 ();
 FILLCELL_X32 FILLER_473_1904 ();
 FILLCELL_X32 FILLER_473_1936 ();
 FILLCELL_X32 FILLER_473_1968 ();
 FILLCELL_X32 FILLER_473_2000 ();
 FILLCELL_X32 FILLER_473_2032 ();
 FILLCELL_X32 FILLER_473_2064 ();
 FILLCELL_X32 FILLER_473_2096 ();
 FILLCELL_X32 FILLER_473_2128 ();
 FILLCELL_X32 FILLER_473_2160 ();
 FILLCELL_X32 FILLER_473_2192 ();
 FILLCELL_X32 FILLER_473_2224 ();
 FILLCELL_X32 FILLER_473_2256 ();
 FILLCELL_X32 FILLER_473_2288 ();
 FILLCELL_X32 FILLER_473_2320 ();
 FILLCELL_X32 FILLER_473_2352 ();
 FILLCELL_X32 FILLER_473_2384 ();
 FILLCELL_X32 FILLER_473_2416 ();
 FILLCELL_X32 FILLER_473_2448 ();
 FILLCELL_X32 FILLER_473_2480 ();
 FILLCELL_X8 FILLER_473_2512 ();
 FILLCELL_X4 FILLER_473_2520 ();
 FILLCELL_X2 FILLER_473_2524 ();
 FILLCELL_X32 FILLER_473_2527 ();
 FILLCELL_X32 FILLER_473_2559 ();
 FILLCELL_X32 FILLER_473_2591 ();
 FILLCELL_X32 FILLER_473_2623 ();
 FILLCELL_X32 FILLER_473_2655 ();
 FILLCELL_X32 FILLER_473_2687 ();
 FILLCELL_X32 FILLER_473_2719 ();
 FILLCELL_X32 FILLER_473_2751 ();
 FILLCELL_X32 FILLER_473_2783 ();
 FILLCELL_X32 FILLER_473_2815 ();
 FILLCELL_X32 FILLER_473_2847 ();
 FILLCELL_X32 FILLER_473_2879 ();
 FILLCELL_X32 FILLER_473_2911 ();
 FILLCELL_X32 FILLER_473_2943 ();
 FILLCELL_X32 FILLER_473_2975 ();
 FILLCELL_X32 FILLER_473_3007 ();
 FILLCELL_X32 FILLER_473_3039 ();
 FILLCELL_X32 FILLER_473_3071 ();
 FILLCELL_X32 FILLER_473_3103 ();
 FILLCELL_X32 FILLER_473_3135 ();
 FILLCELL_X32 FILLER_473_3167 ();
 FILLCELL_X32 FILLER_473_3199 ();
 FILLCELL_X32 FILLER_473_3231 ();
 FILLCELL_X32 FILLER_473_3263 ();
 FILLCELL_X32 FILLER_473_3295 ();
 FILLCELL_X32 FILLER_473_3327 ();
 FILLCELL_X32 FILLER_473_3359 ();
 FILLCELL_X32 FILLER_473_3391 ();
 FILLCELL_X32 FILLER_473_3423 ();
 FILLCELL_X32 FILLER_473_3455 ();
 FILLCELL_X32 FILLER_473_3487 ();
 FILLCELL_X32 FILLER_473_3519 ();
 FILLCELL_X32 FILLER_473_3551 ();
 FILLCELL_X32 FILLER_473_3583 ();
 FILLCELL_X32 FILLER_473_3615 ();
 FILLCELL_X32 FILLER_473_3647 ();
 FILLCELL_X32 FILLER_473_3679 ();
 FILLCELL_X16 FILLER_473_3711 ();
 FILLCELL_X8 FILLER_473_3727 ();
 FILLCELL_X2 FILLER_473_3735 ();
 FILLCELL_X1 FILLER_473_3737 ();
 FILLCELL_X32 FILLER_474_1 ();
 FILLCELL_X32 FILLER_474_33 ();
 FILLCELL_X32 FILLER_474_65 ();
 FILLCELL_X32 FILLER_474_97 ();
 FILLCELL_X32 FILLER_474_129 ();
 FILLCELL_X32 FILLER_474_161 ();
 FILLCELL_X32 FILLER_474_193 ();
 FILLCELL_X32 FILLER_474_225 ();
 FILLCELL_X32 FILLER_474_257 ();
 FILLCELL_X32 FILLER_474_289 ();
 FILLCELL_X32 FILLER_474_321 ();
 FILLCELL_X32 FILLER_474_353 ();
 FILLCELL_X32 FILLER_474_385 ();
 FILLCELL_X32 FILLER_474_417 ();
 FILLCELL_X32 FILLER_474_449 ();
 FILLCELL_X32 FILLER_474_481 ();
 FILLCELL_X32 FILLER_474_513 ();
 FILLCELL_X32 FILLER_474_545 ();
 FILLCELL_X32 FILLER_474_577 ();
 FILLCELL_X16 FILLER_474_609 ();
 FILLCELL_X4 FILLER_474_625 ();
 FILLCELL_X2 FILLER_474_629 ();
 FILLCELL_X32 FILLER_474_632 ();
 FILLCELL_X32 FILLER_474_664 ();
 FILLCELL_X32 FILLER_474_696 ();
 FILLCELL_X32 FILLER_474_728 ();
 FILLCELL_X32 FILLER_474_760 ();
 FILLCELL_X32 FILLER_474_792 ();
 FILLCELL_X32 FILLER_474_824 ();
 FILLCELL_X32 FILLER_474_856 ();
 FILLCELL_X32 FILLER_474_888 ();
 FILLCELL_X32 FILLER_474_920 ();
 FILLCELL_X32 FILLER_474_952 ();
 FILLCELL_X32 FILLER_474_984 ();
 FILLCELL_X32 FILLER_474_1016 ();
 FILLCELL_X32 FILLER_474_1048 ();
 FILLCELL_X32 FILLER_474_1080 ();
 FILLCELL_X32 FILLER_474_1112 ();
 FILLCELL_X32 FILLER_474_1144 ();
 FILLCELL_X32 FILLER_474_1176 ();
 FILLCELL_X32 FILLER_474_1208 ();
 FILLCELL_X32 FILLER_474_1240 ();
 FILLCELL_X32 FILLER_474_1272 ();
 FILLCELL_X32 FILLER_474_1304 ();
 FILLCELL_X32 FILLER_474_1336 ();
 FILLCELL_X32 FILLER_474_1368 ();
 FILLCELL_X32 FILLER_474_1400 ();
 FILLCELL_X32 FILLER_474_1432 ();
 FILLCELL_X32 FILLER_474_1464 ();
 FILLCELL_X32 FILLER_474_1496 ();
 FILLCELL_X32 FILLER_474_1528 ();
 FILLCELL_X32 FILLER_474_1560 ();
 FILLCELL_X32 FILLER_474_1592 ();
 FILLCELL_X32 FILLER_474_1624 ();
 FILLCELL_X32 FILLER_474_1656 ();
 FILLCELL_X32 FILLER_474_1688 ();
 FILLCELL_X32 FILLER_474_1720 ();
 FILLCELL_X32 FILLER_474_1752 ();
 FILLCELL_X32 FILLER_474_1784 ();
 FILLCELL_X32 FILLER_474_1816 ();
 FILLCELL_X32 FILLER_474_1848 ();
 FILLCELL_X8 FILLER_474_1880 ();
 FILLCELL_X4 FILLER_474_1888 ();
 FILLCELL_X2 FILLER_474_1892 ();
 FILLCELL_X32 FILLER_474_1895 ();
 FILLCELL_X32 FILLER_474_1927 ();
 FILLCELL_X32 FILLER_474_1959 ();
 FILLCELL_X32 FILLER_474_1991 ();
 FILLCELL_X32 FILLER_474_2023 ();
 FILLCELL_X32 FILLER_474_2055 ();
 FILLCELL_X32 FILLER_474_2087 ();
 FILLCELL_X32 FILLER_474_2119 ();
 FILLCELL_X32 FILLER_474_2151 ();
 FILLCELL_X32 FILLER_474_2183 ();
 FILLCELL_X32 FILLER_474_2215 ();
 FILLCELL_X32 FILLER_474_2247 ();
 FILLCELL_X32 FILLER_474_2279 ();
 FILLCELL_X32 FILLER_474_2311 ();
 FILLCELL_X32 FILLER_474_2343 ();
 FILLCELL_X32 FILLER_474_2375 ();
 FILLCELL_X32 FILLER_474_2407 ();
 FILLCELL_X32 FILLER_474_2439 ();
 FILLCELL_X32 FILLER_474_2471 ();
 FILLCELL_X32 FILLER_474_2503 ();
 FILLCELL_X32 FILLER_474_2535 ();
 FILLCELL_X32 FILLER_474_2567 ();
 FILLCELL_X32 FILLER_474_2599 ();
 FILLCELL_X32 FILLER_474_2631 ();
 FILLCELL_X32 FILLER_474_2663 ();
 FILLCELL_X32 FILLER_474_2695 ();
 FILLCELL_X32 FILLER_474_2727 ();
 FILLCELL_X32 FILLER_474_2759 ();
 FILLCELL_X32 FILLER_474_2791 ();
 FILLCELL_X32 FILLER_474_2823 ();
 FILLCELL_X32 FILLER_474_2855 ();
 FILLCELL_X32 FILLER_474_2887 ();
 FILLCELL_X32 FILLER_474_2919 ();
 FILLCELL_X32 FILLER_474_2951 ();
 FILLCELL_X32 FILLER_474_2983 ();
 FILLCELL_X32 FILLER_474_3015 ();
 FILLCELL_X32 FILLER_474_3047 ();
 FILLCELL_X32 FILLER_474_3079 ();
 FILLCELL_X32 FILLER_474_3111 ();
 FILLCELL_X8 FILLER_474_3143 ();
 FILLCELL_X4 FILLER_474_3151 ();
 FILLCELL_X2 FILLER_474_3155 ();
 FILLCELL_X32 FILLER_474_3158 ();
 FILLCELL_X32 FILLER_474_3190 ();
 FILLCELL_X32 FILLER_474_3222 ();
 FILLCELL_X32 FILLER_474_3254 ();
 FILLCELL_X32 FILLER_474_3286 ();
 FILLCELL_X32 FILLER_474_3318 ();
 FILLCELL_X32 FILLER_474_3350 ();
 FILLCELL_X32 FILLER_474_3382 ();
 FILLCELL_X32 FILLER_474_3414 ();
 FILLCELL_X32 FILLER_474_3446 ();
 FILLCELL_X32 FILLER_474_3478 ();
 FILLCELL_X32 FILLER_474_3510 ();
 FILLCELL_X32 FILLER_474_3542 ();
 FILLCELL_X32 FILLER_474_3574 ();
 FILLCELL_X32 FILLER_474_3606 ();
 FILLCELL_X32 FILLER_474_3638 ();
 FILLCELL_X32 FILLER_474_3670 ();
 FILLCELL_X32 FILLER_474_3702 ();
 FILLCELL_X4 FILLER_474_3734 ();
 FILLCELL_X32 FILLER_475_1 ();
 FILLCELL_X32 FILLER_475_33 ();
 FILLCELL_X32 FILLER_475_65 ();
 FILLCELL_X32 FILLER_475_97 ();
 FILLCELL_X32 FILLER_475_129 ();
 FILLCELL_X32 FILLER_475_161 ();
 FILLCELL_X32 FILLER_475_193 ();
 FILLCELL_X32 FILLER_475_225 ();
 FILLCELL_X32 FILLER_475_257 ();
 FILLCELL_X32 FILLER_475_289 ();
 FILLCELL_X32 FILLER_475_321 ();
 FILLCELL_X32 FILLER_475_353 ();
 FILLCELL_X32 FILLER_475_385 ();
 FILLCELL_X32 FILLER_475_417 ();
 FILLCELL_X32 FILLER_475_449 ();
 FILLCELL_X32 FILLER_475_481 ();
 FILLCELL_X32 FILLER_475_513 ();
 FILLCELL_X32 FILLER_475_545 ();
 FILLCELL_X32 FILLER_475_577 ();
 FILLCELL_X32 FILLER_475_609 ();
 FILLCELL_X32 FILLER_475_641 ();
 FILLCELL_X32 FILLER_475_673 ();
 FILLCELL_X32 FILLER_475_705 ();
 FILLCELL_X32 FILLER_475_737 ();
 FILLCELL_X32 FILLER_475_769 ();
 FILLCELL_X32 FILLER_475_801 ();
 FILLCELL_X32 FILLER_475_833 ();
 FILLCELL_X32 FILLER_475_865 ();
 FILLCELL_X32 FILLER_475_897 ();
 FILLCELL_X32 FILLER_475_929 ();
 FILLCELL_X32 FILLER_475_961 ();
 FILLCELL_X32 FILLER_475_993 ();
 FILLCELL_X32 FILLER_475_1025 ();
 FILLCELL_X32 FILLER_475_1057 ();
 FILLCELL_X32 FILLER_475_1089 ();
 FILLCELL_X32 FILLER_475_1121 ();
 FILLCELL_X32 FILLER_475_1153 ();
 FILLCELL_X32 FILLER_475_1185 ();
 FILLCELL_X32 FILLER_475_1217 ();
 FILLCELL_X8 FILLER_475_1249 ();
 FILLCELL_X4 FILLER_475_1257 ();
 FILLCELL_X2 FILLER_475_1261 ();
 FILLCELL_X32 FILLER_475_1264 ();
 FILLCELL_X32 FILLER_475_1296 ();
 FILLCELL_X32 FILLER_475_1328 ();
 FILLCELL_X32 FILLER_475_1360 ();
 FILLCELL_X32 FILLER_475_1392 ();
 FILLCELL_X32 FILLER_475_1424 ();
 FILLCELL_X32 FILLER_475_1456 ();
 FILLCELL_X32 FILLER_475_1488 ();
 FILLCELL_X32 FILLER_475_1520 ();
 FILLCELL_X32 FILLER_475_1552 ();
 FILLCELL_X32 FILLER_475_1584 ();
 FILLCELL_X32 FILLER_475_1616 ();
 FILLCELL_X32 FILLER_475_1648 ();
 FILLCELL_X32 FILLER_475_1680 ();
 FILLCELL_X32 FILLER_475_1712 ();
 FILLCELL_X32 FILLER_475_1744 ();
 FILLCELL_X32 FILLER_475_1776 ();
 FILLCELL_X32 FILLER_475_1808 ();
 FILLCELL_X32 FILLER_475_1840 ();
 FILLCELL_X32 FILLER_475_1872 ();
 FILLCELL_X32 FILLER_475_1904 ();
 FILLCELL_X32 FILLER_475_1936 ();
 FILLCELL_X32 FILLER_475_1968 ();
 FILLCELL_X32 FILLER_475_2000 ();
 FILLCELL_X32 FILLER_475_2032 ();
 FILLCELL_X32 FILLER_475_2064 ();
 FILLCELL_X32 FILLER_475_2096 ();
 FILLCELL_X32 FILLER_475_2128 ();
 FILLCELL_X32 FILLER_475_2160 ();
 FILLCELL_X32 FILLER_475_2192 ();
 FILLCELL_X32 FILLER_475_2224 ();
 FILLCELL_X32 FILLER_475_2256 ();
 FILLCELL_X32 FILLER_475_2288 ();
 FILLCELL_X32 FILLER_475_2320 ();
 FILLCELL_X32 FILLER_475_2352 ();
 FILLCELL_X32 FILLER_475_2384 ();
 FILLCELL_X32 FILLER_475_2416 ();
 FILLCELL_X32 FILLER_475_2448 ();
 FILLCELL_X32 FILLER_475_2480 ();
 FILLCELL_X8 FILLER_475_2512 ();
 FILLCELL_X4 FILLER_475_2520 ();
 FILLCELL_X2 FILLER_475_2524 ();
 FILLCELL_X32 FILLER_475_2527 ();
 FILLCELL_X32 FILLER_475_2559 ();
 FILLCELL_X32 FILLER_475_2591 ();
 FILLCELL_X32 FILLER_475_2623 ();
 FILLCELL_X32 FILLER_475_2655 ();
 FILLCELL_X32 FILLER_475_2687 ();
 FILLCELL_X32 FILLER_475_2719 ();
 FILLCELL_X32 FILLER_475_2751 ();
 FILLCELL_X32 FILLER_475_2783 ();
 FILLCELL_X32 FILLER_475_2815 ();
 FILLCELL_X32 FILLER_475_2847 ();
 FILLCELL_X32 FILLER_475_2879 ();
 FILLCELL_X32 FILLER_475_2911 ();
 FILLCELL_X32 FILLER_475_2943 ();
 FILLCELL_X32 FILLER_475_2975 ();
 FILLCELL_X32 FILLER_475_3007 ();
 FILLCELL_X32 FILLER_475_3039 ();
 FILLCELL_X32 FILLER_475_3071 ();
 FILLCELL_X32 FILLER_475_3103 ();
 FILLCELL_X32 FILLER_475_3135 ();
 FILLCELL_X32 FILLER_475_3167 ();
 FILLCELL_X32 FILLER_475_3199 ();
 FILLCELL_X32 FILLER_475_3231 ();
 FILLCELL_X32 FILLER_475_3263 ();
 FILLCELL_X32 FILLER_475_3295 ();
 FILLCELL_X32 FILLER_475_3327 ();
 FILLCELL_X32 FILLER_475_3359 ();
 FILLCELL_X32 FILLER_475_3391 ();
 FILLCELL_X32 FILLER_475_3423 ();
 FILLCELL_X32 FILLER_475_3455 ();
 FILLCELL_X32 FILLER_475_3487 ();
 FILLCELL_X32 FILLER_475_3519 ();
 FILLCELL_X32 FILLER_475_3551 ();
 FILLCELL_X32 FILLER_475_3583 ();
 FILLCELL_X32 FILLER_475_3615 ();
 FILLCELL_X32 FILLER_475_3647 ();
 FILLCELL_X32 FILLER_475_3679 ();
 FILLCELL_X16 FILLER_475_3711 ();
 FILLCELL_X8 FILLER_475_3727 ();
 FILLCELL_X2 FILLER_475_3735 ();
 FILLCELL_X1 FILLER_475_3737 ();
 FILLCELL_X32 FILLER_476_1 ();
 FILLCELL_X32 FILLER_476_33 ();
 FILLCELL_X32 FILLER_476_65 ();
 FILLCELL_X32 FILLER_476_97 ();
 FILLCELL_X32 FILLER_476_129 ();
 FILLCELL_X32 FILLER_476_161 ();
 FILLCELL_X32 FILLER_476_193 ();
 FILLCELL_X32 FILLER_476_225 ();
 FILLCELL_X32 FILLER_476_257 ();
 FILLCELL_X32 FILLER_476_289 ();
 FILLCELL_X32 FILLER_476_321 ();
 FILLCELL_X32 FILLER_476_353 ();
 FILLCELL_X32 FILLER_476_385 ();
 FILLCELL_X32 FILLER_476_417 ();
 FILLCELL_X32 FILLER_476_449 ();
 FILLCELL_X32 FILLER_476_481 ();
 FILLCELL_X32 FILLER_476_513 ();
 FILLCELL_X32 FILLER_476_545 ();
 FILLCELL_X32 FILLER_476_577 ();
 FILLCELL_X16 FILLER_476_609 ();
 FILLCELL_X4 FILLER_476_625 ();
 FILLCELL_X2 FILLER_476_629 ();
 FILLCELL_X32 FILLER_476_632 ();
 FILLCELL_X32 FILLER_476_664 ();
 FILLCELL_X32 FILLER_476_696 ();
 FILLCELL_X32 FILLER_476_728 ();
 FILLCELL_X32 FILLER_476_760 ();
 FILLCELL_X32 FILLER_476_792 ();
 FILLCELL_X32 FILLER_476_824 ();
 FILLCELL_X32 FILLER_476_856 ();
 FILLCELL_X32 FILLER_476_888 ();
 FILLCELL_X32 FILLER_476_920 ();
 FILLCELL_X32 FILLER_476_952 ();
 FILLCELL_X32 FILLER_476_984 ();
 FILLCELL_X32 FILLER_476_1016 ();
 FILLCELL_X32 FILLER_476_1048 ();
 FILLCELL_X32 FILLER_476_1080 ();
 FILLCELL_X32 FILLER_476_1112 ();
 FILLCELL_X32 FILLER_476_1144 ();
 FILLCELL_X32 FILLER_476_1176 ();
 FILLCELL_X32 FILLER_476_1208 ();
 FILLCELL_X32 FILLER_476_1240 ();
 FILLCELL_X32 FILLER_476_1272 ();
 FILLCELL_X32 FILLER_476_1304 ();
 FILLCELL_X32 FILLER_476_1336 ();
 FILLCELL_X32 FILLER_476_1368 ();
 FILLCELL_X32 FILLER_476_1400 ();
 FILLCELL_X32 FILLER_476_1432 ();
 FILLCELL_X32 FILLER_476_1464 ();
 FILLCELL_X32 FILLER_476_1496 ();
 FILLCELL_X32 FILLER_476_1528 ();
 FILLCELL_X32 FILLER_476_1560 ();
 FILLCELL_X32 FILLER_476_1592 ();
 FILLCELL_X32 FILLER_476_1624 ();
 FILLCELL_X32 FILLER_476_1656 ();
 FILLCELL_X32 FILLER_476_1688 ();
 FILLCELL_X32 FILLER_476_1720 ();
 FILLCELL_X32 FILLER_476_1752 ();
 FILLCELL_X32 FILLER_476_1784 ();
 FILLCELL_X32 FILLER_476_1816 ();
 FILLCELL_X32 FILLER_476_1848 ();
 FILLCELL_X8 FILLER_476_1880 ();
 FILLCELL_X4 FILLER_476_1888 ();
 FILLCELL_X2 FILLER_476_1892 ();
 FILLCELL_X32 FILLER_476_1895 ();
 FILLCELL_X32 FILLER_476_1927 ();
 FILLCELL_X32 FILLER_476_1959 ();
 FILLCELL_X32 FILLER_476_1991 ();
 FILLCELL_X32 FILLER_476_2023 ();
 FILLCELL_X32 FILLER_476_2055 ();
 FILLCELL_X32 FILLER_476_2087 ();
 FILLCELL_X32 FILLER_476_2119 ();
 FILLCELL_X32 FILLER_476_2151 ();
 FILLCELL_X32 FILLER_476_2183 ();
 FILLCELL_X32 FILLER_476_2215 ();
 FILLCELL_X32 FILLER_476_2247 ();
 FILLCELL_X32 FILLER_476_2279 ();
 FILLCELL_X32 FILLER_476_2311 ();
 FILLCELL_X32 FILLER_476_2343 ();
 FILLCELL_X32 FILLER_476_2375 ();
 FILLCELL_X32 FILLER_476_2407 ();
 FILLCELL_X32 FILLER_476_2439 ();
 FILLCELL_X32 FILLER_476_2471 ();
 FILLCELL_X32 FILLER_476_2503 ();
 FILLCELL_X32 FILLER_476_2535 ();
 FILLCELL_X32 FILLER_476_2567 ();
 FILLCELL_X32 FILLER_476_2599 ();
 FILLCELL_X32 FILLER_476_2631 ();
 FILLCELL_X32 FILLER_476_2663 ();
 FILLCELL_X32 FILLER_476_2695 ();
 FILLCELL_X32 FILLER_476_2727 ();
 FILLCELL_X32 FILLER_476_2759 ();
 FILLCELL_X32 FILLER_476_2791 ();
 FILLCELL_X32 FILLER_476_2823 ();
 FILLCELL_X32 FILLER_476_2855 ();
 FILLCELL_X32 FILLER_476_2887 ();
 FILLCELL_X32 FILLER_476_2919 ();
 FILLCELL_X32 FILLER_476_2951 ();
 FILLCELL_X32 FILLER_476_2983 ();
 FILLCELL_X32 FILLER_476_3015 ();
 FILLCELL_X32 FILLER_476_3047 ();
 FILLCELL_X32 FILLER_476_3079 ();
 FILLCELL_X32 FILLER_476_3111 ();
 FILLCELL_X8 FILLER_476_3143 ();
 FILLCELL_X4 FILLER_476_3151 ();
 FILLCELL_X2 FILLER_476_3155 ();
 FILLCELL_X32 FILLER_476_3158 ();
 FILLCELL_X32 FILLER_476_3190 ();
 FILLCELL_X32 FILLER_476_3222 ();
 FILLCELL_X32 FILLER_476_3254 ();
 FILLCELL_X32 FILLER_476_3286 ();
 FILLCELL_X32 FILLER_476_3318 ();
 FILLCELL_X32 FILLER_476_3350 ();
 FILLCELL_X32 FILLER_476_3382 ();
 FILLCELL_X32 FILLER_476_3414 ();
 FILLCELL_X32 FILLER_476_3446 ();
 FILLCELL_X32 FILLER_476_3478 ();
 FILLCELL_X32 FILLER_476_3510 ();
 FILLCELL_X32 FILLER_476_3542 ();
 FILLCELL_X32 FILLER_476_3574 ();
 FILLCELL_X32 FILLER_476_3606 ();
 FILLCELL_X32 FILLER_476_3638 ();
 FILLCELL_X32 FILLER_476_3670 ();
 FILLCELL_X32 FILLER_476_3702 ();
 FILLCELL_X4 FILLER_476_3734 ();
 FILLCELL_X32 FILLER_477_1 ();
 FILLCELL_X32 FILLER_477_33 ();
 FILLCELL_X32 FILLER_477_65 ();
 FILLCELL_X32 FILLER_477_97 ();
 FILLCELL_X32 FILLER_477_129 ();
 FILLCELL_X32 FILLER_477_161 ();
 FILLCELL_X32 FILLER_477_193 ();
 FILLCELL_X32 FILLER_477_225 ();
 FILLCELL_X32 FILLER_477_257 ();
 FILLCELL_X32 FILLER_477_289 ();
 FILLCELL_X32 FILLER_477_321 ();
 FILLCELL_X32 FILLER_477_353 ();
 FILLCELL_X32 FILLER_477_385 ();
 FILLCELL_X32 FILLER_477_417 ();
 FILLCELL_X32 FILLER_477_449 ();
 FILLCELL_X32 FILLER_477_481 ();
 FILLCELL_X32 FILLER_477_513 ();
 FILLCELL_X32 FILLER_477_545 ();
 FILLCELL_X32 FILLER_477_577 ();
 FILLCELL_X32 FILLER_477_609 ();
 FILLCELL_X32 FILLER_477_641 ();
 FILLCELL_X32 FILLER_477_673 ();
 FILLCELL_X32 FILLER_477_705 ();
 FILLCELL_X32 FILLER_477_737 ();
 FILLCELL_X32 FILLER_477_769 ();
 FILLCELL_X32 FILLER_477_801 ();
 FILLCELL_X32 FILLER_477_833 ();
 FILLCELL_X32 FILLER_477_865 ();
 FILLCELL_X32 FILLER_477_897 ();
 FILLCELL_X32 FILLER_477_929 ();
 FILLCELL_X32 FILLER_477_961 ();
 FILLCELL_X32 FILLER_477_993 ();
 FILLCELL_X32 FILLER_477_1025 ();
 FILLCELL_X32 FILLER_477_1057 ();
 FILLCELL_X32 FILLER_477_1089 ();
 FILLCELL_X32 FILLER_477_1121 ();
 FILLCELL_X32 FILLER_477_1153 ();
 FILLCELL_X32 FILLER_477_1185 ();
 FILLCELL_X32 FILLER_477_1217 ();
 FILLCELL_X8 FILLER_477_1249 ();
 FILLCELL_X4 FILLER_477_1257 ();
 FILLCELL_X2 FILLER_477_1261 ();
 FILLCELL_X32 FILLER_477_1264 ();
 FILLCELL_X32 FILLER_477_1296 ();
 FILLCELL_X32 FILLER_477_1328 ();
 FILLCELL_X32 FILLER_477_1360 ();
 FILLCELL_X32 FILLER_477_1392 ();
 FILLCELL_X32 FILLER_477_1424 ();
 FILLCELL_X32 FILLER_477_1456 ();
 FILLCELL_X32 FILLER_477_1488 ();
 FILLCELL_X32 FILLER_477_1520 ();
 FILLCELL_X32 FILLER_477_1552 ();
 FILLCELL_X32 FILLER_477_1584 ();
 FILLCELL_X32 FILLER_477_1616 ();
 FILLCELL_X32 FILLER_477_1648 ();
 FILLCELL_X32 FILLER_477_1680 ();
 FILLCELL_X32 FILLER_477_1712 ();
 FILLCELL_X32 FILLER_477_1744 ();
 FILLCELL_X32 FILLER_477_1776 ();
 FILLCELL_X32 FILLER_477_1808 ();
 FILLCELL_X32 FILLER_477_1840 ();
 FILLCELL_X32 FILLER_477_1872 ();
 FILLCELL_X32 FILLER_477_1904 ();
 FILLCELL_X32 FILLER_477_1936 ();
 FILLCELL_X32 FILLER_477_1968 ();
 FILLCELL_X32 FILLER_477_2000 ();
 FILLCELL_X32 FILLER_477_2032 ();
 FILLCELL_X32 FILLER_477_2064 ();
 FILLCELL_X32 FILLER_477_2096 ();
 FILLCELL_X32 FILLER_477_2128 ();
 FILLCELL_X32 FILLER_477_2160 ();
 FILLCELL_X32 FILLER_477_2192 ();
 FILLCELL_X32 FILLER_477_2224 ();
 FILLCELL_X32 FILLER_477_2256 ();
 FILLCELL_X32 FILLER_477_2288 ();
 FILLCELL_X32 FILLER_477_2320 ();
 FILLCELL_X32 FILLER_477_2352 ();
 FILLCELL_X32 FILLER_477_2384 ();
 FILLCELL_X32 FILLER_477_2416 ();
 FILLCELL_X32 FILLER_477_2448 ();
 FILLCELL_X32 FILLER_477_2480 ();
 FILLCELL_X8 FILLER_477_2512 ();
 FILLCELL_X4 FILLER_477_2520 ();
 FILLCELL_X2 FILLER_477_2524 ();
 FILLCELL_X32 FILLER_477_2527 ();
 FILLCELL_X32 FILLER_477_2559 ();
 FILLCELL_X32 FILLER_477_2591 ();
 FILLCELL_X32 FILLER_477_2623 ();
 FILLCELL_X32 FILLER_477_2655 ();
 FILLCELL_X32 FILLER_477_2687 ();
 FILLCELL_X32 FILLER_477_2719 ();
 FILLCELL_X32 FILLER_477_2751 ();
 FILLCELL_X32 FILLER_477_2783 ();
 FILLCELL_X32 FILLER_477_2815 ();
 FILLCELL_X32 FILLER_477_2847 ();
 FILLCELL_X32 FILLER_477_2879 ();
 FILLCELL_X32 FILLER_477_2911 ();
 FILLCELL_X32 FILLER_477_2943 ();
 FILLCELL_X32 FILLER_477_2975 ();
 FILLCELL_X32 FILLER_477_3007 ();
 FILLCELL_X32 FILLER_477_3039 ();
 FILLCELL_X32 FILLER_477_3071 ();
 FILLCELL_X32 FILLER_477_3103 ();
 FILLCELL_X32 FILLER_477_3135 ();
 FILLCELL_X32 FILLER_477_3167 ();
 FILLCELL_X32 FILLER_477_3199 ();
 FILLCELL_X32 FILLER_477_3231 ();
 FILLCELL_X32 FILLER_477_3263 ();
 FILLCELL_X32 FILLER_477_3295 ();
 FILLCELL_X32 FILLER_477_3327 ();
 FILLCELL_X32 FILLER_477_3359 ();
 FILLCELL_X32 FILLER_477_3391 ();
 FILLCELL_X32 FILLER_477_3423 ();
 FILLCELL_X32 FILLER_477_3455 ();
 FILLCELL_X32 FILLER_477_3487 ();
 FILLCELL_X32 FILLER_477_3519 ();
 FILLCELL_X32 FILLER_477_3551 ();
 FILLCELL_X32 FILLER_477_3583 ();
 FILLCELL_X32 FILLER_477_3615 ();
 FILLCELL_X32 FILLER_477_3647 ();
 FILLCELL_X32 FILLER_477_3679 ();
 FILLCELL_X16 FILLER_477_3711 ();
 FILLCELL_X8 FILLER_477_3727 ();
 FILLCELL_X2 FILLER_477_3735 ();
 FILLCELL_X1 FILLER_477_3737 ();
 FILLCELL_X32 FILLER_478_1 ();
 FILLCELL_X32 FILLER_478_33 ();
 FILLCELL_X32 FILLER_478_65 ();
 FILLCELL_X32 FILLER_478_97 ();
 FILLCELL_X32 FILLER_478_129 ();
 FILLCELL_X32 FILLER_478_161 ();
 FILLCELL_X32 FILLER_478_193 ();
 FILLCELL_X32 FILLER_478_225 ();
 FILLCELL_X32 FILLER_478_257 ();
 FILLCELL_X32 FILLER_478_289 ();
 FILLCELL_X32 FILLER_478_321 ();
 FILLCELL_X32 FILLER_478_353 ();
 FILLCELL_X32 FILLER_478_385 ();
 FILLCELL_X32 FILLER_478_417 ();
 FILLCELL_X32 FILLER_478_449 ();
 FILLCELL_X32 FILLER_478_481 ();
 FILLCELL_X32 FILLER_478_513 ();
 FILLCELL_X32 FILLER_478_545 ();
 FILLCELL_X32 FILLER_478_577 ();
 FILLCELL_X16 FILLER_478_609 ();
 FILLCELL_X4 FILLER_478_625 ();
 FILLCELL_X2 FILLER_478_629 ();
 FILLCELL_X32 FILLER_478_632 ();
 FILLCELL_X32 FILLER_478_664 ();
 FILLCELL_X32 FILLER_478_696 ();
 FILLCELL_X32 FILLER_478_728 ();
 FILLCELL_X32 FILLER_478_760 ();
 FILLCELL_X32 FILLER_478_792 ();
 FILLCELL_X32 FILLER_478_824 ();
 FILLCELL_X32 FILLER_478_856 ();
 FILLCELL_X32 FILLER_478_888 ();
 FILLCELL_X32 FILLER_478_920 ();
 FILLCELL_X32 FILLER_478_952 ();
 FILLCELL_X32 FILLER_478_984 ();
 FILLCELL_X32 FILLER_478_1016 ();
 FILLCELL_X32 FILLER_478_1048 ();
 FILLCELL_X32 FILLER_478_1080 ();
 FILLCELL_X32 FILLER_478_1112 ();
 FILLCELL_X32 FILLER_478_1144 ();
 FILLCELL_X32 FILLER_478_1176 ();
 FILLCELL_X32 FILLER_478_1208 ();
 FILLCELL_X32 FILLER_478_1240 ();
 FILLCELL_X32 FILLER_478_1272 ();
 FILLCELL_X32 FILLER_478_1304 ();
 FILLCELL_X32 FILLER_478_1336 ();
 FILLCELL_X32 FILLER_478_1368 ();
 FILLCELL_X32 FILLER_478_1400 ();
 FILLCELL_X32 FILLER_478_1432 ();
 FILLCELL_X32 FILLER_478_1464 ();
 FILLCELL_X32 FILLER_478_1496 ();
 FILLCELL_X32 FILLER_478_1528 ();
 FILLCELL_X32 FILLER_478_1560 ();
 FILLCELL_X32 FILLER_478_1592 ();
 FILLCELL_X32 FILLER_478_1624 ();
 FILLCELL_X32 FILLER_478_1656 ();
 FILLCELL_X32 FILLER_478_1688 ();
 FILLCELL_X32 FILLER_478_1720 ();
 FILLCELL_X32 FILLER_478_1752 ();
 FILLCELL_X32 FILLER_478_1784 ();
 FILLCELL_X32 FILLER_478_1816 ();
 FILLCELL_X32 FILLER_478_1848 ();
 FILLCELL_X8 FILLER_478_1880 ();
 FILLCELL_X4 FILLER_478_1888 ();
 FILLCELL_X2 FILLER_478_1892 ();
 FILLCELL_X32 FILLER_478_1895 ();
 FILLCELL_X32 FILLER_478_1927 ();
 FILLCELL_X32 FILLER_478_1959 ();
 FILLCELL_X32 FILLER_478_1991 ();
 FILLCELL_X32 FILLER_478_2023 ();
 FILLCELL_X32 FILLER_478_2055 ();
 FILLCELL_X32 FILLER_478_2087 ();
 FILLCELL_X32 FILLER_478_2119 ();
 FILLCELL_X32 FILLER_478_2151 ();
 FILLCELL_X32 FILLER_478_2183 ();
 FILLCELL_X32 FILLER_478_2215 ();
 FILLCELL_X32 FILLER_478_2247 ();
 FILLCELL_X32 FILLER_478_2279 ();
 FILLCELL_X32 FILLER_478_2311 ();
 FILLCELL_X32 FILLER_478_2343 ();
 FILLCELL_X32 FILLER_478_2375 ();
 FILLCELL_X32 FILLER_478_2407 ();
 FILLCELL_X32 FILLER_478_2439 ();
 FILLCELL_X32 FILLER_478_2471 ();
 FILLCELL_X32 FILLER_478_2503 ();
 FILLCELL_X32 FILLER_478_2535 ();
 FILLCELL_X32 FILLER_478_2567 ();
 FILLCELL_X32 FILLER_478_2599 ();
 FILLCELL_X32 FILLER_478_2631 ();
 FILLCELL_X32 FILLER_478_2663 ();
 FILLCELL_X32 FILLER_478_2695 ();
 FILLCELL_X32 FILLER_478_2727 ();
 FILLCELL_X32 FILLER_478_2759 ();
 FILLCELL_X32 FILLER_478_2791 ();
 FILLCELL_X32 FILLER_478_2823 ();
 FILLCELL_X32 FILLER_478_2855 ();
 FILLCELL_X32 FILLER_478_2887 ();
 FILLCELL_X32 FILLER_478_2919 ();
 FILLCELL_X32 FILLER_478_2951 ();
 FILLCELL_X32 FILLER_478_2983 ();
 FILLCELL_X32 FILLER_478_3015 ();
 FILLCELL_X32 FILLER_478_3047 ();
 FILLCELL_X32 FILLER_478_3079 ();
 FILLCELL_X32 FILLER_478_3111 ();
 FILLCELL_X8 FILLER_478_3143 ();
 FILLCELL_X4 FILLER_478_3151 ();
 FILLCELL_X2 FILLER_478_3155 ();
 FILLCELL_X32 FILLER_478_3158 ();
 FILLCELL_X32 FILLER_478_3190 ();
 FILLCELL_X32 FILLER_478_3222 ();
 FILLCELL_X32 FILLER_478_3254 ();
 FILLCELL_X32 FILLER_478_3286 ();
 FILLCELL_X32 FILLER_478_3318 ();
 FILLCELL_X32 FILLER_478_3350 ();
 FILLCELL_X32 FILLER_478_3382 ();
 FILLCELL_X32 FILLER_478_3414 ();
 FILLCELL_X32 FILLER_478_3446 ();
 FILLCELL_X32 FILLER_478_3478 ();
 FILLCELL_X32 FILLER_478_3510 ();
 FILLCELL_X32 FILLER_478_3542 ();
 FILLCELL_X32 FILLER_478_3574 ();
 FILLCELL_X32 FILLER_478_3606 ();
 FILLCELL_X32 FILLER_478_3638 ();
 FILLCELL_X32 FILLER_478_3670 ();
 FILLCELL_X32 FILLER_478_3702 ();
 FILLCELL_X4 FILLER_478_3734 ();
 FILLCELL_X32 FILLER_479_1 ();
 FILLCELL_X32 FILLER_479_33 ();
 FILLCELL_X32 FILLER_479_65 ();
 FILLCELL_X32 FILLER_479_97 ();
 FILLCELL_X32 FILLER_479_129 ();
 FILLCELL_X32 FILLER_479_161 ();
 FILLCELL_X32 FILLER_479_193 ();
 FILLCELL_X32 FILLER_479_225 ();
 FILLCELL_X32 FILLER_479_257 ();
 FILLCELL_X32 FILLER_479_289 ();
 FILLCELL_X32 FILLER_479_321 ();
 FILLCELL_X32 FILLER_479_353 ();
 FILLCELL_X32 FILLER_479_385 ();
 FILLCELL_X32 FILLER_479_417 ();
 FILLCELL_X32 FILLER_479_449 ();
 FILLCELL_X32 FILLER_479_481 ();
 FILLCELL_X32 FILLER_479_513 ();
 FILLCELL_X32 FILLER_479_545 ();
 FILLCELL_X32 FILLER_479_577 ();
 FILLCELL_X32 FILLER_479_609 ();
 FILLCELL_X32 FILLER_479_641 ();
 FILLCELL_X32 FILLER_479_673 ();
 FILLCELL_X32 FILLER_479_705 ();
 FILLCELL_X32 FILLER_479_737 ();
 FILLCELL_X32 FILLER_479_769 ();
 FILLCELL_X32 FILLER_479_801 ();
 FILLCELL_X32 FILLER_479_833 ();
 FILLCELL_X32 FILLER_479_865 ();
 FILLCELL_X32 FILLER_479_897 ();
 FILLCELL_X32 FILLER_479_929 ();
 FILLCELL_X32 FILLER_479_961 ();
 FILLCELL_X32 FILLER_479_993 ();
 FILLCELL_X32 FILLER_479_1025 ();
 FILLCELL_X32 FILLER_479_1057 ();
 FILLCELL_X32 FILLER_479_1089 ();
 FILLCELL_X32 FILLER_479_1121 ();
 FILLCELL_X32 FILLER_479_1153 ();
 FILLCELL_X32 FILLER_479_1185 ();
 FILLCELL_X32 FILLER_479_1217 ();
 FILLCELL_X8 FILLER_479_1249 ();
 FILLCELL_X4 FILLER_479_1257 ();
 FILLCELL_X2 FILLER_479_1261 ();
 FILLCELL_X32 FILLER_479_1264 ();
 FILLCELL_X32 FILLER_479_1296 ();
 FILLCELL_X32 FILLER_479_1328 ();
 FILLCELL_X32 FILLER_479_1360 ();
 FILLCELL_X32 FILLER_479_1392 ();
 FILLCELL_X32 FILLER_479_1424 ();
 FILLCELL_X32 FILLER_479_1456 ();
 FILLCELL_X32 FILLER_479_1488 ();
 FILLCELL_X32 FILLER_479_1520 ();
 FILLCELL_X32 FILLER_479_1552 ();
 FILLCELL_X32 FILLER_479_1584 ();
 FILLCELL_X32 FILLER_479_1616 ();
 FILLCELL_X32 FILLER_479_1648 ();
 FILLCELL_X32 FILLER_479_1680 ();
 FILLCELL_X32 FILLER_479_1712 ();
 FILLCELL_X32 FILLER_479_1744 ();
 FILLCELL_X32 FILLER_479_1776 ();
 FILLCELL_X32 FILLER_479_1808 ();
 FILLCELL_X32 FILLER_479_1840 ();
 FILLCELL_X32 FILLER_479_1872 ();
 FILLCELL_X32 FILLER_479_1904 ();
 FILLCELL_X32 FILLER_479_1936 ();
 FILLCELL_X32 FILLER_479_1968 ();
 FILLCELL_X32 FILLER_479_2000 ();
 FILLCELL_X32 FILLER_479_2032 ();
 FILLCELL_X32 FILLER_479_2064 ();
 FILLCELL_X32 FILLER_479_2096 ();
 FILLCELL_X32 FILLER_479_2128 ();
 FILLCELL_X32 FILLER_479_2160 ();
 FILLCELL_X32 FILLER_479_2192 ();
 FILLCELL_X32 FILLER_479_2224 ();
 FILLCELL_X32 FILLER_479_2256 ();
 FILLCELL_X32 FILLER_479_2288 ();
 FILLCELL_X32 FILLER_479_2320 ();
 FILLCELL_X32 FILLER_479_2352 ();
 FILLCELL_X32 FILLER_479_2384 ();
 FILLCELL_X32 FILLER_479_2416 ();
 FILLCELL_X32 FILLER_479_2448 ();
 FILLCELL_X32 FILLER_479_2480 ();
 FILLCELL_X8 FILLER_479_2512 ();
 FILLCELL_X4 FILLER_479_2520 ();
 FILLCELL_X2 FILLER_479_2524 ();
 FILLCELL_X32 FILLER_479_2527 ();
 FILLCELL_X32 FILLER_479_2559 ();
 FILLCELL_X32 FILLER_479_2591 ();
 FILLCELL_X32 FILLER_479_2623 ();
 FILLCELL_X32 FILLER_479_2655 ();
 FILLCELL_X32 FILLER_479_2687 ();
 FILLCELL_X32 FILLER_479_2719 ();
 FILLCELL_X32 FILLER_479_2751 ();
 FILLCELL_X32 FILLER_479_2783 ();
 FILLCELL_X32 FILLER_479_2815 ();
 FILLCELL_X32 FILLER_479_2847 ();
 FILLCELL_X32 FILLER_479_2879 ();
 FILLCELL_X32 FILLER_479_2911 ();
 FILLCELL_X32 FILLER_479_2943 ();
 FILLCELL_X32 FILLER_479_2975 ();
 FILLCELL_X32 FILLER_479_3007 ();
 FILLCELL_X32 FILLER_479_3039 ();
 FILLCELL_X32 FILLER_479_3071 ();
 FILLCELL_X32 FILLER_479_3103 ();
 FILLCELL_X32 FILLER_479_3135 ();
 FILLCELL_X32 FILLER_479_3167 ();
 FILLCELL_X32 FILLER_479_3199 ();
 FILLCELL_X32 FILLER_479_3231 ();
 FILLCELL_X32 FILLER_479_3263 ();
 FILLCELL_X32 FILLER_479_3295 ();
 FILLCELL_X32 FILLER_479_3327 ();
 FILLCELL_X32 FILLER_479_3359 ();
 FILLCELL_X32 FILLER_479_3391 ();
 FILLCELL_X32 FILLER_479_3423 ();
 FILLCELL_X32 FILLER_479_3455 ();
 FILLCELL_X32 FILLER_479_3487 ();
 FILLCELL_X32 FILLER_479_3519 ();
 FILLCELL_X32 FILLER_479_3551 ();
 FILLCELL_X32 FILLER_479_3583 ();
 FILLCELL_X32 FILLER_479_3615 ();
 FILLCELL_X32 FILLER_479_3647 ();
 FILLCELL_X32 FILLER_479_3679 ();
 FILLCELL_X16 FILLER_479_3711 ();
 FILLCELL_X8 FILLER_479_3727 ();
 FILLCELL_X2 FILLER_479_3735 ();
 FILLCELL_X1 FILLER_479_3737 ();
 FILLCELL_X32 FILLER_480_1 ();
 FILLCELL_X32 FILLER_480_33 ();
 FILLCELL_X32 FILLER_480_65 ();
 FILLCELL_X32 FILLER_480_97 ();
 FILLCELL_X32 FILLER_480_129 ();
 FILLCELL_X32 FILLER_480_161 ();
 FILLCELL_X32 FILLER_480_193 ();
 FILLCELL_X32 FILLER_480_225 ();
 FILLCELL_X32 FILLER_480_257 ();
 FILLCELL_X32 FILLER_480_289 ();
 FILLCELL_X32 FILLER_480_321 ();
 FILLCELL_X32 FILLER_480_353 ();
 FILLCELL_X32 FILLER_480_385 ();
 FILLCELL_X32 FILLER_480_417 ();
 FILLCELL_X32 FILLER_480_449 ();
 FILLCELL_X32 FILLER_480_481 ();
 FILLCELL_X32 FILLER_480_513 ();
 FILLCELL_X32 FILLER_480_545 ();
 FILLCELL_X32 FILLER_480_577 ();
 FILLCELL_X16 FILLER_480_609 ();
 FILLCELL_X4 FILLER_480_625 ();
 FILLCELL_X2 FILLER_480_629 ();
 FILLCELL_X32 FILLER_480_632 ();
 FILLCELL_X32 FILLER_480_664 ();
 FILLCELL_X32 FILLER_480_696 ();
 FILLCELL_X32 FILLER_480_728 ();
 FILLCELL_X32 FILLER_480_760 ();
 FILLCELL_X32 FILLER_480_792 ();
 FILLCELL_X32 FILLER_480_824 ();
 FILLCELL_X32 FILLER_480_856 ();
 FILLCELL_X32 FILLER_480_888 ();
 FILLCELL_X32 FILLER_480_920 ();
 FILLCELL_X32 FILLER_480_952 ();
 FILLCELL_X32 FILLER_480_984 ();
 FILLCELL_X32 FILLER_480_1016 ();
 FILLCELL_X32 FILLER_480_1048 ();
 FILLCELL_X32 FILLER_480_1080 ();
 FILLCELL_X32 FILLER_480_1112 ();
 FILLCELL_X32 FILLER_480_1144 ();
 FILLCELL_X32 FILLER_480_1176 ();
 FILLCELL_X32 FILLER_480_1208 ();
 FILLCELL_X32 FILLER_480_1240 ();
 FILLCELL_X32 FILLER_480_1272 ();
 FILLCELL_X32 FILLER_480_1304 ();
 FILLCELL_X32 FILLER_480_1336 ();
 FILLCELL_X32 FILLER_480_1368 ();
 FILLCELL_X32 FILLER_480_1400 ();
 FILLCELL_X32 FILLER_480_1432 ();
 FILLCELL_X32 FILLER_480_1464 ();
 FILLCELL_X32 FILLER_480_1496 ();
 FILLCELL_X32 FILLER_480_1528 ();
 FILLCELL_X32 FILLER_480_1560 ();
 FILLCELL_X32 FILLER_480_1592 ();
 FILLCELL_X32 FILLER_480_1624 ();
 FILLCELL_X32 FILLER_480_1656 ();
 FILLCELL_X32 FILLER_480_1688 ();
 FILLCELL_X32 FILLER_480_1720 ();
 FILLCELL_X32 FILLER_480_1752 ();
 FILLCELL_X32 FILLER_480_1784 ();
 FILLCELL_X32 FILLER_480_1816 ();
 FILLCELL_X32 FILLER_480_1848 ();
 FILLCELL_X8 FILLER_480_1880 ();
 FILLCELL_X4 FILLER_480_1888 ();
 FILLCELL_X2 FILLER_480_1892 ();
 FILLCELL_X32 FILLER_480_1895 ();
 FILLCELL_X32 FILLER_480_1927 ();
 FILLCELL_X32 FILLER_480_1959 ();
 FILLCELL_X32 FILLER_480_1991 ();
 FILLCELL_X32 FILLER_480_2023 ();
 FILLCELL_X32 FILLER_480_2055 ();
 FILLCELL_X32 FILLER_480_2087 ();
 FILLCELL_X32 FILLER_480_2119 ();
 FILLCELL_X32 FILLER_480_2151 ();
 FILLCELL_X32 FILLER_480_2183 ();
 FILLCELL_X32 FILLER_480_2215 ();
 FILLCELL_X32 FILLER_480_2247 ();
 FILLCELL_X32 FILLER_480_2279 ();
 FILLCELL_X32 FILLER_480_2311 ();
 FILLCELL_X32 FILLER_480_2343 ();
 FILLCELL_X32 FILLER_480_2375 ();
 FILLCELL_X32 FILLER_480_2407 ();
 FILLCELL_X32 FILLER_480_2439 ();
 FILLCELL_X32 FILLER_480_2471 ();
 FILLCELL_X32 FILLER_480_2503 ();
 FILLCELL_X32 FILLER_480_2535 ();
 FILLCELL_X32 FILLER_480_2567 ();
 FILLCELL_X32 FILLER_480_2599 ();
 FILLCELL_X32 FILLER_480_2631 ();
 FILLCELL_X32 FILLER_480_2663 ();
 FILLCELL_X32 FILLER_480_2695 ();
 FILLCELL_X32 FILLER_480_2727 ();
 FILLCELL_X32 FILLER_480_2759 ();
 FILLCELL_X32 FILLER_480_2791 ();
 FILLCELL_X32 FILLER_480_2823 ();
 FILLCELL_X32 FILLER_480_2855 ();
 FILLCELL_X32 FILLER_480_2887 ();
 FILLCELL_X32 FILLER_480_2919 ();
 FILLCELL_X32 FILLER_480_2951 ();
 FILLCELL_X32 FILLER_480_2983 ();
 FILLCELL_X32 FILLER_480_3015 ();
 FILLCELL_X32 FILLER_480_3047 ();
 FILLCELL_X32 FILLER_480_3079 ();
 FILLCELL_X32 FILLER_480_3111 ();
 FILLCELL_X8 FILLER_480_3143 ();
 FILLCELL_X4 FILLER_480_3151 ();
 FILLCELL_X2 FILLER_480_3155 ();
 FILLCELL_X32 FILLER_480_3158 ();
 FILLCELL_X32 FILLER_480_3190 ();
 FILLCELL_X32 FILLER_480_3222 ();
 FILLCELL_X32 FILLER_480_3254 ();
 FILLCELL_X32 FILLER_480_3286 ();
 FILLCELL_X32 FILLER_480_3318 ();
 FILLCELL_X32 FILLER_480_3350 ();
 FILLCELL_X32 FILLER_480_3382 ();
 FILLCELL_X32 FILLER_480_3414 ();
 FILLCELL_X32 FILLER_480_3446 ();
 FILLCELL_X32 FILLER_480_3478 ();
 FILLCELL_X32 FILLER_480_3510 ();
 FILLCELL_X32 FILLER_480_3542 ();
 FILLCELL_X32 FILLER_480_3574 ();
 FILLCELL_X32 FILLER_480_3606 ();
 FILLCELL_X32 FILLER_480_3638 ();
 FILLCELL_X32 FILLER_480_3670 ();
 FILLCELL_X32 FILLER_480_3702 ();
 FILLCELL_X4 FILLER_480_3734 ();
 FILLCELL_X32 FILLER_481_1 ();
 FILLCELL_X32 FILLER_481_33 ();
 FILLCELL_X32 FILLER_481_65 ();
 FILLCELL_X32 FILLER_481_97 ();
 FILLCELL_X32 FILLER_481_129 ();
 FILLCELL_X32 FILLER_481_161 ();
 FILLCELL_X32 FILLER_481_193 ();
 FILLCELL_X32 FILLER_481_225 ();
 FILLCELL_X32 FILLER_481_257 ();
 FILLCELL_X32 FILLER_481_289 ();
 FILLCELL_X32 FILLER_481_321 ();
 FILLCELL_X32 FILLER_481_353 ();
 FILLCELL_X32 FILLER_481_385 ();
 FILLCELL_X32 FILLER_481_417 ();
 FILLCELL_X32 FILLER_481_449 ();
 FILLCELL_X32 FILLER_481_481 ();
 FILLCELL_X32 FILLER_481_513 ();
 FILLCELL_X32 FILLER_481_545 ();
 FILLCELL_X32 FILLER_481_577 ();
 FILLCELL_X32 FILLER_481_609 ();
 FILLCELL_X32 FILLER_481_641 ();
 FILLCELL_X32 FILLER_481_673 ();
 FILLCELL_X32 FILLER_481_705 ();
 FILLCELL_X32 FILLER_481_737 ();
 FILLCELL_X32 FILLER_481_769 ();
 FILLCELL_X32 FILLER_481_801 ();
 FILLCELL_X32 FILLER_481_833 ();
 FILLCELL_X32 FILLER_481_865 ();
 FILLCELL_X32 FILLER_481_897 ();
 FILLCELL_X32 FILLER_481_929 ();
 FILLCELL_X32 FILLER_481_961 ();
 FILLCELL_X32 FILLER_481_993 ();
 FILLCELL_X32 FILLER_481_1025 ();
 FILLCELL_X32 FILLER_481_1057 ();
 FILLCELL_X32 FILLER_481_1089 ();
 FILLCELL_X32 FILLER_481_1121 ();
 FILLCELL_X32 FILLER_481_1153 ();
 FILLCELL_X32 FILLER_481_1185 ();
 FILLCELL_X32 FILLER_481_1217 ();
 FILLCELL_X8 FILLER_481_1249 ();
 FILLCELL_X4 FILLER_481_1257 ();
 FILLCELL_X2 FILLER_481_1261 ();
 FILLCELL_X32 FILLER_481_1264 ();
 FILLCELL_X32 FILLER_481_1296 ();
 FILLCELL_X32 FILLER_481_1328 ();
 FILLCELL_X32 FILLER_481_1360 ();
 FILLCELL_X32 FILLER_481_1392 ();
 FILLCELL_X32 FILLER_481_1424 ();
 FILLCELL_X32 FILLER_481_1456 ();
 FILLCELL_X32 FILLER_481_1488 ();
 FILLCELL_X32 FILLER_481_1520 ();
 FILLCELL_X32 FILLER_481_1552 ();
 FILLCELL_X32 FILLER_481_1584 ();
 FILLCELL_X32 FILLER_481_1616 ();
 FILLCELL_X32 FILLER_481_1648 ();
 FILLCELL_X32 FILLER_481_1680 ();
 FILLCELL_X32 FILLER_481_1712 ();
 FILLCELL_X32 FILLER_481_1744 ();
 FILLCELL_X32 FILLER_481_1776 ();
 FILLCELL_X32 FILLER_481_1808 ();
 FILLCELL_X32 FILLER_481_1840 ();
 FILLCELL_X32 FILLER_481_1872 ();
 FILLCELL_X32 FILLER_481_1904 ();
 FILLCELL_X32 FILLER_481_1936 ();
 FILLCELL_X32 FILLER_481_1968 ();
 FILLCELL_X32 FILLER_481_2000 ();
 FILLCELL_X32 FILLER_481_2032 ();
 FILLCELL_X32 FILLER_481_2064 ();
 FILLCELL_X32 FILLER_481_2096 ();
 FILLCELL_X32 FILLER_481_2128 ();
 FILLCELL_X32 FILLER_481_2160 ();
 FILLCELL_X32 FILLER_481_2192 ();
 FILLCELL_X32 FILLER_481_2224 ();
 FILLCELL_X32 FILLER_481_2256 ();
 FILLCELL_X32 FILLER_481_2288 ();
 FILLCELL_X32 FILLER_481_2320 ();
 FILLCELL_X32 FILLER_481_2352 ();
 FILLCELL_X32 FILLER_481_2384 ();
 FILLCELL_X32 FILLER_481_2416 ();
 FILLCELL_X32 FILLER_481_2448 ();
 FILLCELL_X32 FILLER_481_2480 ();
 FILLCELL_X8 FILLER_481_2512 ();
 FILLCELL_X4 FILLER_481_2520 ();
 FILLCELL_X2 FILLER_481_2524 ();
 FILLCELL_X32 FILLER_481_2527 ();
 FILLCELL_X32 FILLER_481_2559 ();
 FILLCELL_X32 FILLER_481_2591 ();
 FILLCELL_X32 FILLER_481_2623 ();
 FILLCELL_X32 FILLER_481_2655 ();
 FILLCELL_X32 FILLER_481_2687 ();
 FILLCELL_X32 FILLER_481_2719 ();
 FILLCELL_X32 FILLER_481_2751 ();
 FILLCELL_X32 FILLER_481_2783 ();
 FILLCELL_X32 FILLER_481_2815 ();
 FILLCELL_X32 FILLER_481_2847 ();
 FILLCELL_X32 FILLER_481_2879 ();
 FILLCELL_X32 FILLER_481_2911 ();
 FILLCELL_X32 FILLER_481_2943 ();
 FILLCELL_X32 FILLER_481_2975 ();
 FILLCELL_X32 FILLER_481_3007 ();
 FILLCELL_X32 FILLER_481_3039 ();
 FILLCELL_X32 FILLER_481_3071 ();
 FILLCELL_X32 FILLER_481_3103 ();
 FILLCELL_X32 FILLER_481_3135 ();
 FILLCELL_X32 FILLER_481_3167 ();
 FILLCELL_X32 FILLER_481_3199 ();
 FILLCELL_X32 FILLER_481_3231 ();
 FILLCELL_X32 FILLER_481_3263 ();
 FILLCELL_X32 FILLER_481_3295 ();
 FILLCELL_X32 FILLER_481_3327 ();
 FILLCELL_X32 FILLER_481_3359 ();
 FILLCELL_X32 FILLER_481_3391 ();
 FILLCELL_X32 FILLER_481_3423 ();
 FILLCELL_X32 FILLER_481_3455 ();
 FILLCELL_X32 FILLER_481_3487 ();
 FILLCELL_X32 FILLER_481_3519 ();
 FILLCELL_X32 FILLER_481_3551 ();
 FILLCELL_X32 FILLER_481_3583 ();
 FILLCELL_X32 FILLER_481_3615 ();
 FILLCELL_X32 FILLER_481_3647 ();
 FILLCELL_X32 FILLER_481_3679 ();
 FILLCELL_X16 FILLER_481_3711 ();
 FILLCELL_X8 FILLER_481_3727 ();
 FILLCELL_X2 FILLER_481_3735 ();
 FILLCELL_X1 FILLER_481_3737 ();
 FILLCELL_X32 FILLER_482_1 ();
 FILLCELL_X32 FILLER_482_33 ();
 FILLCELL_X32 FILLER_482_65 ();
 FILLCELL_X32 FILLER_482_97 ();
 FILLCELL_X32 FILLER_482_129 ();
 FILLCELL_X32 FILLER_482_161 ();
 FILLCELL_X32 FILLER_482_193 ();
 FILLCELL_X32 FILLER_482_225 ();
 FILLCELL_X32 FILLER_482_257 ();
 FILLCELL_X32 FILLER_482_289 ();
 FILLCELL_X32 FILLER_482_321 ();
 FILLCELL_X32 FILLER_482_353 ();
 FILLCELL_X32 FILLER_482_385 ();
 FILLCELL_X32 FILLER_482_417 ();
 FILLCELL_X32 FILLER_482_449 ();
 FILLCELL_X32 FILLER_482_481 ();
 FILLCELL_X32 FILLER_482_513 ();
 FILLCELL_X32 FILLER_482_545 ();
 FILLCELL_X32 FILLER_482_577 ();
 FILLCELL_X16 FILLER_482_609 ();
 FILLCELL_X4 FILLER_482_625 ();
 FILLCELL_X2 FILLER_482_629 ();
 FILLCELL_X32 FILLER_482_632 ();
 FILLCELL_X32 FILLER_482_664 ();
 FILLCELL_X32 FILLER_482_696 ();
 FILLCELL_X32 FILLER_482_728 ();
 FILLCELL_X32 FILLER_482_760 ();
 FILLCELL_X32 FILLER_482_792 ();
 FILLCELL_X32 FILLER_482_824 ();
 FILLCELL_X32 FILLER_482_856 ();
 FILLCELL_X32 FILLER_482_888 ();
 FILLCELL_X32 FILLER_482_920 ();
 FILLCELL_X32 FILLER_482_952 ();
 FILLCELL_X32 FILLER_482_984 ();
 FILLCELL_X32 FILLER_482_1016 ();
 FILLCELL_X32 FILLER_482_1048 ();
 FILLCELL_X32 FILLER_482_1080 ();
 FILLCELL_X32 FILLER_482_1112 ();
 FILLCELL_X32 FILLER_482_1144 ();
 FILLCELL_X32 FILLER_482_1176 ();
 FILLCELL_X32 FILLER_482_1208 ();
 FILLCELL_X32 FILLER_482_1240 ();
 FILLCELL_X32 FILLER_482_1272 ();
 FILLCELL_X32 FILLER_482_1304 ();
 FILLCELL_X32 FILLER_482_1336 ();
 FILLCELL_X32 FILLER_482_1368 ();
 FILLCELL_X32 FILLER_482_1400 ();
 FILLCELL_X32 FILLER_482_1432 ();
 FILLCELL_X32 FILLER_482_1464 ();
 FILLCELL_X32 FILLER_482_1496 ();
 FILLCELL_X32 FILLER_482_1528 ();
 FILLCELL_X32 FILLER_482_1560 ();
 FILLCELL_X32 FILLER_482_1592 ();
 FILLCELL_X32 FILLER_482_1624 ();
 FILLCELL_X32 FILLER_482_1656 ();
 FILLCELL_X32 FILLER_482_1688 ();
 FILLCELL_X32 FILLER_482_1720 ();
 FILLCELL_X32 FILLER_482_1752 ();
 FILLCELL_X32 FILLER_482_1784 ();
 FILLCELL_X32 FILLER_482_1816 ();
 FILLCELL_X32 FILLER_482_1848 ();
 FILLCELL_X8 FILLER_482_1880 ();
 FILLCELL_X4 FILLER_482_1888 ();
 FILLCELL_X2 FILLER_482_1892 ();
 FILLCELL_X32 FILLER_482_1895 ();
 FILLCELL_X32 FILLER_482_1927 ();
 FILLCELL_X32 FILLER_482_1959 ();
 FILLCELL_X32 FILLER_482_1991 ();
 FILLCELL_X32 FILLER_482_2023 ();
 FILLCELL_X32 FILLER_482_2055 ();
 FILLCELL_X32 FILLER_482_2087 ();
 FILLCELL_X32 FILLER_482_2119 ();
 FILLCELL_X32 FILLER_482_2151 ();
 FILLCELL_X32 FILLER_482_2183 ();
 FILLCELL_X32 FILLER_482_2215 ();
 FILLCELL_X32 FILLER_482_2247 ();
 FILLCELL_X32 FILLER_482_2279 ();
 FILLCELL_X32 FILLER_482_2311 ();
 FILLCELL_X32 FILLER_482_2343 ();
 FILLCELL_X32 FILLER_482_2375 ();
 FILLCELL_X32 FILLER_482_2407 ();
 FILLCELL_X32 FILLER_482_2439 ();
 FILLCELL_X32 FILLER_482_2471 ();
 FILLCELL_X32 FILLER_482_2503 ();
 FILLCELL_X32 FILLER_482_2535 ();
 FILLCELL_X32 FILLER_482_2567 ();
 FILLCELL_X32 FILLER_482_2599 ();
 FILLCELL_X32 FILLER_482_2631 ();
 FILLCELL_X32 FILLER_482_2663 ();
 FILLCELL_X32 FILLER_482_2695 ();
 FILLCELL_X32 FILLER_482_2727 ();
 FILLCELL_X32 FILLER_482_2759 ();
 FILLCELL_X32 FILLER_482_2791 ();
 FILLCELL_X32 FILLER_482_2823 ();
 FILLCELL_X32 FILLER_482_2855 ();
 FILLCELL_X32 FILLER_482_2887 ();
 FILLCELL_X32 FILLER_482_2919 ();
 FILLCELL_X32 FILLER_482_2951 ();
 FILLCELL_X32 FILLER_482_2983 ();
 FILLCELL_X32 FILLER_482_3015 ();
 FILLCELL_X32 FILLER_482_3047 ();
 FILLCELL_X32 FILLER_482_3079 ();
 FILLCELL_X32 FILLER_482_3111 ();
 FILLCELL_X8 FILLER_482_3143 ();
 FILLCELL_X4 FILLER_482_3151 ();
 FILLCELL_X2 FILLER_482_3155 ();
 FILLCELL_X32 FILLER_482_3158 ();
 FILLCELL_X32 FILLER_482_3190 ();
 FILLCELL_X32 FILLER_482_3222 ();
 FILLCELL_X32 FILLER_482_3254 ();
 FILLCELL_X32 FILLER_482_3286 ();
 FILLCELL_X32 FILLER_482_3318 ();
 FILLCELL_X32 FILLER_482_3350 ();
 FILLCELL_X32 FILLER_482_3382 ();
 FILLCELL_X32 FILLER_482_3414 ();
 FILLCELL_X32 FILLER_482_3446 ();
 FILLCELL_X32 FILLER_482_3478 ();
 FILLCELL_X32 FILLER_482_3510 ();
 FILLCELL_X32 FILLER_482_3542 ();
 FILLCELL_X32 FILLER_482_3574 ();
 FILLCELL_X32 FILLER_482_3606 ();
 FILLCELL_X32 FILLER_482_3638 ();
 FILLCELL_X32 FILLER_482_3670 ();
 FILLCELL_X32 FILLER_482_3702 ();
 FILLCELL_X4 FILLER_482_3734 ();
 FILLCELL_X32 FILLER_483_1 ();
 FILLCELL_X32 FILLER_483_33 ();
 FILLCELL_X32 FILLER_483_65 ();
 FILLCELL_X32 FILLER_483_97 ();
 FILLCELL_X32 FILLER_483_129 ();
 FILLCELL_X32 FILLER_483_161 ();
 FILLCELL_X32 FILLER_483_193 ();
 FILLCELL_X32 FILLER_483_225 ();
 FILLCELL_X32 FILLER_483_257 ();
 FILLCELL_X32 FILLER_483_289 ();
 FILLCELL_X32 FILLER_483_321 ();
 FILLCELL_X32 FILLER_483_353 ();
 FILLCELL_X32 FILLER_483_385 ();
 FILLCELL_X32 FILLER_483_417 ();
 FILLCELL_X32 FILLER_483_449 ();
 FILLCELL_X32 FILLER_483_481 ();
 FILLCELL_X32 FILLER_483_513 ();
 FILLCELL_X32 FILLER_483_545 ();
 FILLCELL_X32 FILLER_483_577 ();
 FILLCELL_X32 FILLER_483_609 ();
 FILLCELL_X32 FILLER_483_641 ();
 FILLCELL_X32 FILLER_483_673 ();
 FILLCELL_X32 FILLER_483_705 ();
 FILLCELL_X32 FILLER_483_737 ();
 FILLCELL_X32 FILLER_483_769 ();
 FILLCELL_X32 FILLER_483_801 ();
 FILLCELL_X32 FILLER_483_833 ();
 FILLCELL_X32 FILLER_483_865 ();
 FILLCELL_X32 FILLER_483_897 ();
 FILLCELL_X32 FILLER_483_929 ();
 FILLCELL_X32 FILLER_483_961 ();
 FILLCELL_X32 FILLER_483_993 ();
 FILLCELL_X32 FILLER_483_1025 ();
 FILLCELL_X32 FILLER_483_1057 ();
 FILLCELL_X32 FILLER_483_1089 ();
 FILLCELL_X32 FILLER_483_1121 ();
 FILLCELL_X32 FILLER_483_1153 ();
 FILLCELL_X32 FILLER_483_1185 ();
 FILLCELL_X32 FILLER_483_1217 ();
 FILLCELL_X8 FILLER_483_1249 ();
 FILLCELL_X4 FILLER_483_1257 ();
 FILLCELL_X2 FILLER_483_1261 ();
 FILLCELL_X32 FILLER_483_1264 ();
 FILLCELL_X32 FILLER_483_1296 ();
 FILLCELL_X32 FILLER_483_1328 ();
 FILLCELL_X32 FILLER_483_1360 ();
 FILLCELL_X32 FILLER_483_1392 ();
 FILLCELL_X32 FILLER_483_1424 ();
 FILLCELL_X32 FILLER_483_1456 ();
 FILLCELL_X32 FILLER_483_1488 ();
 FILLCELL_X32 FILLER_483_1520 ();
 FILLCELL_X32 FILLER_483_1552 ();
 FILLCELL_X32 FILLER_483_1584 ();
 FILLCELL_X32 FILLER_483_1616 ();
 FILLCELL_X32 FILLER_483_1648 ();
 FILLCELL_X32 FILLER_483_1680 ();
 FILLCELL_X32 FILLER_483_1712 ();
 FILLCELL_X32 FILLER_483_1744 ();
 FILLCELL_X32 FILLER_483_1776 ();
 FILLCELL_X32 FILLER_483_1808 ();
 FILLCELL_X32 FILLER_483_1840 ();
 FILLCELL_X32 FILLER_483_1872 ();
 FILLCELL_X32 FILLER_483_1904 ();
 FILLCELL_X32 FILLER_483_1936 ();
 FILLCELL_X32 FILLER_483_1968 ();
 FILLCELL_X32 FILLER_483_2000 ();
 FILLCELL_X32 FILLER_483_2032 ();
 FILLCELL_X32 FILLER_483_2064 ();
 FILLCELL_X32 FILLER_483_2096 ();
 FILLCELL_X32 FILLER_483_2128 ();
 FILLCELL_X32 FILLER_483_2160 ();
 FILLCELL_X32 FILLER_483_2192 ();
 FILLCELL_X32 FILLER_483_2224 ();
 FILLCELL_X32 FILLER_483_2256 ();
 FILLCELL_X32 FILLER_483_2288 ();
 FILLCELL_X32 FILLER_483_2320 ();
 FILLCELL_X32 FILLER_483_2352 ();
 FILLCELL_X32 FILLER_483_2384 ();
 FILLCELL_X32 FILLER_483_2416 ();
 FILLCELL_X32 FILLER_483_2448 ();
 FILLCELL_X32 FILLER_483_2480 ();
 FILLCELL_X8 FILLER_483_2512 ();
 FILLCELL_X4 FILLER_483_2520 ();
 FILLCELL_X2 FILLER_483_2524 ();
 FILLCELL_X32 FILLER_483_2527 ();
 FILLCELL_X32 FILLER_483_2559 ();
 FILLCELL_X32 FILLER_483_2591 ();
 FILLCELL_X32 FILLER_483_2623 ();
 FILLCELL_X32 FILLER_483_2655 ();
 FILLCELL_X32 FILLER_483_2687 ();
 FILLCELL_X32 FILLER_483_2719 ();
 FILLCELL_X32 FILLER_483_2751 ();
 FILLCELL_X32 FILLER_483_2783 ();
 FILLCELL_X32 FILLER_483_2815 ();
 FILLCELL_X32 FILLER_483_2847 ();
 FILLCELL_X32 FILLER_483_2879 ();
 FILLCELL_X32 FILLER_483_2911 ();
 FILLCELL_X32 FILLER_483_2943 ();
 FILLCELL_X32 FILLER_483_2975 ();
 FILLCELL_X32 FILLER_483_3007 ();
 FILLCELL_X32 FILLER_483_3039 ();
 FILLCELL_X32 FILLER_483_3071 ();
 FILLCELL_X32 FILLER_483_3103 ();
 FILLCELL_X32 FILLER_483_3135 ();
 FILLCELL_X32 FILLER_483_3167 ();
 FILLCELL_X32 FILLER_483_3199 ();
 FILLCELL_X32 FILLER_483_3231 ();
 FILLCELL_X32 FILLER_483_3263 ();
 FILLCELL_X32 FILLER_483_3295 ();
 FILLCELL_X32 FILLER_483_3327 ();
 FILLCELL_X32 FILLER_483_3359 ();
 FILLCELL_X32 FILLER_483_3391 ();
 FILLCELL_X32 FILLER_483_3423 ();
 FILLCELL_X32 FILLER_483_3455 ();
 FILLCELL_X32 FILLER_483_3487 ();
 FILLCELL_X32 FILLER_483_3519 ();
 FILLCELL_X32 FILLER_483_3551 ();
 FILLCELL_X32 FILLER_483_3583 ();
 FILLCELL_X32 FILLER_483_3615 ();
 FILLCELL_X32 FILLER_483_3647 ();
 FILLCELL_X32 FILLER_483_3679 ();
 FILLCELL_X16 FILLER_483_3711 ();
 FILLCELL_X8 FILLER_483_3727 ();
 FILLCELL_X2 FILLER_483_3735 ();
 FILLCELL_X1 FILLER_483_3737 ();
 FILLCELL_X32 FILLER_484_1 ();
 FILLCELL_X32 FILLER_484_33 ();
 FILLCELL_X32 FILLER_484_65 ();
 FILLCELL_X32 FILLER_484_97 ();
 FILLCELL_X32 FILLER_484_129 ();
 FILLCELL_X32 FILLER_484_161 ();
 FILLCELL_X32 FILLER_484_193 ();
 FILLCELL_X32 FILLER_484_225 ();
 FILLCELL_X32 FILLER_484_257 ();
 FILLCELL_X32 FILLER_484_289 ();
 FILLCELL_X32 FILLER_484_321 ();
 FILLCELL_X32 FILLER_484_353 ();
 FILLCELL_X32 FILLER_484_385 ();
 FILLCELL_X32 FILLER_484_417 ();
 FILLCELL_X32 FILLER_484_449 ();
 FILLCELL_X32 FILLER_484_481 ();
 FILLCELL_X32 FILLER_484_513 ();
 FILLCELL_X32 FILLER_484_545 ();
 FILLCELL_X32 FILLER_484_577 ();
 FILLCELL_X16 FILLER_484_609 ();
 FILLCELL_X4 FILLER_484_625 ();
 FILLCELL_X2 FILLER_484_629 ();
 FILLCELL_X32 FILLER_484_632 ();
 FILLCELL_X32 FILLER_484_664 ();
 FILLCELL_X32 FILLER_484_696 ();
 FILLCELL_X32 FILLER_484_728 ();
 FILLCELL_X32 FILLER_484_760 ();
 FILLCELL_X32 FILLER_484_792 ();
 FILLCELL_X32 FILLER_484_824 ();
 FILLCELL_X32 FILLER_484_856 ();
 FILLCELL_X32 FILLER_484_888 ();
 FILLCELL_X32 FILLER_484_920 ();
 FILLCELL_X32 FILLER_484_952 ();
 FILLCELL_X32 FILLER_484_984 ();
 FILLCELL_X32 FILLER_484_1016 ();
 FILLCELL_X32 FILLER_484_1048 ();
 FILLCELL_X32 FILLER_484_1080 ();
 FILLCELL_X32 FILLER_484_1112 ();
 FILLCELL_X32 FILLER_484_1144 ();
 FILLCELL_X32 FILLER_484_1176 ();
 FILLCELL_X32 FILLER_484_1208 ();
 FILLCELL_X32 FILLER_484_1240 ();
 FILLCELL_X32 FILLER_484_1272 ();
 FILLCELL_X32 FILLER_484_1304 ();
 FILLCELL_X32 FILLER_484_1336 ();
 FILLCELL_X32 FILLER_484_1368 ();
 FILLCELL_X32 FILLER_484_1400 ();
 FILLCELL_X32 FILLER_484_1432 ();
 FILLCELL_X32 FILLER_484_1464 ();
 FILLCELL_X32 FILLER_484_1496 ();
 FILLCELL_X32 FILLER_484_1528 ();
 FILLCELL_X32 FILLER_484_1560 ();
 FILLCELL_X32 FILLER_484_1592 ();
 FILLCELL_X32 FILLER_484_1624 ();
 FILLCELL_X32 FILLER_484_1656 ();
 FILLCELL_X32 FILLER_484_1688 ();
 FILLCELL_X32 FILLER_484_1720 ();
 FILLCELL_X32 FILLER_484_1752 ();
 FILLCELL_X32 FILLER_484_1784 ();
 FILLCELL_X32 FILLER_484_1816 ();
 FILLCELL_X32 FILLER_484_1848 ();
 FILLCELL_X8 FILLER_484_1880 ();
 FILLCELL_X4 FILLER_484_1888 ();
 FILLCELL_X2 FILLER_484_1892 ();
 FILLCELL_X32 FILLER_484_1895 ();
 FILLCELL_X32 FILLER_484_1927 ();
 FILLCELL_X32 FILLER_484_1959 ();
 FILLCELL_X32 FILLER_484_1991 ();
 FILLCELL_X32 FILLER_484_2023 ();
 FILLCELL_X32 FILLER_484_2055 ();
 FILLCELL_X32 FILLER_484_2087 ();
 FILLCELL_X32 FILLER_484_2119 ();
 FILLCELL_X32 FILLER_484_2151 ();
 FILLCELL_X32 FILLER_484_2183 ();
 FILLCELL_X32 FILLER_484_2215 ();
 FILLCELL_X32 FILLER_484_2247 ();
 FILLCELL_X32 FILLER_484_2279 ();
 FILLCELL_X32 FILLER_484_2311 ();
 FILLCELL_X32 FILLER_484_2343 ();
 FILLCELL_X32 FILLER_484_2375 ();
 FILLCELL_X32 FILLER_484_2407 ();
 FILLCELL_X32 FILLER_484_2439 ();
 FILLCELL_X32 FILLER_484_2471 ();
 FILLCELL_X32 FILLER_484_2503 ();
 FILLCELL_X32 FILLER_484_2535 ();
 FILLCELL_X32 FILLER_484_2567 ();
 FILLCELL_X32 FILLER_484_2599 ();
 FILLCELL_X32 FILLER_484_2631 ();
 FILLCELL_X32 FILLER_484_2663 ();
 FILLCELL_X32 FILLER_484_2695 ();
 FILLCELL_X32 FILLER_484_2727 ();
 FILLCELL_X32 FILLER_484_2759 ();
 FILLCELL_X32 FILLER_484_2791 ();
 FILLCELL_X32 FILLER_484_2823 ();
 FILLCELL_X32 FILLER_484_2855 ();
 FILLCELL_X32 FILLER_484_2887 ();
 FILLCELL_X32 FILLER_484_2919 ();
 FILLCELL_X32 FILLER_484_2951 ();
 FILLCELL_X32 FILLER_484_2983 ();
 FILLCELL_X32 FILLER_484_3015 ();
 FILLCELL_X32 FILLER_484_3047 ();
 FILLCELL_X32 FILLER_484_3079 ();
 FILLCELL_X32 FILLER_484_3111 ();
 FILLCELL_X8 FILLER_484_3143 ();
 FILLCELL_X4 FILLER_484_3151 ();
 FILLCELL_X2 FILLER_484_3155 ();
 FILLCELL_X32 FILLER_484_3158 ();
 FILLCELL_X32 FILLER_484_3190 ();
 FILLCELL_X32 FILLER_484_3222 ();
 FILLCELL_X32 FILLER_484_3254 ();
 FILLCELL_X32 FILLER_484_3286 ();
 FILLCELL_X32 FILLER_484_3318 ();
 FILLCELL_X32 FILLER_484_3350 ();
 FILLCELL_X32 FILLER_484_3382 ();
 FILLCELL_X32 FILLER_484_3414 ();
 FILLCELL_X32 FILLER_484_3446 ();
 FILLCELL_X32 FILLER_484_3478 ();
 FILLCELL_X32 FILLER_484_3510 ();
 FILLCELL_X32 FILLER_484_3542 ();
 FILLCELL_X32 FILLER_484_3574 ();
 FILLCELL_X32 FILLER_484_3606 ();
 FILLCELL_X32 FILLER_484_3638 ();
 FILLCELL_X32 FILLER_484_3670 ();
 FILLCELL_X32 FILLER_484_3702 ();
 FILLCELL_X4 FILLER_484_3734 ();
 FILLCELL_X32 FILLER_485_1 ();
 FILLCELL_X32 FILLER_485_33 ();
 FILLCELL_X32 FILLER_485_65 ();
 FILLCELL_X32 FILLER_485_97 ();
 FILLCELL_X32 FILLER_485_129 ();
 FILLCELL_X32 FILLER_485_161 ();
 FILLCELL_X32 FILLER_485_193 ();
 FILLCELL_X32 FILLER_485_225 ();
 FILLCELL_X32 FILLER_485_257 ();
 FILLCELL_X32 FILLER_485_289 ();
 FILLCELL_X32 FILLER_485_321 ();
 FILLCELL_X32 FILLER_485_353 ();
 FILLCELL_X32 FILLER_485_385 ();
 FILLCELL_X32 FILLER_485_417 ();
 FILLCELL_X32 FILLER_485_449 ();
 FILLCELL_X32 FILLER_485_481 ();
 FILLCELL_X32 FILLER_485_513 ();
 FILLCELL_X32 FILLER_485_545 ();
 FILLCELL_X32 FILLER_485_577 ();
 FILLCELL_X32 FILLER_485_609 ();
 FILLCELL_X32 FILLER_485_641 ();
 FILLCELL_X32 FILLER_485_673 ();
 FILLCELL_X32 FILLER_485_705 ();
 FILLCELL_X32 FILLER_485_737 ();
 FILLCELL_X32 FILLER_485_769 ();
 FILLCELL_X32 FILLER_485_801 ();
 FILLCELL_X32 FILLER_485_833 ();
 FILLCELL_X32 FILLER_485_865 ();
 FILLCELL_X32 FILLER_485_897 ();
 FILLCELL_X32 FILLER_485_929 ();
 FILLCELL_X32 FILLER_485_961 ();
 FILLCELL_X32 FILLER_485_993 ();
 FILLCELL_X32 FILLER_485_1025 ();
 FILLCELL_X32 FILLER_485_1057 ();
 FILLCELL_X32 FILLER_485_1089 ();
 FILLCELL_X32 FILLER_485_1121 ();
 FILLCELL_X32 FILLER_485_1153 ();
 FILLCELL_X32 FILLER_485_1185 ();
 FILLCELL_X32 FILLER_485_1217 ();
 FILLCELL_X8 FILLER_485_1249 ();
 FILLCELL_X4 FILLER_485_1257 ();
 FILLCELL_X2 FILLER_485_1261 ();
 FILLCELL_X32 FILLER_485_1264 ();
 FILLCELL_X32 FILLER_485_1296 ();
 FILLCELL_X32 FILLER_485_1328 ();
 FILLCELL_X32 FILLER_485_1360 ();
 FILLCELL_X32 FILLER_485_1392 ();
 FILLCELL_X32 FILLER_485_1424 ();
 FILLCELL_X32 FILLER_485_1456 ();
 FILLCELL_X32 FILLER_485_1488 ();
 FILLCELL_X32 FILLER_485_1520 ();
 FILLCELL_X32 FILLER_485_1552 ();
 FILLCELL_X32 FILLER_485_1584 ();
 FILLCELL_X32 FILLER_485_1616 ();
 FILLCELL_X32 FILLER_485_1648 ();
 FILLCELL_X32 FILLER_485_1680 ();
 FILLCELL_X32 FILLER_485_1712 ();
 FILLCELL_X32 FILLER_485_1744 ();
 FILLCELL_X32 FILLER_485_1776 ();
 FILLCELL_X32 FILLER_485_1808 ();
 FILLCELL_X32 FILLER_485_1840 ();
 FILLCELL_X32 FILLER_485_1872 ();
 FILLCELL_X32 FILLER_485_1904 ();
 FILLCELL_X32 FILLER_485_1936 ();
 FILLCELL_X32 FILLER_485_1968 ();
 FILLCELL_X32 FILLER_485_2000 ();
 FILLCELL_X32 FILLER_485_2032 ();
 FILLCELL_X32 FILLER_485_2064 ();
 FILLCELL_X32 FILLER_485_2096 ();
 FILLCELL_X32 FILLER_485_2128 ();
 FILLCELL_X32 FILLER_485_2160 ();
 FILLCELL_X32 FILLER_485_2192 ();
 FILLCELL_X32 FILLER_485_2224 ();
 FILLCELL_X32 FILLER_485_2256 ();
 FILLCELL_X32 FILLER_485_2288 ();
 FILLCELL_X32 FILLER_485_2320 ();
 FILLCELL_X32 FILLER_485_2352 ();
 FILLCELL_X32 FILLER_485_2384 ();
 FILLCELL_X32 FILLER_485_2416 ();
 FILLCELL_X32 FILLER_485_2448 ();
 FILLCELL_X32 FILLER_485_2480 ();
 FILLCELL_X8 FILLER_485_2512 ();
 FILLCELL_X4 FILLER_485_2520 ();
 FILLCELL_X2 FILLER_485_2524 ();
 FILLCELL_X32 FILLER_485_2527 ();
 FILLCELL_X32 FILLER_485_2559 ();
 FILLCELL_X32 FILLER_485_2591 ();
 FILLCELL_X32 FILLER_485_2623 ();
 FILLCELL_X32 FILLER_485_2655 ();
 FILLCELL_X32 FILLER_485_2687 ();
 FILLCELL_X32 FILLER_485_2719 ();
 FILLCELL_X32 FILLER_485_2751 ();
 FILLCELL_X32 FILLER_485_2783 ();
 FILLCELL_X32 FILLER_485_2815 ();
 FILLCELL_X32 FILLER_485_2847 ();
 FILLCELL_X32 FILLER_485_2879 ();
 FILLCELL_X32 FILLER_485_2911 ();
 FILLCELL_X32 FILLER_485_2943 ();
 FILLCELL_X32 FILLER_485_2975 ();
 FILLCELL_X32 FILLER_485_3007 ();
 FILLCELL_X32 FILLER_485_3039 ();
 FILLCELL_X32 FILLER_485_3071 ();
 FILLCELL_X32 FILLER_485_3103 ();
 FILLCELL_X32 FILLER_485_3135 ();
 FILLCELL_X32 FILLER_485_3167 ();
 FILLCELL_X32 FILLER_485_3199 ();
 FILLCELL_X32 FILLER_485_3231 ();
 FILLCELL_X32 FILLER_485_3263 ();
 FILLCELL_X32 FILLER_485_3295 ();
 FILLCELL_X32 FILLER_485_3327 ();
 FILLCELL_X32 FILLER_485_3359 ();
 FILLCELL_X32 FILLER_485_3391 ();
 FILLCELL_X32 FILLER_485_3423 ();
 FILLCELL_X32 FILLER_485_3455 ();
 FILLCELL_X32 FILLER_485_3487 ();
 FILLCELL_X32 FILLER_485_3519 ();
 FILLCELL_X32 FILLER_485_3551 ();
 FILLCELL_X32 FILLER_485_3583 ();
 FILLCELL_X32 FILLER_485_3615 ();
 FILLCELL_X32 FILLER_485_3647 ();
 FILLCELL_X32 FILLER_485_3679 ();
 FILLCELL_X16 FILLER_485_3711 ();
 FILLCELL_X8 FILLER_485_3727 ();
 FILLCELL_X2 FILLER_485_3735 ();
 FILLCELL_X1 FILLER_485_3737 ();
 FILLCELL_X32 FILLER_486_1 ();
 FILLCELL_X32 FILLER_486_33 ();
 FILLCELL_X32 FILLER_486_65 ();
 FILLCELL_X32 FILLER_486_97 ();
 FILLCELL_X32 FILLER_486_129 ();
 FILLCELL_X32 FILLER_486_161 ();
 FILLCELL_X32 FILLER_486_193 ();
 FILLCELL_X32 FILLER_486_225 ();
 FILLCELL_X32 FILLER_486_257 ();
 FILLCELL_X32 FILLER_486_289 ();
 FILLCELL_X32 FILLER_486_321 ();
 FILLCELL_X32 FILLER_486_353 ();
 FILLCELL_X32 FILLER_486_385 ();
 FILLCELL_X32 FILLER_486_417 ();
 FILLCELL_X32 FILLER_486_449 ();
 FILLCELL_X32 FILLER_486_481 ();
 FILLCELL_X32 FILLER_486_513 ();
 FILLCELL_X32 FILLER_486_545 ();
 FILLCELL_X32 FILLER_486_577 ();
 FILLCELL_X16 FILLER_486_609 ();
 FILLCELL_X4 FILLER_486_625 ();
 FILLCELL_X2 FILLER_486_629 ();
 FILLCELL_X32 FILLER_486_632 ();
 FILLCELL_X32 FILLER_486_664 ();
 FILLCELL_X32 FILLER_486_696 ();
 FILLCELL_X32 FILLER_486_728 ();
 FILLCELL_X32 FILLER_486_760 ();
 FILLCELL_X32 FILLER_486_792 ();
 FILLCELL_X32 FILLER_486_824 ();
 FILLCELL_X32 FILLER_486_856 ();
 FILLCELL_X32 FILLER_486_888 ();
 FILLCELL_X32 FILLER_486_920 ();
 FILLCELL_X32 FILLER_486_952 ();
 FILLCELL_X32 FILLER_486_984 ();
 FILLCELL_X32 FILLER_486_1016 ();
 FILLCELL_X32 FILLER_486_1048 ();
 FILLCELL_X32 FILLER_486_1080 ();
 FILLCELL_X32 FILLER_486_1112 ();
 FILLCELL_X32 FILLER_486_1144 ();
 FILLCELL_X32 FILLER_486_1176 ();
 FILLCELL_X32 FILLER_486_1208 ();
 FILLCELL_X32 FILLER_486_1240 ();
 FILLCELL_X32 FILLER_486_1272 ();
 FILLCELL_X32 FILLER_486_1304 ();
 FILLCELL_X32 FILLER_486_1336 ();
 FILLCELL_X32 FILLER_486_1368 ();
 FILLCELL_X32 FILLER_486_1400 ();
 FILLCELL_X32 FILLER_486_1432 ();
 FILLCELL_X32 FILLER_486_1464 ();
 FILLCELL_X32 FILLER_486_1496 ();
 FILLCELL_X32 FILLER_486_1528 ();
 FILLCELL_X32 FILLER_486_1560 ();
 FILLCELL_X32 FILLER_486_1592 ();
 FILLCELL_X32 FILLER_486_1624 ();
 FILLCELL_X32 FILLER_486_1656 ();
 FILLCELL_X32 FILLER_486_1688 ();
 FILLCELL_X32 FILLER_486_1720 ();
 FILLCELL_X32 FILLER_486_1752 ();
 FILLCELL_X32 FILLER_486_1784 ();
 FILLCELL_X32 FILLER_486_1816 ();
 FILLCELL_X32 FILLER_486_1848 ();
 FILLCELL_X8 FILLER_486_1880 ();
 FILLCELL_X4 FILLER_486_1888 ();
 FILLCELL_X2 FILLER_486_1892 ();
 FILLCELL_X32 FILLER_486_1895 ();
 FILLCELL_X32 FILLER_486_1927 ();
 FILLCELL_X32 FILLER_486_1959 ();
 FILLCELL_X32 FILLER_486_1991 ();
 FILLCELL_X32 FILLER_486_2023 ();
 FILLCELL_X32 FILLER_486_2055 ();
 FILLCELL_X32 FILLER_486_2087 ();
 FILLCELL_X32 FILLER_486_2119 ();
 FILLCELL_X32 FILLER_486_2151 ();
 FILLCELL_X32 FILLER_486_2183 ();
 FILLCELL_X32 FILLER_486_2215 ();
 FILLCELL_X32 FILLER_486_2247 ();
 FILLCELL_X32 FILLER_486_2279 ();
 FILLCELL_X32 FILLER_486_2311 ();
 FILLCELL_X32 FILLER_486_2343 ();
 FILLCELL_X32 FILLER_486_2375 ();
 FILLCELL_X32 FILLER_486_2407 ();
 FILLCELL_X32 FILLER_486_2439 ();
 FILLCELL_X32 FILLER_486_2471 ();
 FILLCELL_X32 FILLER_486_2503 ();
 FILLCELL_X32 FILLER_486_2535 ();
 FILLCELL_X32 FILLER_486_2567 ();
 FILLCELL_X32 FILLER_486_2599 ();
 FILLCELL_X32 FILLER_486_2631 ();
 FILLCELL_X32 FILLER_486_2663 ();
 FILLCELL_X32 FILLER_486_2695 ();
 FILLCELL_X32 FILLER_486_2727 ();
 FILLCELL_X32 FILLER_486_2759 ();
 FILLCELL_X32 FILLER_486_2791 ();
 FILLCELL_X32 FILLER_486_2823 ();
 FILLCELL_X32 FILLER_486_2855 ();
 FILLCELL_X32 FILLER_486_2887 ();
 FILLCELL_X32 FILLER_486_2919 ();
 FILLCELL_X32 FILLER_486_2951 ();
 FILLCELL_X32 FILLER_486_2983 ();
 FILLCELL_X32 FILLER_486_3015 ();
 FILLCELL_X32 FILLER_486_3047 ();
 FILLCELL_X32 FILLER_486_3079 ();
 FILLCELL_X32 FILLER_486_3111 ();
 FILLCELL_X8 FILLER_486_3143 ();
 FILLCELL_X4 FILLER_486_3151 ();
 FILLCELL_X2 FILLER_486_3155 ();
 FILLCELL_X32 FILLER_486_3158 ();
 FILLCELL_X32 FILLER_486_3190 ();
 FILLCELL_X32 FILLER_486_3222 ();
 FILLCELL_X32 FILLER_486_3254 ();
 FILLCELL_X32 FILLER_486_3286 ();
 FILLCELL_X32 FILLER_486_3318 ();
 FILLCELL_X32 FILLER_486_3350 ();
 FILLCELL_X32 FILLER_486_3382 ();
 FILLCELL_X32 FILLER_486_3414 ();
 FILLCELL_X32 FILLER_486_3446 ();
 FILLCELL_X32 FILLER_486_3478 ();
 FILLCELL_X32 FILLER_486_3510 ();
 FILLCELL_X32 FILLER_486_3542 ();
 FILLCELL_X32 FILLER_486_3574 ();
 FILLCELL_X32 FILLER_486_3606 ();
 FILLCELL_X32 FILLER_486_3638 ();
 FILLCELL_X32 FILLER_486_3670 ();
 FILLCELL_X32 FILLER_486_3702 ();
 FILLCELL_X4 FILLER_486_3734 ();
 FILLCELL_X32 FILLER_487_1 ();
 FILLCELL_X32 FILLER_487_33 ();
 FILLCELL_X32 FILLER_487_65 ();
 FILLCELL_X32 FILLER_487_97 ();
 FILLCELL_X32 FILLER_487_129 ();
 FILLCELL_X32 FILLER_487_161 ();
 FILLCELL_X32 FILLER_487_193 ();
 FILLCELL_X32 FILLER_487_225 ();
 FILLCELL_X32 FILLER_487_257 ();
 FILLCELL_X32 FILLER_487_289 ();
 FILLCELL_X32 FILLER_487_321 ();
 FILLCELL_X32 FILLER_487_353 ();
 FILLCELL_X32 FILLER_487_385 ();
 FILLCELL_X32 FILLER_487_417 ();
 FILLCELL_X32 FILLER_487_449 ();
 FILLCELL_X32 FILLER_487_481 ();
 FILLCELL_X32 FILLER_487_513 ();
 FILLCELL_X32 FILLER_487_545 ();
 FILLCELL_X32 FILLER_487_577 ();
 FILLCELL_X32 FILLER_487_609 ();
 FILLCELL_X32 FILLER_487_641 ();
 FILLCELL_X32 FILLER_487_673 ();
 FILLCELL_X32 FILLER_487_705 ();
 FILLCELL_X32 FILLER_487_737 ();
 FILLCELL_X32 FILLER_487_769 ();
 FILLCELL_X32 FILLER_487_801 ();
 FILLCELL_X32 FILLER_487_833 ();
 FILLCELL_X32 FILLER_487_865 ();
 FILLCELL_X32 FILLER_487_897 ();
 FILLCELL_X32 FILLER_487_929 ();
 FILLCELL_X32 FILLER_487_961 ();
 FILLCELL_X32 FILLER_487_993 ();
 FILLCELL_X32 FILLER_487_1025 ();
 FILLCELL_X32 FILLER_487_1057 ();
 FILLCELL_X32 FILLER_487_1089 ();
 FILLCELL_X32 FILLER_487_1121 ();
 FILLCELL_X32 FILLER_487_1153 ();
 FILLCELL_X32 FILLER_487_1185 ();
 FILLCELL_X32 FILLER_487_1217 ();
 FILLCELL_X8 FILLER_487_1249 ();
 FILLCELL_X4 FILLER_487_1257 ();
 FILLCELL_X2 FILLER_487_1261 ();
 FILLCELL_X32 FILLER_487_1264 ();
 FILLCELL_X32 FILLER_487_1296 ();
 FILLCELL_X32 FILLER_487_1328 ();
 FILLCELL_X32 FILLER_487_1360 ();
 FILLCELL_X32 FILLER_487_1392 ();
 FILLCELL_X32 FILLER_487_1424 ();
 FILLCELL_X32 FILLER_487_1456 ();
 FILLCELL_X32 FILLER_487_1488 ();
 FILLCELL_X32 FILLER_487_1520 ();
 FILLCELL_X32 FILLER_487_1552 ();
 FILLCELL_X32 FILLER_487_1584 ();
 FILLCELL_X32 FILLER_487_1616 ();
 FILLCELL_X32 FILLER_487_1648 ();
 FILLCELL_X32 FILLER_487_1680 ();
 FILLCELL_X32 FILLER_487_1712 ();
 FILLCELL_X32 FILLER_487_1744 ();
 FILLCELL_X32 FILLER_487_1776 ();
 FILLCELL_X32 FILLER_487_1808 ();
 FILLCELL_X32 FILLER_487_1840 ();
 FILLCELL_X32 FILLER_487_1872 ();
 FILLCELL_X32 FILLER_487_1904 ();
 FILLCELL_X32 FILLER_487_1936 ();
 FILLCELL_X32 FILLER_487_1968 ();
 FILLCELL_X32 FILLER_487_2000 ();
 FILLCELL_X32 FILLER_487_2032 ();
 FILLCELL_X32 FILLER_487_2064 ();
 FILLCELL_X32 FILLER_487_2096 ();
 FILLCELL_X32 FILLER_487_2128 ();
 FILLCELL_X32 FILLER_487_2160 ();
 FILLCELL_X32 FILLER_487_2192 ();
 FILLCELL_X32 FILLER_487_2224 ();
 FILLCELL_X32 FILLER_487_2256 ();
 FILLCELL_X32 FILLER_487_2288 ();
 FILLCELL_X32 FILLER_487_2320 ();
 FILLCELL_X32 FILLER_487_2352 ();
 FILLCELL_X32 FILLER_487_2384 ();
 FILLCELL_X32 FILLER_487_2416 ();
 FILLCELL_X32 FILLER_487_2448 ();
 FILLCELL_X32 FILLER_487_2480 ();
 FILLCELL_X8 FILLER_487_2512 ();
 FILLCELL_X4 FILLER_487_2520 ();
 FILLCELL_X2 FILLER_487_2524 ();
 FILLCELL_X32 FILLER_487_2527 ();
 FILLCELL_X32 FILLER_487_2559 ();
 FILLCELL_X32 FILLER_487_2591 ();
 FILLCELL_X32 FILLER_487_2623 ();
 FILLCELL_X32 FILLER_487_2655 ();
 FILLCELL_X32 FILLER_487_2687 ();
 FILLCELL_X32 FILLER_487_2719 ();
 FILLCELL_X32 FILLER_487_2751 ();
 FILLCELL_X32 FILLER_487_2783 ();
 FILLCELL_X32 FILLER_487_2815 ();
 FILLCELL_X32 FILLER_487_2847 ();
 FILLCELL_X32 FILLER_487_2879 ();
 FILLCELL_X32 FILLER_487_2911 ();
 FILLCELL_X32 FILLER_487_2943 ();
 FILLCELL_X32 FILLER_487_2975 ();
 FILLCELL_X32 FILLER_487_3007 ();
 FILLCELL_X32 FILLER_487_3039 ();
 FILLCELL_X32 FILLER_487_3071 ();
 FILLCELL_X32 FILLER_487_3103 ();
 FILLCELL_X32 FILLER_487_3135 ();
 FILLCELL_X32 FILLER_487_3167 ();
 FILLCELL_X32 FILLER_487_3199 ();
 FILLCELL_X32 FILLER_487_3231 ();
 FILLCELL_X32 FILLER_487_3263 ();
 FILLCELL_X32 FILLER_487_3295 ();
 FILLCELL_X32 FILLER_487_3327 ();
 FILLCELL_X32 FILLER_487_3359 ();
 FILLCELL_X32 FILLER_487_3391 ();
 FILLCELL_X32 FILLER_487_3423 ();
 FILLCELL_X32 FILLER_487_3455 ();
 FILLCELL_X32 FILLER_487_3487 ();
 FILLCELL_X32 FILLER_487_3519 ();
 FILLCELL_X32 FILLER_487_3551 ();
 FILLCELL_X32 FILLER_487_3583 ();
 FILLCELL_X32 FILLER_487_3615 ();
 FILLCELL_X32 FILLER_487_3647 ();
 FILLCELL_X32 FILLER_487_3679 ();
 FILLCELL_X16 FILLER_487_3711 ();
 FILLCELL_X8 FILLER_487_3727 ();
 FILLCELL_X2 FILLER_487_3735 ();
 FILLCELL_X1 FILLER_487_3737 ();
 FILLCELL_X32 FILLER_488_1 ();
 FILLCELL_X32 FILLER_488_33 ();
 FILLCELL_X32 FILLER_488_65 ();
 FILLCELL_X32 FILLER_488_97 ();
 FILLCELL_X32 FILLER_488_129 ();
 FILLCELL_X32 FILLER_488_161 ();
 FILLCELL_X32 FILLER_488_193 ();
 FILLCELL_X32 FILLER_488_225 ();
 FILLCELL_X32 FILLER_488_257 ();
 FILLCELL_X32 FILLER_488_289 ();
 FILLCELL_X32 FILLER_488_321 ();
 FILLCELL_X32 FILLER_488_353 ();
 FILLCELL_X32 FILLER_488_385 ();
 FILLCELL_X32 FILLER_488_417 ();
 FILLCELL_X32 FILLER_488_449 ();
 FILLCELL_X32 FILLER_488_481 ();
 FILLCELL_X32 FILLER_488_513 ();
 FILLCELL_X32 FILLER_488_545 ();
 FILLCELL_X32 FILLER_488_577 ();
 FILLCELL_X16 FILLER_488_609 ();
 FILLCELL_X4 FILLER_488_625 ();
 FILLCELL_X2 FILLER_488_629 ();
 FILLCELL_X32 FILLER_488_632 ();
 FILLCELL_X32 FILLER_488_664 ();
 FILLCELL_X32 FILLER_488_696 ();
 FILLCELL_X32 FILLER_488_728 ();
 FILLCELL_X32 FILLER_488_760 ();
 FILLCELL_X32 FILLER_488_792 ();
 FILLCELL_X32 FILLER_488_824 ();
 FILLCELL_X32 FILLER_488_856 ();
 FILLCELL_X32 FILLER_488_888 ();
 FILLCELL_X32 FILLER_488_920 ();
 FILLCELL_X32 FILLER_488_952 ();
 FILLCELL_X32 FILLER_488_984 ();
 FILLCELL_X32 FILLER_488_1016 ();
 FILLCELL_X32 FILLER_488_1048 ();
 FILLCELL_X32 FILLER_488_1080 ();
 FILLCELL_X32 FILLER_488_1112 ();
 FILLCELL_X32 FILLER_488_1144 ();
 FILLCELL_X32 FILLER_488_1176 ();
 FILLCELL_X32 FILLER_488_1208 ();
 FILLCELL_X32 FILLER_488_1240 ();
 FILLCELL_X32 FILLER_488_1272 ();
 FILLCELL_X32 FILLER_488_1304 ();
 FILLCELL_X32 FILLER_488_1336 ();
 FILLCELL_X32 FILLER_488_1368 ();
 FILLCELL_X32 FILLER_488_1400 ();
 FILLCELL_X32 FILLER_488_1432 ();
 FILLCELL_X32 FILLER_488_1464 ();
 FILLCELL_X32 FILLER_488_1496 ();
 FILLCELL_X32 FILLER_488_1528 ();
 FILLCELL_X32 FILLER_488_1560 ();
 FILLCELL_X32 FILLER_488_1592 ();
 FILLCELL_X32 FILLER_488_1624 ();
 FILLCELL_X32 FILLER_488_1656 ();
 FILLCELL_X32 FILLER_488_1688 ();
 FILLCELL_X32 FILLER_488_1720 ();
 FILLCELL_X32 FILLER_488_1752 ();
 FILLCELL_X32 FILLER_488_1784 ();
 FILLCELL_X32 FILLER_488_1816 ();
 FILLCELL_X32 FILLER_488_1848 ();
 FILLCELL_X8 FILLER_488_1880 ();
 FILLCELL_X4 FILLER_488_1888 ();
 FILLCELL_X2 FILLER_488_1892 ();
 FILLCELL_X32 FILLER_488_1895 ();
 FILLCELL_X32 FILLER_488_1927 ();
 FILLCELL_X32 FILLER_488_1959 ();
 FILLCELL_X32 FILLER_488_1991 ();
 FILLCELL_X32 FILLER_488_2023 ();
 FILLCELL_X32 FILLER_488_2055 ();
 FILLCELL_X32 FILLER_488_2087 ();
 FILLCELL_X32 FILLER_488_2119 ();
 FILLCELL_X32 FILLER_488_2151 ();
 FILLCELL_X32 FILLER_488_2183 ();
 FILLCELL_X32 FILLER_488_2215 ();
 FILLCELL_X32 FILLER_488_2247 ();
 FILLCELL_X32 FILLER_488_2279 ();
 FILLCELL_X32 FILLER_488_2311 ();
 FILLCELL_X32 FILLER_488_2343 ();
 FILLCELL_X32 FILLER_488_2375 ();
 FILLCELL_X32 FILLER_488_2407 ();
 FILLCELL_X32 FILLER_488_2439 ();
 FILLCELL_X32 FILLER_488_2471 ();
 FILLCELL_X32 FILLER_488_2503 ();
 FILLCELL_X32 FILLER_488_2535 ();
 FILLCELL_X32 FILLER_488_2567 ();
 FILLCELL_X32 FILLER_488_2599 ();
 FILLCELL_X32 FILLER_488_2631 ();
 FILLCELL_X32 FILLER_488_2663 ();
 FILLCELL_X32 FILLER_488_2695 ();
 FILLCELL_X32 FILLER_488_2727 ();
 FILLCELL_X32 FILLER_488_2759 ();
 FILLCELL_X32 FILLER_488_2791 ();
 FILLCELL_X32 FILLER_488_2823 ();
 FILLCELL_X32 FILLER_488_2855 ();
 FILLCELL_X32 FILLER_488_2887 ();
 FILLCELL_X32 FILLER_488_2919 ();
 FILLCELL_X32 FILLER_488_2951 ();
 FILLCELL_X32 FILLER_488_2983 ();
 FILLCELL_X32 FILLER_488_3015 ();
 FILLCELL_X32 FILLER_488_3047 ();
 FILLCELL_X32 FILLER_488_3079 ();
 FILLCELL_X32 FILLER_488_3111 ();
 FILLCELL_X8 FILLER_488_3143 ();
 FILLCELL_X4 FILLER_488_3151 ();
 FILLCELL_X2 FILLER_488_3155 ();
 FILLCELL_X32 FILLER_488_3158 ();
 FILLCELL_X32 FILLER_488_3190 ();
 FILLCELL_X32 FILLER_488_3222 ();
 FILLCELL_X32 FILLER_488_3254 ();
 FILLCELL_X32 FILLER_488_3286 ();
 FILLCELL_X32 FILLER_488_3318 ();
 FILLCELL_X32 FILLER_488_3350 ();
 FILLCELL_X32 FILLER_488_3382 ();
 FILLCELL_X32 FILLER_488_3414 ();
 FILLCELL_X32 FILLER_488_3446 ();
 FILLCELL_X32 FILLER_488_3478 ();
 FILLCELL_X32 FILLER_488_3510 ();
 FILLCELL_X32 FILLER_488_3542 ();
 FILLCELL_X32 FILLER_488_3574 ();
 FILLCELL_X32 FILLER_488_3606 ();
 FILLCELL_X32 FILLER_488_3638 ();
 FILLCELL_X32 FILLER_488_3670 ();
 FILLCELL_X32 FILLER_488_3702 ();
 FILLCELL_X4 FILLER_488_3734 ();
 FILLCELL_X32 FILLER_489_1 ();
 FILLCELL_X32 FILLER_489_33 ();
 FILLCELL_X32 FILLER_489_65 ();
 FILLCELL_X32 FILLER_489_97 ();
 FILLCELL_X32 FILLER_489_129 ();
 FILLCELL_X32 FILLER_489_161 ();
 FILLCELL_X32 FILLER_489_193 ();
 FILLCELL_X32 FILLER_489_225 ();
 FILLCELL_X32 FILLER_489_257 ();
 FILLCELL_X32 FILLER_489_289 ();
 FILLCELL_X32 FILLER_489_321 ();
 FILLCELL_X32 FILLER_489_353 ();
 FILLCELL_X32 FILLER_489_385 ();
 FILLCELL_X32 FILLER_489_417 ();
 FILLCELL_X32 FILLER_489_449 ();
 FILLCELL_X32 FILLER_489_481 ();
 FILLCELL_X32 FILLER_489_513 ();
 FILLCELL_X32 FILLER_489_545 ();
 FILLCELL_X32 FILLER_489_577 ();
 FILLCELL_X32 FILLER_489_609 ();
 FILLCELL_X32 FILLER_489_641 ();
 FILLCELL_X32 FILLER_489_673 ();
 FILLCELL_X32 FILLER_489_705 ();
 FILLCELL_X32 FILLER_489_737 ();
 FILLCELL_X32 FILLER_489_769 ();
 FILLCELL_X32 FILLER_489_801 ();
 FILLCELL_X32 FILLER_489_833 ();
 FILLCELL_X32 FILLER_489_865 ();
 FILLCELL_X32 FILLER_489_897 ();
 FILLCELL_X32 FILLER_489_929 ();
 FILLCELL_X32 FILLER_489_961 ();
 FILLCELL_X32 FILLER_489_993 ();
 FILLCELL_X32 FILLER_489_1025 ();
 FILLCELL_X32 FILLER_489_1057 ();
 FILLCELL_X32 FILLER_489_1089 ();
 FILLCELL_X32 FILLER_489_1121 ();
 FILLCELL_X32 FILLER_489_1153 ();
 FILLCELL_X32 FILLER_489_1185 ();
 FILLCELL_X32 FILLER_489_1217 ();
 FILLCELL_X8 FILLER_489_1249 ();
 FILLCELL_X4 FILLER_489_1257 ();
 FILLCELL_X2 FILLER_489_1261 ();
 FILLCELL_X32 FILLER_489_1264 ();
 FILLCELL_X32 FILLER_489_1296 ();
 FILLCELL_X32 FILLER_489_1328 ();
 FILLCELL_X32 FILLER_489_1360 ();
 FILLCELL_X32 FILLER_489_1392 ();
 FILLCELL_X32 FILLER_489_1424 ();
 FILLCELL_X32 FILLER_489_1456 ();
 FILLCELL_X32 FILLER_489_1488 ();
 FILLCELL_X32 FILLER_489_1520 ();
 FILLCELL_X32 FILLER_489_1552 ();
 FILLCELL_X32 FILLER_489_1584 ();
 FILLCELL_X32 FILLER_489_1616 ();
 FILLCELL_X32 FILLER_489_1648 ();
 FILLCELL_X32 FILLER_489_1680 ();
 FILLCELL_X32 FILLER_489_1712 ();
 FILLCELL_X32 FILLER_489_1744 ();
 FILLCELL_X32 FILLER_489_1776 ();
 FILLCELL_X32 FILLER_489_1808 ();
 FILLCELL_X32 FILLER_489_1840 ();
 FILLCELL_X32 FILLER_489_1872 ();
 FILLCELL_X32 FILLER_489_1904 ();
 FILLCELL_X32 FILLER_489_1936 ();
 FILLCELL_X32 FILLER_489_1968 ();
 FILLCELL_X32 FILLER_489_2000 ();
 FILLCELL_X32 FILLER_489_2032 ();
 FILLCELL_X32 FILLER_489_2064 ();
 FILLCELL_X32 FILLER_489_2096 ();
 FILLCELL_X32 FILLER_489_2128 ();
 FILLCELL_X32 FILLER_489_2160 ();
 FILLCELL_X32 FILLER_489_2192 ();
 FILLCELL_X32 FILLER_489_2224 ();
 FILLCELL_X32 FILLER_489_2256 ();
 FILLCELL_X32 FILLER_489_2288 ();
 FILLCELL_X32 FILLER_489_2320 ();
 FILLCELL_X32 FILLER_489_2352 ();
 FILLCELL_X32 FILLER_489_2384 ();
 FILLCELL_X32 FILLER_489_2416 ();
 FILLCELL_X32 FILLER_489_2448 ();
 FILLCELL_X32 FILLER_489_2480 ();
 FILLCELL_X8 FILLER_489_2512 ();
 FILLCELL_X4 FILLER_489_2520 ();
 FILLCELL_X2 FILLER_489_2524 ();
 FILLCELL_X32 FILLER_489_2527 ();
 FILLCELL_X32 FILLER_489_2559 ();
 FILLCELL_X32 FILLER_489_2591 ();
 FILLCELL_X32 FILLER_489_2623 ();
 FILLCELL_X32 FILLER_489_2655 ();
 FILLCELL_X32 FILLER_489_2687 ();
 FILLCELL_X32 FILLER_489_2719 ();
 FILLCELL_X32 FILLER_489_2751 ();
 FILLCELL_X32 FILLER_489_2783 ();
 FILLCELL_X32 FILLER_489_2815 ();
 FILLCELL_X32 FILLER_489_2847 ();
 FILLCELL_X32 FILLER_489_2879 ();
 FILLCELL_X32 FILLER_489_2911 ();
 FILLCELL_X32 FILLER_489_2943 ();
 FILLCELL_X32 FILLER_489_2975 ();
 FILLCELL_X32 FILLER_489_3007 ();
 FILLCELL_X32 FILLER_489_3039 ();
 FILLCELL_X32 FILLER_489_3071 ();
 FILLCELL_X32 FILLER_489_3103 ();
 FILLCELL_X32 FILLER_489_3135 ();
 FILLCELL_X32 FILLER_489_3167 ();
 FILLCELL_X32 FILLER_489_3199 ();
 FILLCELL_X32 FILLER_489_3231 ();
 FILLCELL_X32 FILLER_489_3263 ();
 FILLCELL_X32 FILLER_489_3295 ();
 FILLCELL_X32 FILLER_489_3327 ();
 FILLCELL_X32 FILLER_489_3359 ();
 FILLCELL_X32 FILLER_489_3391 ();
 FILLCELL_X32 FILLER_489_3423 ();
 FILLCELL_X32 FILLER_489_3455 ();
 FILLCELL_X32 FILLER_489_3487 ();
 FILLCELL_X32 FILLER_489_3519 ();
 FILLCELL_X32 FILLER_489_3551 ();
 FILLCELL_X32 FILLER_489_3583 ();
 FILLCELL_X32 FILLER_489_3615 ();
 FILLCELL_X32 FILLER_489_3647 ();
 FILLCELL_X32 FILLER_489_3679 ();
 FILLCELL_X16 FILLER_489_3711 ();
 FILLCELL_X8 FILLER_489_3727 ();
 FILLCELL_X2 FILLER_489_3735 ();
 FILLCELL_X1 FILLER_489_3737 ();
 FILLCELL_X32 FILLER_490_1 ();
 FILLCELL_X32 FILLER_490_33 ();
 FILLCELL_X32 FILLER_490_65 ();
 FILLCELL_X32 FILLER_490_97 ();
 FILLCELL_X32 FILLER_490_129 ();
 FILLCELL_X32 FILLER_490_161 ();
 FILLCELL_X32 FILLER_490_193 ();
 FILLCELL_X32 FILLER_490_225 ();
 FILLCELL_X32 FILLER_490_257 ();
 FILLCELL_X32 FILLER_490_289 ();
 FILLCELL_X32 FILLER_490_321 ();
 FILLCELL_X32 FILLER_490_353 ();
 FILLCELL_X32 FILLER_490_385 ();
 FILLCELL_X32 FILLER_490_417 ();
 FILLCELL_X32 FILLER_490_449 ();
 FILLCELL_X32 FILLER_490_481 ();
 FILLCELL_X32 FILLER_490_513 ();
 FILLCELL_X32 FILLER_490_545 ();
 FILLCELL_X32 FILLER_490_577 ();
 FILLCELL_X16 FILLER_490_609 ();
 FILLCELL_X4 FILLER_490_625 ();
 FILLCELL_X2 FILLER_490_629 ();
 FILLCELL_X32 FILLER_490_632 ();
 FILLCELL_X32 FILLER_490_664 ();
 FILLCELL_X32 FILLER_490_696 ();
 FILLCELL_X32 FILLER_490_728 ();
 FILLCELL_X32 FILLER_490_760 ();
 FILLCELL_X32 FILLER_490_792 ();
 FILLCELL_X32 FILLER_490_824 ();
 FILLCELL_X32 FILLER_490_856 ();
 FILLCELL_X32 FILLER_490_888 ();
 FILLCELL_X32 FILLER_490_920 ();
 FILLCELL_X32 FILLER_490_952 ();
 FILLCELL_X32 FILLER_490_984 ();
 FILLCELL_X32 FILLER_490_1016 ();
 FILLCELL_X32 FILLER_490_1048 ();
 FILLCELL_X32 FILLER_490_1080 ();
 FILLCELL_X32 FILLER_490_1112 ();
 FILLCELL_X32 FILLER_490_1144 ();
 FILLCELL_X32 FILLER_490_1176 ();
 FILLCELL_X32 FILLER_490_1208 ();
 FILLCELL_X32 FILLER_490_1240 ();
 FILLCELL_X32 FILLER_490_1272 ();
 FILLCELL_X32 FILLER_490_1304 ();
 FILLCELL_X32 FILLER_490_1336 ();
 FILLCELL_X32 FILLER_490_1368 ();
 FILLCELL_X32 FILLER_490_1400 ();
 FILLCELL_X32 FILLER_490_1432 ();
 FILLCELL_X32 FILLER_490_1464 ();
 FILLCELL_X32 FILLER_490_1496 ();
 FILLCELL_X32 FILLER_490_1528 ();
 FILLCELL_X32 FILLER_490_1560 ();
 FILLCELL_X32 FILLER_490_1592 ();
 FILLCELL_X32 FILLER_490_1624 ();
 FILLCELL_X32 FILLER_490_1656 ();
 FILLCELL_X32 FILLER_490_1688 ();
 FILLCELL_X32 FILLER_490_1720 ();
 FILLCELL_X32 FILLER_490_1752 ();
 FILLCELL_X32 FILLER_490_1784 ();
 FILLCELL_X32 FILLER_490_1816 ();
 FILLCELL_X32 FILLER_490_1848 ();
 FILLCELL_X8 FILLER_490_1880 ();
 FILLCELL_X4 FILLER_490_1888 ();
 FILLCELL_X2 FILLER_490_1892 ();
 FILLCELL_X32 FILLER_490_1895 ();
 FILLCELL_X32 FILLER_490_1927 ();
 FILLCELL_X32 FILLER_490_1959 ();
 FILLCELL_X32 FILLER_490_1991 ();
 FILLCELL_X32 FILLER_490_2023 ();
 FILLCELL_X32 FILLER_490_2055 ();
 FILLCELL_X32 FILLER_490_2087 ();
 FILLCELL_X32 FILLER_490_2119 ();
 FILLCELL_X32 FILLER_490_2151 ();
 FILLCELL_X32 FILLER_490_2183 ();
 FILLCELL_X32 FILLER_490_2215 ();
 FILLCELL_X32 FILLER_490_2247 ();
 FILLCELL_X32 FILLER_490_2279 ();
 FILLCELL_X32 FILLER_490_2311 ();
 FILLCELL_X32 FILLER_490_2343 ();
 FILLCELL_X32 FILLER_490_2375 ();
 FILLCELL_X32 FILLER_490_2407 ();
 FILLCELL_X32 FILLER_490_2439 ();
 FILLCELL_X32 FILLER_490_2471 ();
 FILLCELL_X32 FILLER_490_2503 ();
 FILLCELL_X32 FILLER_490_2535 ();
 FILLCELL_X32 FILLER_490_2567 ();
 FILLCELL_X32 FILLER_490_2599 ();
 FILLCELL_X32 FILLER_490_2631 ();
 FILLCELL_X32 FILLER_490_2663 ();
 FILLCELL_X32 FILLER_490_2695 ();
 FILLCELL_X32 FILLER_490_2727 ();
 FILLCELL_X32 FILLER_490_2759 ();
 FILLCELL_X32 FILLER_490_2791 ();
 FILLCELL_X32 FILLER_490_2823 ();
 FILLCELL_X32 FILLER_490_2855 ();
 FILLCELL_X32 FILLER_490_2887 ();
 FILLCELL_X32 FILLER_490_2919 ();
 FILLCELL_X32 FILLER_490_2951 ();
 FILLCELL_X32 FILLER_490_2983 ();
 FILLCELL_X32 FILLER_490_3015 ();
 FILLCELL_X32 FILLER_490_3047 ();
 FILLCELL_X32 FILLER_490_3079 ();
 FILLCELL_X32 FILLER_490_3111 ();
 FILLCELL_X8 FILLER_490_3143 ();
 FILLCELL_X4 FILLER_490_3151 ();
 FILLCELL_X2 FILLER_490_3155 ();
 FILLCELL_X32 FILLER_490_3158 ();
 FILLCELL_X32 FILLER_490_3190 ();
 FILLCELL_X32 FILLER_490_3222 ();
 FILLCELL_X32 FILLER_490_3254 ();
 FILLCELL_X32 FILLER_490_3286 ();
 FILLCELL_X32 FILLER_490_3318 ();
 FILLCELL_X32 FILLER_490_3350 ();
 FILLCELL_X32 FILLER_490_3382 ();
 FILLCELL_X32 FILLER_490_3414 ();
 FILLCELL_X32 FILLER_490_3446 ();
 FILLCELL_X32 FILLER_490_3478 ();
 FILLCELL_X32 FILLER_490_3510 ();
 FILLCELL_X32 FILLER_490_3542 ();
 FILLCELL_X32 FILLER_490_3574 ();
 FILLCELL_X32 FILLER_490_3606 ();
 FILLCELL_X32 FILLER_490_3638 ();
 FILLCELL_X32 FILLER_490_3670 ();
 FILLCELL_X32 FILLER_490_3702 ();
 FILLCELL_X4 FILLER_490_3734 ();
 FILLCELL_X32 FILLER_491_1 ();
 FILLCELL_X32 FILLER_491_33 ();
 FILLCELL_X32 FILLER_491_65 ();
 FILLCELL_X32 FILLER_491_97 ();
 FILLCELL_X32 FILLER_491_129 ();
 FILLCELL_X32 FILLER_491_161 ();
 FILLCELL_X32 FILLER_491_193 ();
 FILLCELL_X32 FILLER_491_225 ();
 FILLCELL_X32 FILLER_491_257 ();
 FILLCELL_X32 FILLER_491_289 ();
 FILLCELL_X32 FILLER_491_321 ();
 FILLCELL_X32 FILLER_491_353 ();
 FILLCELL_X32 FILLER_491_385 ();
 FILLCELL_X32 FILLER_491_417 ();
 FILLCELL_X32 FILLER_491_449 ();
 FILLCELL_X32 FILLER_491_481 ();
 FILLCELL_X32 FILLER_491_513 ();
 FILLCELL_X32 FILLER_491_545 ();
 FILLCELL_X32 FILLER_491_577 ();
 FILLCELL_X32 FILLER_491_609 ();
 FILLCELL_X32 FILLER_491_641 ();
 FILLCELL_X32 FILLER_491_673 ();
 FILLCELL_X32 FILLER_491_705 ();
 FILLCELL_X32 FILLER_491_737 ();
 FILLCELL_X32 FILLER_491_769 ();
 FILLCELL_X32 FILLER_491_801 ();
 FILLCELL_X32 FILLER_491_833 ();
 FILLCELL_X32 FILLER_491_865 ();
 FILLCELL_X32 FILLER_491_897 ();
 FILLCELL_X32 FILLER_491_929 ();
 FILLCELL_X32 FILLER_491_961 ();
 FILLCELL_X32 FILLER_491_993 ();
 FILLCELL_X32 FILLER_491_1025 ();
 FILLCELL_X32 FILLER_491_1057 ();
 FILLCELL_X32 FILLER_491_1089 ();
 FILLCELL_X32 FILLER_491_1121 ();
 FILLCELL_X32 FILLER_491_1153 ();
 FILLCELL_X32 FILLER_491_1185 ();
 FILLCELL_X32 FILLER_491_1217 ();
 FILLCELL_X8 FILLER_491_1249 ();
 FILLCELL_X4 FILLER_491_1257 ();
 FILLCELL_X2 FILLER_491_1261 ();
 FILLCELL_X32 FILLER_491_1264 ();
 FILLCELL_X32 FILLER_491_1296 ();
 FILLCELL_X32 FILLER_491_1328 ();
 FILLCELL_X32 FILLER_491_1360 ();
 FILLCELL_X32 FILLER_491_1392 ();
 FILLCELL_X32 FILLER_491_1424 ();
 FILLCELL_X32 FILLER_491_1456 ();
 FILLCELL_X32 FILLER_491_1488 ();
 FILLCELL_X32 FILLER_491_1520 ();
 FILLCELL_X32 FILLER_491_1552 ();
 FILLCELL_X32 FILLER_491_1584 ();
 FILLCELL_X32 FILLER_491_1616 ();
 FILLCELL_X32 FILLER_491_1648 ();
 FILLCELL_X32 FILLER_491_1680 ();
 FILLCELL_X32 FILLER_491_1712 ();
 FILLCELL_X32 FILLER_491_1744 ();
 FILLCELL_X32 FILLER_491_1776 ();
 FILLCELL_X32 FILLER_491_1808 ();
 FILLCELL_X32 FILLER_491_1840 ();
 FILLCELL_X32 FILLER_491_1872 ();
 FILLCELL_X32 FILLER_491_1904 ();
 FILLCELL_X32 FILLER_491_1936 ();
 FILLCELL_X32 FILLER_491_1968 ();
 FILLCELL_X32 FILLER_491_2000 ();
 FILLCELL_X32 FILLER_491_2032 ();
 FILLCELL_X32 FILLER_491_2064 ();
 FILLCELL_X32 FILLER_491_2096 ();
 FILLCELL_X32 FILLER_491_2128 ();
 FILLCELL_X32 FILLER_491_2160 ();
 FILLCELL_X32 FILLER_491_2192 ();
 FILLCELL_X32 FILLER_491_2224 ();
 FILLCELL_X32 FILLER_491_2256 ();
 FILLCELL_X32 FILLER_491_2288 ();
 FILLCELL_X32 FILLER_491_2320 ();
 FILLCELL_X32 FILLER_491_2352 ();
 FILLCELL_X32 FILLER_491_2384 ();
 FILLCELL_X32 FILLER_491_2416 ();
 FILLCELL_X32 FILLER_491_2448 ();
 FILLCELL_X32 FILLER_491_2480 ();
 FILLCELL_X8 FILLER_491_2512 ();
 FILLCELL_X4 FILLER_491_2520 ();
 FILLCELL_X2 FILLER_491_2524 ();
 FILLCELL_X32 FILLER_491_2527 ();
 FILLCELL_X32 FILLER_491_2559 ();
 FILLCELL_X32 FILLER_491_2591 ();
 FILLCELL_X32 FILLER_491_2623 ();
 FILLCELL_X32 FILLER_491_2655 ();
 FILLCELL_X32 FILLER_491_2687 ();
 FILLCELL_X32 FILLER_491_2719 ();
 FILLCELL_X32 FILLER_491_2751 ();
 FILLCELL_X32 FILLER_491_2783 ();
 FILLCELL_X32 FILLER_491_2815 ();
 FILLCELL_X32 FILLER_491_2847 ();
 FILLCELL_X32 FILLER_491_2879 ();
 FILLCELL_X32 FILLER_491_2911 ();
 FILLCELL_X32 FILLER_491_2943 ();
 FILLCELL_X32 FILLER_491_2975 ();
 FILLCELL_X32 FILLER_491_3007 ();
 FILLCELL_X32 FILLER_491_3039 ();
 FILLCELL_X32 FILLER_491_3071 ();
 FILLCELL_X32 FILLER_491_3103 ();
 FILLCELL_X32 FILLER_491_3135 ();
 FILLCELL_X32 FILLER_491_3167 ();
 FILLCELL_X32 FILLER_491_3199 ();
 FILLCELL_X32 FILLER_491_3231 ();
 FILLCELL_X32 FILLER_491_3263 ();
 FILLCELL_X32 FILLER_491_3295 ();
 FILLCELL_X32 FILLER_491_3327 ();
 FILLCELL_X32 FILLER_491_3359 ();
 FILLCELL_X32 FILLER_491_3391 ();
 FILLCELL_X32 FILLER_491_3423 ();
 FILLCELL_X32 FILLER_491_3455 ();
 FILLCELL_X32 FILLER_491_3487 ();
 FILLCELL_X32 FILLER_491_3519 ();
 FILLCELL_X32 FILLER_491_3551 ();
 FILLCELL_X32 FILLER_491_3583 ();
 FILLCELL_X32 FILLER_491_3615 ();
 FILLCELL_X32 FILLER_491_3647 ();
 FILLCELL_X32 FILLER_491_3679 ();
 FILLCELL_X16 FILLER_491_3711 ();
 FILLCELL_X8 FILLER_491_3727 ();
 FILLCELL_X2 FILLER_491_3735 ();
 FILLCELL_X1 FILLER_491_3737 ();
 FILLCELL_X32 FILLER_492_1 ();
 FILLCELL_X32 FILLER_492_33 ();
 FILLCELL_X32 FILLER_492_65 ();
 FILLCELL_X32 FILLER_492_97 ();
 FILLCELL_X32 FILLER_492_129 ();
 FILLCELL_X32 FILLER_492_161 ();
 FILLCELL_X32 FILLER_492_193 ();
 FILLCELL_X32 FILLER_492_225 ();
 FILLCELL_X32 FILLER_492_257 ();
 FILLCELL_X32 FILLER_492_289 ();
 FILLCELL_X32 FILLER_492_321 ();
 FILLCELL_X32 FILLER_492_353 ();
 FILLCELL_X32 FILLER_492_385 ();
 FILLCELL_X32 FILLER_492_417 ();
 FILLCELL_X32 FILLER_492_449 ();
 FILLCELL_X32 FILLER_492_481 ();
 FILLCELL_X32 FILLER_492_513 ();
 FILLCELL_X32 FILLER_492_545 ();
 FILLCELL_X32 FILLER_492_577 ();
 FILLCELL_X16 FILLER_492_609 ();
 FILLCELL_X4 FILLER_492_625 ();
 FILLCELL_X2 FILLER_492_629 ();
 FILLCELL_X32 FILLER_492_632 ();
 FILLCELL_X32 FILLER_492_664 ();
 FILLCELL_X32 FILLER_492_696 ();
 FILLCELL_X32 FILLER_492_728 ();
 FILLCELL_X32 FILLER_492_760 ();
 FILLCELL_X32 FILLER_492_792 ();
 FILLCELL_X32 FILLER_492_824 ();
 FILLCELL_X32 FILLER_492_856 ();
 FILLCELL_X32 FILLER_492_888 ();
 FILLCELL_X32 FILLER_492_920 ();
 FILLCELL_X32 FILLER_492_952 ();
 FILLCELL_X32 FILLER_492_984 ();
 FILLCELL_X32 FILLER_492_1016 ();
 FILLCELL_X32 FILLER_492_1048 ();
 FILLCELL_X32 FILLER_492_1080 ();
 FILLCELL_X32 FILLER_492_1112 ();
 FILLCELL_X32 FILLER_492_1144 ();
 FILLCELL_X32 FILLER_492_1176 ();
 FILLCELL_X32 FILLER_492_1208 ();
 FILLCELL_X32 FILLER_492_1240 ();
 FILLCELL_X32 FILLER_492_1272 ();
 FILLCELL_X32 FILLER_492_1304 ();
 FILLCELL_X32 FILLER_492_1336 ();
 FILLCELL_X32 FILLER_492_1368 ();
 FILLCELL_X32 FILLER_492_1400 ();
 FILLCELL_X32 FILLER_492_1432 ();
 FILLCELL_X32 FILLER_492_1464 ();
 FILLCELL_X32 FILLER_492_1496 ();
 FILLCELL_X32 FILLER_492_1528 ();
 FILLCELL_X32 FILLER_492_1560 ();
 FILLCELL_X32 FILLER_492_1592 ();
 FILLCELL_X32 FILLER_492_1624 ();
 FILLCELL_X32 FILLER_492_1656 ();
 FILLCELL_X32 FILLER_492_1688 ();
 FILLCELL_X32 FILLER_492_1720 ();
 FILLCELL_X32 FILLER_492_1752 ();
 FILLCELL_X32 FILLER_492_1784 ();
 FILLCELL_X32 FILLER_492_1816 ();
 FILLCELL_X32 FILLER_492_1848 ();
 FILLCELL_X8 FILLER_492_1880 ();
 FILLCELL_X4 FILLER_492_1888 ();
 FILLCELL_X2 FILLER_492_1892 ();
 FILLCELL_X32 FILLER_492_1895 ();
 FILLCELL_X32 FILLER_492_1927 ();
 FILLCELL_X32 FILLER_492_1959 ();
 FILLCELL_X32 FILLER_492_1991 ();
 FILLCELL_X32 FILLER_492_2023 ();
 FILLCELL_X32 FILLER_492_2055 ();
 FILLCELL_X32 FILLER_492_2087 ();
 FILLCELL_X32 FILLER_492_2119 ();
 FILLCELL_X32 FILLER_492_2151 ();
 FILLCELL_X32 FILLER_492_2183 ();
 FILLCELL_X32 FILLER_492_2215 ();
 FILLCELL_X32 FILLER_492_2247 ();
 FILLCELL_X32 FILLER_492_2279 ();
 FILLCELL_X32 FILLER_492_2311 ();
 FILLCELL_X32 FILLER_492_2343 ();
 FILLCELL_X32 FILLER_492_2375 ();
 FILLCELL_X32 FILLER_492_2407 ();
 FILLCELL_X32 FILLER_492_2439 ();
 FILLCELL_X32 FILLER_492_2471 ();
 FILLCELL_X32 FILLER_492_2503 ();
 FILLCELL_X32 FILLER_492_2535 ();
 FILLCELL_X32 FILLER_492_2567 ();
 FILLCELL_X32 FILLER_492_2599 ();
 FILLCELL_X32 FILLER_492_2631 ();
 FILLCELL_X32 FILLER_492_2663 ();
 FILLCELL_X32 FILLER_492_2695 ();
 FILLCELL_X32 FILLER_492_2727 ();
 FILLCELL_X32 FILLER_492_2759 ();
 FILLCELL_X32 FILLER_492_2791 ();
 FILLCELL_X32 FILLER_492_2823 ();
 FILLCELL_X32 FILLER_492_2855 ();
 FILLCELL_X32 FILLER_492_2887 ();
 FILLCELL_X32 FILLER_492_2919 ();
 FILLCELL_X32 FILLER_492_2951 ();
 FILLCELL_X32 FILLER_492_2983 ();
 FILLCELL_X32 FILLER_492_3015 ();
 FILLCELL_X32 FILLER_492_3047 ();
 FILLCELL_X32 FILLER_492_3079 ();
 FILLCELL_X32 FILLER_492_3111 ();
 FILLCELL_X8 FILLER_492_3143 ();
 FILLCELL_X4 FILLER_492_3151 ();
 FILLCELL_X2 FILLER_492_3155 ();
 FILLCELL_X32 FILLER_492_3158 ();
 FILLCELL_X32 FILLER_492_3190 ();
 FILLCELL_X32 FILLER_492_3222 ();
 FILLCELL_X32 FILLER_492_3254 ();
 FILLCELL_X32 FILLER_492_3286 ();
 FILLCELL_X32 FILLER_492_3318 ();
 FILLCELL_X32 FILLER_492_3350 ();
 FILLCELL_X32 FILLER_492_3382 ();
 FILLCELL_X32 FILLER_492_3414 ();
 FILLCELL_X32 FILLER_492_3446 ();
 FILLCELL_X32 FILLER_492_3478 ();
 FILLCELL_X32 FILLER_492_3510 ();
 FILLCELL_X32 FILLER_492_3542 ();
 FILLCELL_X32 FILLER_492_3574 ();
 FILLCELL_X32 FILLER_492_3606 ();
 FILLCELL_X32 FILLER_492_3638 ();
 FILLCELL_X32 FILLER_492_3670 ();
 FILLCELL_X32 FILLER_492_3702 ();
 FILLCELL_X4 FILLER_492_3734 ();
 FILLCELL_X32 FILLER_493_1 ();
 FILLCELL_X32 FILLER_493_33 ();
 FILLCELL_X32 FILLER_493_65 ();
 FILLCELL_X32 FILLER_493_97 ();
 FILLCELL_X32 FILLER_493_129 ();
 FILLCELL_X32 FILLER_493_161 ();
 FILLCELL_X32 FILLER_493_193 ();
 FILLCELL_X32 FILLER_493_225 ();
 FILLCELL_X32 FILLER_493_257 ();
 FILLCELL_X32 FILLER_493_289 ();
 FILLCELL_X32 FILLER_493_321 ();
 FILLCELL_X32 FILLER_493_353 ();
 FILLCELL_X32 FILLER_493_385 ();
 FILLCELL_X32 FILLER_493_417 ();
 FILLCELL_X32 FILLER_493_449 ();
 FILLCELL_X32 FILLER_493_481 ();
 FILLCELL_X32 FILLER_493_513 ();
 FILLCELL_X32 FILLER_493_545 ();
 FILLCELL_X32 FILLER_493_577 ();
 FILLCELL_X32 FILLER_493_609 ();
 FILLCELL_X32 FILLER_493_641 ();
 FILLCELL_X32 FILLER_493_673 ();
 FILLCELL_X32 FILLER_493_705 ();
 FILLCELL_X32 FILLER_493_737 ();
 FILLCELL_X32 FILLER_493_769 ();
 FILLCELL_X32 FILLER_493_801 ();
 FILLCELL_X32 FILLER_493_833 ();
 FILLCELL_X32 FILLER_493_865 ();
 FILLCELL_X32 FILLER_493_897 ();
 FILLCELL_X32 FILLER_493_929 ();
 FILLCELL_X32 FILLER_493_961 ();
 FILLCELL_X32 FILLER_493_993 ();
 FILLCELL_X32 FILLER_493_1025 ();
 FILLCELL_X32 FILLER_493_1057 ();
 FILLCELL_X32 FILLER_493_1089 ();
 FILLCELL_X32 FILLER_493_1121 ();
 FILLCELL_X32 FILLER_493_1153 ();
 FILLCELL_X32 FILLER_493_1185 ();
 FILLCELL_X32 FILLER_493_1217 ();
 FILLCELL_X8 FILLER_493_1249 ();
 FILLCELL_X4 FILLER_493_1257 ();
 FILLCELL_X2 FILLER_493_1261 ();
 FILLCELL_X32 FILLER_493_1264 ();
 FILLCELL_X32 FILLER_493_1296 ();
 FILLCELL_X32 FILLER_493_1328 ();
 FILLCELL_X32 FILLER_493_1360 ();
 FILLCELL_X32 FILLER_493_1392 ();
 FILLCELL_X32 FILLER_493_1424 ();
 FILLCELL_X32 FILLER_493_1456 ();
 FILLCELL_X32 FILLER_493_1488 ();
 FILLCELL_X32 FILLER_493_1520 ();
 FILLCELL_X32 FILLER_493_1552 ();
 FILLCELL_X32 FILLER_493_1584 ();
 FILLCELL_X32 FILLER_493_1616 ();
 FILLCELL_X32 FILLER_493_1648 ();
 FILLCELL_X32 FILLER_493_1680 ();
 FILLCELL_X32 FILLER_493_1712 ();
 FILLCELL_X32 FILLER_493_1744 ();
 FILLCELL_X32 FILLER_493_1776 ();
 FILLCELL_X32 FILLER_493_1808 ();
 FILLCELL_X32 FILLER_493_1840 ();
 FILLCELL_X32 FILLER_493_1872 ();
 FILLCELL_X32 FILLER_493_1904 ();
 FILLCELL_X32 FILLER_493_1936 ();
 FILLCELL_X32 FILLER_493_1968 ();
 FILLCELL_X32 FILLER_493_2000 ();
 FILLCELL_X32 FILLER_493_2032 ();
 FILLCELL_X32 FILLER_493_2064 ();
 FILLCELL_X32 FILLER_493_2096 ();
 FILLCELL_X32 FILLER_493_2128 ();
 FILLCELL_X32 FILLER_493_2160 ();
 FILLCELL_X32 FILLER_493_2192 ();
 FILLCELL_X32 FILLER_493_2224 ();
 FILLCELL_X32 FILLER_493_2256 ();
 FILLCELL_X32 FILLER_493_2288 ();
 FILLCELL_X32 FILLER_493_2320 ();
 FILLCELL_X32 FILLER_493_2352 ();
 FILLCELL_X32 FILLER_493_2384 ();
 FILLCELL_X32 FILLER_493_2416 ();
 FILLCELL_X32 FILLER_493_2448 ();
 FILLCELL_X32 FILLER_493_2480 ();
 FILLCELL_X8 FILLER_493_2512 ();
 FILLCELL_X4 FILLER_493_2520 ();
 FILLCELL_X2 FILLER_493_2524 ();
 FILLCELL_X32 FILLER_493_2527 ();
 FILLCELL_X32 FILLER_493_2559 ();
 FILLCELL_X32 FILLER_493_2591 ();
 FILLCELL_X32 FILLER_493_2623 ();
 FILLCELL_X32 FILLER_493_2655 ();
 FILLCELL_X32 FILLER_493_2687 ();
 FILLCELL_X32 FILLER_493_2719 ();
 FILLCELL_X32 FILLER_493_2751 ();
 FILLCELL_X32 FILLER_493_2783 ();
 FILLCELL_X32 FILLER_493_2815 ();
 FILLCELL_X32 FILLER_493_2847 ();
 FILLCELL_X32 FILLER_493_2879 ();
 FILLCELL_X32 FILLER_493_2911 ();
 FILLCELL_X32 FILLER_493_2943 ();
 FILLCELL_X32 FILLER_493_2975 ();
 FILLCELL_X32 FILLER_493_3007 ();
 FILLCELL_X32 FILLER_493_3039 ();
 FILLCELL_X32 FILLER_493_3071 ();
 FILLCELL_X32 FILLER_493_3103 ();
 FILLCELL_X32 FILLER_493_3135 ();
 FILLCELL_X32 FILLER_493_3167 ();
 FILLCELL_X32 FILLER_493_3199 ();
 FILLCELL_X32 FILLER_493_3231 ();
 FILLCELL_X32 FILLER_493_3263 ();
 FILLCELL_X32 FILLER_493_3295 ();
 FILLCELL_X32 FILLER_493_3327 ();
 FILLCELL_X32 FILLER_493_3359 ();
 FILLCELL_X32 FILLER_493_3391 ();
 FILLCELL_X32 FILLER_493_3423 ();
 FILLCELL_X32 FILLER_493_3455 ();
 FILLCELL_X32 FILLER_493_3487 ();
 FILLCELL_X32 FILLER_493_3519 ();
 FILLCELL_X32 FILLER_493_3551 ();
 FILLCELL_X32 FILLER_493_3583 ();
 FILLCELL_X32 FILLER_493_3615 ();
 FILLCELL_X32 FILLER_493_3647 ();
 FILLCELL_X32 FILLER_493_3679 ();
 FILLCELL_X16 FILLER_493_3711 ();
 FILLCELL_X8 FILLER_493_3727 ();
 FILLCELL_X2 FILLER_493_3735 ();
 FILLCELL_X1 FILLER_493_3737 ();
 FILLCELL_X32 FILLER_494_1 ();
 FILLCELL_X32 FILLER_494_33 ();
 FILLCELL_X32 FILLER_494_65 ();
 FILLCELL_X32 FILLER_494_97 ();
 FILLCELL_X32 FILLER_494_129 ();
 FILLCELL_X32 FILLER_494_161 ();
 FILLCELL_X32 FILLER_494_193 ();
 FILLCELL_X32 FILLER_494_225 ();
 FILLCELL_X32 FILLER_494_257 ();
 FILLCELL_X32 FILLER_494_289 ();
 FILLCELL_X32 FILLER_494_321 ();
 FILLCELL_X32 FILLER_494_353 ();
 FILLCELL_X32 FILLER_494_385 ();
 FILLCELL_X32 FILLER_494_417 ();
 FILLCELL_X32 FILLER_494_449 ();
 FILLCELL_X32 FILLER_494_481 ();
 FILLCELL_X32 FILLER_494_513 ();
 FILLCELL_X32 FILLER_494_545 ();
 FILLCELL_X32 FILLER_494_577 ();
 FILLCELL_X16 FILLER_494_609 ();
 FILLCELL_X4 FILLER_494_625 ();
 FILLCELL_X2 FILLER_494_629 ();
 FILLCELL_X32 FILLER_494_632 ();
 FILLCELL_X32 FILLER_494_664 ();
 FILLCELL_X32 FILLER_494_696 ();
 FILLCELL_X32 FILLER_494_728 ();
 FILLCELL_X32 FILLER_494_760 ();
 FILLCELL_X32 FILLER_494_792 ();
 FILLCELL_X32 FILLER_494_824 ();
 FILLCELL_X32 FILLER_494_856 ();
 FILLCELL_X32 FILLER_494_888 ();
 FILLCELL_X32 FILLER_494_920 ();
 FILLCELL_X32 FILLER_494_952 ();
 FILLCELL_X32 FILLER_494_984 ();
 FILLCELL_X32 FILLER_494_1016 ();
 FILLCELL_X32 FILLER_494_1048 ();
 FILLCELL_X32 FILLER_494_1080 ();
 FILLCELL_X32 FILLER_494_1112 ();
 FILLCELL_X32 FILLER_494_1144 ();
 FILLCELL_X32 FILLER_494_1176 ();
 FILLCELL_X32 FILLER_494_1208 ();
 FILLCELL_X32 FILLER_494_1240 ();
 FILLCELL_X32 FILLER_494_1272 ();
 FILLCELL_X32 FILLER_494_1304 ();
 FILLCELL_X32 FILLER_494_1336 ();
 FILLCELL_X32 FILLER_494_1368 ();
 FILLCELL_X32 FILLER_494_1400 ();
 FILLCELL_X32 FILLER_494_1432 ();
 FILLCELL_X32 FILLER_494_1464 ();
 FILLCELL_X32 FILLER_494_1496 ();
 FILLCELL_X32 FILLER_494_1528 ();
 FILLCELL_X32 FILLER_494_1560 ();
 FILLCELL_X32 FILLER_494_1592 ();
 FILLCELL_X32 FILLER_494_1624 ();
 FILLCELL_X32 FILLER_494_1656 ();
 FILLCELL_X32 FILLER_494_1688 ();
 FILLCELL_X32 FILLER_494_1720 ();
 FILLCELL_X32 FILLER_494_1752 ();
 FILLCELL_X32 FILLER_494_1784 ();
 FILLCELL_X32 FILLER_494_1816 ();
 FILLCELL_X32 FILLER_494_1848 ();
 FILLCELL_X8 FILLER_494_1880 ();
 FILLCELL_X4 FILLER_494_1888 ();
 FILLCELL_X2 FILLER_494_1892 ();
 FILLCELL_X32 FILLER_494_1895 ();
 FILLCELL_X32 FILLER_494_1927 ();
 FILLCELL_X32 FILLER_494_1959 ();
 FILLCELL_X32 FILLER_494_1991 ();
 FILLCELL_X32 FILLER_494_2023 ();
 FILLCELL_X32 FILLER_494_2055 ();
 FILLCELL_X32 FILLER_494_2087 ();
 FILLCELL_X32 FILLER_494_2119 ();
 FILLCELL_X32 FILLER_494_2151 ();
 FILLCELL_X32 FILLER_494_2183 ();
 FILLCELL_X32 FILLER_494_2215 ();
 FILLCELL_X32 FILLER_494_2247 ();
 FILLCELL_X32 FILLER_494_2279 ();
 FILLCELL_X32 FILLER_494_2311 ();
 FILLCELL_X32 FILLER_494_2343 ();
 FILLCELL_X32 FILLER_494_2375 ();
 FILLCELL_X32 FILLER_494_2407 ();
 FILLCELL_X32 FILLER_494_2439 ();
 FILLCELL_X32 FILLER_494_2471 ();
 FILLCELL_X32 FILLER_494_2503 ();
 FILLCELL_X32 FILLER_494_2535 ();
 FILLCELL_X32 FILLER_494_2567 ();
 FILLCELL_X32 FILLER_494_2599 ();
 FILLCELL_X32 FILLER_494_2631 ();
 FILLCELL_X32 FILLER_494_2663 ();
 FILLCELL_X32 FILLER_494_2695 ();
 FILLCELL_X32 FILLER_494_2727 ();
 FILLCELL_X32 FILLER_494_2759 ();
 FILLCELL_X32 FILLER_494_2791 ();
 FILLCELL_X32 FILLER_494_2823 ();
 FILLCELL_X32 FILLER_494_2855 ();
 FILLCELL_X32 FILLER_494_2887 ();
 FILLCELL_X32 FILLER_494_2919 ();
 FILLCELL_X32 FILLER_494_2951 ();
 FILLCELL_X32 FILLER_494_2983 ();
 FILLCELL_X32 FILLER_494_3015 ();
 FILLCELL_X32 FILLER_494_3047 ();
 FILLCELL_X32 FILLER_494_3079 ();
 FILLCELL_X32 FILLER_494_3111 ();
 FILLCELL_X8 FILLER_494_3143 ();
 FILLCELL_X4 FILLER_494_3151 ();
 FILLCELL_X2 FILLER_494_3155 ();
 FILLCELL_X32 FILLER_494_3158 ();
 FILLCELL_X32 FILLER_494_3190 ();
 FILLCELL_X32 FILLER_494_3222 ();
 FILLCELL_X32 FILLER_494_3254 ();
 FILLCELL_X32 FILLER_494_3286 ();
 FILLCELL_X32 FILLER_494_3318 ();
 FILLCELL_X32 FILLER_494_3350 ();
 FILLCELL_X32 FILLER_494_3382 ();
 FILLCELL_X32 FILLER_494_3414 ();
 FILLCELL_X32 FILLER_494_3446 ();
 FILLCELL_X32 FILLER_494_3478 ();
 FILLCELL_X32 FILLER_494_3510 ();
 FILLCELL_X32 FILLER_494_3542 ();
 FILLCELL_X32 FILLER_494_3574 ();
 FILLCELL_X32 FILLER_494_3606 ();
 FILLCELL_X32 FILLER_494_3638 ();
 FILLCELL_X32 FILLER_494_3670 ();
 FILLCELL_X32 FILLER_494_3702 ();
 FILLCELL_X4 FILLER_494_3734 ();
 FILLCELL_X32 FILLER_495_1 ();
 FILLCELL_X32 FILLER_495_33 ();
 FILLCELL_X32 FILLER_495_65 ();
 FILLCELL_X32 FILLER_495_97 ();
 FILLCELL_X32 FILLER_495_129 ();
 FILLCELL_X32 FILLER_495_161 ();
 FILLCELL_X32 FILLER_495_193 ();
 FILLCELL_X32 FILLER_495_225 ();
 FILLCELL_X32 FILLER_495_257 ();
 FILLCELL_X32 FILLER_495_289 ();
 FILLCELL_X32 FILLER_495_321 ();
 FILLCELL_X32 FILLER_495_353 ();
 FILLCELL_X32 FILLER_495_385 ();
 FILLCELL_X32 FILLER_495_417 ();
 FILLCELL_X32 FILLER_495_449 ();
 FILLCELL_X32 FILLER_495_481 ();
 FILLCELL_X32 FILLER_495_513 ();
 FILLCELL_X32 FILLER_495_545 ();
 FILLCELL_X32 FILLER_495_577 ();
 FILLCELL_X32 FILLER_495_609 ();
 FILLCELL_X32 FILLER_495_641 ();
 FILLCELL_X32 FILLER_495_673 ();
 FILLCELL_X32 FILLER_495_705 ();
 FILLCELL_X32 FILLER_495_737 ();
 FILLCELL_X32 FILLER_495_769 ();
 FILLCELL_X32 FILLER_495_801 ();
 FILLCELL_X32 FILLER_495_833 ();
 FILLCELL_X32 FILLER_495_865 ();
 FILLCELL_X32 FILLER_495_897 ();
 FILLCELL_X32 FILLER_495_929 ();
 FILLCELL_X32 FILLER_495_961 ();
 FILLCELL_X32 FILLER_495_993 ();
 FILLCELL_X32 FILLER_495_1025 ();
 FILLCELL_X32 FILLER_495_1057 ();
 FILLCELL_X32 FILLER_495_1089 ();
 FILLCELL_X32 FILLER_495_1121 ();
 FILLCELL_X32 FILLER_495_1153 ();
 FILLCELL_X32 FILLER_495_1185 ();
 FILLCELL_X32 FILLER_495_1217 ();
 FILLCELL_X8 FILLER_495_1249 ();
 FILLCELL_X4 FILLER_495_1257 ();
 FILLCELL_X2 FILLER_495_1261 ();
 FILLCELL_X32 FILLER_495_1264 ();
 FILLCELL_X32 FILLER_495_1296 ();
 FILLCELL_X32 FILLER_495_1328 ();
 FILLCELL_X32 FILLER_495_1360 ();
 FILLCELL_X32 FILLER_495_1392 ();
 FILLCELL_X32 FILLER_495_1424 ();
 FILLCELL_X32 FILLER_495_1456 ();
 FILLCELL_X32 FILLER_495_1488 ();
 FILLCELL_X32 FILLER_495_1520 ();
 FILLCELL_X32 FILLER_495_1552 ();
 FILLCELL_X32 FILLER_495_1584 ();
 FILLCELL_X32 FILLER_495_1616 ();
 FILLCELL_X32 FILLER_495_1648 ();
 FILLCELL_X32 FILLER_495_1680 ();
 FILLCELL_X32 FILLER_495_1712 ();
 FILLCELL_X32 FILLER_495_1744 ();
 FILLCELL_X32 FILLER_495_1776 ();
 FILLCELL_X32 FILLER_495_1808 ();
 FILLCELL_X32 FILLER_495_1840 ();
 FILLCELL_X32 FILLER_495_1872 ();
 FILLCELL_X32 FILLER_495_1904 ();
 FILLCELL_X32 FILLER_495_1936 ();
 FILLCELL_X32 FILLER_495_1968 ();
 FILLCELL_X32 FILLER_495_2000 ();
 FILLCELL_X32 FILLER_495_2032 ();
 FILLCELL_X32 FILLER_495_2064 ();
 FILLCELL_X32 FILLER_495_2096 ();
 FILLCELL_X32 FILLER_495_2128 ();
 FILLCELL_X32 FILLER_495_2160 ();
 FILLCELL_X32 FILLER_495_2192 ();
 FILLCELL_X32 FILLER_495_2224 ();
 FILLCELL_X32 FILLER_495_2256 ();
 FILLCELL_X32 FILLER_495_2288 ();
 FILLCELL_X32 FILLER_495_2320 ();
 FILLCELL_X32 FILLER_495_2352 ();
 FILLCELL_X32 FILLER_495_2384 ();
 FILLCELL_X32 FILLER_495_2416 ();
 FILLCELL_X32 FILLER_495_2448 ();
 FILLCELL_X32 FILLER_495_2480 ();
 FILLCELL_X8 FILLER_495_2512 ();
 FILLCELL_X4 FILLER_495_2520 ();
 FILLCELL_X2 FILLER_495_2524 ();
 FILLCELL_X32 FILLER_495_2527 ();
 FILLCELL_X32 FILLER_495_2559 ();
 FILLCELL_X32 FILLER_495_2591 ();
 FILLCELL_X32 FILLER_495_2623 ();
 FILLCELL_X32 FILLER_495_2655 ();
 FILLCELL_X32 FILLER_495_2687 ();
 FILLCELL_X32 FILLER_495_2719 ();
 FILLCELL_X32 FILLER_495_2751 ();
 FILLCELL_X32 FILLER_495_2783 ();
 FILLCELL_X32 FILLER_495_2815 ();
 FILLCELL_X32 FILLER_495_2847 ();
 FILLCELL_X32 FILLER_495_2879 ();
 FILLCELL_X32 FILLER_495_2911 ();
 FILLCELL_X32 FILLER_495_2943 ();
 FILLCELL_X32 FILLER_495_2975 ();
 FILLCELL_X32 FILLER_495_3007 ();
 FILLCELL_X32 FILLER_495_3039 ();
 FILLCELL_X32 FILLER_495_3071 ();
 FILLCELL_X32 FILLER_495_3103 ();
 FILLCELL_X32 FILLER_495_3135 ();
 FILLCELL_X32 FILLER_495_3167 ();
 FILLCELL_X32 FILLER_495_3199 ();
 FILLCELL_X32 FILLER_495_3231 ();
 FILLCELL_X32 FILLER_495_3263 ();
 FILLCELL_X32 FILLER_495_3295 ();
 FILLCELL_X32 FILLER_495_3327 ();
 FILLCELL_X32 FILLER_495_3359 ();
 FILLCELL_X32 FILLER_495_3391 ();
 FILLCELL_X32 FILLER_495_3423 ();
 FILLCELL_X32 FILLER_495_3455 ();
 FILLCELL_X32 FILLER_495_3487 ();
 FILLCELL_X32 FILLER_495_3519 ();
 FILLCELL_X32 FILLER_495_3551 ();
 FILLCELL_X32 FILLER_495_3583 ();
 FILLCELL_X32 FILLER_495_3615 ();
 FILLCELL_X32 FILLER_495_3647 ();
 FILLCELL_X32 FILLER_495_3679 ();
 FILLCELL_X16 FILLER_495_3711 ();
 FILLCELL_X8 FILLER_495_3727 ();
 FILLCELL_X2 FILLER_495_3735 ();
 FILLCELL_X1 FILLER_495_3737 ();
 FILLCELL_X32 FILLER_496_1 ();
 FILLCELL_X32 FILLER_496_33 ();
 FILLCELL_X32 FILLER_496_65 ();
 FILLCELL_X32 FILLER_496_97 ();
 FILLCELL_X32 FILLER_496_129 ();
 FILLCELL_X32 FILLER_496_161 ();
 FILLCELL_X32 FILLER_496_193 ();
 FILLCELL_X32 FILLER_496_225 ();
 FILLCELL_X32 FILLER_496_257 ();
 FILLCELL_X32 FILLER_496_289 ();
 FILLCELL_X32 FILLER_496_321 ();
 FILLCELL_X32 FILLER_496_353 ();
 FILLCELL_X32 FILLER_496_385 ();
 FILLCELL_X32 FILLER_496_417 ();
 FILLCELL_X32 FILLER_496_449 ();
 FILLCELL_X32 FILLER_496_481 ();
 FILLCELL_X32 FILLER_496_513 ();
 FILLCELL_X32 FILLER_496_545 ();
 FILLCELL_X32 FILLER_496_577 ();
 FILLCELL_X16 FILLER_496_609 ();
 FILLCELL_X4 FILLER_496_625 ();
 FILLCELL_X2 FILLER_496_629 ();
 FILLCELL_X32 FILLER_496_632 ();
 FILLCELL_X32 FILLER_496_664 ();
 FILLCELL_X32 FILLER_496_696 ();
 FILLCELL_X32 FILLER_496_728 ();
 FILLCELL_X32 FILLER_496_760 ();
 FILLCELL_X32 FILLER_496_792 ();
 FILLCELL_X32 FILLER_496_824 ();
 FILLCELL_X32 FILLER_496_856 ();
 FILLCELL_X32 FILLER_496_888 ();
 FILLCELL_X32 FILLER_496_920 ();
 FILLCELL_X32 FILLER_496_952 ();
 FILLCELL_X32 FILLER_496_984 ();
 FILLCELL_X32 FILLER_496_1016 ();
 FILLCELL_X32 FILLER_496_1048 ();
 FILLCELL_X32 FILLER_496_1080 ();
 FILLCELL_X32 FILLER_496_1112 ();
 FILLCELL_X32 FILLER_496_1144 ();
 FILLCELL_X32 FILLER_496_1176 ();
 FILLCELL_X32 FILLER_496_1208 ();
 FILLCELL_X32 FILLER_496_1240 ();
 FILLCELL_X32 FILLER_496_1272 ();
 FILLCELL_X32 FILLER_496_1304 ();
 FILLCELL_X32 FILLER_496_1336 ();
 FILLCELL_X32 FILLER_496_1368 ();
 FILLCELL_X32 FILLER_496_1400 ();
 FILLCELL_X32 FILLER_496_1432 ();
 FILLCELL_X32 FILLER_496_1464 ();
 FILLCELL_X32 FILLER_496_1496 ();
 FILLCELL_X32 FILLER_496_1528 ();
 FILLCELL_X32 FILLER_496_1560 ();
 FILLCELL_X32 FILLER_496_1592 ();
 FILLCELL_X32 FILLER_496_1624 ();
 FILLCELL_X32 FILLER_496_1656 ();
 FILLCELL_X32 FILLER_496_1688 ();
 FILLCELL_X32 FILLER_496_1720 ();
 FILLCELL_X32 FILLER_496_1752 ();
 FILLCELL_X32 FILLER_496_1784 ();
 FILLCELL_X32 FILLER_496_1816 ();
 FILLCELL_X32 FILLER_496_1848 ();
 FILLCELL_X8 FILLER_496_1880 ();
 FILLCELL_X4 FILLER_496_1888 ();
 FILLCELL_X2 FILLER_496_1892 ();
 FILLCELL_X32 FILLER_496_1895 ();
 FILLCELL_X32 FILLER_496_1927 ();
 FILLCELL_X32 FILLER_496_1959 ();
 FILLCELL_X32 FILLER_496_1991 ();
 FILLCELL_X32 FILLER_496_2023 ();
 FILLCELL_X32 FILLER_496_2055 ();
 FILLCELL_X32 FILLER_496_2087 ();
 FILLCELL_X32 FILLER_496_2119 ();
 FILLCELL_X32 FILLER_496_2151 ();
 FILLCELL_X32 FILLER_496_2183 ();
 FILLCELL_X32 FILLER_496_2215 ();
 FILLCELL_X32 FILLER_496_2247 ();
 FILLCELL_X32 FILLER_496_2279 ();
 FILLCELL_X32 FILLER_496_2311 ();
 FILLCELL_X32 FILLER_496_2343 ();
 FILLCELL_X32 FILLER_496_2375 ();
 FILLCELL_X32 FILLER_496_2407 ();
 FILLCELL_X32 FILLER_496_2439 ();
 FILLCELL_X32 FILLER_496_2471 ();
 FILLCELL_X32 FILLER_496_2503 ();
 FILLCELL_X32 FILLER_496_2535 ();
 FILLCELL_X32 FILLER_496_2567 ();
 FILLCELL_X32 FILLER_496_2599 ();
 FILLCELL_X32 FILLER_496_2631 ();
 FILLCELL_X32 FILLER_496_2663 ();
 FILLCELL_X32 FILLER_496_2695 ();
 FILLCELL_X32 FILLER_496_2727 ();
 FILLCELL_X32 FILLER_496_2759 ();
 FILLCELL_X32 FILLER_496_2791 ();
 FILLCELL_X32 FILLER_496_2823 ();
 FILLCELL_X32 FILLER_496_2855 ();
 FILLCELL_X32 FILLER_496_2887 ();
 FILLCELL_X32 FILLER_496_2919 ();
 FILLCELL_X32 FILLER_496_2951 ();
 FILLCELL_X32 FILLER_496_2983 ();
 FILLCELL_X32 FILLER_496_3015 ();
 FILLCELL_X32 FILLER_496_3047 ();
 FILLCELL_X32 FILLER_496_3079 ();
 FILLCELL_X32 FILLER_496_3111 ();
 FILLCELL_X8 FILLER_496_3143 ();
 FILLCELL_X4 FILLER_496_3151 ();
 FILLCELL_X2 FILLER_496_3155 ();
 FILLCELL_X32 FILLER_496_3158 ();
 FILLCELL_X32 FILLER_496_3190 ();
 FILLCELL_X32 FILLER_496_3222 ();
 FILLCELL_X32 FILLER_496_3254 ();
 FILLCELL_X32 FILLER_496_3286 ();
 FILLCELL_X32 FILLER_496_3318 ();
 FILLCELL_X32 FILLER_496_3350 ();
 FILLCELL_X32 FILLER_496_3382 ();
 FILLCELL_X32 FILLER_496_3414 ();
 FILLCELL_X32 FILLER_496_3446 ();
 FILLCELL_X32 FILLER_496_3478 ();
 FILLCELL_X32 FILLER_496_3510 ();
 FILLCELL_X32 FILLER_496_3542 ();
 FILLCELL_X32 FILLER_496_3574 ();
 FILLCELL_X32 FILLER_496_3606 ();
 FILLCELL_X32 FILLER_496_3638 ();
 FILLCELL_X32 FILLER_496_3670 ();
 FILLCELL_X32 FILLER_496_3702 ();
 FILLCELL_X4 FILLER_496_3734 ();
 FILLCELL_X32 FILLER_497_1 ();
 FILLCELL_X32 FILLER_497_33 ();
 FILLCELL_X32 FILLER_497_65 ();
 FILLCELL_X32 FILLER_497_97 ();
 FILLCELL_X32 FILLER_497_129 ();
 FILLCELL_X32 FILLER_497_161 ();
 FILLCELL_X32 FILLER_497_193 ();
 FILLCELL_X32 FILLER_497_225 ();
 FILLCELL_X32 FILLER_497_257 ();
 FILLCELL_X32 FILLER_497_289 ();
 FILLCELL_X32 FILLER_497_321 ();
 FILLCELL_X32 FILLER_497_353 ();
 FILLCELL_X32 FILLER_497_385 ();
 FILLCELL_X32 FILLER_497_417 ();
 FILLCELL_X32 FILLER_497_449 ();
 FILLCELL_X32 FILLER_497_481 ();
 FILLCELL_X32 FILLER_497_513 ();
 FILLCELL_X32 FILLER_497_545 ();
 FILLCELL_X32 FILLER_497_577 ();
 FILLCELL_X32 FILLER_497_609 ();
 FILLCELL_X32 FILLER_497_641 ();
 FILLCELL_X32 FILLER_497_673 ();
 FILLCELL_X32 FILLER_497_705 ();
 FILLCELL_X32 FILLER_497_737 ();
 FILLCELL_X32 FILLER_497_769 ();
 FILLCELL_X32 FILLER_497_801 ();
 FILLCELL_X32 FILLER_497_833 ();
 FILLCELL_X32 FILLER_497_865 ();
 FILLCELL_X32 FILLER_497_897 ();
 FILLCELL_X32 FILLER_497_929 ();
 FILLCELL_X32 FILLER_497_961 ();
 FILLCELL_X32 FILLER_497_993 ();
 FILLCELL_X32 FILLER_497_1025 ();
 FILLCELL_X32 FILLER_497_1057 ();
 FILLCELL_X32 FILLER_497_1089 ();
 FILLCELL_X32 FILLER_497_1121 ();
 FILLCELL_X32 FILLER_497_1153 ();
 FILLCELL_X32 FILLER_497_1185 ();
 FILLCELL_X32 FILLER_497_1217 ();
 FILLCELL_X8 FILLER_497_1249 ();
 FILLCELL_X4 FILLER_497_1257 ();
 FILLCELL_X2 FILLER_497_1261 ();
 FILLCELL_X32 FILLER_497_1264 ();
 FILLCELL_X32 FILLER_497_1296 ();
 FILLCELL_X32 FILLER_497_1328 ();
 FILLCELL_X32 FILLER_497_1360 ();
 FILLCELL_X32 FILLER_497_1392 ();
 FILLCELL_X32 FILLER_497_1424 ();
 FILLCELL_X32 FILLER_497_1456 ();
 FILLCELL_X32 FILLER_497_1488 ();
 FILLCELL_X32 FILLER_497_1520 ();
 FILLCELL_X32 FILLER_497_1552 ();
 FILLCELL_X32 FILLER_497_1584 ();
 FILLCELL_X32 FILLER_497_1616 ();
 FILLCELL_X32 FILLER_497_1648 ();
 FILLCELL_X32 FILLER_497_1680 ();
 FILLCELL_X32 FILLER_497_1712 ();
 FILLCELL_X32 FILLER_497_1744 ();
 FILLCELL_X32 FILLER_497_1776 ();
 FILLCELL_X32 FILLER_497_1808 ();
 FILLCELL_X32 FILLER_497_1840 ();
 FILLCELL_X32 FILLER_497_1872 ();
 FILLCELL_X32 FILLER_497_1904 ();
 FILLCELL_X32 FILLER_497_1936 ();
 FILLCELL_X32 FILLER_497_1968 ();
 FILLCELL_X32 FILLER_497_2000 ();
 FILLCELL_X32 FILLER_497_2032 ();
 FILLCELL_X32 FILLER_497_2064 ();
 FILLCELL_X32 FILLER_497_2096 ();
 FILLCELL_X32 FILLER_497_2128 ();
 FILLCELL_X32 FILLER_497_2160 ();
 FILLCELL_X32 FILLER_497_2192 ();
 FILLCELL_X32 FILLER_497_2224 ();
 FILLCELL_X32 FILLER_497_2256 ();
 FILLCELL_X32 FILLER_497_2288 ();
 FILLCELL_X32 FILLER_497_2320 ();
 FILLCELL_X32 FILLER_497_2352 ();
 FILLCELL_X32 FILLER_497_2384 ();
 FILLCELL_X32 FILLER_497_2416 ();
 FILLCELL_X32 FILLER_497_2448 ();
 FILLCELL_X32 FILLER_497_2480 ();
 FILLCELL_X8 FILLER_497_2512 ();
 FILLCELL_X4 FILLER_497_2520 ();
 FILLCELL_X2 FILLER_497_2524 ();
 FILLCELL_X32 FILLER_497_2527 ();
 FILLCELL_X32 FILLER_497_2559 ();
 FILLCELL_X32 FILLER_497_2591 ();
 FILLCELL_X32 FILLER_497_2623 ();
 FILLCELL_X32 FILLER_497_2655 ();
 FILLCELL_X32 FILLER_497_2687 ();
 FILLCELL_X32 FILLER_497_2719 ();
 FILLCELL_X32 FILLER_497_2751 ();
 FILLCELL_X32 FILLER_497_2783 ();
 FILLCELL_X32 FILLER_497_2815 ();
 FILLCELL_X32 FILLER_497_2847 ();
 FILLCELL_X32 FILLER_497_2879 ();
 FILLCELL_X32 FILLER_497_2911 ();
 FILLCELL_X32 FILLER_497_2943 ();
 FILLCELL_X32 FILLER_497_2975 ();
 FILLCELL_X32 FILLER_497_3007 ();
 FILLCELL_X32 FILLER_497_3039 ();
 FILLCELL_X32 FILLER_497_3071 ();
 FILLCELL_X32 FILLER_497_3103 ();
 FILLCELL_X32 FILLER_497_3135 ();
 FILLCELL_X32 FILLER_497_3167 ();
 FILLCELL_X32 FILLER_497_3199 ();
 FILLCELL_X32 FILLER_497_3231 ();
 FILLCELL_X32 FILLER_497_3263 ();
 FILLCELL_X32 FILLER_497_3295 ();
 FILLCELL_X32 FILLER_497_3327 ();
 FILLCELL_X32 FILLER_497_3359 ();
 FILLCELL_X32 FILLER_497_3391 ();
 FILLCELL_X32 FILLER_497_3423 ();
 FILLCELL_X32 FILLER_497_3455 ();
 FILLCELL_X32 FILLER_497_3487 ();
 FILLCELL_X32 FILLER_497_3519 ();
 FILLCELL_X32 FILLER_497_3551 ();
 FILLCELL_X32 FILLER_497_3583 ();
 FILLCELL_X32 FILLER_497_3615 ();
 FILLCELL_X32 FILLER_497_3647 ();
 FILLCELL_X32 FILLER_497_3679 ();
 FILLCELL_X16 FILLER_497_3711 ();
 FILLCELL_X8 FILLER_497_3727 ();
 FILLCELL_X2 FILLER_497_3735 ();
 FILLCELL_X1 FILLER_497_3737 ();
 FILLCELL_X32 FILLER_498_1 ();
 FILLCELL_X32 FILLER_498_33 ();
 FILLCELL_X32 FILLER_498_65 ();
 FILLCELL_X32 FILLER_498_97 ();
 FILLCELL_X32 FILLER_498_129 ();
 FILLCELL_X32 FILLER_498_161 ();
 FILLCELL_X32 FILLER_498_193 ();
 FILLCELL_X32 FILLER_498_225 ();
 FILLCELL_X32 FILLER_498_257 ();
 FILLCELL_X32 FILLER_498_289 ();
 FILLCELL_X32 FILLER_498_321 ();
 FILLCELL_X32 FILLER_498_353 ();
 FILLCELL_X32 FILLER_498_385 ();
 FILLCELL_X32 FILLER_498_417 ();
 FILLCELL_X32 FILLER_498_449 ();
 FILLCELL_X32 FILLER_498_481 ();
 FILLCELL_X32 FILLER_498_513 ();
 FILLCELL_X32 FILLER_498_545 ();
 FILLCELL_X32 FILLER_498_577 ();
 FILLCELL_X16 FILLER_498_609 ();
 FILLCELL_X4 FILLER_498_625 ();
 FILLCELL_X2 FILLER_498_629 ();
 FILLCELL_X32 FILLER_498_632 ();
 FILLCELL_X32 FILLER_498_664 ();
 FILLCELL_X32 FILLER_498_696 ();
 FILLCELL_X32 FILLER_498_728 ();
 FILLCELL_X32 FILLER_498_760 ();
 FILLCELL_X32 FILLER_498_792 ();
 FILLCELL_X32 FILLER_498_824 ();
 FILLCELL_X32 FILLER_498_856 ();
 FILLCELL_X32 FILLER_498_888 ();
 FILLCELL_X32 FILLER_498_920 ();
 FILLCELL_X32 FILLER_498_952 ();
 FILLCELL_X32 FILLER_498_984 ();
 FILLCELL_X32 FILLER_498_1016 ();
 FILLCELL_X32 FILLER_498_1048 ();
 FILLCELL_X32 FILLER_498_1080 ();
 FILLCELL_X32 FILLER_498_1112 ();
 FILLCELL_X32 FILLER_498_1144 ();
 FILLCELL_X32 FILLER_498_1176 ();
 FILLCELL_X32 FILLER_498_1208 ();
 FILLCELL_X32 FILLER_498_1240 ();
 FILLCELL_X32 FILLER_498_1272 ();
 FILLCELL_X32 FILLER_498_1304 ();
 FILLCELL_X32 FILLER_498_1336 ();
 FILLCELL_X32 FILLER_498_1368 ();
 FILLCELL_X32 FILLER_498_1400 ();
 FILLCELL_X32 FILLER_498_1432 ();
 FILLCELL_X32 FILLER_498_1464 ();
 FILLCELL_X32 FILLER_498_1496 ();
 FILLCELL_X32 FILLER_498_1528 ();
 FILLCELL_X32 FILLER_498_1560 ();
 FILLCELL_X32 FILLER_498_1592 ();
 FILLCELL_X32 FILLER_498_1624 ();
 FILLCELL_X32 FILLER_498_1656 ();
 FILLCELL_X32 FILLER_498_1688 ();
 FILLCELL_X32 FILLER_498_1720 ();
 FILLCELL_X32 FILLER_498_1752 ();
 FILLCELL_X32 FILLER_498_1784 ();
 FILLCELL_X32 FILLER_498_1816 ();
 FILLCELL_X32 FILLER_498_1848 ();
 FILLCELL_X8 FILLER_498_1880 ();
 FILLCELL_X4 FILLER_498_1888 ();
 FILLCELL_X2 FILLER_498_1892 ();
 FILLCELL_X32 FILLER_498_1895 ();
 FILLCELL_X32 FILLER_498_1927 ();
 FILLCELL_X32 FILLER_498_1959 ();
 FILLCELL_X32 FILLER_498_1991 ();
 FILLCELL_X32 FILLER_498_2023 ();
 FILLCELL_X32 FILLER_498_2055 ();
 FILLCELL_X32 FILLER_498_2087 ();
 FILLCELL_X32 FILLER_498_2119 ();
 FILLCELL_X32 FILLER_498_2151 ();
 FILLCELL_X32 FILLER_498_2183 ();
 FILLCELL_X32 FILLER_498_2215 ();
 FILLCELL_X32 FILLER_498_2247 ();
 FILLCELL_X32 FILLER_498_2279 ();
 FILLCELL_X32 FILLER_498_2311 ();
 FILLCELL_X32 FILLER_498_2343 ();
 FILLCELL_X32 FILLER_498_2375 ();
 FILLCELL_X32 FILLER_498_2407 ();
 FILLCELL_X32 FILLER_498_2439 ();
 FILLCELL_X32 FILLER_498_2471 ();
 FILLCELL_X32 FILLER_498_2503 ();
 FILLCELL_X32 FILLER_498_2535 ();
 FILLCELL_X32 FILLER_498_2567 ();
 FILLCELL_X32 FILLER_498_2599 ();
 FILLCELL_X32 FILLER_498_2631 ();
 FILLCELL_X32 FILLER_498_2663 ();
 FILLCELL_X32 FILLER_498_2695 ();
 FILLCELL_X32 FILLER_498_2727 ();
 FILLCELL_X32 FILLER_498_2759 ();
 FILLCELL_X32 FILLER_498_2791 ();
 FILLCELL_X32 FILLER_498_2823 ();
 FILLCELL_X32 FILLER_498_2855 ();
 FILLCELL_X32 FILLER_498_2887 ();
 FILLCELL_X32 FILLER_498_2919 ();
 FILLCELL_X32 FILLER_498_2951 ();
 FILLCELL_X32 FILLER_498_2983 ();
 FILLCELL_X32 FILLER_498_3015 ();
 FILLCELL_X32 FILLER_498_3047 ();
 FILLCELL_X32 FILLER_498_3079 ();
 FILLCELL_X32 FILLER_498_3111 ();
 FILLCELL_X8 FILLER_498_3143 ();
 FILLCELL_X4 FILLER_498_3151 ();
 FILLCELL_X2 FILLER_498_3155 ();
 FILLCELL_X32 FILLER_498_3158 ();
 FILLCELL_X32 FILLER_498_3190 ();
 FILLCELL_X32 FILLER_498_3222 ();
 FILLCELL_X32 FILLER_498_3254 ();
 FILLCELL_X32 FILLER_498_3286 ();
 FILLCELL_X32 FILLER_498_3318 ();
 FILLCELL_X32 FILLER_498_3350 ();
 FILLCELL_X32 FILLER_498_3382 ();
 FILLCELL_X32 FILLER_498_3414 ();
 FILLCELL_X32 FILLER_498_3446 ();
 FILLCELL_X32 FILLER_498_3478 ();
 FILLCELL_X32 FILLER_498_3510 ();
 FILLCELL_X32 FILLER_498_3542 ();
 FILLCELL_X32 FILLER_498_3574 ();
 FILLCELL_X32 FILLER_498_3606 ();
 FILLCELL_X32 FILLER_498_3638 ();
 FILLCELL_X32 FILLER_498_3670 ();
 FILLCELL_X32 FILLER_498_3702 ();
 FILLCELL_X4 FILLER_498_3734 ();
 FILLCELL_X32 FILLER_499_1 ();
 FILLCELL_X32 FILLER_499_33 ();
 FILLCELL_X32 FILLER_499_65 ();
 FILLCELL_X32 FILLER_499_97 ();
 FILLCELL_X32 FILLER_499_129 ();
 FILLCELL_X32 FILLER_499_161 ();
 FILLCELL_X32 FILLER_499_193 ();
 FILLCELL_X32 FILLER_499_225 ();
 FILLCELL_X32 FILLER_499_257 ();
 FILLCELL_X32 FILLER_499_289 ();
 FILLCELL_X32 FILLER_499_321 ();
 FILLCELL_X32 FILLER_499_353 ();
 FILLCELL_X32 FILLER_499_385 ();
 FILLCELL_X32 FILLER_499_417 ();
 FILLCELL_X32 FILLER_499_449 ();
 FILLCELL_X32 FILLER_499_481 ();
 FILLCELL_X32 FILLER_499_513 ();
 FILLCELL_X32 FILLER_499_545 ();
 FILLCELL_X32 FILLER_499_577 ();
 FILLCELL_X32 FILLER_499_609 ();
 FILLCELL_X32 FILLER_499_641 ();
 FILLCELL_X32 FILLER_499_673 ();
 FILLCELL_X32 FILLER_499_705 ();
 FILLCELL_X32 FILLER_499_737 ();
 FILLCELL_X32 FILLER_499_769 ();
 FILLCELL_X32 FILLER_499_801 ();
 FILLCELL_X32 FILLER_499_833 ();
 FILLCELL_X32 FILLER_499_865 ();
 FILLCELL_X32 FILLER_499_897 ();
 FILLCELL_X32 FILLER_499_929 ();
 FILLCELL_X32 FILLER_499_961 ();
 FILLCELL_X32 FILLER_499_993 ();
 FILLCELL_X32 FILLER_499_1025 ();
 FILLCELL_X32 FILLER_499_1057 ();
 FILLCELL_X32 FILLER_499_1089 ();
 FILLCELL_X32 FILLER_499_1121 ();
 FILLCELL_X32 FILLER_499_1153 ();
 FILLCELL_X32 FILLER_499_1185 ();
 FILLCELL_X32 FILLER_499_1217 ();
 FILLCELL_X8 FILLER_499_1249 ();
 FILLCELL_X4 FILLER_499_1257 ();
 FILLCELL_X2 FILLER_499_1261 ();
 FILLCELL_X32 FILLER_499_1264 ();
 FILLCELL_X32 FILLER_499_1296 ();
 FILLCELL_X32 FILLER_499_1328 ();
 FILLCELL_X32 FILLER_499_1360 ();
 FILLCELL_X32 FILLER_499_1392 ();
 FILLCELL_X32 FILLER_499_1424 ();
 FILLCELL_X32 FILLER_499_1456 ();
 FILLCELL_X32 FILLER_499_1488 ();
 FILLCELL_X32 FILLER_499_1520 ();
 FILLCELL_X32 FILLER_499_1552 ();
 FILLCELL_X32 FILLER_499_1584 ();
 FILLCELL_X32 FILLER_499_1616 ();
 FILLCELL_X32 FILLER_499_1648 ();
 FILLCELL_X32 FILLER_499_1680 ();
 FILLCELL_X32 FILLER_499_1712 ();
 FILLCELL_X32 FILLER_499_1744 ();
 FILLCELL_X32 FILLER_499_1776 ();
 FILLCELL_X32 FILLER_499_1808 ();
 FILLCELL_X32 FILLER_499_1840 ();
 FILLCELL_X32 FILLER_499_1872 ();
 FILLCELL_X32 FILLER_499_1904 ();
 FILLCELL_X32 FILLER_499_1936 ();
 FILLCELL_X32 FILLER_499_1968 ();
 FILLCELL_X32 FILLER_499_2000 ();
 FILLCELL_X32 FILLER_499_2032 ();
 FILLCELL_X32 FILLER_499_2064 ();
 FILLCELL_X32 FILLER_499_2096 ();
 FILLCELL_X32 FILLER_499_2128 ();
 FILLCELL_X32 FILLER_499_2160 ();
 FILLCELL_X32 FILLER_499_2192 ();
 FILLCELL_X32 FILLER_499_2224 ();
 FILLCELL_X32 FILLER_499_2256 ();
 FILLCELL_X32 FILLER_499_2288 ();
 FILLCELL_X32 FILLER_499_2320 ();
 FILLCELL_X32 FILLER_499_2352 ();
 FILLCELL_X32 FILLER_499_2384 ();
 FILLCELL_X32 FILLER_499_2416 ();
 FILLCELL_X32 FILLER_499_2448 ();
 FILLCELL_X32 FILLER_499_2480 ();
 FILLCELL_X8 FILLER_499_2512 ();
 FILLCELL_X4 FILLER_499_2520 ();
 FILLCELL_X2 FILLER_499_2524 ();
 FILLCELL_X32 FILLER_499_2527 ();
 FILLCELL_X32 FILLER_499_2559 ();
 FILLCELL_X32 FILLER_499_2591 ();
 FILLCELL_X32 FILLER_499_2623 ();
 FILLCELL_X32 FILLER_499_2655 ();
 FILLCELL_X32 FILLER_499_2687 ();
 FILLCELL_X32 FILLER_499_2719 ();
 FILLCELL_X32 FILLER_499_2751 ();
 FILLCELL_X32 FILLER_499_2783 ();
 FILLCELL_X32 FILLER_499_2815 ();
 FILLCELL_X32 FILLER_499_2847 ();
 FILLCELL_X32 FILLER_499_2879 ();
 FILLCELL_X32 FILLER_499_2911 ();
 FILLCELL_X32 FILLER_499_2943 ();
 FILLCELL_X32 FILLER_499_2975 ();
 FILLCELL_X32 FILLER_499_3007 ();
 FILLCELL_X32 FILLER_499_3039 ();
 FILLCELL_X32 FILLER_499_3071 ();
 FILLCELL_X32 FILLER_499_3103 ();
 FILLCELL_X32 FILLER_499_3135 ();
 FILLCELL_X32 FILLER_499_3167 ();
 FILLCELL_X32 FILLER_499_3199 ();
 FILLCELL_X32 FILLER_499_3231 ();
 FILLCELL_X32 FILLER_499_3263 ();
 FILLCELL_X32 FILLER_499_3295 ();
 FILLCELL_X32 FILLER_499_3327 ();
 FILLCELL_X32 FILLER_499_3359 ();
 FILLCELL_X32 FILLER_499_3391 ();
 FILLCELL_X32 FILLER_499_3423 ();
 FILLCELL_X32 FILLER_499_3455 ();
 FILLCELL_X32 FILLER_499_3487 ();
 FILLCELL_X32 FILLER_499_3519 ();
 FILLCELL_X32 FILLER_499_3551 ();
 FILLCELL_X32 FILLER_499_3583 ();
 FILLCELL_X32 FILLER_499_3615 ();
 FILLCELL_X32 FILLER_499_3647 ();
 FILLCELL_X32 FILLER_499_3679 ();
 FILLCELL_X16 FILLER_499_3711 ();
 FILLCELL_X8 FILLER_499_3727 ();
 FILLCELL_X2 FILLER_499_3735 ();
 FILLCELL_X1 FILLER_499_3737 ();
 FILLCELL_X32 FILLER_500_1 ();
 FILLCELL_X32 FILLER_500_33 ();
 FILLCELL_X32 FILLER_500_65 ();
 FILLCELL_X32 FILLER_500_97 ();
 FILLCELL_X32 FILLER_500_129 ();
 FILLCELL_X32 FILLER_500_161 ();
 FILLCELL_X32 FILLER_500_193 ();
 FILLCELL_X32 FILLER_500_225 ();
 FILLCELL_X32 FILLER_500_257 ();
 FILLCELL_X32 FILLER_500_289 ();
 FILLCELL_X32 FILLER_500_321 ();
 FILLCELL_X32 FILLER_500_353 ();
 FILLCELL_X32 FILLER_500_385 ();
 FILLCELL_X32 FILLER_500_417 ();
 FILLCELL_X32 FILLER_500_449 ();
 FILLCELL_X32 FILLER_500_481 ();
 FILLCELL_X32 FILLER_500_513 ();
 FILLCELL_X32 FILLER_500_545 ();
 FILLCELL_X32 FILLER_500_577 ();
 FILLCELL_X16 FILLER_500_609 ();
 FILLCELL_X4 FILLER_500_625 ();
 FILLCELL_X2 FILLER_500_629 ();
 FILLCELL_X32 FILLER_500_632 ();
 FILLCELL_X32 FILLER_500_664 ();
 FILLCELL_X32 FILLER_500_696 ();
 FILLCELL_X32 FILLER_500_728 ();
 FILLCELL_X32 FILLER_500_760 ();
 FILLCELL_X32 FILLER_500_792 ();
 FILLCELL_X32 FILLER_500_824 ();
 FILLCELL_X32 FILLER_500_856 ();
 FILLCELL_X32 FILLER_500_888 ();
 FILLCELL_X32 FILLER_500_920 ();
 FILLCELL_X32 FILLER_500_952 ();
 FILLCELL_X32 FILLER_500_984 ();
 FILLCELL_X32 FILLER_500_1016 ();
 FILLCELL_X32 FILLER_500_1048 ();
 FILLCELL_X32 FILLER_500_1080 ();
 FILLCELL_X32 FILLER_500_1112 ();
 FILLCELL_X32 FILLER_500_1144 ();
 FILLCELL_X32 FILLER_500_1176 ();
 FILLCELL_X32 FILLER_500_1208 ();
 FILLCELL_X32 FILLER_500_1240 ();
 FILLCELL_X32 FILLER_500_1272 ();
 FILLCELL_X32 FILLER_500_1304 ();
 FILLCELL_X32 FILLER_500_1336 ();
 FILLCELL_X32 FILLER_500_1368 ();
 FILLCELL_X32 FILLER_500_1400 ();
 FILLCELL_X32 FILLER_500_1432 ();
 FILLCELL_X32 FILLER_500_1464 ();
 FILLCELL_X32 FILLER_500_1496 ();
 FILLCELL_X32 FILLER_500_1528 ();
 FILLCELL_X32 FILLER_500_1560 ();
 FILLCELL_X32 FILLER_500_1592 ();
 FILLCELL_X32 FILLER_500_1624 ();
 FILLCELL_X32 FILLER_500_1656 ();
 FILLCELL_X32 FILLER_500_1688 ();
 FILLCELL_X32 FILLER_500_1720 ();
 FILLCELL_X32 FILLER_500_1752 ();
 FILLCELL_X32 FILLER_500_1784 ();
 FILLCELL_X32 FILLER_500_1816 ();
 FILLCELL_X32 FILLER_500_1848 ();
 FILLCELL_X8 FILLER_500_1880 ();
 FILLCELL_X4 FILLER_500_1888 ();
 FILLCELL_X2 FILLER_500_1892 ();
 FILLCELL_X32 FILLER_500_1895 ();
 FILLCELL_X32 FILLER_500_1927 ();
 FILLCELL_X32 FILLER_500_1959 ();
 FILLCELL_X32 FILLER_500_1991 ();
 FILLCELL_X32 FILLER_500_2023 ();
 FILLCELL_X32 FILLER_500_2055 ();
 FILLCELL_X32 FILLER_500_2087 ();
 FILLCELL_X32 FILLER_500_2119 ();
 FILLCELL_X32 FILLER_500_2151 ();
 FILLCELL_X32 FILLER_500_2183 ();
 FILLCELL_X32 FILLER_500_2215 ();
 FILLCELL_X32 FILLER_500_2247 ();
 FILLCELL_X32 FILLER_500_2279 ();
 FILLCELL_X32 FILLER_500_2311 ();
 FILLCELL_X32 FILLER_500_2343 ();
 FILLCELL_X32 FILLER_500_2375 ();
 FILLCELL_X32 FILLER_500_2407 ();
 FILLCELL_X32 FILLER_500_2439 ();
 FILLCELL_X32 FILLER_500_2471 ();
 FILLCELL_X32 FILLER_500_2503 ();
 FILLCELL_X32 FILLER_500_2535 ();
 FILLCELL_X32 FILLER_500_2567 ();
 FILLCELL_X32 FILLER_500_2599 ();
 FILLCELL_X32 FILLER_500_2631 ();
 FILLCELL_X32 FILLER_500_2663 ();
 FILLCELL_X32 FILLER_500_2695 ();
 FILLCELL_X32 FILLER_500_2727 ();
 FILLCELL_X32 FILLER_500_2759 ();
 FILLCELL_X32 FILLER_500_2791 ();
 FILLCELL_X32 FILLER_500_2823 ();
 FILLCELL_X32 FILLER_500_2855 ();
 FILLCELL_X32 FILLER_500_2887 ();
 FILLCELL_X32 FILLER_500_2919 ();
 FILLCELL_X32 FILLER_500_2951 ();
 FILLCELL_X32 FILLER_500_2983 ();
 FILLCELL_X32 FILLER_500_3015 ();
 FILLCELL_X32 FILLER_500_3047 ();
 FILLCELL_X32 FILLER_500_3079 ();
 FILLCELL_X32 FILLER_500_3111 ();
 FILLCELL_X8 FILLER_500_3143 ();
 FILLCELL_X4 FILLER_500_3151 ();
 FILLCELL_X2 FILLER_500_3155 ();
 FILLCELL_X32 FILLER_500_3158 ();
 FILLCELL_X32 FILLER_500_3190 ();
 FILLCELL_X32 FILLER_500_3222 ();
 FILLCELL_X32 FILLER_500_3254 ();
 FILLCELL_X32 FILLER_500_3286 ();
 FILLCELL_X32 FILLER_500_3318 ();
 FILLCELL_X32 FILLER_500_3350 ();
 FILLCELL_X32 FILLER_500_3382 ();
 FILLCELL_X32 FILLER_500_3414 ();
 FILLCELL_X32 FILLER_500_3446 ();
 FILLCELL_X32 FILLER_500_3478 ();
 FILLCELL_X32 FILLER_500_3510 ();
 FILLCELL_X32 FILLER_500_3542 ();
 FILLCELL_X32 FILLER_500_3574 ();
 FILLCELL_X32 FILLER_500_3606 ();
 FILLCELL_X32 FILLER_500_3638 ();
 FILLCELL_X32 FILLER_500_3670 ();
 FILLCELL_X32 FILLER_500_3702 ();
 FILLCELL_X4 FILLER_500_3734 ();
 FILLCELL_X32 FILLER_501_1 ();
 FILLCELL_X32 FILLER_501_33 ();
 FILLCELL_X32 FILLER_501_65 ();
 FILLCELL_X32 FILLER_501_97 ();
 FILLCELL_X32 FILLER_501_129 ();
 FILLCELL_X32 FILLER_501_161 ();
 FILLCELL_X32 FILLER_501_193 ();
 FILLCELL_X32 FILLER_501_225 ();
 FILLCELL_X32 FILLER_501_257 ();
 FILLCELL_X32 FILLER_501_289 ();
 FILLCELL_X32 FILLER_501_321 ();
 FILLCELL_X32 FILLER_501_353 ();
 FILLCELL_X32 FILLER_501_385 ();
 FILLCELL_X32 FILLER_501_417 ();
 FILLCELL_X32 FILLER_501_449 ();
 FILLCELL_X32 FILLER_501_481 ();
 FILLCELL_X32 FILLER_501_513 ();
 FILLCELL_X32 FILLER_501_545 ();
 FILLCELL_X32 FILLER_501_577 ();
 FILLCELL_X32 FILLER_501_609 ();
 FILLCELL_X32 FILLER_501_641 ();
 FILLCELL_X32 FILLER_501_673 ();
 FILLCELL_X32 FILLER_501_705 ();
 FILLCELL_X32 FILLER_501_737 ();
 FILLCELL_X32 FILLER_501_769 ();
 FILLCELL_X32 FILLER_501_801 ();
 FILLCELL_X32 FILLER_501_833 ();
 FILLCELL_X32 FILLER_501_865 ();
 FILLCELL_X32 FILLER_501_897 ();
 FILLCELL_X32 FILLER_501_929 ();
 FILLCELL_X32 FILLER_501_961 ();
 FILLCELL_X32 FILLER_501_993 ();
 FILLCELL_X32 FILLER_501_1025 ();
 FILLCELL_X32 FILLER_501_1057 ();
 FILLCELL_X32 FILLER_501_1089 ();
 FILLCELL_X32 FILLER_501_1121 ();
 FILLCELL_X32 FILLER_501_1153 ();
 FILLCELL_X32 FILLER_501_1185 ();
 FILLCELL_X32 FILLER_501_1217 ();
 FILLCELL_X8 FILLER_501_1249 ();
 FILLCELL_X4 FILLER_501_1257 ();
 FILLCELL_X2 FILLER_501_1261 ();
 FILLCELL_X32 FILLER_501_1264 ();
 FILLCELL_X32 FILLER_501_1296 ();
 FILLCELL_X32 FILLER_501_1328 ();
 FILLCELL_X32 FILLER_501_1360 ();
 FILLCELL_X32 FILLER_501_1392 ();
 FILLCELL_X32 FILLER_501_1424 ();
 FILLCELL_X32 FILLER_501_1456 ();
 FILLCELL_X32 FILLER_501_1488 ();
 FILLCELL_X32 FILLER_501_1520 ();
 FILLCELL_X32 FILLER_501_1552 ();
 FILLCELL_X32 FILLER_501_1584 ();
 FILLCELL_X32 FILLER_501_1616 ();
 FILLCELL_X32 FILLER_501_1648 ();
 FILLCELL_X32 FILLER_501_1680 ();
 FILLCELL_X32 FILLER_501_1712 ();
 FILLCELL_X32 FILLER_501_1744 ();
 FILLCELL_X32 FILLER_501_1776 ();
 FILLCELL_X32 FILLER_501_1808 ();
 FILLCELL_X32 FILLER_501_1840 ();
 FILLCELL_X32 FILLER_501_1872 ();
 FILLCELL_X32 FILLER_501_1904 ();
 FILLCELL_X32 FILLER_501_1936 ();
 FILLCELL_X32 FILLER_501_1968 ();
 FILLCELL_X32 FILLER_501_2000 ();
 FILLCELL_X32 FILLER_501_2032 ();
 FILLCELL_X32 FILLER_501_2064 ();
 FILLCELL_X32 FILLER_501_2096 ();
 FILLCELL_X32 FILLER_501_2128 ();
 FILLCELL_X32 FILLER_501_2160 ();
 FILLCELL_X32 FILLER_501_2192 ();
 FILLCELL_X32 FILLER_501_2224 ();
 FILLCELL_X32 FILLER_501_2256 ();
 FILLCELL_X32 FILLER_501_2288 ();
 FILLCELL_X32 FILLER_501_2320 ();
 FILLCELL_X32 FILLER_501_2352 ();
 FILLCELL_X32 FILLER_501_2384 ();
 FILLCELL_X32 FILLER_501_2416 ();
 FILLCELL_X32 FILLER_501_2448 ();
 FILLCELL_X32 FILLER_501_2480 ();
 FILLCELL_X8 FILLER_501_2512 ();
 FILLCELL_X4 FILLER_501_2520 ();
 FILLCELL_X2 FILLER_501_2524 ();
 FILLCELL_X32 FILLER_501_2527 ();
 FILLCELL_X32 FILLER_501_2559 ();
 FILLCELL_X32 FILLER_501_2591 ();
 FILLCELL_X32 FILLER_501_2623 ();
 FILLCELL_X32 FILLER_501_2655 ();
 FILLCELL_X32 FILLER_501_2687 ();
 FILLCELL_X32 FILLER_501_2719 ();
 FILLCELL_X32 FILLER_501_2751 ();
 FILLCELL_X32 FILLER_501_2783 ();
 FILLCELL_X32 FILLER_501_2815 ();
 FILLCELL_X32 FILLER_501_2847 ();
 FILLCELL_X32 FILLER_501_2879 ();
 FILLCELL_X32 FILLER_501_2911 ();
 FILLCELL_X32 FILLER_501_2943 ();
 FILLCELL_X32 FILLER_501_2975 ();
 FILLCELL_X32 FILLER_501_3007 ();
 FILLCELL_X32 FILLER_501_3039 ();
 FILLCELL_X32 FILLER_501_3071 ();
 FILLCELL_X32 FILLER_501_3103 ();
 FILLCELL_X32 FILLER_501_3135 ();
 FILLCELL_X32 FILLER_501_3167 ();
 FILLCELL_X32 FILLER_501_3199 ();
 FILLCELL_X32 FILLER_501_3231 ();
 FILLCELL_X32 FILLER_501_3263 ();
 FILLCELL_X32 FILLER_501_3295 ();
 FILLCELL_X32 FILLER_501_3327 ();
 FILLCELL_X32 FILLER_501_3359 ();
 FILLCELL_X32 FILLER_501_3391 ();
 FILLCELL_X32 FILLER_501_3423 ();
 FILLCELL_X32 FILLER_501_3455 ();
 FILLCELL_X32 FILLER_501_3487 ();
 FILLCELL_X32 FILLER_501_3519 ();
 FILLCELL_X32 FILLER_501_3551 ();
 FILLCELL_X32 FILLER_501_3583 ();
 FILLCELL_X32 FILLER_501_3615 ();
 FILLCELL_X32 FILLER_501_3647 ();
 FILLCELL_X32 FILLER_501_3679 ();
 FILLCELL_X16 FILLER_501_3711 ();
 FILLCELL_X8 FILLER_501_3727 ();
 FILLCELL_X2 FILLER_501_3735 ();
 FILLCELL_X1 FILLER_501_3737 ();
 FILLCELL_X32 FILLER_502_1 ();
 FILLCELL_X32 FILLER_502_33 ();
 FILLCELL_X32 FILLER_502_65 ();
 FILLCELL_X32 FILLER_502_97 ();
 FILLCELL_X32 FILLER_502_129 ();
 FILLCELL_X32 FILLER_502_161 ();
 FILLCELL_X32 FILLER_502_193 ();
 FILLCELL_X32 FILLER_502_225 ();
 FILLCELL_X32 FILLER_502_257 ();
 FILLCELL_X32 FILLER_502_289 ();
 FILLCELL_X32 FILLER_502_321 ();
 FILLCELL_X32 FILLER_502_353 ();
 FILLCELL_X32 FILLER_502_385 ();
 FILLCELL_X32 FILLER_502_417 ();
 FILLCELL_X32 FILLER_502_449 ();
 FILLCELL_X32 FILLER_502_481 ();
 FILLCELL_X32 FILLER_502_513 ();
 FILLCELL_X32 FILLER_502_545 ();
 FILLCELL_X32 FILLER_502_577 ();
 FILLCELL_X16 FILLER_502_609 ();
 FILLCELL_X4 FILLER_502_625 ();
 FILLCELL_X2 FILLER_502_629 ();
 FILLCELL_X32 FILLER_502_632 ();
 FILLCELL_X32 FILLER_502_664 ();
 FILLCELL_X32 FILLER_502_696 ();
 FILLCELL_X32 FILLER_502_728 ();
 FILLCELL_X32 FILLER_502_760 ();
 FILLCELL_X32 FILLER_502_792 ();
 FILLCELL_X32 FILLER_502_824 ();
 FILLCELL_X32 FILLER_502_856 ();
 FILLCELL_X32 FILLER_502_888 ();
 FILLCELL_X32 FILLER_502_920 ();
 FILLCELL_X32 FILLER_502_952 ();
 FILLCELL_X32 FILLER_502_984 ();
 FILLCELL_X32 FILLER_502_1016 ();
 FILLCELL_X32 FILLER_502_1048 ();
 FILLCELL_X32 FILLER_502_1080 ();
 FILLCELL_X32 FILLER_502_1112 ();
 FILLCELL_X32 FILLER_502_1144 ();
 FILLCELL_X32 FILLER_502_1176 ();
 FILLCELL_X32 FILLER_502_1208 ();
 FILLCELL_X32 FILLER_502_1240 ();
 FILLCELL_X32 FILLER_502_1272 ();
 FILLCELL_X32 FILLER_502_1304 ();
 FILLCELL_X32 FILLER_502_1336 ();
 FILLCELL_X32 FILLER_502_1368 ();
 FILLCELL_X32 FILLER_502_1400 ();
 FILLCELL_X32 FILLER_502_1432 ();
 FILLCELL_X32 FILLER_502_1464 ();
 FILLCELL_X32 FILLER_502_1496 ();
 FILLCELL_X32 FILLER_502_1528 ();
 FILLCELL_X32 FILLER_502_1560 ();
 FILLCELL_X32 FILLER_502_1592 ();
 FILLCELL_X32 FILLER_502_1624 ();
 FILLCELL_X32 FILLER_502_1656 ();
 FILLCELL_X32 FILLER_502_1688 ();
 FILLCELL_X32 FILLER_502_1720 ();
 FILLCELL_X32 FILLER_502_1752 ();
 FILLCELL_X32 FILLER_502_1784 ();
 FILLCELL_X32 FILLER_502_1816 ();
 FILLCELL_X32 FILLER_502_1848 ();
 FILLCELL_X8 FILLER_502_1880 ();
 FILLCELL_X4 FILLER_502_1888 ();
 FILLCELL_X2 FILLER_502_1892 ();
 FILLCELL_X32 FILLER_502_1895 ();
 FILLCELL_X32 FILLER_502_1927 ();
 FILLCELL_X32 FILLER_502_1959 ();
 FILLCELL_X32 FILLER_502_1991 ();
 FILLCELL_X32 FILLER_502_2023 ();
 FILLCELL_X32 FILLER_502_2055 ();
 FILLCELL_X32 FILLER_502_2087 ();
 FILLCELL_X32 FILLER_502_2119 ();
 FILLCELL_X32 FILLER_502_2151 ();
 FILLCELL_X32 FILLER_502_2183 ();
 FILLCELL_X32 FILLER_502_2215 ();
 FILLCELL_X32 FILLER_502_2247 ();
 FILLCELL_X32 FILLER_502_2279 ();
 FILLCELL_X32 FILLER_502_2311 ();
 FILLCELL_X32 FILLER_502_2343 ();
 FILLCELL_X32 FILLER_502_2375 ();
 FILLCELL_X32 FILLER_502_2407 ();
 FILLCELL_X32 FILLER_502_2439 ();
 FILLCELL_X32 FILLER_502_2471 ();
 FILLCELL_X32 FILLER_502_2503 ();
 FILLCELL_X32 FILLER_502_2535 ();
 FILLCELL_X32 FILLER_502_2567 ();
 FILLCELL_X32 FILLER_502_2599 ();
 FILLCELL_X32 FILLER_502_2631 ();
 FILLCELL_X32 FILLER_502_2663 ();
 FILLCELL_X32 FILLER_502_2695 ();
 FILLCELL_X32 FILLER_502_2727 ();
 FILLCELL_X32 FILLER_502_2759 ();
 FILLCELL_X32 FILLER_502_2791 ();
 FILLCELL_X32 FILLER_502_2823 ();
 FILLCELL_X32 FILLER_502_2855 ();
 FILLCELL_X32 FILLER_502_2887 ();
 FILLCELL_X32 FILLER_502_2919 ();
 FILLCELL_X32 FILLER_502_2951 ();
 FILLCELL_X32 FILLER_502_2983 ();
 FILLCELL_X32 FILLER_502_3015 ();
 FILLCELL_X32 FILLER_502_3047 ();
 FILLCELL_X32 FILLER_502_3079 ();
 FILLCELL_X32 FILLER_502_3111 ();
 FILLCELL_X8 FILLER_502_3143 ();
 FILLCELL_X4 FILLER_502_3151 ();
 FILLCELL_X2 FILLER_502_3155 ();
 FILLCELL_X32 FILLER_502_3158 ();
 FILLCELL_X32 FILLER_502_3190 ();
 FILLCELL_X32 FILLER_502_3222 ();
 FILLCELL_X32 FILLER_502_3254 ();
 FILLCELL_X32 FILLER_502_3286 ();
 FILLCELL_X32 FILLER_502_3318 ();
 FILLCELL_X32 FILLER_502_3350 ();
 FILLCELL_X32 FILLER_502_3382 ();
 FILLCELL_X32 FILLER_502_3414 ();
 FILLCELL_X32 FILLER_502_3446 ();
 FILLCELL_X32 FILLER_502_3478 ();
 FILLCELL_X32 FILLER_502_3510 ();
 FILLCELL_X32 FILLER_502_3542 ();
 FILLCELL_X32 FILLER_502_3574 ();
 FILLCELL_X32 FILLER_502_3606 ();
 FILLCELL_X32 FILLER_502_3638 ();
 FILLCELL_X32 FILLER_502_3670 ();
 FILLCELL_X32 FILLER_502_3702 ();
 FILLCELL_X4 FILLER_502_3734 ();
 FILLCELL_X32 FILLER_503_1 ();
 FILLCELL_X32 FILLER_503_33 ();
 FILLCELL_X32 FILLER_503_65 ();
 FILLCELL_X32 FILLER_503_97 ();
 FILLCELL_X32 FILLER_503_129 ();
 FILLCELL_X32 FILLER_503_161 ();
 FILLCELL_X32 FILLER_503_193 ();
 FILLCELL_X32 FILLER_503_225 ();
 FILLCELL_X32 FILLER_503_257 ();
 FILLCELL_X32 FILLER_503_289 ();
 FILLCELL_X32 FILLER_503_321 ();
 FILLCELL_X32 FILLER_503_353 ();
 FILLCELL_X32 FILLER_503_385 ();
 FILLCELL_X32 FILLER_503_417 ();
 FILLCELL_X32 FILLER_503_449 ();
 FILLCELL_X32 FILLER_503_481 ();
 FILLCELL_X32 FILLER_503_513 ();
 FILLCELL_X32 FILLER_503_545 ();
 FILLCELL_X32 FILLER_503_577 ();
 FILLCELL_X32 FILLER_503_609 ();
 FILLCELL_X32 FILLER_503_641 ();
 FILLCELL_X32 FILLER_503_673 ();
 FILLCELL_X32 FILLER_503_705 ();
 FILLCELL_X32 FILLER_503_737 ();
 FILLCELL_X32 FILLER_503_769 ();
 FILLCELL_X32 FILLER_503_801 ();
 FILLCELL_X32 FILLER_503_833 ();
 FILLCELL_X32 FILLER_503_865 ();
 FILLCELL_X32 FILLER_503_897 ();
 FILLCELL_X32 FILLER_503_929 ();
 FILLCELL_X32 FILLER_503_961 ();
 FILLCELL_X32 FILLER_503_993 ();
 FILLCELL_X32 FILLER_503_1025 ();
 FILLCELL_X32 FILLER_503_1057 ();
 FILLCELL_X32 FILLER_503_1089 ();
 FILLCELL_X32 FILLER_503_1121 ();
 FILLCELL_X32 FILLER_503_1153 ();
 FILLCELL_X32 FILLER_503_1185 ();
 FILLCELL_X32 FILLER_503_1217 ();
 FILLCELL_X8 FILLER_503_1249 ();
 FILLCELL_X4 FILLER_503_1257 ();
 FILLCELL_X2 FILLER_503_1261 ();
 FILLCELL_X32 FILLER_503_1264 ();
 FILLCELL_X32 FILLER_503_1296 ();
 FILLCELL_X32 FILLER_503_1328 ();
 FILLCELL_X32 FILLER_503_1360 ();
 FILLCELL_X32 FILLER_503_1392 ();
 FILLCELL_X32 FILLER_503_1424 ();
 FILLCELL_X32 FILLER_503_1456 ();
 FILLCELL_X32 FILLER_503_1488 ();
 FILLCELL_X32 FILLER_503_1520 ();
 FILLCELL_X32 FILLER_503_1552 ();
 FILLCELL_X32 FILLER_503_1584 ();
 FILLCELL_X32 FILLER_503_1616 ();
 FILLCELL_X32 FILLER_503_1648 ();
 FILLCELL_X32 FILLER_503_1680 ();
 FILLCELL_X32 FILLER_503_1712 ();
 FILLCELL_X32 FILLER_503_1744 ();
 FILLCELL_X32 FILLER_503_1776 ();
 FILLCELL_X32 FILLER_503_1808 ();
 FILLCELL_X32 FILLER_503_1840 ();
 FILLCELL_X32 FILLER_503_1872 ();
 FILLCELL_X32 FILLER_503_1904 ();
 FILLCELL_X32 FILLER_503_1936 ();
 FILLCELL_X32 FILLER_503_1968 ();
 FILLCELL_X32 FILLER_503_2000 ();
 FILLCELL_X32 FILLER_503_2032 ();
 FILLCELL_X32 FILLER_503_2064 ();
 FILLCELL_X32 FILLER_503_2096 ();
 FILLCELL_X32 FILLER_503_2128 ();
 FILLCELL_X32 FILLER_503_2160 ();
 FILLCELL_X32 FILLER_503_2192 ();
 FILLCELL_X32 FILLER_503_2224 ();
 FILLCELL_X32 FILLER_503_2256 ();
 FILLCELL_X32 FILLER_503_2288 ();
 FILLCELL_X32 FILLER_503_2320 ();
 FILLCELL_X32 FILLER_503_2352 ();
 FILLCELL_X32 FILLER_503_2384 ();
 FILLCELL_X32 FILLER_503_2416 ();
 FILLCELL_X32 FILLER_503_2448 ();
 FILLCELL_X32 FILLER_503_2480 ();
 FILLCELL_X8 FILLER_503_2512 ();
 FILLCELL_X4 FILLER_503_2520 ();
 FILLCELL_X2 FILLER_503_2524 ();
 FILLCELL_X32 FILLER_503_2527 ();
 FILLCELL_X32 FILLER_503_2559 ();
 FILLCELL_X32 FILLER_503_2591 ();
 FILLCELL_X32 FILLER_503_2623 ();
 FILLCELL_X32 FILLER_503_2655 ();
 FILLCELL_X32 FILLER_503_2687 ();
 FILLCELL_X32 FILLER_503_2719 ();
 FILLCELL_X32 FILLER_503_2751 ();
 FILLCELL_X32 FILLER_503_2783 ();
 FILLCELL_X32 FILLER_503_2815 ();
 FILLCELL_X32 FILLER_503_2847 ();
 FILLCELL_X32 FILLER_503_2879 ();
 FILLCELL_X32 FILLER_503_2911 ();
 FILLCELL_X32 FILLER_503_2943 ();
 FILLCELL_X32 FILLER_503_2975 ();
 FILLCELL_X32 FILLER_503_3007 ();
 FILLCELL_X32 FILLER_503_3039 ();
 FILLCELL_X32 FILLER_503_3071 ();
 FILLCELL_X32 FILLER_503_3103 ();
 FILLCELL_X32 FILLER_503_3135 ();
 FILLCELL_X32 FILLER_503_3167 ();
 FILLCELL_X32 FILLER_503_3199 ();
 FILLCELL_X32 FILLER_503_3231 ();
 FILLCELL_X32 FILLER_503_3263 ();
 FILLCELL_X32 FILLER_503_3295 ();
 FILLCELL_X32 FILLER_503_3327 ();
 FILLCELL_X32 FILLER_503_3359 ();
 FILLCELL_X32 FILLER_503_3391 ();
 FILLCELL_X32 FILLER_503_3423 ();
 FILLCELL_X32 FILLER_503_3455 ();
 FILLCELL_X32 FILLER_503_3487 ();
 FILLCELL_X32 FILLER_503_3519 ();
 FILLCELL_X32 FILLER_503_3551 ();
 FILLCELL_X32 FILLER_503_3583 ();
 FILLCELL_X32 FILLER_503_3615 ();
 FILLCELL_X32 FILLER_503_3647 ();
 FILLCELL_X32 FILLER_503_3679 ();
 FILLCELL_X16 FILLER_503_3711 ();
 FILLCELL_X8 FILLER_503_3727 ();
 FILLCELL_X2 FILLER_503_3735 ();
 FILLCELL_X1 FILLER_503_3737 ();
 FILLCELL_X32 FILLER_504_1 ();
 FILLCELL_X32 FILLER_504_33 ();
 FILLCELL_X32 FILLER_504_65 ();
 FILLCELL_X32 FILLER_504_97 ();
 FILLCELL_X32 FILLER_504_129 ();
 FILLCELL_X32 FILLER_504_161 ();
 FILLCELL_X32 FILLER_504_193 ();
 FILLCELL_X32 FILLER_504_225 ();
 FILLCELL_X32 FILLER_504_257 ();
 FILLCELL_X32 FILLER_504_289 ();
 FILLCELL_X32 FILLER_504_321 ();
 FILLCELL_X32 FILLER_504_353 ();
 FILLCELL_X32 FILLER_504_385 ();
 FILLCELL_X32 FILLER_504_417 ();
 FILLCELL_X32 FILLER_504_449 ();
 FILLCELL_X32 FILLER_504_481 ();
 FILLCELL_X32 FILLER_504_513 ();
 FILLCELL_X32 FILLER_504_545 ();
 FILLCELL_X32 FILLER_504_577 ();
 FILLCELL_X16 FILLER_504_609 ();
 FILLCELL_X4 FILLER_504_625 ();
 FILLCELL_X2 FILLER_504_629 ();
 FILLCELL_X32 FILLER_504_632 ();
 FILLCELL_X32 FILLER_504_664 ();
 FILLCELL_X32 FILLER_504_696 ();
 FILLCELL_X32 FILLER_504_728 ();
 FILLCELL_X32 FILLER_504_760 ();
 FILLCELL_X32 FILLER_504_792 ();
 FILLCELL_X32 FILLER_504_824 ();
 FILLCELL_X32 FILLER_504_856 ();
 FILLCELL_X32 FILLER_504_888 ();
 FILLCELL_X32 FILLER_504_920 ();
 FILLCELL_X32 FILLER_504_952 ();
 FILLCELL_X32 FILLER_504_984 ();
 FILLCELL_X32 FILLER_504_1016 ();
 FILLCELL_X32 FILLER_504_1048 ();
 FILLCELL_X32 FILLER_504_1080 ();
 FILLCELL_X32 FILLER_504_1112 ();
 FILLCELL_X32 FILLER_504_1144 ();
 FILLCELL_X32 FILLER_504_1176 ();
 FILLCELL_X32 FILLER_504_1208 ();
 FILLCELL_X32 FILLER_504_1240 ();
 FILLCELL_X32 FILLER_504_1272 ();
 FILLCELL_X32 FILLER_504_1304 ();
 FILLCELL_X32 FILLER_504_1336 ();
 FILLCELL_X32 FILLER_504_1368 ();
 FILLCELL_X32 FILLER_504_1400 ();
 FILLCELL_X32 FILLER_504_1432 ();
 FILLCELL_X32 FILLER_504_1464 ();
 FILLCELL_X32 FILLER_504_1496 ();
 FILLCELL_X32 FILLER_504_1528 ();
 FILLCELL_X32 FILLER_504_1560 ();
 FILLCELL_X32 FILLER_504_1592 ();
 FILLCELL_X32 FILLER_504_1624 ();
 FILLCELL_X32 FILLER_504_1656 ();
 FILLCELL_X32 FILLER_504_1688 ();
 FILLCELL_X32 FILLER_504_1720 ();
 FILLCELL_X32 FILLER_504_1752 ();
 FILLCELL_X32 FILLER_504_1784 ();
 FILLCELL_X32 FILLER_504_1816 ();
 FILLCELL_X32 FILLER_504_1848 ();
 FILLCELL_X8 FILLER_504_1880 ();
 FILLCELL_X4 FILLER_504_1888 ();
 FILLCELL_X2 FILLER_504_1892 ();
 FILLCELL_X32 FILLER_504_1895 ();
 FILLCELL_X32 FILLER_504_1927 ();
 FILLCELL_X32 FILLER_504_1959 ();
 FILLCELL_X32 FILLER_504_1991 ();
 FILLCELL_X32 FILLER_504_2023 ();
 FILLCELL_X32 FILLER_504_2055 ();
 FILLCELL_X32 FILLER_504_2087 ();
 FILLCELL_X32 FILLER_504_2119 ();
 FILLCELL_X32 FILLER_504_2151 ();
 FILLCELL_X32 FILLER_504_2183 ();
 FILLCELL_X32 FILLER_504_2215 ();
 FILLCELL_X32 FILLER_504_2247 ();
 FILLCELL_X32 FILLER_504_2279 ();
 FILLCELL_X32 FILLER_504_2311 ();
 FILLCELL_X32 FILLER_504_2343 ();
 FILLCELL_X32 FILLER_504_2375 ();
 FILLCELL_X32 FILLER_504_2407 ();
 FILLCELL_X32 FILLER_504_2439 ();
 FILLCELL_X32 FILLER_504_2471 ();
 FILLCELL_X32 FILLER_504_2503 ();
 FILLCELL_X32 FILLER_504_2535 ();
 FILLCELL_X32 FILLER_504_2567 ();
 FILLCELL_X32 FILLER_504_2599 ();
 FILLCELL_X32 FILLER_504_2631 ();
 FILLCELL_X32 FILLER_504_2663 ();
 FILLCELL_X32 FILLER_504_2695 ();
 FILLCELL_X32 FILLER_504_2727 ();
 FILLCELL_X32 FILLER_504_2759 ();
 FILLCELL_X32 FILLER_504_2791 ();
 FILLCELL_X32 FILLER_504_2823 ();
 FILLCELL_X32 FILLER_504_2855 ();
 FILLCELL_X32 FILLER_504_2887 ();
 FILLCELL_X32 FILLER_504_2919 ();
 FILLCELL_X32 FILLER_504_2951 ();
 FILLCELL_X32 FILLER_504_2983 ();
 FILLCELL_X32 FILLER_504_3015 ();
 FILLCELL_X32 FILLER_504_3047 ();
 FILLCELL_X32 FILLER_504_3079 ();
 FILLCELL_X32 FILLER_504_3111 ();
 FILLCELL_X8 FILLER_504_3143 ();
 FILLCELL_X4 FILLER_504_3151 ();
 FILLCELL_X2 FILLER_504_3155 ();
 FILLCELL_X32 FILLER_504_3158 ();
 FILLCELL_X32 FILLER_504_3190 ();
 FILLCELL_X32 FILLER_504_3222 ();
 FILLCELL_X32 FILLER_504_3254 ();
 FILLCELL_X32 FILLER_504_3286 ();
 FILLCELL_X32 FILLER_504_3318 ();
 FILLCELL_X32 FILLER_504_3350 ();
 FILLCELL_X32 FILLER_504_3382 ();
 FILLCELL_X32 FILLER_504_3414 ();
 FILLCELL_X32 FILLER_504_3446 ();
 FILLCELL_X32 FILLER_504_3478 ();
 FILLCELL_X32 FILLER_504_3510 ();
 FILLCELL_X32 FILLER_504_3542 ();
 FILLCELL_X32 FILLER_504_3574 ();
 FILLCELL_X32 FILLER_504_3606 ();
 FILLCELL_X32 FILLER_504_3638 ();
 FILLCELL_X32 FILLER_504_3670 ();
 FILLCELL_X32 FILLER_504_3702 ();
 FILLCELL_X4 FILLER_504_3734 ();
 FILLCELL_X32 FILLER_505_1 ();
 FILLCELL_X32 FILLER_505_33 ();
 FILLCELL_X32 FILLER_505_65 ();
 FILLCELL_X32 FILLER_505_97 ();
 FILLCELL_X32 FILLER_505_129 ();
 FILLCELL_X32 FILLER_505_161 ();
 FILLCELL_X32 FILLER_505_193 ();
 FILLCELL_X32 FILLER_505_225 ();
 FILLCELL_X32 FILLER_505_257 ();
 FILLCELL_X32 FILLER_505_289 ();
 FILLCELL_X32 FILLER_505_321 ();
 FILLCELL_X32 FILLER_505_353 ();
 FILLCELL_X32 FILLER_505_385 ();
 FILLCELL_X32 FILLER_505_417 ();
 FILLCELL_X32 FILLER_505_449 ();
 FILLCELL_X32 FILLER_505_481 ();
 FILLCELL_X32 FILLER_505_513 ();
 FILLCELL_X32 FILLER_505_545 ();
 FILLCELL_X32 FILLER_505_577 ();
 FILLCELL_X32 FILLER_505_609 ();
 FILLCELL_X32 FILLER_505_641 ();
 FILLCELL_X32 FILLER_505_673 ();
 FILLCELL_X32 FILLER_505_705 ();
 FILLCELL_X32 FILLER_505_737 ();
 FILLCELL_X32 FILLER_505_769 ();
 FILLCELL_X32 FILLER_505_801 ();
 FILLCELL_X32 FILLER_505_833 ();
 FILLCELL_X32 FILLER_505_865 ();
 FILLCELL_X32 FILLER_505_897 ();
 FILLCELL_X32 FILLER_505_929 ();
 FILLCELL_X32 FILLER_505_961 ();
 FILLCELL_X32 FILLER_505_993 ();
 FILLCELL_X32 FILLER_505_1025 ();
 FILLCELL_X32 FILLER_505_1057 ();
 FILLCELL_X32 FILLER_505_1089 ();
 FILLCELL_X32 FILLER_505_1121 ();
 FILLCELL_X32 FILLER_505_1153 ();
 FILLCELL_X32 FILLER_505_1185 ();
 FILLCELL_X32 FILLER_505_1217 ();
 FILLCELL_X8 FILLER_505_1249 ();
 FILLCELL_X4 FILLER_505_1257 ();
 FILLCELL_X2 FILLER_505_1261 ();
 FILLCELL_X32 FILLER_505_1264 ();
 FILLCELL_X32 FILLER_505_1296 ();
 FILLCELL_X32 FILLER_505_1328 ();
 FILLCELL_X32 FILLER_505_1360 ();
 FILLCELL_X32 FILLER_505_1392 ();
 FILLCELL_X32 FILLER_505_1424 ();
 FILLCELL_X32 FILLER_505_1456 ();
 FILLCELL_X32 FILLER_505_1488 ();
 FILLCELL_X32 FILLER_505_1520 ();
 FILLCELL_X32 FILLER_505_1552 ();
 FILLCELL_X32 FILLER_505_1584 ();
 FILLCELL_X32 FILLER_505_1616 ();
 FILLCELL_X16 FILLER_505_1648 ();
 FILLCELL_X8 FILLER_505_1664 ();
 FILLCELL_X4 FILLER_505_1672 ();
 FILLCELL_X1 FILLER_505_1676 ();
 FILLCELL_X32 FILLER_505_1680 ();
 FILLCELL_X32 FILLER_505_1712 ();
 FILLCELL_X16 FILLER_505_1744 ();
 FILLCELL_X4 FILLER_505_1760 ();
 FILLCELL_X32 FILLER_505_1767 ();
 FILLCELL_X32 FILLER_505_1799 ();
 FILLCELL_X32 FILLER_505_1831 ();
 FILLCELL_X32 FILLER_505_1863 ();
 FILLCELL_X32 FILLER_505_1895 ();
 FILLCELL_X32 FILLER_505_1927 ();
 FILLCELL_X32 FILLER_505_1959 ();
 FILLCELL_X32 FILLER_505_1991 ();
 FILLCELL_X32 FILLER_505_2023 ();
 FILLCELL_X32 FILLER_505_2055 ();
 FILLCELL_X32 FILLER_505_2087 ();
 FILLCELL_X32 FILLER_505_2119 ();
 FILLCELL_X32 FILLER_505_2151 ();
 FILLCELL_X32 FILLER_505_2183 ();
 FILLCELL_X32 FILLER_505_2215 ();
 FILLCELL_X32 FILLER_505_2247 ();
 FILLCELL_X32 FILLER_505_2279 ();
 FILLCELL_X32 FILLER_505_2311 ();
 FILLCELL_X32 FILLER_505_2343 ();
 FILLCELL_X32 FILLER_505_2375 ();
 FILLCELL_X32 FILLER_505_2407 ();
 FILLCELL_X32 FILLER_505_2439 ();
 FILLCELL_X32 FILLER_505_2471 ();
 FILLCELL_X16 FILLER_505_2503 ();
 FILLCELL_X4 FILLER_505_2519 ();
 FILLCELL_X2 FILLER_505_2523 ();
 FILLCELL_X1 FILLER_505_2525 ();
 FILLCELL_X32 FILLER_505_2527 ();
 FILLCELL_X32 FILLER_505_2559 ();
 FILLCELL_X32 FILLER_505_2591 ();
 FILLCELL_X32 FILLER_505_2623 ();
 FILLCELL_X32 FILLER_505_2655 ();
 FILLCELL_X32 FILLER_505_2687 ();
 FILLCELL_X32 FILLER_505_2719 ();
 FILLCELL_X32 FILLER_505_2751 ();
 FILLCELL_X32 FILLER_505_2783 ();
 FILLCELL_X32 FILLER_505_2815 ();
 FILLCELL_X32 FILLER_505_2847 ();
 FILLCELL_X32 FILLER_505_2879 ();
 FILLCELL_X32 FILLER_505_2911 ();
 FILLCELL_X32 FILLER_505_2943 ();
 FILLCELL_X32 FILLER_505_2975 ();
 FILLCELL_X32 FILLER_505_3007 ();
 FILLCELL_X32 FILLER_505_3039 ();
 FILLCELL_X32 FILLER_505_3071 ();
 FILLCELL_X32 FILLER_505_3103 ();
 FILLCELL_X32 FILLER_505_3135 ();
 FILLCELL_X32 FILLER_505_3167 ();
 FILLCELL_X32 FILLER_505_3199 ();
 FILLCELL_X32 FILLER_505_3231 ();
 FILLCELL_X32 FILLER_505_3263 ();
 FILLCELL_X32 FILLER_505_3295 ();
 FILLCELL_X32 FILLER_505_3327 ();
 FILLCELL_X32 FILLER_505_3359 ();
 FILLCELL_X32 FILLER_505_3391 ();
 FILLCELL_X32 FILLER_505_3423 ();
 FILLCELL_X32 FILLER_505_3455 ();
 FILLCELL_X32 FILLER_505_3487 ();
 FILLCELL_X32 FILLER_505_3519 ();
 FILLCELL_X32 FILLER_505_3551 ();
 FILLCELL_X32 FILLER_505_3583 ();
 FILLCELL_X32 FILLER_505_3615 ();
 FILLCELL_X32 FILLER_505_3647 ();
 FILLCELL_X32 FILLER_505_3679 ();
 FILLCELL_X16 FILLER_505_3711 ();
 FILLCELL_X8 FILLER_505_3727 ();
 FILLCELL_X2 FILLER_505_3735 ();
 FILLCELL_X1 FILLER_505_3737 ();
 FILLCELL_X32 FILLER_506_1 ();
 FILLCELL_X32 FILLER_506_33 ();
 FILLCELL_X32 FILLER_506_65 ();
 FILLCELL_X32 FILLER_506_97 ();
 FILLCELL_X32 FILLER_506_129 ();
 FILLCELL_X32 FILLER_506_161 ();
 FILLCELL_X32 FILLER_506_193 ();
 FILLCELL_X32 FILLER_506_225 ();
 FILLCELL_X32 FILLER_506_257 ();
 FILLCELL_X32 FILLER_506_289 ();
 FILLCELL_X32 FILLER_506_321 ();
 FILLCELL_X32 FILLER_506_353 ();
 FILLCELL_X32 FILLER_506_385 ();
 FILLCELL_X32 FILLER_506_417 ();
 FILLCELL_X32 FILLER_506_449 ();
 FILLCELL_X32 FILLER_506_481 ();
 FILLCELL_X32 FILLER_506_513 ();
 FILLCELL_X32 FILLER_506_545 ();
 FILLCELL_X32 FILLER_506_577 ();
 FILLCELL_X16 FILLER_506_609 ();
 FILLCELL_X4 FILLER_506_625 ();
 FILLCELL_X2 FILLER_506_629 ();
 FILLCELL_X32 FILLER_506_632 ();
 FILLCELL_X32 FILLER_506_664 ();
 FILLCELL_X32 FILLER_506_696 ();
 FILLCELL_X32 FILLER_506_728 ();
 FILLCELL_X32 FILLER_506_760 ();
 FILLCELL_X32 FILLER_506_792 ();
 FILLCELL_X32 FILLER_506_824 ();
 FILLCELL_X32 FILLER_506_856 ();
 FILLCELL_X32 FILLER_506_888 ();
 FILLCELL_X32 FILLER_506_920 ();
 FILLCELL_X32 FILLER_506_952 ();
 FILLCELL_X32 FILLER_506_984 ();
 FILLCELL_X32 FILLER_506_1016 ();
 FILLCELL_X32 FILLER_506_1048 ();
 FILLCELL_X32 FILLER_506_1080 ();
 FILLCELL_X32 FILLER_506_1112 ();
 FILLCELL_X32 FILLER_506_1144 ();
 FILLCELL_X32 FILLER_506_1176 ();
 FILLCELL_X32 FILLER_506_1208 ();
 FILLCELL_X16 FILLER_506_1240 ();
 FILLCELL_X4 FILLER_506_1256 ();
 FILLCELL_X2 FILLER_506_1260 ();
 FILLCELL_X32 FILLER_506_1263 ();
 FILLCELL_X32 FILLER_506_1295 ();
 FILLCELL_X32 FILLER_506_1327 ();
 FILLCELL_X32 FILLER_506_1359 ();
 FILLCELL_X32 FILLER_506_1391 ();
 FILLCELL_X32 FILLER_506_1423 ();
 FILLCELL_X32 FILLER_506_1455 ();
 FILLCELL_X32 FILLER_506_1487 ();
 FILLCELL_X32 FILLER_506_1519 ();
 FILLCELL_X32 FILLER_506_1551 ();
 FILLCELL_X32 FILLER_506_1583 ();
 FILLCELL_X32 FILLER_506_1615 ();
 FILLCELL_X16 FILLER_506_1647 ();
 FILLCELL_X8 FILLER_506_1663 ();
 FILLCELL_X4 FILLER_506_1671 ();
 FILLCELL_X2 FILLER_506_1675 ();
 FILLCELL_X32 FILLER_506_1680 ();
 FILLCELL_X32 FILLER_506_1712 ();
 FILLCELL_X16 FILLER_506_1744 ();
 FILLCELL_X8 FILLER_506_1760 ();
 FILLCELL_X32 FILLER_506_1771 ();
 FILLCELL_X32 FILLER_506_1803 ();
 FILLCELL_X32 FILLER_506_1835 ();
 FILLCELL_X16 FILLER_506_1867 ();
 FILLCELL_X4 FILLER_506_1883 ();
 FILLCELL_X2 FILLER_506_1890 ();
 FILLCELL_X1 FILLER_506_1892 ();
 FILLCELL_X32 FILLER_506_1894 ();
 FILLCELL_X32 FILLER_506_1926 ();
 FILLCELL_X32 FILLER_506_1958 ();
 FILLCELL_X32 FILLER_506_1990 ();
 FILLCELL_X32 FILLER_506_2022 ();
 FILLCELL_X32 FILLER_506_2054 ();
 FILLCELL_X32 FILLER_506_2086 ();
 FILLCELL_X32 FILLER_506_2118 ();
 FILLCELL_X32 FILLER_506_2150 ();
 FILLCELL_X32 FILLER_506_2182 ();
 FILLCELL_X32 FILLER_506_2214 ();
 FILLCELL_X32 FILLER_506_2246 ();
 FILLCELL_X32 FILLER_506_2278 ();
 FILLCELL_X32 FILLER_506_2310 ();
 FILLCELL_X32 FILLER_506_2342 ();
 FILLCELL_X32 FILLER_506_2374 ();
 FILLCELL_X32 FILLER_506_2406 ();
 FILLCELL_X32 FILLER_506_2438 ();
 FILLCELL_X32 FILLER_506_2470 ();
 FILLCELL_X16 FILLER_506_2502 ();
 FILLCELL_X4 FILLER_506_2518 ();
 FILLCELL_X2 FILLER_506_2522 ();
 FILLCELL_X32 FILLER_506_2525 ();
 FILLCELL_X32 FILLER_506_2557 ();
 FILLCELL_X32 FILLER_506_2589 ();
 FILLCELL_X32 FILLER_506_2621 ();
 FILLCELL_X32 FILLER_506_2653 ();
 FILLCELL_X32 FILLER_506_2685 ();
 FILLCELL_X32 FILLER_506_2717 ();
 FILLCELL_X32 FILLER_506_2749 ();
 FILLCELL_X32 FILLER_506_2781 ();
 FILLCELL_X32 FILLER_506_2813 ();
 FILLCELL_X32 FILLER_506_2845 ();
 FILLCELL_X32 FILLER_506_2877 ();
 FILLCELL_X32 FILLER_506_2909 ();
 FILLCELL_X32 FILLER_506_2941 ();
 FILLCELL_X32 FILLER_506_2973 ();
 FILLCELL_X32 FILLER_506_3005 ();
 FILLCELL_X32 FILLER_506_3037 ();
 FILLCELL_X32 FILLER_506_3069 ();
 FILLCELL_X32 FILLER_506_3101 ();
 FILLCELL_X16 FILLER_506_3133 ();
 FILLCELL_X4 FILLER_506_3149 ();
 FILLCELL_X2 FILLER_506_3153 ();
 FILLCELL_X32 FILLER_506_3156 ();
 FILLCELL_X32 FILLER_506_3188 ();
 FILLCELL_X32 FILLER_506_3220 ();
 FILLCELL_X32 FILLER_506_3252 ();
 FILLCELL_X32 FILLER_506_3284 ();
 FILLCELL_X32 FILLER_506_3316 ();
 FILLCELL_X32 FILLER_506_3348 ();
 FILLCELL_X32 FILLER_506_3380 ();
 FILLCELL_X32 FILLER_506_3412 ();
 FILLCELL_X32 FILLER_506_3444 ();
 FILLCELL_X32 FILLER_506_3476 ();
 FILLCELL_X32 FILLER_506_3508 ();
 FILLCELL_X32 FILLER_506_3540 ();
 FILLCELL_X32 FILLER_506_3572 ();
 FILLCELL_X32 FILLER_506_3604 ();
 FILLCELL_X32 FILLER_506_3636 ();
 FILLCELL_X32 FILLER_506_3668 ();
 FILLCELL_X32 FILLER_506_3700 ();
 FILLCELL_X4 FILLER_506_3732 ();
 FILLCELL_X2 FILLER_506_3736 ();
endmodule
