module configurable_brent_kung_adder (cin,
    cout,
    a,
    b,
    sum);
 input cin;
 output cout;
 input [31:0] a;
 input [31:0] b;
 output [31:0] sum;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _070_ (.I(net1),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _071_ (.I(net25),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_8 _072_ (.I(net33),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _073_ (.I(net57),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _074_ (.I(net65),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _075_ (.I(_006_),
    .ZN(net68));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _076_ (.I(_008_),
    .ZN(net69));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _077_ (.I(_010_),
    .ZN(net70));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _078_ (.I(_012_),
    .ZN(net71));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _079_ (.I(_014_),
    .ZN(net72));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _080_ (.I(_016_),
    .ZN(net73));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _081_ (.I(_018_),
    .ZN(net74));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _082_ (.I(_020_),
    .ZN(net75));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _083_ (.I(_022_),
    .ZN(net76));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _084_ (.I(_024_),
    .ZN(net77));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _085_ (.I(_027_),
    .ZN(net78));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _086_ (.I(_029_),
    .ZN(net79));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _087_ (.I(_031_),
    .ZN(net80));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _088_ (.I(_033_),
    .ZN(net81));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _089_ (.I(_035_),
    .ZN(net82));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _090_ (.I(_037_),
    .ZN(net83));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _091_ (.I(_039_),
    .ZN(net84));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 _092_ (.I(_041_),
    .ZN(net85));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _093_ (.I(_043_),
    .ZN(net86));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _094_ (.I(_045_),
    .ZN(net87));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _095_ (.I(_047_),
    .ZN(net88));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _096_ (.I(_049_),
    .ZN(net89));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _097_ (.I(_051_),
    .ZN(net90));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _098_ (.I(_056_),
    .ZN(net91));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _099_ (.I(_058_),
    .ZN(net92));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _100_ (.I(_060_),
    .ZN(net93));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _101_ (.I(_062_),
    .ZN(net94));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _102_ (.I(_064_),
    .ZN(net95));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _103_ (.I(_066_),
    .ZN(net96));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _104_ (.I(_068_),
    .ZN(net97));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _105_ (.I(_069_),
    .ZN(net98));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _106_ (.I(_050_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _107_ (.I(_055_),
    .ZN(net66));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _108_ (.I(_003_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _109_ (.A(_000_),
    .B(_001_),
    .CI(_002_),
    .CO(_003_),
    .S(net67));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _110_ (.A(net2),
    .B(net34),
    .CI(_004_),
    .CO(_005_),
    .S(_006_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _111_ (.A(net3),
    .B(net35),
    .CI(_005_),
    .CO(_007_),
    .S(_008_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _112_ (.A(net4),
    .B(net36),
    .CI(_007_),
    .CO(_009_),
    .S(_010_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _113_ (.A(net5),
    .B(net37),
    .CI(_009_),
    .CO(_011_),
    .S(_012_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _114_ (.A(net6),
    .B(net38),
    .CI(_011_),
    .CO(_013_),
    .S(_014_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _115_ (.A(net7),
    .B(net39),
    .CI(_013_),
    .CO(_015_),
    .S(_016_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _116_ (.A(net8),
    .B(net40),
    .CI(_015_),
    .CO(_017_),
    .S(_018_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _117_ (.A(net9),
    .B(net41),
    .CI(_017_),
    .CO(_019_),
    .S(_020_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _118_ (.A(net10),
    .B(net42),
    .CI(_019_),
    .CO(_021_),
    .S(_022_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _119_ (.A(net11),
    .B(net43),
    .CI(_021_),
    .CO(_023_),
    .S(_024_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _120_ (.A(net12),
    .B(net44),
    .CI(_025_),
    .CO(_026_),
    .S(_027_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _121_ (.A(net13),
    .B(net45),
    .CI(_023_),
    .CO(_028_),
    .S(_029_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _122_ (.A(net14),
    .B(net46),
    .CI(_028_),
    .CO(_030_),
    .S(_031_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _123_ (.A(net15),
    .B(net47),
    .CI(_030_),
    .CO(_032_),
    .S(_033_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _124_ (.A(net16),
    .B(net48),
    .CI(_032_),
    .CO(_034_),
    .S(_035_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _125_ (.A(net17),
    .B(net49),
    .CI(_034_),
    .CO(_036_),
    .S(_037_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _126_ (.A(net18),
    .B(net50),
    .CI(_036_),
    .CO(_038_),
    .S(_039_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _127_ (.A(net19),
    .B(net51),
    .CI(_038_),
    .CO(_040_),
    .S(_041_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _128_ (.A(net20),
    .B(net52),
    .CI(_040_),
    .CO(_042_),
    .S(_043_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _129_ (.A(net21),
    .B(net53),
    .CI(_042_),
    .CO(_044_),
    .S(_045_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _130_ (.A(net22),
    .B(net54),
    .CI(_044_),
    .CO(_046_),
    .S(_047_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _131_ (.A(net23),
    .B(net55),
    .CI(_026_),
    .CO(_048_),
    .S(_049_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _132_ (.A(net24),
    .B(net56),
    .CI(_046_),
    .CO(_050_),
    .S(_051_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _133_ (.A(_052_),
    .B(_053_),
    .CI(_054_),
    .CO(_055_),
    .S(_056_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _134_ (.A(net26),
    .B(net58),
    .CI(_048_),
    .CO(_057_),
    .S(_058_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _135_ (.A(net27),
    .B(net59),
    .CI(_057_),
    .CO(_059_),
    .S(_060_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _136_ (.A(net28),
    .B(net60),
    .CI(_059_),
    .CO(_061_),
    .S(_062_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _137_ (.A(net29),
    .B(net61),
    .CI(_061_),
    .CO(_063_),
    .S(_064_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _138_ (.A(net30),
    .B(net62),
    .CI(_063_),
    .CO(_065_),
    .S(_066_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _139_ (.A(net31),
    .B(net63),
    .CI(_065_),
    .CO(_067_),
    .S(_068_));
 gf180mcu_fd_sc_mcu9t5v0__addf_2 _140_ (.A(net32),
    .B(net64),
    .CI(_067_),
    .CO(_004_),
    .S(_069_));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_65 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_66 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_67 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_68 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_69 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_70 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_71 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_72 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_73 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_74 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_75 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_76 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_77 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_78 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_79 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_80 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_81 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_82 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_83 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_84 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_85 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_86 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_87 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_88 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_89 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_90 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_91 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_27_Left_92 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_28_Left_93 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_29_Left_94 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_30_Left_95 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_31_Left_96 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_32_Left_97 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_33_Left_98 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_34_Left_99 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_35_Left_100 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_36_Left_101 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_37_Left_102 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_38_Left_103 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_39_Left_104 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_40_Left_105 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_41_Left_106 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_42_Left_107 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_43_Left_108 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_44_Left_109 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_45_Left_110 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_46_Left_111 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_47_Left_112 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_48_Left_113 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_49_Left_114 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_50_Left_115 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_51_Left_116 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_52_Left_117 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_53_Left_118 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_54_Left_119 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_55_Left_120 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_56_Left_121 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_57_Left_122 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_58_Left_123 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_59_Left_124 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_60_Left_125 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_61_Left_126 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_62_Left_127 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_63_Left_128 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_64_Left_129 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_131 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_132 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_1_133 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_134 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_135 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_3_136 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_137 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_138 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_5_139 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_140 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_141 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_7_142 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_143 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_144 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_9_145 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_146 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_147 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_11_148 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_149 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_150 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_13_151 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_152 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_153 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_15_154 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_155 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_156 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_17_157 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_158 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_159 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_19_160 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_161 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_21_163 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_164 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_165 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_23_166 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_167 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_168 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_169 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_170 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_171 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_27_172 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_173 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_28_174 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_29_175 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_176 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_30_177 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_31_178 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_179 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_33_181 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_182 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_34_183 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_35_184 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_185 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_36_186 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_37_187 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_188 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_38_189 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_39_190 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_191 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_40_192 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_41_193 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_194 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_42_195 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_43_196 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_197 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_44_198 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_45_199 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_200 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_46_201 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_47_202 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_203 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_48_204 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_49_205 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_206 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_50_207 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_51_208 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_209 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_52_210 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_53_211 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_212 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_54_213 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_55_214 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_215 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_56_216 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_57_217 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_218 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_58_219 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_59_220 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_221 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_60_222 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_61_223 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_224 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_62_225 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_63_226 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_227 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_228 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_64_229 ();
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 input1 (.I(a[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(a[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(a[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(a[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(a[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(a[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input7 (.I(a[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlya_2 input8 (.I(a[16]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(a[17]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(a[18]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input11 (.I(a[19]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input12 (.I(a[1]),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input13 (.I(a[20]),
    .Z(net13));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input14 (.I(a[21]),
    .Z(net14));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input15 (.I(a[22]),
    .Z(net15));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input16 (.I(a[23]),
    .Z(net16));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input17 (.I(a[24]),
    .Z(net17));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input18 (.I(a[25]),
    .Z(net18));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input19 (.I(a[26]),
    .Z(net19));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input20 (.I(a[27]),
    .Z(net20));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input21 (.I(a[28]),
    .Z(net21));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input22 (.I(a[29]),
    .Z(net22));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input23 (.I(a[2]),
    .Z(net23));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input24 (.I(a[30]),
    .Z(net24));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input25 (.I(a[31]),
    .Z(net25));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input26 (.I(a[3]),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input27 (.I(a[4]),
    .Z(net27));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input28 (.I(a[5]),
    .Z(net28));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input29 (.I(a[6]),
    .Z(net29));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input30 (.I(a[7]),
    .Z(net30));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input31 (.I(a[8]),
    .Z(net31));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input32 (.I(a[9]),
    .Z(net32));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 input33 (.I(b[0]),
    .Z(net33));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input34 (.I(b[10]),
    .Z(net34));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input35 (.I(b[11]),
    .Z(net35));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input36 (.I(b[12]),
    .Z(net36));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input37 (.I(b[13]),
    .Z(net37));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input38 (.I(b[14]),
    .Z(net38));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input39 (.I(b[15]),
    .Z(net39));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input40 (.I(b[16]),
    .Z(net40));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input41 (.I(b[17]),
    .Z(net41));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input42 (.I(b[18]),
    .Z(net42));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input43 (.I(b[19]),
    .Z(net43));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input44 (.I(b[1]),
    .Z(net44));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input45 (.I(b[20]),
    .Z(net45));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input46 (.I(b[21]),
    .Z(net46));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input47 (.I(b[22]),
    .Z(net47));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input48 (.I(b[23]),
    .Z(net48));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input49 (.I(b[24]),
    .Z(net49));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input50 (.I(b[25]),
    .Z(net50));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input51 (.I(b[26]),
    .Z(net51));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input52 (.I(b[27]),
    .Z(net52));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input53 (.I(b[28]),
    .Z(net53));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input54 (.I(b[29]),
    .Z(net54));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input55 (.I(b[2]),
    .Z(net55));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input56 (.I(b[30]),
    .Z(net56));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input57 (.I(b[31]),
    .Z(net57));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input58 (.I(b[3]),
    .Z(net58));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input59 (.I(b[4]),
    .Z(net59));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input60 (.I(b[5]),
    .Z(net60));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input61 (.I(b[6]),
    .Z(net61));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input62 (.I(b[7]),
    .Z(net62));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input63 (.I(b[8]),
    .Z(net63));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input64 (.I(b[9]),
    .Z(net64));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 input65 (.I(cin),
    .Z(net65));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 output66 (.I(net66),
    .Z(cout));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output67 (.I(net67),
    .Z(sum[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output68 (.I(net68),
    .Z(sum[10]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output69 (.I(net69),
    .Z(sum[11]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output70 (.I(net70),
    .Z(sum[12]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output71 (.I(net71),
    .Z(sum[13]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output72 (.I(net72),
    .Z(sum[14]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output73 (.I(net73),
    .Z(sum[15]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output74 (.I(net74),
    .Z(sum[16]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output75 (.I(net75),
    .Z(sum[17]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output76 (.I(net76),
    .Z(sum[18]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output77 (.I(net77),
    .Z(sum[19]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output78 (.I(net78),
    .Z(sum[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output79 (.I(net79),
    .Z(sum[20]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output80 (.I(net80),
    .Z(sum[21]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output81 (.I(net81),
    .Z(sum[22]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output82 (.I(net82),
    .Z(sum[23]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output83 (.I(net83),
    .Z(sum[24]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output84 (.I(net84),
    .Z(sum[25]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output85 (.I(net85),
    .Z(sum[26]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output86 (.I(net86),
    .Z(sum[27]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output87 (.I(net87),
    .Z(sum[28]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 output88 (.I(net88),
    .Z(sum[29]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output89 (.I(net89),
    .Z(sum[2]));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 output90 (.I(net90),
    .Z(sum[30]));
 gf180mcu_fd_sc_mcu9t5v0__buf_2 output91 (.I(net91),
    .Z(sum[31]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output92 (.I(net92),
    .Z(sum[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output93 (.I(net93),
    .Z(sum[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output94 (.I(net94),
    .Z(sum[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output95 (.I(net95),
    .Z(sum[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output96 (.I(net96),
    .Z(sum[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output97 (.I(net97),
    .Z(sum[8]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output98 (.I(net98),
    .Z(sum[9]));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_342 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_154 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_299 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_331 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_347 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_293 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_357 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_421 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_485 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_218 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_222 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_262 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_313 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_345 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_261 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_453 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_517 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_269 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_349 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_417 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_481 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_529 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_7_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_8_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_9_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_10_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_14_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_15_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_16_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_18_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_19_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_22_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_24_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_13 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_25 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_26_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_27_338 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_27_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_27_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_27_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_27_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_27_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_28_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_28_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_28_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_28_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_28_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_28_560 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_28_564 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_29_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_302 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_334 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_29_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_29_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_29_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_29_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_29_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_29_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_30_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_30_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_30_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_30_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_30_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_30_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_30_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_57 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_272 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_336 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_31_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_31_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_31_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_31_534 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_31_538 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_31_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_32_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_32_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_32_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_32_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_32_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_32_561 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_33_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_33_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_312 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_344 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_33_352 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_33_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_33_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_33_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_33_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_34_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_287 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_34_415 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_479 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_487 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_34_491 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_493 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_34_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_34_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_34_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_548 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_34_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_35_348 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_35_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_35_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_35_518 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_35_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_35_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_35_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_8 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_17 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_41 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_45 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_36_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_310 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_374 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_36_438 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_36_502 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_36_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_544 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_559 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_563 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_565 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_36_581 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_36_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_36_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_33 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_289 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_353 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_37_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_37_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_558 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_37_574 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_37_578 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_37_580 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_38_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_38_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_38_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_552 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_569 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_38_589 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_38_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_38_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_39_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_39_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_39_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_39_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_39_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_40_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_40_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_40_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_40_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_40_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_40_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_41_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_41_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_41_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_41_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_41_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_42_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_42_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_42_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_42_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_42_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_42_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_43_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_43_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_43_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_43_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_43_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_44_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_44_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_44_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_44_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_44_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_44_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_45_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_45_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_45_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_45_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_45_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_46_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_46_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_46_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_46_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_46_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_47_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_47_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_47_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_47_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_47_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_48_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_48_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_48_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_48_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_48_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_48_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_49_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_49_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_49_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_49_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_49_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_50_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_50_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_50_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_50_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_50_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_50_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_51_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_51_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_51_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_51_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_51_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_52_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_52_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_52_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_52_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_52_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_53_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_53_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_53_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_53_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_53_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_54_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_54_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_54_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_54_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_54_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_55_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_55_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_55_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_55_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_55_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_56_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_56_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_56_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_56_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_56_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_56_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_57_486 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_57_550 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_57_582 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_57_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_57_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_58_436 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_500 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_58_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_58_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_58_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_58_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_58_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_322 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_59_373 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_389 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_59_391 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_398 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_462 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_59_526 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_59_590 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_59_594 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_308 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_325 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_333 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_337 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_423 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_431 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_60_433 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_60_468 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_60_532 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_60_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_60_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_60_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_60_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_61_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_324 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_61_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_358 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_61_409 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_426 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_440 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_61_504 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_61_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_61_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_61_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_372 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_412 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_420 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_62_455 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_519 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_62_533 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_62_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_62_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_62_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_62_592 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_258 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_63_274 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_282 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_316 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_63_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_449 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_63_513 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_63_577 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_63_593 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_63_595 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_276 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_284 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_311 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_351 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_64_355 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_448 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_64_470 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_64_536 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_64_568 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_64_584 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_64_592 ();
endmodule
