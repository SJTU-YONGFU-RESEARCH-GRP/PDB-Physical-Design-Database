module configurable_comparator (result,
    signed_mode,
    a,
    b,
    op_sel);
 output result;
 input signed_mode;
 input [15:0] a;
 input [15:0] b;
 input [2:0] op_sel;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;

 INV_X1 _086_ (.A(net1),
    .ZN(_083_));
 INV_X1 _087_ (.A(net23),
    .ZN(_038_));
 INV_X1 _088_ (.A(net22),
    .ZN(_041_));
 INV_X1 _089_ (.A(net21),
    .ZN(_044_));
 INV_X1 _090_ (.A(net20),
    .ZN(_047_));
 INV_X1 _091_ (.A(net19),
    .ZN(_050_));
 INV_X1 _092_ (.A(net18),
    .ZN(_053_));
 INV_X1 _093_ (.A(net32),
    .ZN(_056_));
 INV_X1 _094_ (.A(net31),
    .ZN(_059_));
 INV_X1 _095_ (.A(net30),
    .ZN(_062_));
 INV_X1 _096_ (.A(net29),
    .ZN(_065_));
 INV_X1 _097_ (.A(net28),
    .ZN(_068_));
 INV_X1 _098_ (.A(net27),
    .ZN(_071_));
 INV_X1 _099_ (.A(net26),
    .ZN(_074_));
 INV_X1 _100_ (.A(net25),
    .ZN(_077_));
 INV_X1 _101_ (.A(net24),
    .ZN(_080_));
 INV_X1 _102_ (.A(net33),
    .ZN(_024_));
 NAND4_X4 _103_ (.A1(_040_),
    .A2(_043_),
    .A3(_046_),
    .A4(_049_),
    .ZN(_025_));
 NAND4_X4 _104_ (.A1(_052_),
    .A2(_058_),
    .A3(_055_),
    .A4(_061_),
    .ZN(_026_));
 NAND4_X2 _105_ (.A1(_064_),
    .A2(_067_),
    .A3(_070_),
    .A4(_073_),
    .ZN(_027_));
 NAND4_X4 _106_ (.A1(_076_),
    .A2(_085_),
    .A3(_082_),
    .A4(_079_),
    .ZN(_028_));
 NOR4_X4 _107_ (.A1(_025_),
    .A2(_026_),
    .A3(_027_),
    .A4(_028_),
    .ZN(_029_));
 XNOR2_X1 _108_ (.A(_024_),
    .B(_029_),
    .ZN(_030_));
 NOR3_X1 _109_ (.A1(net35),
    .A2(net34),
    .A3(_030_),
    .ZN(_031_));
 AOI21_X1 _110_ (.A(_031_),
    .B1(net34),
    .B2(net35),
    .ZN(_032_));
 NAND2_X1 _111_ (.A1(net33),
    .A2(_029_),
    .ZN(_033_));
 NAND2_X1 _112_ (.A1(net34),
    .A2(_033_),
    .ZN(_034_));
 NOR2_X1 _113_ (.A1(_025_),
    .A2(_026_),
    .ZN(_035_));
 AOI21_X2 _114_ (.A(_063_),
    .B1(_066_),
    .B2(_064_),
    .ZN(_036_));
 AOI21_X2 _115_ (.A(_069_),
    .B1(_072_),
    .B2(_070_),
    .ZN(_037_));
 NAND2_X1 _116_ (.A1(_064_),
    .A2(_067_),
    .ZN(_000_));
 OAI21_X1 _117_ (.A(_036_),
    .B1(_037_),
    .B2(_000_),
    .ZN(_001_));
 NAND3_X1 _118_ (.A1(_043_),
    .A2(_046_),
    .A3(_048_),
    .ZN(_002_));
 AOI21_X2 _119_ (.A(_042_),
    .B1(_045_),
    .B2(_043_),
    .ZN(_003_));
 NAND2_X1 _120_ (.A1(_002_),
    .A2(_003_),
    .ZN(_004_));
 AOI221_X2 _121_ (.A(_039_),
    .B1(_035_),
    .B2(_001_),
    .C1(_004_),
    .C2(_040_),
    .ZN(_005_));
 INV_X1 _122_ (.A(_025_),
    .ZN(_006_));
 AOI21_X1 _123_ (.A(_051_),
    .B1(_054_),
    .B2(_052_),
    .ZN(_007_));
 NAND2_X1 _124_ (.A1(_052_),
    .A2(_055_),
    .ZN(_008_));
 AOI21_X1 _125_ (.A(_057_),
    .B1(_060_),
    .B2(_058_),
    .ZN(_009_));
 OAI21_X2 _126_ (.A(_007_),
    .B1(_008_),
    .B2(_009_),
    .ZN(_010_));
 NAND2_X1 _127_ (.A1(_006_),
    .A2(_010_),
    .ZN(_011_));
 AND2_X1 _128_ (.A1(_076_),
    .A2(_079_),
    .ZN(_012_));
 INV_X1 _129_ (.A(_081_),
    .ZN(_013_));
 INV_X1 _130_ (.A(_082_),
    .ZN(_014_));
 OAI21_X1 _131_ (.A(_013_),
    .B1(_084_),
    .B2(_014_),
    .ZN(_015_));
 AOI221_X2 _132_ (.A(_075_),
    .B1(_012_),
    .B2(_015_),
    .C1(_078_),
    .C2(_076_),
    .ZN(_016_));
 OR3_X1 _133_ (.A1(_025_),
    .A2(_026_),
    .A3(_027_),
    .ZN(_017_));
 OAI211_X2 _134_ (.A(_005_),
    .B(_011_),
    .C1(_016_),
    .C2(_017_),
    .ZN(_018_));
 INV_X1 _135_ (.A(net36),
    .ZN(_019_));
 NOR2_X1 _136_ (.A1(_040_),
    .A2(_019_),
    .ZN(_020_));
 XNOR2_X2 _137_ (.A(_018_),
    .B(_020_),
    .ZN(_021_));
 OAI21_X1 _138_ (.A(_032_),
    .B1(_034_),
    .B2(_021_),
    .ZN(_022_));
 MUX2_X1 _139_ (.A(_021_),
    .B(_024_),
    .S(_029_),
    .Z(_023_));
 AOI21_X1 _140_ (.A(_022_),
    .B1(_023_),
    .B2(net35),
    .ZN(net37));
 HA_X1 _141_ (.A(net7),
    .B(_038_),
    .CO(_039_),
    .S(_040_));
 HA_X1 _142_ (.A(net6),
    .B(_041_),
    .CO(_042_),
    .S(_043_));
 HA_X1 _143_ (.A(net5),
    .B(_044_),
    .CO(_045_),
    .S(_046_));
 HA_X1 _144_ (.A(net4),
    .B(_047_),
    .CO(_048_),
    .S(_049_));
 HA_X1 _145_ (.A(net3),
    .B(_050_),
    .CO(_051_),
    .S(_052_));
 HA_X1 _146_ (.A(net2),
    .B(_053_),
    .CO(_054_),
    .S(_055_));
 HA_X1 _147_ (.A(net16),
    .B(_056_),
    .CO(_057_),
    .S(_058_));
 HA_X1 _148_ (.A(net15),
    .B(_059_),
    .CO(_060_),
    .S(_061_));
 HA_X1 _149_ (.A(net14),
    .B(_062_),
    .CO(_063_),
    .S(_064_));
 HA_X1 _150_ (.A(net13),
    .B(_065_),
    .CO(_066_),
    .S(_067_));
 HA_X1 _151_ (.A(net12),
    .B(_068_),
    .CO(_069_),
    .S(_070_));
 HA_X1 _152_ (.A(net11),
    .B(_071_),
    .CO(_072_),
    .S(_073_));
 HA_X1 _153_ (.A(net10),
    .B(_074_),
    .CO(_075_),
    .S(_076_));
 HA_X1 _154_ (.A(net9),
    .B(_077_),
    .CO(_078_),
    .S(_079_));
 HA_X1 _155_ (.A(net8),
    .B(_080_),
    .CO(_081_),
    .S(_082_));
 HA_X1 _156_ (.A(_083_),
    .B(net17),
    .CO(_084_),
    .S(_085_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_213 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_214 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_215 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_216 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_217 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_218 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_219 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_220 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_221 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_222 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_223 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_224 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_225 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_226 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_227 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_228 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_229 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_230 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_231 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_232 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_233 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_234 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_235 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_236 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_237 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_238 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_239 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_240 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_241 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_242 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_243 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_244 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_245 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_246 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_247 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_248 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_249 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_250 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_251 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_252 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_253 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_254 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_255 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_256 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_257 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_258 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_259 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_260 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_261 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_262 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_263 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_264 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_265 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_266 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_267 ();
 BUF_X1 input1 (.A(a[0]),
    .Z(net1));
 BUF_X1 input2 (.A(a[10]),
    .Z(net2));
 BUF_X1 input3 (.A(a[11]),
    .Z(net3));
 BUF_X1 input4 (.A(a[12]),
    .Z(net4));
 BUF_X1 input5 (.A(a[13]),
    .Z(net5));
 BUF_X1 input6 (.A(a[14]),
    .Z(net6));
 BUF_X1 input7 (.A(a[15]),
    .Z(net7));
 BUF_X1 input8 (.A(a[1]),
    .Z(net8));
 BUF_X1 input9 (.A(a[2]),
    .Z(net9));
 BUF_X2 input10 (.A(a[3]),
    .Z(net10));
 BUF_X1 input11 (.A(a[4]),
    .Z(net11));
 BUF_X1 input12 (.A(a[5]),
    .Z(net12));
 BUF_X1 input13 (.A(a[6]),
    .Z(net13));
 BUF_X1 input14 (.A(a[7]),
    .Z(net14));
 BUF_X2 input15 (.A(a[8]),
    .Z(net15));
 BUF_X1 input16 (.A(a[9]),
    .Z(net16));
 BUF_X1 input17 (.A(b[0]),
    .Z(net17));
 BUF_X1 input18 (.A(b[10]),
    .Z(net18));
 BUF_X1 input19 (.A(b[11]),
    .Z(net19));
 BUF_X1 input20 (.A(b[12]),
    .Z(net20));
 BUF_X1 input21 (.A(b[13]),
    .Z(net21));
 BUF_X1 input22 (.A(b[14]),
    .Z(net22));
 BUF_X1 input23 (.A(b[15]),
    .Z(net23));
 BUF_X1 input24 (.A(b[1]),
    .Z(net24));
 BUF_X1 input25 (.A(b[2]),
    .Z(net25));
 BUF_X1 input26 (.A(b[3]),
    .Z(net26));
 BUF_X1 input27 (.A(b[4]),
    .Z(net27));
 BUF_X1 input28 (.A(b[5]),
    .Z(net28));
 BUF_X1 input29 (.A(b[6]),
    .Z(net29));
 BUF_X1 input30 (.A(b[7]),
    .Z(net30));
 BUF_X1 input31 (.A(b[8]),
    .Z(net31));
 BUF_X1 input32 (.A(b[9]),
    .Z(net32));
 BUF_X1 input33 (.A(op_sel[0]),
    .Z(net33));
 BUF_X1 input34 (.A(op_sel[1]),
    .Z(net34));
 BUF_X1 input35 (.A(op_sel[2]),
    .Z(net35));
 BUF_X1 input36 (.A(signed_mode),
    .Z(net36));
 BUF_X1 output37 (.A(net37),
    .Z(result));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X32 FILLER_0_257 ();
 FILLCELL_X32 FILLER_0_289 ();
 FILLCELL_X16 FILLER_0_321 ();
 FILLCELL_X8 FILLER_0_337 ();
 FILLCELL_X2 FILLER_0_350 ();
 FILLCELL_X1 FILLER_0_352 ();
 FILLCELL_X1 FILLER_0_356 ();
 FILLCELL_X2 FILLER_0_360 ();
 FILLCELL_X1 FILLER_0_362 ();
 FILLCELL_X1 FILLER_0_366 ();
 FILLCELL_X1 FILLER_0_370 ();
 FILLCELL_X1 FILLER_0_377 ();
 FILLCELL_X8 FILLER_0_381 ();
 FILLCELL_X2 FILLER_0_392 ();
 FILLCELL_X1 FILLER_0_394 ();
 FILLCELL_X32 FILLER_0_398 ();
 FILLCELL_X32 FILLER_0_430 ();
 FILLCELL_X32 FILLER_0_462 ();
 FILLCELL_X32 FILLER_0_494 ();
 FILLCELL_X32 FILLER_0_526 ();
 FILLCELL_X32 FILLER_0_558 ();
 FILLCELL_X32 FILLER_0_590 ();
 FILLCELL_X8 FILLER_0_622 ();
 FILLCELL_X1 FILLER_0_630 ();
 FILLCELL_X32 FILLER_0_632 ();
 FILLCELL_X32 FILLER_0_664 ();
 FILLCELL_X32 FILLER_0_696 ();
 FILLCELL_X32 FILLER_0_728 ();
 FILLCELL_X16 FILLER_0_760 ();
 FILLCELL_X8 FILLER_0_776 ();
 FILLCELL_X4 FILLER_0_784 ();
 FILLCELL_X2 FILLER_0_788 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X16 FILLER_1_321 ();
 FILLCELL_X4 FILLER_1_337 ();
 FILLCELL_X1 FILLER_1_341 ();
 FILLCELL_X4 FILLER_1_364 ();
 FILLCELL_X2 FILLER_1_368 ();
 FILLCELL_X1 FILLER_1_370 ();
 FILLCELL_X2 FILLER_1_373 ();
 FILLCELL_X4 FILLER_1_387 ();
 FILLCELL_X32 FILLER_1_403 ();
 FILLCELL_X32 FILLER_1_435 ();
 FILLCELL_X32 FILLER_1_467 ();
 FILLCELL_X32 FILLER_1_499 ();
 FILLCELL_X32 FILLER_1_531 ();
 FILLCELL_X32 FILLER_1_563 ();
 FILLCELL_X32 FILLER_1_595 ();
 FILLCELL_X32 FILLER_1_627 ();
 FILLCELL_X32 FILLER_1_659 ();
 FILLCELL_X32 FILLER_1_691 ();
 FILLCELL_X32 FILLER_1_723 ();
 FILLCELL_X32 FILLER_1_755 ();
 FILLCELL_X2 FILLER_1_787 ();
 FILLCELL_X1 FILLER_1_789 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X16 FILLER_2_321 ();
 FILLCELL_X8 FILLER_2_337 ();
 FILLCELL_X4 FILLER_2_345 ();
 FILLCELL_X2 FILLER_2_349 ();
 FILLCELL_X8 FILLER_2_358 ();
 FILLCELL_X4 FILLER_2_366 ();
 FILLCELL_X32 FILLER_2_380 ();
 FILLCELL_X32 FILLER_2_412 ();
 FILLCELL_X32 FILLER_2_444 ();
 FILLCELL_X32 FILLER_2_476 ();
 FILLCELL_X32 FILLER_2_508 ();
 FILLCELL_X32 FILLER_2_540 ();
 FILLCELL_X32 FILLER_2_572 ();
 FILLCELL_X16 FILLER_2_604 ();
 FILLCELL_X8 FILLER_2_620 ();
 FILLCELL_X2 FILLER_2_628 ();
 FILLCELL_X1 FILLER_2_630 ();
 FILLCELL_X32 FILLER_2_632 ();
 FILLCELL_X32 FILLER_2_664 ();
 FILLCELL_X32 FILLER_2_696 ();
 FILLCELL_X32 FILLER_2_728 ();
 FILLCELL_X16 FILLER_2_760 ();
 FILLCELL_X8 FILLER_2_776 ();
 FILLCELL_X4 FILLER_2_784 ();
 FILLCELL_X2 FILLER_2_788 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X16 FILLER_3_353 ();
 FILLCELL_X8 FILLER_3_369 ();
 FILLCELL_X1 FILLER_3_377 ();
 FILLCELL_X32 FILLER_3_385 ();
 FILLCELL_X32 FILLER_3_417 ();
 FILLCELL_X32 FILLER_3_449 ();
 FILLCELL_X32 FILLER_3_481 ();
 FILLCELL_X32 FILLER_3_513 ();
 FILLCELL_X32 FILLER_3_545 ();
 FILLCELL_X32 FILLER_3_577 ();
 FILLCELL_X32 FILLER_3_609 ();
 FILLCELL_X32 FILLER_3_641 ();
 FILLCELL_X32 FILLER_3_673 ();
 FILLCELL_X32 FILLER_3_705 ();
 FILLCELL_X32 FILLER_3_737 ();
 FILLCELL_X16 FILLER_3_769 ();
 FILLCELL_X4 FILLER_3_785 ();
 FILLCELL_X1 FILLER_3_789 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X16 FILLER_4_353 ();
 FILLCELL_X8 FILLER_4_369 ();
 FILLCELL_X2 FILLER_4_377 ();
 FILLCELL_X8 FILLER_4_386 ();
 FILLCELL_X32 FILLER_4_398 ();
 FILLCELL_X32 FILLER_4_430 ();
 FILLCELL_X32 FILLER_4_462 ();
 FILLCELL_X32 FILLER_4_494 ();
 FILLCELL_X32 FILLER_4_526 ();
 FILLCELL_X32 FILLER_4_558 ();
 FILLCELL_X32 FILLER_4_590 ();
 FILLCELL_X8 FILLER_4_622 ();
 FILLCELL_X1 FILLER_4_630 ();
 FILLCELL_X32 FILLER_4_632 ();
 FILLCELL_X32 FILLER_4_664 ();
 FILLCELL_X32 FILLER_4_696 ();
 FILLCELL_X32 FILLER_4_728 ();
 FILLCELL_X16 FILLER_4_760 ();
 FILLCELL_X8 FILLER_4_776 ();
 FILLCELL_X4 FILLER_4_784 ();
 FILLCELL_X2 FILLER_4_788 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X32 FILLER_5_321 ();
 FILLCELL_X32 FILLER_5_353 ();
 FILLCELL_X32 FILLER_5_403 ();
 FILLCELL_X32 FILLER_5_435 ();
 FILLCELL_X32 FILLER_5_467 ();
 FILLCELL_X32 FILLER_5_499 ();
 FILLCELL_X32 FILLER_5_531 ();
 FILLCELL_X32 FILLER_5_563 ();
 FILLCELL_X32 FILLER_5_595 ();
 FILLCELL_X32 FILLER_5_627 ();
 FILLCELL_X32 FILLER_5_659 ();
 FILLCELL_X32 FILLER_5_691 ();
 FILLCELL_X32 FILLER_5_723 ();
 FILLCELL_X32 FILLER_5_755 ();
 FILLCELL_X2 FILLER_5_787 ();
 FILLCELL_X1 FILLER_5_789 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X32 FILLER_6_257 ();
 FILLCELL_X32 FILLER_6_289 ();
 FILLCELL_X32 FILLER_6_321 ();
 FILLCELL_X32 FILLER_6_353 ();
 FILLCELL_X32 FILLER_6_385 ();
 FILLCELL_X4 FILLER_6_417 ();
 FILLCELL_X32 FILLER_6_431 ();
 FILLCELL_X32 FILLER_6_463 ();
 FILLCELL_X32 FILLER_6_495 ();
 FILLCELL_X32 FILLER_6_527 ();
 FILLCELL_X32 FILLER_6_559 ();
 FILLCELL_X32 FILLER_6_591 ();
 FILLCELL_X8 FILLER_6_623 ();
 FILLCELL_X32 FILLER_6_632 ();
 FILLCELL_X32 FILLER_6_664 ();
 FILLCELL_X32 FILLER_6_696 ();
 FILLCELL_X32 FILLER_6_728 ();
 FILLCELL_X16 FILLER_6_760 ();
 FILLCELL_X8 FILLER_6_776 ();
 FILLCELL_X4 FILLER_6_784 ();
 FILLCELL_X2 FILLER_6_788 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X32 FILLER_7_257 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X32 FILLER_7_321 ();
 FILLCELL_X32 FILLER_7_353 ();
 FILLCELL_X32 FILLER_7_385 ();
 FILLCELL_X32 FILLER_7_417 ();
 FILLCELL_X32 FILLER_7_449 ();
 FILLCELL_X32 FILLER_7_481 ();
 FILLCELL_X32 FILLER_7_513 ();
 FILLCELL_X32 FILLER_7_545 ();
 FILLCELL_X32 FILLER_7_577 ();
 FILLCELL_X32 FILLER_7_609 ();
 FILLCELL_X32 FILLER_7_641 ();
 FILLCELL_X32 FILLER_7_673 ();
 FILLCELL_X32 FILLER_7_705 ();
 FILLCELL_X32 FILLER_7_737 ();
 FILLCELL_X16 FILLER_7_769 ();
 FILLCELL_X4 FILLER_7_785 ();
 FILLCELL_X1 FILLER_7_789 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X32 FILLER_8_257 ();
 FILLCELL_X32 FILLER_8_289 ();
 FILLCELL_X32 FILLER_8_321 ();
 FILLCELL_X32 FILLER_8_353 ();
 FILLCELL_X32 FILLER_8_385 ();
 FILLCELL_X32 FILLER_8_417 ();
 FILLCELL_X32 FILLER_8_449 ();
 FILLCELL_X32 FILLER_8_481 ();
 FILLCELL_X32 FILLER_8_513 ();
 FILLCELL_X32 FILLER_8_545 ();
 FILLCELL_X32 FILLER_8_577 ();
 FILLCELL_X16 FILLER_8_609 ();
 FILLCELL_X4 FILLER_8_625 ();
 FILLCELL_X2 FILLER_8_629 ();
 FILLCELL_X32 FILLER_8_632 ();
 FILLCELL_X32 FILLER_8_664 ();
 FILLCELL_X32 FILLER_8_696 ();
 FILLCELL_X32 FILLER_8_728 ();
 FILLCELL_X16 FILLER_8_760 ();
 FILLCELL_X8 FILLER_8_776 ();
 FILLCELL_X4 FILLER_8_784 ();
 FILLCELL_X2 FILLER_8_788 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X32 FILLER_9_257 ();
 FILLCELL_X32 FILLER_9_289 ();
 FILLCELL_X32 FILLER_9_321 ();
 FILLCELL_X32 FILLER_9_353 ();
 FILLCELL_X32 FILLER_9_385 ();
 FILLCELL_X32 FILLER_9_417 ();
 FILLCELL_X32 FILLER_9_449 ();
 FILLCELL_X32 FILLER_9_481 ();
 FILLCELL_X32 FILLER_9_513 ();
 FILLCELL_X32 FILLER_9_545 ();
 FILLCELL_X32 FILLER_9_577 ();
 FILLCELL_X32 FILLER_9_609 ();
 FILLCELL_X32 FILLER_9_641 ();
 FILLCELL_X32 FILLER_9_673 ();
 FILLCELL_X32 FILLER_9_705 ();
 FILLCELL_X32 FILLER_9_737 ();
 FILLCELL_X16 FILLER_9_769 ();
 FILLCELL_X4 FILLER_9_785 ();
 FILLCELL_X1 FILLER_9_789 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X32 FILLER_10_257 ();
 FILLCELL_X32 FILLER_10_289 ();
 FILLCELL_X32 FILLER_10_321 ();
 FILLCELL_X32 FILLER_10_353 ();
 FILLCELL_X32 FILLER_10_385 ();
 FILLCELL_X32 FILLER_10_417 ();
 FILLCELL_X32 FILLER_10_449 ();
 FILLCELL_X32 FILLER_10_481 ();
 FILLCELL_X32 FILLER_10_513 ();
 FILLCELL_X32 FILLER_10_545 ();
 FILLCELL_X32 FILLER_10_577 ();
 FILLCELL_X16 FILLER_10_609 ();
 FILLCELL_X4 FILLER_10_625 ();
 FILLCELL_X2 FILLER_10_629 ();
 FILLCELL_X32 FILLER_10_632 ();
 FILLCELL_X32 FILLER_10_664 ();
 FILLCELL_X32 FILLER_10_696 ();
 FILLCELL_X32 FILLER_10_728 ();
 FILLCELL_X16 FILLER_10_760 ();
 FILLCELL_X8 FILLER_10_776 ();
 FILLCELL_X4 FILLER_10_784 ();
 FILLCELL_X2 FILLER_10_788 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_257 ();
 FILLCELL_X32 FILLER_11_289 ();
 FILLCELL_X32 FILLER_11_321 ();
 FILLCELL_X32 FILLER_11_353 ();
 FILLCELL_X32 FILLER_11_385 ();
 FILLCELL_X32 FILLER_11_417 ();
 FILLCELL_X32 FILLER_11_449 ();
 FILLCELL_X32 FILLER_11_481 ();
 FILLCELL_X32 FILLER_11_513 ();
 FILLCELL_X32 FILLER_11_545 ();
 FILLCELL_X32 FILLER_11_577 ();
 FILLCELL_X32 FILLER_11_609 ();
 FILLCELL_X32 FILLER_11_641 ();
 FILLCELL_X32 FILLER_11_673 ();
 FILLCELL_X32 FILLER_11_705 ();
 FILLCELL_X32 FILLER_11_737 ();
 FILLCELL_X16 FILLER_11_769 ();
 FILLCELL_X4 FILLER_11_785 ();
 FILLCELL_X1 FILLER_11_789 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X32 FILLER_12_257 ();
 FILLCELL_X32 FILLER_12_289 ();
 FILLCELL_X32 FILLER_12_321 ();
 FILLCELL_X32 FILLER_12_353 ();
 FILLCELL_X32 FILLER_12_385 ();
 FILLCELL_X32 FILLER_12_417 ();
 FILLCELL_X32 FILLER_12_449 ();
 FILLCELL_X32 FILLER_12_481 ();
 FILLCELL_X32 FILLER_12_513 ();
 FILLCELL_X32 FILLER_12_545 ();
 FILLCELL_X32 FILLER_12_577 ();
 FILLCELL_X16 FILLER_12_609 ();
 FILLCELL_X4 FILLER_12_625 ();
 FILLCELL_X2 FILLER_12_629 ();
 FILLCELL_X32 FILLER_12_632 ();
 FILLCELL_X32 FILLER_12_664 ();
 FILLCELL_X32 FILLER_12_696 ();
 FILLCELL_X32 FILLER_12_728 ();
 FILLCELL_X16 FILLER_12_760 ();
 FILLCELL_X8 FILLER_12_776 ();
 FILLCELL_X4 FILLER_12_784 ();
 FILLCELL_X2 FILLER_12_788 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X32 FILLER_13_257 ();
 FILLCELL_X32 FILLER_13_289 ();
 FILLCELL_X32 FILLER_13_321 ();
 FILLCELL_X32 FILLER_13_353 ();
 FILLCELL_X32 FILLER_13_385 ();
 FILLCELL_X32 FILLER_13_417 ();
 FILLCELL_X32 FILLER_13_449 ();
 FILLCELL_X32 FILLER_13_481 ();
 FILLCELL_X32 FILLER_13_513 ();
 FILLCELL_X32 FILLER_13_545 ();
 FILLCELL_X32 FILLER_13_577 ();
 FILLCELL_X32 FILLER_13_609 ();
 FILLCELL_X32 FILLER_13_641 ();
 FILLCELL_X32 FILLER_13_673 ();
 FILLCELL_X32 FILLER_13_705 ();
 FILLCELL_X32 FILLER_13_737 ();
 FILLCELL_X16 FILLER_13_769 ();
 FILLCELL_X4 FILLER_13_785 ();
 FILLCELL_X1 FILLER_13_789 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X32 FILLER_14_257 ();
 FILLCELL_X32 FILLER_14_289 ();
 FILLCELL_X32 FILLER_14_321 ();
 FILLCELL_X32 FILLER_14_353 ();
 FILLCELL_X32 FILLER_14_385 ();
 FILLCELL_X32 FILLER_14_417 ();
 FILLCELL_X32 FILLER_14_449 ();
 FILLCELL_X32 FILLER_14_481 ();
 FILLCELL_X32 FILLER_14_513 ();
 FILLCELL_X32 FILLER_14_545 ();
 FILLCELL_X32 FILLER_14_577 ();
 FILLCELL_X16 FILLER_14_609 ();
 FILLCELL_X4 FILLER_14_625 ();
 FILLCELL_X2 FILLER_14_629 ();
 FILLCELL_X32 FILLER_14_632 ();
 FILLCELL_X32 FILLER_14_664 ();
 FILLCELL_X32 FILLER_14_696 ();
 FILLCELL_X32 FILLER_14_728 ();
 FILLCELL_X16 FILLER_14_760 ();
 FILLCELL_X8 FILLER_14_776 ();
 FILLCELL_X4 FILLER_14_784 ();
 FILLCELL_X2 FILLER_14_788 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X32 FILLER_15_257 ();
 FILLCELL_X32 FILLER_15_289 ();
 FILLCELL_X32 FILLER_15_321 ();
 FILLCELL_X32 FILLER_15_353 ();
 FILLCELL_X32 FILLER_15_385 ();
 FILLCELL_X32 FILLER_15_417 ();
 FILLCELL_X32 FILLER_15_449 ();
 FILLCELL_X32 FILLER_15_481 ();
 FILLCELL_X32 FILLER_15_513 ();
 FILLCELL_X32 FILLER_15_545 ();
 FILLCELL_X32 FILLER_15_577 ();
 FILLCELL_X32 FILLER_15_609 ();
 FILLCELL_X32 FILLER_15_641 ();
 FILLCELL_X32 FILLER_15_673 ();
 FILLCELL_X32 FILLER_15_705 ();
 FILLCELL_X32 FILLER_15_737 ();
 FILLCELL_X16 FILLER_15_769 ();
 FILLCELL_X4 FILLER_15_785 ();
 FILLCELL_X1 FILLER_15_789 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X32 FILLER_16_257 ();
 FILLCELL_X32 FILLER_16_289 ();
 FILLCELL_X32 FILLER_16_321 ();
 FILLCELL_X32 FILLER_16_353 ();
 FILLCELL_X32 FILLER_16_385 ();
 FILLCELL_X32 FILLER_16_417 ();
 FILLCELL_X32 FILLER_16_449 ();
 FILLCELL_X32 FILLER_16_481 ();
 FILLCELL_X32 FILLER_16_513 ();
 FILLCELL_X32 FILLER_16_545 ();
 FILLCELL_X32 FILLER_16_577 ();
 FILLCELL_X16 FILLER_16_609 ();
 FILLCELL_X4 FILLER_16_625 ();
 FILLCELL_X2 FILLER_16_629 ();
 FILLCELL_X32 FILLER_16_632 ();
 FILLCELL_X32 FILLER_16_664 ();
 FILLCELL_X32 FILLER_16_696 ();
 FILLCELL_X32 FILLER_16_728 ();
 FILLCELL_X16 FILLER_16_760 ();
 FILLCELL_X8 FILLER_16_776 ();
 FILLCELL_X4 FILLER_16_784 ();
 FILLCELL_X2 FILLER_16_788 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X32 FILLER_17_193 ();
 FILLCELL_X32 FILLER_17_225 ();
 FILLCELL_X32 FILLER_17_257 ();
 FILLCELL_X32 FILLER_17_289 ();
 FILLCELL_X32 FILLER_17_321 ();
 FILLCELL_X32 FILLER_17_353 ();
 FILLCELL_X32 FILLER_17_385 ();
 FILLCELL_X32 FILLER_17_417 ();
 FILLCELL_X32 FILLER_17_449 ();
 FILLCELL_X32 FILLER_17_481 ();
 FILLCELL_X32 FILLER_17_513 ();
 FILLCELL_X32 FILLER_17_545 ();
 FILLCELL_X32 FILLER_17_577 ();
 FILLCELL_X32 FILLER_17_609 ();
 FILLCELL_X32 FILLER_17_641 ();
 FILLCELL_X32 FILLER_17_673 ();
 FILLCELL_X32 FILLER_17_705 ();
 FILLCELL_X32 FILLER_17_737 ();
 FILLCELL_X16 FILLER_17_769 ();
 FILLCELL_X4 FILLER_17_785 ();
 FILLCELL_X1 FILLER_17_789 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X32 FILLER_18_225 ();
 FILLCELL_X32 FILLER_18_257 ();
 FILLCELL_X32 FILLER_18_289 ();
 FILLCELL_X32 FILLER_18_321 ();
 FILLCELL_X32 FILLER_18_353 ();
 FILLCELL_X32 FILLER_18_385 ();
 FILLCELL_X32 FILLER_18_417 ();
 FILLCELL_X32 FILLER_18_449 ();
 FILLCELL_X32 FILLER_18_481 ();
 FILLCELL_X32 FILLER_18_513 ();
 FILLCELL_X32 FILLER_18_545 ();
 FILLCELL_X32 FILLER_18_577 ();
 FILLCELL_X16 FILLER_18_609 ();
 FILLCELL_X4 FILLER_18_625 ();
 FILLCELL_X2 FILLER_18_629 ();
 FILLCELL_X32 FILLER_18_632 ();
 FILLCELL_X32 FILLER_18_664 ();
 FILLCELL_X32 FILLER_18_696 ();
 FILLCELL_X32 FILLER_18_728 ();
 FILLCELL_X16 FILLER_18_760 ();
 FILLCELL_X8 FILLER_18_776 ();
 FILLCELL_X4 FILLER_18_784 ();
 FILLCELL_X2 FILLER_18_788 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X32 FILLER_19_257 ();
 FILLCELL_X32 FILLER_19_289 ();
 FILLCELL_X32 FILLER_19_321 ();
 FILLCELL_X32 FILLER_19_353 ();
 FILLCELL_X32 FILLER_19_385 ();
 FILLCELL_X32 FILLER_19_417 ();
 FILLCELL_X32 FILLER_19_449 ();
 FILLCELL_X32 FILLER_19_481 ();
 FILLCELL_X32 FILLER_19_513 ();
 FILLCELL_X32 FILLER_19_545 ();
 FILLCELL_X32 FILLER_19_577 ();
 FILLCELL_X32 FILLER_19_609 ();
 FILLCELL_X32 FILLER_19_641 ();
 FILLCELL_X32 FILLER_19_673 ();
 FILLCELL_X32 FILLER_19_705 ();
 FILLCELL_X32 FILLER_19_737 ();
 FILLCELL_X16 FILLER_19_769 ();
 FILLCELL_X4 FILLER_19_785 ();
 FILLCELL_X1 FILLER_19_789 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X32 FILLER_20_225 ();
 FILLCELL_X32 FILLER_20_257 ();
 FILLCELL_X32 FILLER_20_289 ();
 FILLCELL_X32 FILLER_20_321 ();
 FILLCELL_X32 FILLER_20_353 ();
 FILLCELL_X32 FILLER_20_385 ();
 FILLCELL_X32 FILLER_20_417 ();
 FILLCELL_X32 FILLER_20_449 ();
 FILLCELL_X32 FILLER_20_481 ();
 FILLCELL_X32 FILLER_20_513 ();
 FILLCELL_X32 FILLER_20_545 ();
 FILLCELL_X32 FILLER_20_577 ();
 FILLCELL_X16 FILLER_20_609 ();
 FILLCELL_X4 FILLER_20_625 ();
 FILLCELL_X2 FILLER_20_629 ();
 FILLCELL_X32 FILLER_20_632 ();
 FILLCELL_X32 FILLER_20_664 ();
 FILLCELL_X32 FILLER_20_696 ();
 FILLCELL_X32 FILLER_20_728 ();
 FILLCELL_X16 FILLER_20_760 ();
 FILLCELL_X8 FILLER_20_776 ();
 FILLCELL_X4 FILLER_20_784 ();
 FILLCELL_X2 FILLER_20_788 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X32 FILLER_21_225 ();
 FILLCELL_X32 FILLER_21_257 ();
 FILLCELL_X32 FILLER_21_289 ();
 FILLCELL_X32 FILLER_21_321 ();
 FILLCELL_X32 FILLER_21_353 ();
 FILLCELL_X32 FILLER_21_385 ();
 FILLCELL_X32 FILLER_21_417 ();
 FILLCELL_X32 FILLER_21_449 ();
 FILLCELL_X32 FILLER_21_481 ();
 FILLCELL_X32 FILLER_21_513 ();
 FILLCELL_X32 FILLER_21_545 ();
 FILLCELL_X32 FILLER_21_577 ();
 FILLCELL_X32 FILLER_21_609 ();
 FILLCELL_X32 FILLER_21_641 ();
 FILLCELL_X32 FILLER_21_673 ();
 FILLCELL_X32 FILLER_21_705 ();
 FILLCELL_X32 FILLER_21_737 ();
 FILLCELL_X16 FILLER_21_769 ();
 FILLCELL_X4 FILLER_21_785 ();
 FILLCELL_X1 FILLER_21_789 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X32 FILLER_22_225 ();
 FILLCELL_X32 FILLER_22_257 ();
 FILLCELL_X32 FILLER_22_289 ();
 FILLCELL_X32 FILLER_22_321 ();
 FILLCELL_X32 FILLER_22_353 ();
 FILLCELL_X32 FILLER_22_385 ();
 FILLCELL_X32 FILLER_22_417 ();
 FILLCELL_X32 FILLER_22_449 ();
 FILLCELL_X32 FILLER_22_481 ();
 FILLCELL_X32 FILLER_22_513 ();
 FILLCELL_X32 FILLER_22_545 ();
 FILLCELL_X32 FILLER_22_577 ();
 FILLCELL_X16 FILLER_22_609 ();
 FILLCELL_X4 FILLER_22_625 ();
 FILLCELL_X2 FILLER_22_629 ();
 FILLCELL_X32 FILLER_22_632 ();
 FILLCELL_X32 FILLER_22_664 ();
 FILLCELL_X32 FILLER_22_696 ();
 FILLCELL_X32 FILLER_22_728 ();
 FILLCELL_X16 FILLER_22_760 ();
 FILLCELL_X8 FILLER_22_776 ();
 FILLCELL_X4 FILLER_22_784 ();
 FILLCELL_X2 FILLER_22_788 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X32 FILLER_23_225 ();
 FILLCELL_X32 FILLER_23_257 ();
 FILLCELL_X32 FILLER_23_289 ();
 FILLCELL_X32 FILLER_23_321 ();
 FILLCELL_X32 FILLER_23_353 ();
 FILLCELL_X32 FILLER_23_385 ();
 FILLCELL_X32 FILLER_23_417 ();
 FILLCELL_X32 FILLER_23_449 ();
 FILLCELL_X32 FILLER_23_481 ();
 FILLCELL_X32 FILLER_23_513 ();
 FILLCELL_X32 FILLER_23_545 ();
 FILLCELL_X32 FILLER_23_577 ();
 FILLCELL_X32 FILLER_23_609 ();
 FILLCELL_X32 FILLER_23_641 ();
 FILLCELL_X32 FILLER_23_673 ();
 FILLCELL_X32 FILLER_23_705 ();
 FILLCELL_X32 FILLER_23_737 ();
 FILLCELL_X16 FILLER_23_769 ();
 FILLCELL_X4 FILLER_23_785 ();
 FILLCELL_X1 FILLER_23_789 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X32 FILLER_24_225 ();
 FILLCELL_X32 FILLER_24_257 ();
 FILLCELL_X32 FILLER_24_289 ();
 FILLCELL_X32 FILLER_24_321 ();
 FILLCELL_X32 FILLER_24_353 ();
 FILLCELL_X32 FILLER_24_385 ();
 FILLCELL_X32 FILLER_24_417 ();
 FILLCELL_X32 FILLER_24_449 ();
 FILLCELL_X32 FILLER_24_481 ();
 FILLCELL_X32 FILLER_24_513 ();
 FILLCELL_X32 FILLER_24_545 ();
 FILLCELL_X32 FILLER_24_577 ();
 FILLCELL_X16 FILLER_24_609 ();
 FILLCELL_X4 FILLER_24_625 ();
 FILLCELL_X2 FILLER_24_629 ();
 FILLCELL_X32 FILLER_24_632 ();
 FILLCELL_X32 FILLER_24_664 ();
 FILLCELL_X32 FILLER_24_696 ();
 FILLCELL_X32 FILLER_24_728 ();
 FILLCELL_X16 FILLER_24_760 ();
 FILLCELL_X8 FILLER_24_776 ();
 FILLCELL_X4 FILLER_24_784 ();
 FILLCELL_X2 FILLER_24_788 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X32 FILLER_25_225 ();
 FILLCELL_X32 FILLER_25_257 ();
 FILLCELL_X32 FILLER_25_289 ();
 FILLCELL_X32 FILLER_25_321 ();
 FILLCELL_X32 FILLER_25_353 ();
 FILLCELL_X32 FILLER_25_385 ();
 FILLCELL_X32 FILLER_25_417 ();
 FILLCELL_X32 FILLER_25_449 ();
 FILLCELL_X32 FILLER_25_481 ();
 FILLCELL_X32 FILLER_25_513 ();
 FILLCELL_X32 FILLER_25_545 ();
 FILLCELL_X32 FILLER_25_577 ();
 FILLCELL_X32 FILLER_25_609 ();
 FILLCELL_X32 FILLER_25_641 ();
 FILLCELL_X32 FILLER_25_673 ();
 FILLCELL_X32 FILLER_25_705 ();
 FILLCELL_X32 FILLER_25_737 ();
 FILLCELL_X16 FILLER_25_769 ();
 FILLCELL_X4 FILLER_25_785 ();
 FILLCELL_X1 FILLER_25_789 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X32 FILLER_26_225 ();
 FILLCELL_X32 FILLER_26_257 ();
 FILLCELL_X32 FILLER_26_289 ();
 FILLCELL_X32 FILLER_26_321 ();
 FILLCELL_X32 FILLER_26_353 ();
 FILLCELL_X32 FILLER_26_385 ();
 FILLCELL_X32 FILLER_26_417 ();
 FILLCELL_X32 FILLER_26_449 ();
 FILLCELL_X32 FILLER_26_481 ();
 FILLCELL_X32 FILLER_26_513 ();
 FILLCELL_X32 FILLER_26_545 ();
 FILLCELL_X32 FILLER_26_577 ();
 FILLCELL_X16 FILLER_26_609 ();
 FILLCELL_X4 FILLER_26_625 ();
 FILLCELL_X2 FILLER_26_629 ();
 FILLCELL_X32 FILLER_26_632 ();
 FILLCELL_X32 FILLER_26_664 ();
 FILLCELL_X32 FILLER_26_696 ();
 FILLCELL_X32 FILLER_26_728 ();
 FILLCELL_X16 FILLER_26_760 ();
 FILLCELL_X8 FILLER_26_776 ();
 FILLCELL_X4 FILLER_26_784 ();
 FILLCELL_X2 FILLER_26_788 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X32 FILLER_27_225 ();
 FILLCELL_X32 FILLER_27_257 ();
 FILLCELL_X32 FILLER_27_289 ();
 FILLCELL_X32 FILLER_27_321 ();
 FILLCELL_X32 FILLER_27_353 ();
 FILLCELL_X32 FILLER_27_385 ();
 FILLCELL_X32 FILLER_27_417 ();
 FILLCELL_X32 FILLER_27_449 ();
 FILLCELL_X32 FILLER_27_481 ();
 FILLCELL_X32 FILLER_27_513 ();
 FILLCELL_X32 FILLER_27_545 ();
 FILLCELL_X32 FILLER_27_577 ();
 FILLCELL_X32 FILLER_27_609 ();
 FILLCELL_X32 FILLER_27_641 ();
 FILLCELL_X32 FILLER_27_673 ();
 FILLCELL_X32 FILLER_27_705 ();
 FILLCELL_X32 FILLER_27_737 ();
 FILLCELL_X16 FILLER_27_769 ();
 FILLCELL_X4 FILLER_27_785 ();
 FILLCELL_X1 FILLER_27_789 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X32 FILLER_28_257 ();
 FILLCELL_X32 FILLER_28_289 ();
 FILLCELL_X32 FILLER_28_321 ();
 FILLCELL_X32 FILLER_28_353 ();
 FILLCELL_X32 FILLER_28_385 ();
 FILLCELL_X32 FILLER_28_417 ();
 FILLCELL_X32 FILLER_28_449 ();
 FILLCELL_X32 FILLER_28_481 ();
 FILLCELL_X32 FILLER_28_513 ();
 FILLCELL_X32 FILLER_28_545 ();
 FILLCELL_X32 FILLER_28_577 ();
 FILLCELL_X16 FILLER_28_609 ();
 FILLCELL_X4 FILLER_28_625 ();
 FILLCELL_X2 FILLER_28_629 ();
 FILLCELL_X32 FILLER_28_632 ();
 FILLCELL_X32 FILLER_28_664 ();
 FILLCELL_X32 FILLER_28_696 ();
 FILLCELL_X32 FILLER_28_728 ();
 FILLCELL_X16 FILLER_28_760 ();
 FILLCELL_X8 FILLER_28_776 ();
 FILLCELL_X4 FILLER_28_784 ();
 FILLCELL_X2 FILLER_28_788 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X32 FILLER_29_257 ();
 FILLCELL_X32 FILLER_29_289 ();
 FILLCELL_X32 FILLER_29_321 ();
 FILLCELL_X32 FILLER_29_353 ();
 FILLCELL_X32 FILLER_29_385 ();
 FILLCELL_X32 FILLER_29_417 ();
 FILLCELL_X32 FILLER_29_449 ();
 FILLCELL_X32 FILLER_29_481 ();
 FILLCELL_X32 FILLER_29_513 ();
 FILLCELL_X32 FILLER_29_545 ();
 FILLCELL_X32 FILLER_29_577 ();
 FILLCELL_X32 FILLER_29_609 ();
 FILLCELL_X32 FILLER_29_641 ();
 FILLCELL_X32 FILLER_29_673 ();
 FILLCELL_X32 FILLER_29_705 ();
 FILLCELL_X32 FILLER_29_737 ();
 FILLCELL_X16 FILLER_29_769 ();
 FILLCELL_X4 FILLER_29_785 ();
 FILLCELL_X1 FILLER_29_789 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X32 FILLER_30_257 ();
 FILLCELL_X32 FILLER_30_289 ();
 FILLCELL_X32 FILLER_30_321 ();
 FILLCELL_X32 FILLER_30_353 ();
 FILLCELL_X32 FILLER_30_385 ();
 FILLCELL_X32 FILLER_30_417 ();
 FILLCELL_X32 FILLER_30_449 ();
 FILLCELL_X32 FILLER_30_481 ();
 FILLCELL_X32 FILLER_30_513 ();
 FILLCELL_X32 FILLER_30_545 ();
 FILLCELL_X32 FILLER_30_577 ();
 FILLCELL_X16 FILLER_30_609 ();
 FILLCELL_X4 FILLER_30_625 ();
 FILLCELL_X2 FILLER_30_629 ();
 FILLCELL_X32 FILLER_30_632 ();
 FILLCELL_X32 FILLER_30_664 ();
 FILLCELL_X32 FILLER_30_696 ();
 FILLCELL_X32 FILLER_30_728 ();
 FILLCELL_X16 FILLER_30_760 ();
 FILLCELL_X8 FILLER_30_776 ();
 FILLCELL_X4 FILLER_30_784 ();
 FILLCELL_X2 FILLER_30_788 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X32 FILLER_31_257 ();
 FILLCELL_X32 FILLER_31_289 ();
 FILLCELL_X32 FILLER_31_321 ();
 FILLCELL_X32 FILLER_31_353 ();
 FILLCELL_X32 FILLER_31_385 ();
 FILLCELL_X32 FILLER_31_417 ();
 FILLCELL_X32 FILLER_31_449 ();
 FILLCELL_X32 FILLER_31_481 ();
 FILLCELL_X32 FILLER_31_513 ();
 FILLCELL_X32 FILLER_31_545 ();
 FILLCELL_X32 FILLER_31_577 ();
 FILLCELL_X32 FILLER_31_609 ();
 FILLCELL_X32 FILLER_31_641 ();
 FILLCELL_X32 FILLER_31_673 ();
 FILLCELL_X32 FILLER_31_705 ();
 FILLCELL_X32 FILLER_31_737 ();
 FILLCELL_X16 FILLER_31_769 ();
 FILLCELL_X4 FILLER_31_785 ();
 FILLCELL_X1 FILLER_31_789 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X32 FILLER_32_289 ();
 FILLCELL_X32 FILLER_32_321 ();
 FILLCELL_X32 FILLER_32_353 ();
 FILLCELL_X32 FILLER_32_385 ();
 FILLCELL_X32 FILLER_32_417 ();
 FILLCELL_X32 FILLER_32_449 ();
 FILLCELL_X32 FILLER_32_481 ();
 FILLCELL_X32 FILLER_32_513 ();
 FILLCELL_X32 FILLER_32_545 ();
 FILLCELL_X32 FILLER_32_577 ();
 FILLCELL_X16 FILLER_32_609 ();
 FILLCELL_X4 FILLER_32_625 ();
 FILLCELL_X2 FILLER_32_629 ();
 FILLCELL_X32 FILLER_32_632 ();
 FILLCELL_X32 FILLER_32_664 ();
 FILLCELL_X32 FILLER_32_696 ();
 FILLCELL_X32 FILLER_32_728 ();
 FILLCELL_X16 FILLER_32_760 ();
 FILLCELL_X8 FILLER_32_776 ();
 FILLCELL_X4 FILLER_32_784 ();
 FILLCELL_X2 FILLER_32_788 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X32 FILLER_33_257 ();
 FILLCELL_X32 FILLER_33_289 ();
 FILLCELL_X32 FILLER_33_321 ();
 FILLCELL_X32 FILLER_33_353 ();
 FILLCELL_X32 FILLER_33_385 ();
 FILLCELL_X32 FILLER_33_417 ();
 FILLCELL_X32 FILLER_33_449 ();
 FILLCELL_X32 FILLER_33_481 ();
 FILLCELL_X32 FILLER_33_513 ();
 FILLCELL_X32 FILLER_33_545 ();
 FILLCELL_X32 FILLER_33_577 ();
 FILLCELL_X32 FILLER_33_609 ();
 FILLCELL_X32 FILLER_33_641 ();
 FILLCELL_X32 FILLER_33_673 ();
 FILLCELL_X32 FILLER_33_705 ();
 FILLCELL_X32 FILLER_33_737 ();
 FILLCELL_X16 FILLER_33_769 ();
 FILLCELL_X4 FILLER_33_785 ();
 FILLCELL_X1 FILLER_33_789 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X32 FILLER_34_257 ();
 FILLCELL_X32 FILLER_34_289 ();
 FILLCELL_X32 FILLER_34_321 ();
 FILLCELL_X32 FILLER_34_353 ();
 FILLCELL_X32 FILLER_34_385 ();
 FILLCELL_X32 FILLER_34_417 ();
 FILLCELL_X32 FILLER_34_449 ();
 FILLCELL_X32 FILLER_34_481 ();
 FILLCELL_X32 FILLER_34_513 ();
 FILLCELL_X32 FILLER_34_545 ();
 FILLCELL_X32 FILLER_34_577 ();
 FILLCELL_X16 FILLER_34_609 ();
 FILLCELL_X4 FILLER_34_625 ();
 FILLCELL_X2 FILLER_34_629 ();
 FILLCELL_X32 FILLER_34_632 ();
 FILLCELL_X32 FILLER_34_664 ();
 FILLCELL_X32 FILLER_34_696 ();
 FILLCELL_X32 FILLER_34_728 ();
 FILLCELL_X16 FILLER_34_760 ();
 FILLCELL_X8 FILLER_34_776 ();
 FILLCELL_X4 FILLER_34_784 ();
 FILLCELL_X2 FILLER_34_788 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X32 FILLER_35_97 ();
 FILLCELL_X32 FILLER_35_129 ();
 FILLCELL_X32 FILLER_35_161 ();
 FILLCELL_X32 FILLER_35_193 ();
 FILLCELL_X32 FILLER_35_225 ();
 FILLCELL_X32 FILLER_35_257 ();
 FILLCELL_X32 FILLER_35_289 ();
 FILLCELL_X32 FILLER_35_321 ();
 FILLCELL_X32 FILLER_35_353 ();
 FILLCELL_X32 FILLER_35_385 ();
 FILLCELL_X32 FILLER_35_417 ();
 FILLCELL_X32 FILLER_35_449 ();
 FILLCELL_X32 FILLER_35_481 ();
 FILLCELL_X32 FILLER_35_513 ();
 FILLCELL_X32 FILLER_35_545 ();
 FILLCELL_X32 FILLER_35_577 ();
 FILLCELL_X32 FILLER_35_609 ();
 FILLCELL_X32 FILLER_35_641 ();
 FILLCELL_X32 FILLER_35_673 ();
 FILLCELL_X32 FILLER_35_705 ();
 FILLCELL_X32 FILLER_35_737 ();
 FILLCELL_X16 FILLER_35_769 ();
 FILLCELL_X4 FILLER_35_785 ();
 FILLCELL_X1 FILLER_35_789 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X32 FILLER_36_65 ();
 FILLCELL_X32 FILLER_36_97 ();
 FILLCELL_X32 FILLER_36_129 ();
 FILLCELL_X32 FILLER_36_161 ();
 FILLCELL_X32 FILLER_36_193 ();
 FILLCELL_X32 FILLER_36_225 ();
 FILLCELL_X32 FILLER_36_257 ();
 FILLCELL_X32 FILLER_36_289 ();
 FILLCELL_X32 FILLER_36_321 ();
 FILLCELL_X32 FILLER_36_353 ();
 FILLCELL_X32 FILLER_36_385 ();
 FILLCELL_X32 FILLER_36_417 ();
 FILLCELL_X32 FILLER_36_449 ();
 FILLCELL_X32 FILLER_36_481 ();
 FILLCELL_X32 FILLER_36_513 ();
 FILLCELL_X32 FILLER_36_545 ();
 FILLCELL_X32 FILLER_36_577 ();
 FILLCELL_X16 FILLER_36_609 ();
 FILLCELL_X4 FILLER_36_625 ();
 FILLCELL_X2 FILLER_36_629 ();
 FILLCELL_X32 FILLER_36_632 ();
 FILLCELL_X32 FILLER_36_664 ();
 FILLCELL_X32 FILLER_36_696 ();
 FILLCELL_X32 FILLER_36_728 ();
 FILLCELL_X16 FILLER_36_760 ();
 FILLCELL_X8 FILLER_36_776 ();
 FILLCELL_X4 FILLER_36_784 ();
 FILLCELL_X2 FILLER_36_788 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X32 FILLER_37_65 ();
 FILLCELL_X32 FILLER_37_97 ();
 FILLCELL_X32 FILLER_37_129 ();
 FILLCELL_X32 FILLER_37_161 ();
 FILLCELL_X32 FILLER_37_193 ();
 FILLCELL_X32 FILLER_37_225 ();
 FILLCELL_X32 FILLER_37_257 ();
 FILLCELL_X32 FILLER_37_289 ();
 FILLCELL_X32 FILLER_37_321 ();
 FILLCELL_X32 FILLER_37_353 ();
 FILLCELL_X32 FILLER_37_385 ();
 FILLCELL_X32 FILLER_37_417 ();
 FILLCELL_X32 FILLER_37_449 ();
 FILLCELL_X32 FILLER_37_481 ();
 FILLCELL_X32 FILLER_37_513 ();
 FILLCELL_X32 FILLER_37_545 ();
 FILLCELL_X32 FILLER_37_577 ();
 FILLCELL_X32 FILLER_37_609 ();
 FILLCELL_X32 FILLER_37_641 ();
 FILLCELL_X32 FILLER_37_673 ();
 FILLCELL_X32 FILLER_37_705 ();
 FILLCELL_X32 FILLER_37_737 ();
 FILLCELL_X16 FILLER_37_769 ();
 FILLCELL_X4 FILLER_37_785 ();
 FILLCELL_X1 FILLER_37_789 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X32 FILLER_38_65 ();
 FILLCELL_X32 FILLER_38_97 ();
 FILLCELL_X32 FILLER_38_129 ();
 FILLCELL_X32 FILLER_38_161 ();
 FILLCELL_X32 FILLER_38_193 ();
 FILLCELL_X32 FILLER_38_225 ();
 FILLCELL_X32 FILLER_38_257 ();
 FILLCELL_X32 FILLER_38_289 ();
 FILLCELL_X32 FILLER_38_321 ();
 FILLCELL_X32 FILLER_38_353 ();
 FILLCELL_X32 FILLER_38_385 ();
 FILLCELL_X32 FILLER_38_417 ();
 FILLCELL_X32 FILLER_38_449 ();
 FILLCELL_X32 FILLER_38_481 ();
 FILLCELL_X32 FILLER_38_513 ();
 FILLCELL_X32 FILLER_38_545 ();
 FILLCELL_X32 FILLER_38_577 ();
 FILLCELL_X16 FILLER_38_609 ();
 FILLCELL_X4 FILLER_38_625 ();
 FILLCELL_X2 FILLER_38_629 ();
 FILLCELL_X32 FILLER_38_632 ();
 FILLCELL_X32 FILLER_38_664 ();
 FILLCELL_X32 FILLER_38_696 ();
 FILLCELL_X32 FILLER_38_728 ();
 FILLCELL_X16 FILLER_38_760 ();
 FILLCELL_X8 FILLER_38_776 ();
 FILLCELL_X4 FILLER_38_784 ();
 FILLCELL_X2 FILLER_38_788 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X32 FILLER_39_65 ();
 FILLCELL_X32 FILLER_39_97 ();
 FILLCELL_X32 FILLER_39_129 ();
 FILLCELL_X32 FILLER_39_161 ();
 FILLCELL_X32 FILLER_39_193 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X32 FILLER_39_257 ();
 FILLCELL_X32 FILLER_39_289 ();
 FILLCELL_X32 FILLER_39_321 ();
 FILLCELL_X32 FILLER_39_353 ();
 FILLCELL_X32 FILLER_39_385 ();
 FILLCELL_X32 FILLER_39_417 ();
 FILLCELL_X32 FILLER_39_449 ();
 FILLCELL_X32 FILLER_39_481 ();
 FILLCELL_X32 FILLER_39_513 ();
 FILLCELL_X32 FILLER_39_545 ();
 FILLCELL_X32 FILLER_39_577 ();
 FILLCELL_X32 FILLER_39_609 ();
 FILLCELL_X32 FILLER_39_641 ();
 FILLCELL_X32 FILLER_39_673 ();
 FILLCELL_X32 FILLER_39_705 ();
 FILLCELL_X32 FILLER_39_737 ();
 FILLCELL_X16 FILLER_39_769 ();
 FILLCELL_X4 FILLER_39_785 ();
 FILLCELL_X1 FILLER_39_789 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X32 FILLER_40_33 ();
 FILLCELL_X32 FILLER_40_65 ();
 FILLCELL_X32 FILLER_40_97 ();
 FILLCELL_X32 FILLER_40_129 ();
 FILLCELL_X32 FILLER_40_161 ();
 FILLCELL_X32 FILLER_40_193 ();
 FILLCELL_X32 FILLER_40_225 ();
 FILLCELL_X32 FILLER_40_257 ();
 FILLCELL_X32 FILLER_40_289 ();
 FILLCELL_X32 FILLER_40_321 ();
 FILLCELL_X32 FILLER_40_353 ();
 FILLCELL_X32 FILLER_40_385 ();
 FILLCELL_X32 FILLER_40_417 ();
 FILLCELL_X32 FILLER_40_449 ();
 FILLCELL_X32 FILLER_40_481 ();
 FILLCELL_X32 FILLER_40_513 ();
 FILLCELL_X32 FILLER_40_545 ();
 FILLCELL_X32 FILLER_40_577 ();
 FILLCELL_X16 FILLER_40_609 ();
 FILLCELL_X4 FILLER_40_625 ();
 FILLCELL_X2 FILLER_40_629 ();
 FILLCELL_X32 FILLER_40_632 ();
 FILLCELL_X32 FILLER_40_664 ();
 FILLCELL_X32 FILLER_40_696 ();
 FILLCELL_X32 FILLER_40_728 ();
 FILLCELL_X16 FILLER_40_760 ();
 FILLCELL_X8 FILLER_40_776 ();
 FILLCELL_X4 FILLER_40_784 ();
 FILLCELL_X2 FILLER_40_788 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X32 FILLER_41_33 ();
 FILLCELL_X32 FILLER_41_65 ();
 FILLCELL_X32 FILLER_41_97 ();
 FILLCELL_X32 FILLER_41_129 ();
 FILLCELL_X32 FILLER_41_161 ();
 FILLCELL_X32 FILLER_41_193 ();
 FILLCELL_X32 FILLER_41_225 ();
 FILLCELL_X32 FILLER_41_257 ();
 FILLCELL_X32 FILLER_41_289 ();
 FILLCELL_X32 FILLER_41_321 ();
 FILLCELL_X32 FILLER_41_353 ();
 FILLCELL_X32 FILLER_41_385 ();
 FILLCELL_X32 FILLER_41_417 ();
 FILLCELL_X32 FILLER_41_449 ();
 FILLCELL_X32 FILLER_41_481 ();
 FILLCELL_X32 FILLER_41_513 ();
 FILLCELL_X32 FILLER_41_545 ();
 FILLCELL_X32 FILLER_41_577 ();
 FILLCELL_X32 FILLER_41_609 ();
 FILLCELL_X32 FILLER_41_641 ();
 FILLCELL_X32 FILLER_41_673 ();
 FILLCELL_X32 FILLER_41_705 ();
 FILLCELL_X32 FILLER_41_737 ();
 FILLCELL_X16 FILLER_41_769 ();
 FILLCELL_X4 FILLER_41_785 ();
 FILLCELL_X1 FILLER_41_789 ();
 FILLCELL_X32 FILLER_42_1 ();
 FILLCELL_X32 FILLER_42_33 ();
 FILLCELL_X32 FILLER_42_65 ();
 FILLCELL_X32 FILLER_42_97 ();
 FILLCELL_X32 FILLER_42_129 ();
 FILLCELL_X32 FILLER_42_161 ();
 FILLCELL_X32 FILLER_42_193 ();
 FILLCELL_X32 FILLER_42_225 ();
 FILLCELL_X32 FILLER_42_257 ();
 FILLCELL_X32 FILLER_42_289 ();
 FILLCELL_X32 FILLER_42_321 ();
 FILLCELL_X32 FILLER_42_353 ();
 FILLCELL_X32 FILLER_42_385 ();
 FILLCELL_X32 FILLER_42_417 ();
 FILLCELL_X32 FILLER_42_449 ();
 FILLCELL_X32 FILLER_42_481 ();
 FILLCELL_X32 FILLER_42_513 ();
 FILLCELL_X32 FILLER_42_545 ();
 FILLCELL_X32 FILLER_42_577 ();
 FILLCELL_X16 FILLER_42_609 ();
 FILLCELL_X4 FILLER_42_625 ();
 FILLCELL_X2 FILLER_42_629 ();
 FILLCELL_X32 FILLER_42_632 ();
 FILLCELL_X32 FILLER_42_664 ();
 FILLCELL_X32 FILLER_42_696 ();
 FILLCELL_X32 FILLER_42_728 ();
 FILLCELL_X16 FILLER_42_760 ();
 FILLCELL_X8 FILLER_42_776 ();
 FILLCELL_X4 FILLER_42_784 ();
 FILLCELL_X2 FILLER_42_788 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X32 FILLER_43_33 ();
 FILLCELL_X32 FILLER_43_65 ();
 FILLCELL_X32 FILLER_43_97 ();
 FILLCELL_X32 FILLER_43_129 ();
 FILLCELL_X32 FILLER_43_161 ();
 FILLCELL_X32 FILLER_43_193 ();
 FILLCELL_X32 FILLER_43_225 ();
 FILLCELL_X32 FILLER_43_257 ();
 FILLCELL_X32 FILLER_43_289 ();
 FILLCELL_X32 FILLER_43_321 ();
 FILLCELL_X32 FILLER_43_353 ();
 FILLCELL_X32 FILLER_43_385 ();
 FILLCELL_X32 FILLER_43_417 ();
 FILLCELL_X32 FILLER_43_449 ();
 FILLCELL_X32 FILLER_43_481 ();
 FILLCELL_X32 FILLER_43_513 ();
 FILLCELL_X32 FILLER_43_545 ();
 FILLCELL_X32 FILLER_43_577 ();
 FILLCELL_X32 FILLER_43_609 ();
 FILLCELL_X32 FILLER_43_641 ();
 FILLCELL_X32 FILLER_43_673 ();
 FILLCELL_X32 FILLER_43_705 ();
 FILLCELL_X32 FILLER_43_737 ();
 FILLCELL_X16 FILLER_43_769 ();
 FILLCELL_X4 FILLER_43_785 ();
 FILLCELL_X1 FILLER_43_789 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X32 FILLER_44_33 ();
 FILLCELL_X32 FILLER_44_65 ();
 FILLCELL_X32 FILLER_44_97 ();
 FILLCELL_X32 FILLER_44_129 ();
 FILLCELL_X32 FILLER_44_161 ();
 FILLCELL_X32 FILLER_44_193 ();
 FILLCELL_X32 FILLER_44_225 ();
 FILLCELL_X32 FILLER_44_257 ();
 FILLCELL_X32 FILLER_44_289 ();
 FILLCELL_X32 FILLER_44_321 ();
 FILLCELL_X32 FILLER_44_353 ();
 FILLCELL_X32 FILLER_44_385 ();
 FILLCELL_X32 FILLER_44_417 ();
 FILLCELL_X32 FILLER_44_449 ();
 FILLCELL_X32 FILLER_44_481 ();
 FILLCELL_X32 FILLER_44_513 ();
 FILLCELL_X32 FILLER_44_545 ();
 FILLCELL_X32 FILLER_44_577 ();
 FILLCELL_X16 FILLER_44_609 ();
 FILLCELL_X4 FILLER_44_625 ();
 FILLCELL_X2 FILLER_44_629 ();
 FILLCELL_X32 FILLER_44_632 ();
 FILLCELL_X32 FILLER_44_664 ();
 FILLCELL_X32 FILLER_44_696 ();
 FILLCELL_X32 FILLER_44_728 ();
 FILLCELL_X16 FILLER_44_760 ();
 FILLCELL_X8 FILLER_44_776 ();
 FILLCELL_X4 FILLER_44_784 ();
 FILLCELL_X2 FILLER_44_788 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X32 FILLER_45_33 ();
 FILLCELL_X32 FILLER_45_65 ();
 FILLCELL_X32 FILLER_45_97 ();
 FILLCELL_X32 FILLER_45_129 ();
 FILLCELL_X32 FILLER_45_161 ();
 FILLCELL_X32 FILLER_45_193 ();
 FILLCELL_X32 FILLER_45_225 ();
 FILLCELL_X32 FILLER_45_257 ();
 FILLCELL_X32 FILLER_45_289 ();
 FILLCELL_X32 FILLER_45_321 ();
 FILLCELL_X32 FILLER_45_353 ();
 FILLCELL_X32 FILLER_45_385 ();
 FILLCELL_X32 FILLER_45_417 ();
 FILLCELL_X32 FILLER_45_449 ();
 FILLCELL_X32 FILLER_45_481 ();
 FILLCELL_X32 FILLER_45_513 ();
 FILLCELL_X32 FILLER_45_545 ();
 FILLCELL_X32 FILLER_45_577 ();
 FILLCELL_X32 FILLER_45_609 ();
 FILLCELL_X32 FILLER_45_641 ();
 FILLCELL_X32 FILLER_45_673 ();
 FILLCELL_X32 FILLER_45_705 ();
 FILLCELL_X32 FILLER_45_737 ();
 FILLCELL_X16 FILLER_45_769 ();
 FILLCELL_X4 FILLER_45_785 ();
 FILLCELL_X1 FILLER_45_789 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X32 FILLER_46_33 ();
 FILLCELL_X32 FILLER_46_65 ();
 FILLCELL_X32 FILLER_46_97 ();
 FILLCELL_X32 FILLER_46_129 ();
 FILLCELL_X32 FILLER_46_161 ();
 FILLCELL_X32 FILLER_46_193 ();
 FILLCELL_X32 FILLER_46_225 ();
 FILLCELL_X32 FILLER_46_257 ();
 FILLCELL_X32 FILLER_46_289 ();
 FILLCELL_X32 FILLER_46_321 ();
 FILLCELL_X32 FILLER_46_353 ();
 FILLCELL_X32 FILLER_46_385 ();
 FILLCELL_X8 FILLER_46_417 ();
 FILLCELL_X1 FILLER_46_425 ();
 FILLCELL_X32 FILLER_46_428 ();
 FILLCELL_X32 FILLER_46_460 ();
 FILLCELL_X32 FILLER_46_492 ();
 FILLCELL_X32 FILLER_46_524 ();
 FILLCELL_X32 FILLER_46_556 ();
 FILLCELL_X32 FILLER_46_588 ();
 FILLCELL_X8 FILLER_46_620 ();
 FILLCELL_X2 FILLER_46_628 ();
 FILLCELL_X1 FILLER_46_630 ();
 FILLCELL_X32 FILLER_46_632 ();
 FILLCELL_X32 FILLER_46_664 ();
 FILLCELL_X32 FILLER_46_696 ();
 FILLCELL_X32 FILLER_46_728 ();
 FILLCELL_X8 FILLER_46_760 ();
 FILLCELL_X4 FILLER_46_768 ();
 FILLCELL_X2 FILLER_46_775 ();
 FILLCELL_X8 FILLER_46_781 ();
 FILLCELL_X1 FILLER_46_789 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X32 FILLER_47_33 ();
 FILLCELL_X32 FILLER_47_65 ();
 FILLCELL_X32 FILLER_47_97 ();
 FILLCELL_X32 FILLER_47_129 ();
 FILLCELL_X32 FILLER_47_161 ();
 FILLCELL_X32 FILLER_47_193 ();
 FILLCELL_X32 FILLER_47_225 ();
 FILLCELL_X32 FILLER_47_257 ();
 FILLCELL_X32 FILLER_47_289 ();
 FILLCELL_X32 FILLER_47_321 ();
 FILLCELL_X32 FILLER_47_353 ();
 FILLCELL_X32 FILLER_47_385 ();
 FILLCELL_X32 FILLER_47_417 ();
 FILLCELL_X32 FILLER_47_449 ();
 FILLCELL_X32 FILLER_47_481 ();
 FILLCELL_X32 FILLER_47_513 ();
 FILLCELL_X32 FILLER_47_545 ();
 FILLCELL_X32 FILLER_47_577 ();
 FILLCELL_X32 FILLER_47_609 ();
 FILLCELL_X32 FILLER_47_641 ();
 FILLCELL_X32 FILLER_47_673 ();
 FILLCELL_X32 FILLER_47_705 ();
 FILLCELL_X32 FILLER_47_737 ();
 FILLCELL_X16 FILLER_47_769 ();
 FILLCELL_X4 FILLER_47_785 ();
 FILLCELL_X1 FILLER_47_789 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X32 FILLER_48_65 ();
 FILLCELL_X32 FILLER_48_97 ();
 FILLCELL_X32 FILLER_48_129 ();
 FILLCELL_X32 FILLER_48_161 ();
 FILLCELL_X32 FILLER_48_193 ();
 FILLCELL_X32 FILLER_48_225 ();
 FILLCELL_X32 FILLER_48_257 ();
 FILLCELL_X32 FILLER_48_289 ();
 FILLCELL_X32 FILLER_48_321 ();
 FILLCELL_X32 FILLER_48_353 ();
 FILLCELL_X32 FILLER_48_385 ();
 FILLCELL_X32 FILLER_48_417 ();
 FILLCELL_X32 FILLER_48_449 ();
 FILLCELL_X32 FILLER_48_481 ();
 FILLCELL_X32 FILLER_48_513 ();
 FILLCELL_X32 FILLER_48_545 ();
 FILLCELL_X32 FILLER_48_577 ();
 FILLCELL_X16 FILLER_48_609 ();
 FILLCELL_X4 FILLER_48_625 ();
 FILLCELL_X2 FILLER_48_629 ();
 FILLCELL_X32 FILLER_48_632 ();
 FILLCELL_X32 FILLER_48_664 ();
 FILLCELL_X32 FILLER_48_696 ();
 FILLCELL_X32 FILLER_48_728 ();
 FILLCELL_X16 FILLER_48_760 ();
 FILLCELL_X8 FILLER_48_776 ();
 FILLCELL_X4 FILLER_48_784 ();
 FILLCELL_X2 FILLER_48_788 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X32 FILLER_49_33 ();
 FILLCELL_X32 FILLER_49_65 ();
 FILLCELL_X32 FILLER_49_97 ();
 FILLCELL_X32 FILLER_49_129 ();
 FILLCELL_X32 FILLER_49_161 ();
 FILLCELL_X32 FILLER_49_193 ();
 FILLCELL_X32 FILLER_49_225 ();
 FILLCELL_X32 FILLER_49_257 ();
 FILLCELL_X32 FILLER_49_289 ();
 FILLCELL_X32 FILLER_49_321 ();
 FILLCELL_X32 FILLER_49_353 ();
 FILLCELL_X32 FILLER_49_385 ();
 FILLCELL_X32 FILLER_49_417 ();
 FILLCELL_X32 FILLER_49_449 ();
 FILLCELL_X32 FILLER_49_481 ();
 FILLCELL_X32 FILLER_49_513 ();
 FILLCELL_X32 FILLER_49_545 ();
 FILLCELL_X32 FILLER_49_577 ();
 FILLCELL_X32 FILLER_49_609 ();
 FILLCELL_X32 FILLER_49_641 ();
 FILLCELL_X32 FILLER_49_673 ();
 FILLCELL_X32 FILLER_49_705 ();
 FILLCELL_X32 FILLER_49_737 ();
 FILLCELL_X4 FILLER_49_769 ();
 FILLCELL_X2 FILLER_49_773 ();
 FILLCELL_X1 FILLER_49_775 ();
 FILLCELL_X8 FILLER_49_779 ();
 FILLCELL_X2 FILLER_49_787 ();
 FILLCELL_X1 FILLER_49_789 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X32 FILLER_50_33 ();
 FILLCELL_X32 FILLER_50_65 ();
 FILLCELL_X32 FILLER_50_97 ();
 FILLCELL_X32 FILLER_50_129 ();
 FILLCELL_X32 FILLER_50_161 ();
 FILLCELL_X32 FILLER_50_193 ();
 FILLCELL_X32 FILLER_50_225 ();
 FILLCELL_X32 FILLER_50_257 ();
 FILLCELL_X32 FILLER_50_289 ();
 FILLCELL_X32 FILLER_50_321 ();
 FILLCELL_X32 FILLER_50_353 ();
 FILLCELL_X32 FILLER_50_385 ();
 FILLCELL_X32 FILLER_50_417 ();
 FILLCELL_X32 FILLER_50_449 ();
 FILLCELL_X32 FILLER_50_481 ();
 FILLCELL_X32 FILLER_50_513 ();
 FILLCELL_X32 FILLER_50_545 ();
 FILLCELL_X32 FILLER_50_577 ();
 FILLCELL_X16 FILLER_50_609 ();
 FILLCELL_X4 FILLER_50_625 ();
 FILLCELL_X2 FILLER_50_629 ();
 FILLCELL_X32 FILLER_50_632 ();
 FILLCELL_X32 FILLER_50_664 ();
 FILLCELL_X32 FILLER_50_696 ();
 FILLCELL_X32 FILLER_50_728 ();
 FILLCELL_X2 FILLER_50_760 ();
 FILLCELL_X2 FILLER_50_772 ();
 FILLCELL_X1 FILLER_50_774 ();
 FILLCELL_X2 FILLER_50_777 ();
 FILLCELL_X1 FILLER_50_779 ();
 FILLCELL_X1 FILLER_50_783 ();
 FILLCELL_X32 FILLER_51_1 ();
 FILLCELL_X32 FILLER_51_33 ();
 FILLCELL_X32 FILLER_51_65 ();
 FILLCELL_X32 FILLER_51_97 ();
 FILLCELL_X32 FILLER_51_129 ();
 FILLCELL_X32 FILLER_51_161 ();
 FILLCELL_X32 FILLER_51_193 ();
 FILLCELL_X32 FILLER_51_225 ();
 FILLCELL_X32 FILLER_51_257 ();
 FILLCELL_X32 FILLER_51_289 ();
 FILLCELL_X32 FILLER_51_321 ();
 FILLCELL_X32 FILLER_51_353 ();
 FILLCELL_X32 FILLER_51_385 ();
 FILLCELL_X32 FILLER_51_417 ();
 FILLCELL_X32 FILLER_51_449 ();
 FILLCELL_X32 FILLER_51_481 ();
 FILLCELL_X32 FILLER_51_513 ();
 FILLCELL_X32 FILLER_51_545 ();
 FILLCELL_X32 FILLER_51_577 ();
 FILLCELL_X32 FILLER_51_609 ();
 FILLCELL_X32 FILLER_51_641 ();
 FILLCELL_X32 FILLER_51_673 ();
 FILLCELL_X32 FILLER_51_705 ();
 FILLCELL_X16 FILLER_51_737 ();
 FILLCELL_X8 FILLER_51_753 ();
 FILLCELL_X4 FILLER_51_761 ();
 FILLCELL_X1 FILLER_51_765 ();
 FILLCELL_X2 FILLER_51_772 ();
 FILLCELL_X1 FILLER_51_774 ();
 FILLCELL_X1 FILLER_51_789 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X32 FILLER_52_33 ();
 FILLCELL_X32 FILLER_52_65 ();
 FILLCELL_X32 FILLER_52_97 ();
 FILLCELL_X32 FILLER_52_129 ();
 FILLCELL_X32 FILLER_52_161 ();
 FILLCELL_X32 FILLER_52_193 ();
 FILLCELL_X32 FILLER_52_225 ();
 FILLCELL_X32 FILLER_52_257 ();
 FILLCELL_X32 FILLER_52_289 ();
 FILLCELL_X32 FILLER_52_321 ();
 FILLCELL_X32 FILLER_52_353 ();
 FILLCELL_X32 FILLER_52_385 ();
 FILLCELL_X32 FILLER_52_417 ();
 FILLCELL_X32 FILLER_52_449 ();
 FILLCELL_X32 FILLER_52_481 ();
 FILLCELL_X32 FILLER_52_513 ();
 FILLCELL_X32 FILLER_52_545 ();
 FILLCELL_X32 FILLER_52_577 ();
 FILLCELL_X16 FILLER_52_609 ();
 FILLCELL_X4 FILLER_52_625 ();
 FILLCELL_X2 FILLER_52_629 ();
 FILLCELL_X32 FILLER_52_632 ();
 FILLCELL_X32 FILLER_52_664 ();
 FILLCELL_X32 FILLER_52_696 ();
 FILLCELL_X32 FILLER_52_728 ();
 FILLCELL_X16 FILLER_52_760 ();
 FILLCELL_X8 FILLER_52_776 ();
 FILLCELL_X4 FILLER_52_784 ();
 FILLCELL_X2 FILLER_52_788 ();
 FILLCELL_X32 FILLER_53_1 ();
 FILLCELL_X32 FILLER_53_33 ();
 FILLCELL_X32 FILLER_53_65 ();
 FILLCELL_X32 FILLER_53_97 ();
 FILLCELL_X32 FILLER_53_129 ();
 FILLCELL_X32 FILLER_53_161 ();
 FILLCELL_X32 FILLER_53_193 ();
 FILLCELL_X32 FILLER_53_225 ();
 FILLCELL_X32 FILLER_53_257 ();
 FILLCELL_X32 FILLER_53_289 ();
 FILLCELL_X16 FILLER_53_321 ();
 FILLCELL_X4 FILLER_53_337 ();
 FILLCELL_X2 FILLER_53_341 ();
 FILLCELL_X32 FILLER_53_352 ();
 FILLCELL_X32 FILLER_53_384 ();
 FILLCELL_X32 FILLER_53_416 ();
 FILLCELL_X32 FILLER_53_448 ();
 FILLCELL_X32 FILLER_53_480 ();
 FILLCELL_X32 FILLER_53_512 ();
 FILLCELL_X32 FILLER_53_544 ();
 FILLCELL_X32 FILLER_53_576 ();
 FILLCELL_X32 FILLER_53_608 ();
 FILLCELL_X32 FILLER_53_640 ();
 FILLCELL_X32 FILLER_53_672 ();
 FILLCELL_X32 FILLER_53_704 ();
 FILLCELL_X8 FILLER_53_736 ();
 FILLCELL_X4 FILLER_53_744 ();
 FILLCELL_X2 FILLER_53_748 ();
 FILLCELL_X2 FILLER_54_6 ();
 FILLCELL_X1 FILLER_54_18 ();
 FILLCELL_X32 FILLER_54_26 ();
 FILLCELL_X32 FILLER_54_58 ();
 FILLCELL_X32 FILLER_54_90 ();
 FILLCELL_X32 FILLER_54_122 ();
 FILLCELL_X32 FILLER_54_154 ();
 FILLCELL_X32 FILLER_54_186 ();
 FILLCELL_X32 FILLER_54_218 ();
 FILLCELL_X32 FILLER_54_250 ();
 FILLCELL_X32 FILLER_54_282 ();
 FILLCELL_X16 FILLER_54_314 ();
 FILLCELL_X8 FILLER_54_330 ();
 FILLCELL_X4 FILLER_54_338 ();
 FILLCELL_X2 FILLER_54_342 ();
 FILLCELL_X8 FILLER_54_351 ();
 FILLCELL_X4 FILLER_54_359 ();
 FILLCELL_X2 FILLER_54_363 ();
 FILLCELL_X1 FILLER_54_365 ();
 FILLCELL_X1 FILLER_54_369 ();
 FILLCELL_X4 FILLER_54_380 ();
 FILLCELL_X2 FILLER_54_384 ();
 FILLCELL_X1 FILLER_54_386 ();
 FILLCELL_X32 FILLER_54_405 ();
 FILLCELL_X32 FILLER_54_437 ();
 FILLCELL_X32 FILLER_54_469 ();
 FILLCELL_X32 FILLER_54_501 ();
 FILLCELL_X32 FILLER_54_533 ();
 FILLCELL_X32 FILLER_54_565 ();
 FILLCELL_X32 FILLER_54_597 ();
 FILLCELL_X2 FILLER_54_629 ();
 FILLCELL_X32 FILLER_54_632 ();
 FILLCELL_X32 FILLER_54_664 ();
 FILLCELL_X32 FILLER_54_696 ();
 FILLCELL_X16 FILLER_54_728 ();
 FILLCELL_X2 FILLER_54_744 ();
 FILLCELL_X1 FILLER_54_746 ();
 FILLCELL_X32 FILLER_54_758 ();
 FILLCELL_X4 FILLER_55_19 ();
 FILLCELL_X1 FILLER_55_23 ();
 FILLCELL_X2 FILLER_55_27 ();
 FILLCELL_X1 FILLER_55_29 ();
 FILLCELL_X32 FILLER_55_33 ();
 FILLCELL_X32 FILLER_55_65 ();
 FILLCELL_X32 FILLER_55_97 ();
 FILLCELL_X32 FILLER_55_129 ();
 FILLCELL_X32 FILLER_55_161 ();
 FILLCELL_X32 FILLER_55_193 ();
 FILLCELL_X32 FILLER_55_225 ();
 FILLCELL_X32 FILLER_55_257 ();
 FILLCELL_X16 FILLER_55_289 ();
 FILLCELL_X8 FILLER_55_305 ();
 FILLCELL_X16 FILLER_55_315 ();
 FILLCELL_X2 FILLER_55_331 ();
 FILLCELL_X1 FILLER_55_333 ();
 FILLCELL_X8 FILLER_55_357 ();
 FILLCELL_X4 FILLER_55_365 ();
 FILLCELL_X1 FILLER_55_369 ();
 FILLCELL_X32 FILLER_55_379 ();
 FILLCELL_X32 FILLER_55_411 ();
 FILLCELL_X32 FILLER_55_443 ();
 FILLCELL_X32 FILLER_55_475 ();
 FILLCELL_X32 FILLER_55_507 ();
 FILLCELL_X32 FILLER_55_539 ();
 FILLCELL_X32 FILLER_55_571 ();
 FILLCELL_X32 FILLER_55_603 ();
 FILLCELL_X32 FILLER_55_635 ();
 FILLCELL_X32 FILLER_55_667 ();
 FILLCELL_X16 FILLER_55_699 ();
 FILLCELL_X8 FILLER_55_715 ();
 FILLCELL_X2 FILLER_55_723 ();
 FILLCELL_X1 FILLER_55_725 ();
 FILLCELL_X32 FILLER_55_736 ();
 FILLCELL_X16 FILLER_55_768 ();
 FILLCELL_X4 FILLER_55_784 ();
 FILLCELL_X2 FILLER_55_788 ();
 FILLCELL_X2 FILLER_56_1 ();
 FILLCELL_X1 FILLER_56_3 ();
 FILLCELL_X4 FILLER_56_7 ();
 FILLCELL_X2 FILLER_56_11 ();
 FILLCELL_X1 FILLER_56_13 ();
 FILLCELL_X32 FILLER_56_17 ();
 FILLCELL_X32 FILLER_56_49 ();
 FILLCELL_X32 FILLER_56_81 ();
 FILLCELL_X32 FILLER_56_113 ();
 FILLCELL_X32 FILLER_56_145 ();
 FILLCELL_X32 FILLER_56_177 ();
 FILLCELL_X32 FILLER_56_209 ();
 FILLCELL_X32 FILLER_56_241 ();
 FILLCELL_X32 FILLER_56_273 ();
 FILLCELL_X32 FILLER_56_305 ();
 FILLCELL_X4 FILLER_56_337 ();
 FILLCELL_X16 FILLER_56_344 ();
 FILLCELL_X8 FILLER_56_360 ();
 FILLCELL_X4 FILLER_56_368 ();
 FILLCELL_X32 FILLER_56_382 ();
 FILLCELL_X32 FILLER_56_414 ();
 FILLCELL_X16 FILLER_56_446 ();
 FILLCELL_X2 FILLER_56_462 ();
 FILLCELL_X1 FILLER_56_464 ();
 FILLCELL_X32 FILLER_56_467 ();
 FILLCELL_X32 FILLER_56_499 ();
 FILLCELL_X32 FILLER_56_531 ();
 FILLCELL_X32 FILLER_56_563 ();
 FILLCELL_X32 FILLER_56_595 ();
 FILLCELL_X4 FILLER_56_627 ();
 FILLCELL_X32 FILLER_56_632 ();
 FILLCELL_X32 FILLER_56_664 ();
 FILLCELL_X32 FILLER_56_696 ();
 FILLCELL_X32 FILLER_56_728 ();
 FILLCELL_X16 FILLER_56_760 ();
 FILLCELL_X8 FILLER_56_776 ();
 FILLCELL_X4 FILLER_56_784 ();
 FILLCELL_X2 FILLER_56_788 ();
 FILLCELL_X32 FILLER_57_1 ();
 FILLCELL_X32 FILLER_57_33 ();
 FILLCELL_X32 FILLER_57_65 ();
 FILLCELL_X32 FILLER_57_97 ();
 FILLCELL_X32 FILLER_57_129 ();
 FILLCELL_X32 FILLER_57_161 ();
 FILLCELL_X32 FILLER_57_193 ();
 FILLCELL_X32 FILLER_57_225 ();
 FILLCELL_X32 FILLER_57_257 ();
 FILLCELL_X32 FILLER_57_289 ();
 FILLCELL_X32 FILLER_57_321 ();
 FILLCELL_X32 FILLER_57_353 ();
 FILLCELL_X32 FILLER_57_385 ();
 FILLCELL_X32 FILLER_57_417 ();
 FILLCELL_X32 FILLER_57_449 ();
 FILLCELL_X32 FILLER_57_481 ();
 FILLCELL_X32 FILLER_57_513 ();
 FILLCELL_X32 FILLER_57_545 ();
 FILLCELL_X32 FILLER_57_577 ();
 FILLCELL_X32 FILLER_57_609 ();
 FILLCELL_X32 FILLER_57_641 ();
 FILLCELL_X32 FILLER_57_673 ();
 FILLCELL_X32 FILLER_57_705 ();
 FILLCELL_X32 FILLER_57_737 ();
 FILLCELL_X16 FILLER_57_769 ();
 FILLCELL_X4 FILLER_57_785 ();
 FILLCELL_X1 FILLER_57_789 ();
 FILLCELL_X32 FILLER_58_1 ();
 FILLCELL_X32 FILLER_58_33 ();
 FILLCELL_X32 FILLER_58_65 ();
 FILLCELL_X32 FILLER_58_97 ();
 FILLCELL_X32 FILLER_58_129 ();
 FILLCELL_X32 FILLER_58_161 ();
 FILLCELL_X32 FILLER_58_193 ();
 FILLCELL_X32 FILLER_58_225 ();
 FILLCELL_X32 FILLER_58_257 ();
 FILLCELL_X32 FILLER_58_289 ();
 FILLCELL_X32 FILLER_58_321 ();
 FILLCELL_X32 FILLER_58_353 ();
 FILLCELL_X32 FILLER_58_385 ();
 FILLCELL_X32 FILLER_58_417 ();
 FILLCELL_X32 FILLER_58_449 ();
 FILLCELL_X32 FILLER_58_481 ();
 FILLCELL_X32 FILLER_58_513 ();
 FILLCELL_X32 FILLER_58_545 ();
 FILLCELL_X32 FILLER_58_577 ();
 FILLCELL_X16 FILLER_58_609 ();
 FILLCELL_X4 FILLER_58_625 ();
 FILLCELL_X2 FILLER_58_629 ();
 FILLCELL_X32 FILLER_58_632 ();
 FILLCELL_X32 FILLER_58_664 ();
 FILLCELL_X32 FILLER_58_696 ();
 FILLCELL_X32 FILLER_58_728 ();
 FILLCELL_X16 FILLER_58_760 ();
 FILLCELL_X8 FILLER_58_776 ();
 FILLCELL_X4 FILLER_58_784 ();
 FILLCELL_X2 FILLER_58_788 ();
 FILLCELL_X32 FILLER_59_1 ();
 FILLCELL_X32 FILLER_59_33 ();
 FILLCELL_X32 FILLER_59_65 ();
 FILLCELL_X32 FILLER_59_97 ();
 FILLCELL_X32 FILLER_59_129 ();
 FILLCELL_X32 FILLER_59_161 ();
 FILLCELL_X32 FILLER_59_193 ();
 FILLCELL_X32 FILLER_59_225 ();
 FILLCELL_X32 FILLER_59_257 ();
 FILLCELL_X32 FILLER_59_289 ();
 FILLCELL_X32 FILLER_59_321 ();
 FILLCELL_X32 FILLER_59_353 ();
 FILLCELL_X32 FILLER_59_385 ();
 FILLCELL_X32 FILLER_59_417 ();
 FILLCELL_X32 FILLER_59_449 ();
 FILLCELL_X32 FILLER_59_481 ();
 FILLCELL_X32 FILLER_59_513 ();
 FILLCELL_X32 FILLER_59_545 ();
 FILLCELL_X32 FILLER_59_577 ();
 FILLCELL_X32 FILLER_59_609 ();
 FILLCELL_X32 FILLER_59_641 ();
 FILLCELL_X32 FILLER_59_673 ();
 FILLCELL_X32 FILLER_59_705 ();
 FILLCELL_X32 FILLER_59_737 ();
 FILLCELL_X16 FILLER_59_769 ();
 FILLCELL_X4 FILLER_59_785 ();
 FILLCELL_X1 FILLER_59_789 ();
 FILLCELL_X2 FILLER_60_1 ();
 FILLCELL_X2 FILLER_60_6 ();
 FILLCELL_X32 FILLER_60_25 ();
 FILLCELL_X32 FILLER_60_57 ();
 FILLCELL_X32 FILLER_60_89 ();
 FILLCELL_X32 FILLER_60_121 ();
 FILLCELL_X32 FILLER_60_153 ();
 FILLCELL_X32 FILLER_60_185 ();
 FILLCELL_X32 FILLER_60_217 ();
 FILLCELL_X32 FILLER_60_249 ();
 FILLCELL_X32 FILLER_60_281 ();
 FILLCELL_X32 FILLER_60_313 ();
 FILLCELL_X2 FILLER_60_345 ();
 FILLCELL_X1 FILLER_60_347 ();
 FILLCELL_X32 FILLER_60_373 ();
 FILLCELL_X32 FILLER_60_405 ();
 FILLCELL_X32 FILLER_60_437 ();
 FILLCELL_X32 FILLER_60_469 ();
 FILLCELL_X32 FILLER_60_501 ();
 FILLCELL_X32 FILLER_60_533 ();
 FILLCELL_X32 FILLER_60_565 ();
 FILLCELL_X32 FILLER_60_597 ();
 FILLCELL_X2 FILLER_60_629 ();
 FILLCELL_X32 FILLER_60_632 ();
 FILLCELL_X32 FILLER_60_664 ();
 FILLCELL_X32 FILLER_60_696 ();
 FILLCELL_X32 FILLER_60_728 ();
 FILLCELL_X16 FILLER_60_760 ();
 FILLCELL_X8 FILLER_60_776 ();
 FILLCELL_X4 FILLER_60_784 ();
 FILLCELL_X2 FILLER_60_788 ();
 FILLCELL_X1 FILLER_61_6 ();
 FILLCELL_X32 FILLER_61_20 ();
 FILLCELL_X32 FILLER_61_52 ();
 FILLCELL_X32 FILLER_61_84 ();
 FILLCELL_X32 FILLER_61_116 ();
 FILLCELL_X32 FILLER_61_148 ();
 FILLCELL_X32 FILLER_61_180 ();
 FILLCELL_X32 FILLER_61_212 ();
 FILLCELL_X32 FILLER_61_244 ();
 FILLCELL_X32 FILLER_61_276 ();
 FILLCELL_X32 FILLER_61_308 ();
 FILLCELL_X32 FILLER_61_340 ();
 FILLCELL_X8 FILLER_61_372 ();
 FILLCELL_X4 FILLER_61_380 ();
 FILLCELL_X1 FILLER_61_384 ();
 FILLCELL_X32 FILLER_61_395 ();
 FILLCELL_X32 FILLER_61_427 ();
 FILLCELL_X32 FILLER_61_459 ();
 FILLCELL_X32 FILLER_61_491 ();
 FILLCELL_X32 FILLER_61_523 ();
 FILLCELL_X32 FILLER_61_555 ();
 FILLCELL_X32 FILLER_61_587 ();
 FILLCELL_X32 FILLER_61_619 ();
 FILLCELL_X32 FILLER_61_651 ();
 FILLCELL_X32 FILLER_61_683 ();
 FILLCELL_X32 FILLER_61_715 ();
 FILLCELL_X32 FILLER_61_747 ();
 FILLCELL_X8 FILLER_61_779 ();
 FILLCELL_X2 FILLER_61_787 ();
 FILLCELL_X1 FILLER_61_789 ();
 FILLCELL_X1 FILLER_62_1 ();
 FILLCELL_X1 FILLER_62_5 ();
 FILLCELL_X32 FILLER_62_8 ();
 FILLCELL_X32 FILLER_62_40 ();
 FILLCELL_X32 FILLER_62_72 ();
 FILLCELL_X32 FILLER_62_104 ();
 FILLCELL_X32 FILLER_62_136 ();
 FILLCELL_X32 FILLER_62_168 ();
 FILLCELL_X32 FILLER_62_200 ();
 FILLCELL_X32 FILLER_62_232 ();
 FILLCELL_X32 FILLER_62_264 ();
 FILLCELL_X32 FILLER_62_296 ();
 FILLCELL_X32 FILLER_62_328 ();
 FILLCELL_X32 FILLER_62_360 ();
 FILLCELL_X32 FILLER_62_392 ();
 FILLCELL_X32 FILLER_62_424 ();
 FILLCELL_X32 FILLER_62_456 ();
 FILLCELL_X32 FILLER_62_488 ();
 FILLCELL_X32 FILLER_62_520 ();
 FILLCELL_X32 FILLER_62_552 ();
 FILLCELL_X32 FILLER_62_584 ();
 FILLCELL_X8 FILLER_62_616 ();
 FILLCELL_X4 FILLER_62_624 ();
 FILLCELL_X2 FILLER_62_628 ();
 FILLCELL_X1 FILLER_62_630 ();
 FILLCELL_X32 FILLER_62_632 ();
 FILLCELL_X32 FILLER_62_664 ();
 FILLCELL_X32 FILLER_62_696 ();
 FILLCELL_X32 FILLER_62_728 ();
 FILLCELL_X16 FILLER_62_760 ();
 FILLCELL_X8 FILLER_62_776 ();
 FILLCELL_X4 FILLER_62_784 ();
 FILLCELL_X2 FILLER_62_788 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X32 FILLER_63_33 ();
 FILLCELL_X32 FILLER_63_65 ();
 FILLCELL_X32 FILLER_63_97 ();
 FILLCELL_X32 FILLER_63_129 ();
 FILLCELL_X32 FILLER_63_161 ();
 FILLCELL_X32 FILLER_63_193 ();
 FILLCELL_X32 FILLER_63_225 ();
 FILLCELL_X32 FILLER_63_257 ();
 FILLCELL_X32 FILLER_63_289 ();
 FILLCELL_X32 FILLER_63_321 ();
 FILLCELL_X32 FILLER_63_353 ();
 FILLCELL_X2 FILLER_63_385 ();
 FILLCELL_X32 FILLER_63_389 ();
 FILLCELL_X32 FILLER_63_421 ();
 FILLCELL_X32 FILLER_63_453 ();
 FILLCELL_X32 FILLER_63_485 ();
 FILLCELL_X32 FILLER_63_517 ();
 FILLCELL_X32 FILLER_63_549 ();
 FILLCELL_X32 FILLER_63_581 ();
 FILLCELL_X32 FILLER_63_613 ();
 FILLCELL_X32 FILLER_63_645 ();
 FILLCELL_X32 FILLER_63_677 ();
 FILLCELL_X32 FILLER_63_709 ();
 FILLCELL_X32 FILLER_63_741 ();
 FILLCELL_X16 FILLER_63_773 ();
 FILLCELL_X1 FILLER_63_789 ();
 FILLCELL_X32 FILLER_64_1 ();
 FILLCELL_X32 FILLER_64_33 ();
 FILLCELL_X32 FILLER_64_65 ();
 FILLCELL_X32 FILLER_64_97 ();
 FILLCELL_X32 FILLER_64_129 ();
 FILLCELL_X32 FILLER_64_161 ();
 FILLCELL_X32 FILLER_64_193 ();
 FILLCELL_X32 FILLER_64_225 ();
 FILLCELL_X32 FILLER_64_257 ();
 FILLCELL_X32 FILLER_64_289 ();
 FILLCELL_X32 FILLER_64_321 ();
 FILLCELL_X32 FILLER_64_353 ();
 FILLCELL_X32 FILLER_64_385 ();
 FILLCELL_X32 FILLER_64_417 ();
 FILLCELL_X32 FILLER_64_449 ();
 FILLCELL_X32 FILLER_64_481 ();
 FILLCELL_X32 FILLER_64_513 ();
 FILLCELL_X32 FILLER_64_545 ();
 FILLCELL_X32 FILLER_64_577 ();
 FILLCELL_X16 FILLER_64_609 ();
 FILLCELL_X4 FILLER_64_625 ();
 FILLCELL_X2 FILLER_64_629 ();
 FILLCELL_X32 FILLER_64_632 ();
 FILLCELL_X32 FILLER_64_664 ();
 FILLCELL_X32 FILLER_64_696 ();
 FILLCELL_X32 FILLER_64_728 ();
 FILLCELL_X16 FILLER_64_760 ();
 FILLCELL_X8 FILLER_64_776 ();
 FILLCELL_X4 FILLER_64_784 ();
 FILLCELL_X2 FILLER_64_788 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X32 FILLER_65_33 ();
 FILLCELL_X32 FILLER_65_65 ();
 FILLCELL_X32 FILLER_65_97 ();
 FILLCELL_X32 FILLER_65_129 ();
 FILLCELL_X32 FILLER_65_161 ();
 FILLCELL_X32 FILLER_65_193 ();
 FILLCELL_X32 FILLER_65_225 ();
 FILLCELL_X32 FILLER_65_257 ();
 FILLCELL_X32 FILLER_65_289 ();
 FILLCELL_X32 FILLER_65_321 ();
 FILLCELL_X32 FILLER_65_353 ();
 FILLCELL_X32 FILLER_65_385 ();
 FILLCELL_X32 FILLER_65_417 ();
 FILLCELL_X32 FILLER_65_449 ();
 FILLCELL_X32 FILLER_65_481 ();
 FILLCELL_X32 FILLER_65_513 ();
 FILLCELL_X32 FILLER_65_545 ();
 FILLCELL_X32 FILLER_65_577 ();
 FILLCELL_X32 FILLER_65_609 ();
 FILLCELL_X32 FILLER_65_641 ();
 FILLCELL_X32 FILLER_65_673 ();
 FILLCELL_X32 FILLER_65_705 ();
 FILLCELL_X32 FILLER_65_737 ();
 FILLCELL_X16 FILLER_65_769 ();
 FILLCELL_X4 FILLER_65_785 ();
 FILLCELL_X1 FILLER_65_789 ();
 FILLCELL_X32 FILLER_66_1 ();
 FILLCELL_X32 FILLER_66_33 ();
 FILLCELL_X32 FILLER_66_65 ();
 FILLCELL_X32 FILLER_66_97 ();
 FILLCELL_X32 FILLER_66_129 ();
 FILLCELL_X32 FILLER_66_161 ();
 FILLCELL_X32 FILLER_66_193 ();
 FILLCELL_X32 FILLER_66_225 ();
 FILLCELL_X32 FILLER_66_257 ();
 FILLCELL_X32 FILLER_66_289 ();
 FILLCELL_X32 FILLER_66_321 ();
 FILLCELL_X32 FILLER_66_353 ();
 FILLCELL_X32 FILLER_66_385 ();
 FILLCELL_X32 FILLER_66_417 ();
 FILLCELL_X32 FILLER_66_449 ();
 FILLCELL_X32 FILLER_66_481 ();
 FILLCELL_X32 FILLER_66_513 ();
 FILLCELL_X32 FILLER_66_545 ();
 FILLCELL_X32 FILLER_66_577 ();
 FILLCELL_X16 FILLER_66_609 ();
 FILLCELL_X4 FILLER_66_625 ();
 FILLCELL_X2 FILLER_66_629 ();
 FILLCELL_X32 FILLER_66_632 ();
 FILLCELL_X32 FILLER_66_664 ();
 FILLCELL_X32 FILLER_66_696 ();
 FILLCELL_X32 FILLER_66_728 ();
 FILLCELL_X16 FILLER_66_760 ();
 FILLCELL_X8 FILLER_66_776 ();
 FILLCELL_X4 FILLER_66_784 ();
 FILLCELL_X2 FILLER_66_788 ();
 FILLCELL_X32 FILLER_67_1 ();
 FILLCELL_X32 FILLER_67_33 ();
 FILLCELL_X32 FILLER_67_65 ();
 FILLCELL_X32 FILLER_67_97 ();
 FILLCELL_X32 FILLER_67_129 ();
 FILLCELL_X32 FILLER_67_161 ();
 FILLCELL_X32 FILLER_67_193 ();
 FILLCELL_X32 FILLER_67_225 ();
 FILLCELL_X32 FILLER_67_257 ();
 FILLCELL_X32 FILLER_67_289 ();
 FILLCELL_X32 FILLER_67_321 ();
 FILLCELL_X32 FILLER_67_353 ();
 FILLCELL_X32 FILLER_67_385 ();
 FILLCELL_X32 FILLER_67_417 ();
 FILLCELL_X32 FILLER_67_449 ();
 FILLCELL_X32 FILLER_67_481 ();
 FILLCELL_X32 FILLER_67_513 ();
 FILLCELL_X32 FILLER_67_545 ();
 FILLCELL_X32 FILLER_67_577 ();
 FILLCELL_X32 FILLER_67_609 ();
 FILLCELL_X32 FILLER_67_641 ();
 FILLCELL_X32 FILLER_67_673 ();
 FILLCELL_X32 FILLER_67_705 ();
 FILLCELL_X32 FILLER_67_737 ();
 FILLCELL_X16 FILLER_67_769 ();
 FILLCELL_X4 FILLER_67_785 ();
 FILLCELL_X1 FILLER_67_789 ();
 FILLCELL_X32 FILLER_68_1 ();
 FILLCELL_X32 FILLER_68_33 ();
 FILLCELL_X32 FILLER_68_65 ();
 FILLCELL_X32 FILLER_68_97 ();
 FILLCELL_X32 FILLER_68_129 ();
 FILLCELL_X32 FILLER_68_161 ();
 FILLCELL_X32 FILLER_68_193 ();
 FILLCELL_X32 FILLER_68_225 ();
 FILLCELL_X32 FILLER_68_257 ();
 FILLCELL_X32 FILLER_68_289 ();
 FILLCELL_X32 FILLER_68_321 ();
 FILLCELL_X32 FILLER_68_353 ();
 FILLCELL_X32 FILLER_68_385 ();
 FILLCELL_X32 FILLER_68_417 ();
 FILLCELL_X32 FILLER_68_449 ();
 FILLCELL_X32 FILLER_68_481 ();
 FILLCELL_X32 FILLER_68_513 ();
 FILLCELL_X32 FILLER_68_545 ();
 FILLCELL_X32 FILLER_68_577 ();
 FILLCELL_X16 FILLER_68_609 ();
 FILLCELL_X4 FILLER_68_625 ();
 FILLCELL_X2 FILLER_68_629 ();
 FILLCELL_X32 FILLER_68_632 ();
 FILLCELL_X32 FILLER_68_664 ();
 FILLCELL_X32 FILLER_68_696 ();
 FILLCELL_X32 FILLER_68_728 ();
 FILLCELL_X16 FILLER_68_760 ();
 FILLCELL_X8 FILLER_68_776 ();
 FILLCELL_X4 FILLER_68_784 ();
 FILLCELL_X2 FILLER_68_788 ();
 FILLCELL_X32 FILLER_69_1 ();
 FILLCELL_X32 FILLER_69_33 ();
 FILLCELL_X32 FILLER_69_65 ();
 FILLCELL_X32 FILLER_69_97 ();
 FILLCELL_X32 FILLER_69_129 ();
 FILLCELL_X32 FILLER_69_161 ();
 FILLCELL_X32 FILLER_69_193 ();
 FILLCELL_X32 FILLER_69_225 ();
 FILLCELL_X32 FILLER_69_257 ();
 FILLCELL_X32 FILLER_69_289 ();
 FILLCELL_X32 FILLER_69_321 ();
 FILLCELL_X32 FILLER_69_353 ();
 FILLCELL_X32 FILLER_69_385 ();
 FILLCELL_X32 FILLER_69_417 ();
 FILLCELL_X32 FILLER_69_449 ();
 FILLCELL_X32 FILLER_69_481 ();
 FILLCELL_X32 FILLER_69_513 ();
 FILLCELL_X32 FILLER_69_545 ();
 FILLCELL_X32 FILLER_69_577 ();
 FILLCELL_X32 FILLER_69_609 ();
 FILLCELL_X32 FILLER_69_641 ();
 FILLCELL_X32 FILLER_69_673 ();
 FILLCELL_X32 FILLER_69_705 ();
 FILLCELL_X32 FILLER_69_737 ();
 FILLCELL_X16 FILLER_69_769 ();
 FILLCELL_X4 FILLER_69_785 ();
 FILLCELL_X1 FILLER_69_789 ();
 FILLCELL_X32 FILLER_70_1 ();
 FILLCELL_X32 FILLER_70_33 ();
 FILLCELL_X32 FILLER_70_65 ();
 FILLCELL_X32 FILLER_70_97 ();
 FILLCELL_X32 FILLER_70_129 ();
 FILLCELL_X32 FILLER_70_161 ();
 FILLCELL_X32 FILLER_70_193 ();
 FILLCELL_X32 FILLER_70_225 ();
 FILLCELL_X32 FILLER_70_257 ();
 FILLCELL_X32 FILLER_70_289 ();
 FILLCELL_X32 FILLER_70_321 ();
 FILLCELL_X32 FILLER_70_353 ();
 FILLCELL_X32 FILLER_70_385 ();
 FILLCELL_X32 FILLER_70_417 ();
 FILLCELL_X32 FILLER_70_449 ();
 FILLCELL_X32 FILLER_70_481 ();
 FILLCELL_X32 FILLER_70_513 ();
 FILLCELL_X32 FILLER_70_545 ();
 FILLCELL_X32 FILLER_70_577 ();
 FILLCELL_X16 FILLER_70_609 ();
 FILLCELL_X4 FILLER_70_625 ();
 FILLCELL_X2 FILLER_70_629 ();
 FILLCELL_X32 FILLER_70_632 ();
 FILLCELL_X32 FILLER_70_664 ();
 FILLCELL_X32 FILLER_70_696 ();
 FILLCELL_X32 FILLER_70_728 ();
 FILLCELL_X16 FILLER_70_760 ();
 FILLCELL_X8 FILLER_70_776 ();
 FILLCELL_X4 FILLER_70_784 ();
 FILLCELL_X2 FILLER_70_788 ();
 FILLCELL_X32 FILLER_71_1 ();
 FILLCELL_X32 FILLER_71_33 ();
 FILLCELL_X32 FILLER_71_65 ();
 FILLCELL_X32 FILLER_71_97 ();
 FILLCELL_X32 FILLER_71_129 ();
 FILLCELL_X32 FILLER_71_161 ();
 FILLCELL_X32 FILLER_71_193 ();
 FILLCELL_X32 FILLER_71_225 ();
 FILLCELL_X32 FILLER_71_257 ();
 FILLCELL_X32 FILLER_71_289 ();
 FILLCELL_X32 FILLER_71_321 ();
 FILLCELL_X32 FILLER_71_353 ();
 FILLCELL_X32 FILLER_71_385 ();
 FILLCELL_X32 FILLER_71_417 ();
 FILLCELL_X32 FILLER_71_449 ();
 FILLCELL_X32 FILLER_71_481 ();
 FILLCELL_X32 FILLER_71_513 ();
 FILLCELL_X32 FILLER_71_545 ();
 FILLCELL_X32 FILLER_71_577 ();
 FILLCELL_X32 FILLER_71_609 ();
 FILLCELL_X32 FILLER_71_641 ();
 FILLCELL_X32 FILLER_71_673 ();
 FILLCELL_X32 FILLER_71_705 ();
 FILLCELL_X32 FILLER_71_737 ();
 FILLCELL_X16 FILLER_71_769 ();
 FILLCELL_X4 FILLER_71_785 ();
 FILLCELL_X1 FILLER_71_789 ();
 FILLCELL_X32 FILLER_72_1 ();
 FILLCELL_X32 FILLER_72_33 ();
 FILLCELL_X32 FILLER_72_65 ();
 FILLCELL_X32 FILLER_72_97 ();
 FILLCELL_X32 FILLER_72_129 ();
 FILLCELL_X32 FILLER_72_161 ();
 FILLCELL_X32 FILLER_72_193 ();
 FILLCELL_X32 FILLER_72_225 ();
 FILLCELL_X32 FILLER_72_257 ();
 FILLCELL_X32 FILLER_72_289 ();
 FILLCELL_X32 FILLER_72_321 ();
 FILLCELL_X32 FILLER_72_353 ();
 FILLCELL_X32 FILLER_72_385 ();
 FILLCELL_X32 FILLER_72_417 ();
 FILLCELL_X32 FILLER_72_449 ();
 FILLCELL_X32 FILLER_72_481 ();
 FILLCELL_X32 FILLER_72_513 ();
 FILLCELL_X32 FILLER_72_545 ();
 FILLCELL_X32 FILLER_72_577 ();
 FILLCELL_X16 FILLER_72_609 ();
 FILLCELL_X4 FILLER_72_625 ();
 FILLCELL_X2 FILLER_72_629 ();
 FILLCELL_X32 FILLER_72_632 ();
 FILLCELL_X32 FILLER_72_664 ();
 FILLCELL_X32 FILLER_72_696 ();
 FILLCELL_X32 FILLER_72_728 ();
 FILLCELL_X16 FILLER_72_760 ();
 FILLCELL_X8 FILLER_72_776 ();
 FILLCELL_X4 FILLER_72_784 ();
 FILLCELL_X2 FILLER_72_788 ();
 FILLCELL_X32 FILLER_73_1 ();
 FILLCELL_X32 FILLER_73_33 ();
 FILLCELL_X32 FILLER_73_65 ();
 FILLCELL_X32 FILLER_73_97 ();
 FILLCELL_X32 FILLER_73_129 ();
 FILLCELL_X32 FILLER_73_161 ();
 FILLCELL_X32 FILLER_73_193 ();
 FILLCELL_X32 FILLER_73_225 ();
 FILLCELL_X32 FILLER_73_257 ();
 FILLCELL_X32 FILLER_73_289 ();
 FILLCELL_X32 FILLER_73_321 ();
 FILLCELL_X32 FILLER_73_353 ();
 FILLCELL_X32 FILLER_73_385 ();
 FILLCELL_X32 FILLER_73_417 ();
 FILLCELL_X32 FILLER_73_449 ();
 FILLCELL_X32 FILLER_73_481 ();
 FILLCELL_X32 FILLER_73_513 ();
 FILLCELL_X32 FILLER_73_545 ();
 FILLCELL_X32 FILLER_73_577 ();
 FILLCELL_X32 FILLER_73_609 ();
 FILLCELL_X32 FILLER_73_641 ();
 FILLCELL_X32 FILLER_73_673 ();
 FILLCELL_X32 FILLER_73_705 ();
 FILLCELL_X32 FILLER_73_737 ();
 FILLCELL_X16 FILLER_73_769 ();
 FILLCELL_X4 FILLER_73_785 ();
 FILLCELL_X1 FILLER_73_789 ();
 FILLCELL_X32 FILLER_74_1 ();
 FILLCELL_X32 FILLER_74_33 ();
 FILLCELL_X32 FILLER_74_65 ();
 FILLCELL_X32 FILLER_74_97 ();
 FILLCELL_X32 FILLER_74_129 ();
 FILLCELL_X32 FILLER_74_161 ();
 FILLCELL_X32 FILLER_74_193 ();
 FILLCELL_X32 FILLER_74_225 ();
 FILLCELL_X32 FILLER_74_257 ();
 FILLCELL_X32 FILLER_74_289 ();
 FILLCELL_X32 FILLER_74_321 ();
 FILLCELL_X32 FILLER_74_353 ();
 FILLCELL_X32 FILLER_74_385 ();
 FILLCELL_X32 FILLER_74_417 ();
 FILLCELL_X32 FILLER_74_449 ();
 FILLCELL_X32 FILLER_74_481 ();
 FILLCELL_X32 FILLER_74_513 ();
 FILLCELL_X32 FILLER_74_545 ();
 FILLCELL_X32 FILLER_74_577 ();
 FILLCELL_X16 FILLER_74_609 ();
 FILLCELL_X4 FILLER_74_625 ();
 FILLCELL_X2 FILLER_74_629 ();
 FILLCELL_X32 FILLER_74_632 ();
 FILLCELL_X32 FILLER_74_664 ();
 FILLCELL_X32 FILLER_74_696 ();
 FILLCELL_X32 FILLER_74_728 ();
 FILLCELL_X16 FILLER_74_760 ();
 FILLCELL_X8 FILLER_74_776 ();
 FILLCELL_X4 FILLER_74_784 ();
 FILLCELL_X2 FILLER_74_788 ();
 FILLCELL_X32 FILLER_75_1 ();
 FILLCELL_X32 FILLER_75_33 ();
 FILLCELL_X32 FILLER_75_65 ();
 FILLCELL_X32 FILLER_75_97 ();
 FILLCELL_X32 FILLER_75_129 ();
 FILLCELL_X32 FILLER_75_161 ();
 FILLCELL_X32 FILLER_75_193 ();
 FILLCELL_X32 FILLER_75_225 ();
 FILLCELL_X32 FILLER_75_257 ();
 FILLCELL_X32 FILLER_75_289 ();
 FILLCELL_X32 FILLER_75_321 ();
 FILLCELL_X32 FILLER_75_353 ();
 FILLCELL_X32 FILLER_75_385 ();
 FILLCELL_X32 FILLER_75_417 ();
 FILLCELL_X32 FILLER_75_449 ();
 FILLCELL_X32 FILLER_75_481 ();
 FILLCELL_X32 FILLER_75_513 ();
 FILLCELL_X32 FILLER_75_545 ();
 FILLCELL_X32 FILLER_75_577 ();
 FILLCELL_X32 FILLER_75_609 ();
 FILLCELL_X32 FILLER_75_641 ();
 FILLCELL_X32 FILLER_75_673 ();
 FILLCELL_X32 FILLER_75_705 ();
 FILLCELL_X32 FILLER_75_737 ();
 FILLCELL_X16 FILLER_75_769 ();
 FILLCELL_X4 FILLER_75_785 ();
 FILLCELL_X1 FILLER_75_789 ();
 FILLCELL_X32 FILLER_76_1 ();
 FILLCELL_X32 FILLER_76_33 ();
 FILLCELL_X32 FILLER_76_65 ();
 FILLCELL_X32 FILLER_76_97 ();
 FILLCELL_X32 FILLER_76_129 ();
 FILLCELL_X32 FILLER_76_161 ();
 FILLCELL_X32 FILLER_76_193 ();
 FILLCELL_X32 FILLER_76_225 ();
 FILLCELL_X32 FILLER_76_257 ();
 FILLCELL_X32 FILLER_76_289 ();
 FILLCELL_X32 FILLER_76_321 ();
 FILLCELL_X32 FILLER_76_353 ();
 FILLCELL_X32 FILLER_76_385 ();
 FILLCELL_X32 FILLER_76_417 ();
 FILLCELL_X32 FILLER_76_449 ();
 FILLCELL_X32 FILLER_76_481 ();
 FILLCELL_X32 FILLER_76_513 ();
 FILLCELL_X32 FILLER_76_545 ();
 FILLCELL_X32 FILLER_76_577 ();
 FILLCELL_X16 FILLER_76_609 ();
 FILLCELL_X4 FILLER_76_625 ();
 FILLCELL_X2 FILLER_76_629 ();
 FILLCELL_X32 FILLER_76_632 ();
 FILLCELL_X32 FILLER_76_664 ();
 FILLCELL_X32 FILLER_76_696 ();
 FILLCELL_X32 FILLER_76_728 ();
 FILLCELL_X16 FILLER_76_760 ();
 FILLCELL_X8 FILLER_76_776 ();
 FILLCELL_X4 FILLER_76_784 ();
 FILLCELL_X2 FILLER_76_788 ();
 FILLCELL_X32 FILLER_77_1 ();
 FILLCELL_X32 FILLER_77_33 ();
 FILLCELL_X32 FILLER_77_65 ();
 FILLCELL_X32 FILLER_77_97 ();
 FILLCELL_X32 FILLER_77_129 ();
 FILLCELL_X32 FILLER_77_161 ();
 FILLCELL_X32 FILLER_77_193 ();
 FILLCELL_X32 FILLER_77_225 ();
 FILLCELL_X32 FILLER_77_257 ();
 FILLCELL_X32 FILLER_77_289 ();
 FILLCELL_X32 FILLER_77_321 ();
 FILLCELL_X32 FILLER_77_353 ();
 FILLCELL_X32 FILLER_77_385 ();
 FILLCELL_X32 FILLER_77_417 ();
 FILLCELL_X32 FILLER_77_449 ();
 FILLCELL_X32 FILLER_77_481 ();
 FILLCELL_X32 FILLER_77_513 ();
 FILLCELL_X32 FILLER_77_545 ();
 FILLCELL_X32 FILLER_77_577 ();
 FILLCELL_X32 FILLER_77_609 ();
 FILLCELL_X32 FILLER_77_641 ();
 FILLCELL_X32 FILLER_77_673 ();
 FILLCELL_X32 FILLER_77_705 ();
 FILLCELL_X32 FILLER_77_737 ();
 FILLCELL_X16 FILLER_77_769 ();
 FILLCELL_X4 FILLER_77_785 ();
 FILLCELL_X1 FILLER_77_789 ();
 FILLCELL_X32 FILLER_78_1 ();
 FILLCELL_X32 FILLER_78_33 ();
 FILLCELL_X32 FILLER_78_65 ();
 FILLCELL_X32 FILLER_78_97 ();
 FILLCELL_X32 FILLER_78_129 ();
 FILLCELL_X32 FILLER_78_161 ();
 FILLCELL_X32 FILLER_78_193 ();
 FILLCELL_X32 FILLER_78_225 ();
 FILLCELL_X32 FILLER_78_257 ();
 FILLCELL_X32 FILLER_78_289 ();
 FILLCELL_X32 FILLER_78_321 ();
 FILLCELL_X32 FILLER_78_353 ();
 FILLCELL_X32 FILLER_78_385 ();
 FILLCELL_X32 FILLER_78_417 ();
 FILLCELL_X32 FILLER_78_449 ();
 FILLCELL_X32 FILLER_78_481 ();
 FILLCELL_X32 FILLER_78_513 ();
 FILLCELL_X32 FILLER_78_545 ();
 FILLCELL_X32 FILLER_78_577 ();
 FILLCELL_X16 FILLER_78_609 ();
 FILLCELL_X4 FILLER_78_625 ();
 FILLCELL_X2 FILLER_78_629 ();
 FILLCELL_X32 FILLER_78_632 ();
 FILLCELL_X32 FILLER_78_664 ();
 FILLCELL_X32 FILLER_78_696 ();
 FILLCELL_X32 FILLER_78_728 ();
 FILLCELL_X16 FILLER_78_760 ();
 FILLCELL_X8 FILLER_78_776 ();
 FILLCELL_X4 FILLER_78_784 ();
 FILLCELL_X2 FILLER_78_788 ();
 FILLCELL_X32 FILLER_79_1 ();
 FILLCELL_X32 FILLER_79_33 ();
 FILLCELL_X32 FILLER_79_65 ();
 FILLCELL_X32 FILLER_79_97 ();
 FILLCELL_X32 FILLER_79_129 ();
 FILLCELL_X32 FILLER_79_161 ();
 FILLCELL_X32 FILLER_79_193 ();
 FILLCELL_X32 FILLER_79_225 ();
 FILLCELL_X32 FILLER_79_257 ();
 FILLCELL_X32 FILLER_79_289 ();
 FILLCELL_X32 FILLER_79_321 ();
 FILLCELL_X32 FILLER_79_353 ();
 FILLCELL_X32 FILLER_79_385 ();
 FILLCELL_X32 FILLER_79_417 ();
 FILLCELL_X32 FILLER_79_449 ();
 FILLCELL_X32 FILLER_79_481 ();
 FILLCELL_X32 FILLER_79_513 ();
 FILLCELL_X32 FILLER_79_545 ();
 FILLCELL_X32 FILLER_79_577 ();
 FILLCELL_X32 FILLER_79_609 ();
 FILLCELL_X32 FILLER_79_641 ();
 FILLCELL_X32 FILLER_79_673 ();
 FILLCELL_X32 FILLER_79_705 ();
 FILLCELL_X32 FILLER_79_737 ();
 FILLCELL_X16 FILLER_79_769 ();
 FILLCELL_X4 FILLER_79_785 ();
 FILLCELL_X1 FILLER_79_789 ();
 FILLCELL_X32 FILLER_80_1 ();
 FILLCELL_X32 FILLER_80_33 ();
 FILLCELL_X32 FILLER_80_65 ();
 FILLCELL_X32 FILLER_80_97 ();
 FILLCELL_X32 FILLER_80_129 ();
 FILLCELL_X32 FILLER_80_161 ();
 FILLCELL_X32 FILLER_80_193 ();
 FILLCELL_X32 FILLER_80_225 ();
 FILLCELL_X32 FILLER_80_257 ();
 FILLCELL_X32 FILLER_80_289 ();
 FILLCELL_X32 FILLER_80_321 ();
 FILLCELL_X32 FILLER_80_353 ();
 FILLCELL_X32 FILLER_80_385 ();
 FILLCELL_X32 FILLER_80_417 ();
 FILLCELL_X32 FILLER_80_449 ();
 FILLCELL_X32 FILLER_80_481 ();
 FILLCELL_X32 FILLER_80_513 ();
 FILLCELL_X32 FILLER_80_545 ();
 FILLCELL_X32 FILLER_80_577 ();
 FILLCELL_X16 FILLER_80_609 ();
 FILLCELL_X4 FILLER_80_625 ();
 FILLCELL_X2 FILLER_80_629 ();
 FILLCELL_X32 FILLER_80_632 ();
 FILLCELL_X32 FILLER_80_664 ();
 FILLCELL_X32 FILLER_80_696 ();
 FILLCELL_X32 FILLER_80_728 ();
 FILLCELL_X16 FILLER_80_760 ();
 FILLCELL_X8 FILLER_80_776 ();
 FILLCELL_X4 FILLER_80_784 ();
 FILLCELL_X2 FILLER_80_788 ();
 FILLCELL_X32 FILLER_81_1 ();
 FILLCELL_X32 FILLER_81_33 ();
 FILLCELL_X32 FILLER_81_65 ();
 FILLCELL_X32 FILLER_81_97 ();
 FILLCELL_X32 FILLER_81_129 ();
 FILLCELL_X32 FILLER_81_161 ();
 FILLCELL_X32 FILLER_81_193 ();
 FILLCELL_X32 FILLER_81_225 ();
 FILLCELL_X32 FILLER_81_257 ();
 FILLCELL_X32 FILLER_81_289 ();
 FILLCELL_X32 FILLER_81_321 ();
 FILLCELL_X32 FILLER_81_353 ();
 FILLCELL_X32 FILLER_81_385 ();
 FILLCELL_X32 FILLER_81_417 ();
 FILLCELL_X32 FILLER_81_449 ();
 FILLCELL_X32 FILLER_81_481 ();
 FILLCELL_X32 FILLER_81_513 ();
 FILLCELL_X32 FILLER_81_545 ();
 FILLCELL_X32 FILLER_81_577 ();
 FILLCELL_X32 FILLER_81_609 ();
 FILLCELL_X32 FILLER_81_641 ();
 FILLCELL_X32 FILLER_81_673 ();
 FILLCELL_X32 FILLER_81_705 ();
 FILLCELL_X32 FILLER_81_737 ();
 FILLCELL_X16 FILLER_81_769 ();
 FILLCELL_X4 FILLER_81_785 ();
 FILLCELL_X1 FILLER_81_789 ();
 FILLCELL_X32 FILLER_82_1 ();
 FILLCELL_X32 FILLER_82_33 ();
 FILLCELL_X32 FILLER_82_65 ();
 FILLCELL_X32 FILLER_82_97 ();
 FILLCELL_X32 FILLER_82_129 ();
 FILLCELL_X32 FILLER_82_161 ();
 FILLCELL_X32 FILLER_82_193 ();
 FILLCELL_X32 FILLER_82_225 ();
 FILLCELL_X32 FILLER_82_257 ();
 FILLCELL_X32 FILLER_82_289 ();
 FILLCELL_X32 FILLER_82_321 ();
 FILLCELL_X32 FILLER_82_353 ();
 FILLCELL_X32 FILLER_82_385 ();
 FILLCELL_X32 FILLER_82_417 ();
 FILLCELL_X32 FILLER_82_449 ();
 FILLCELL_X32 FILLER_82_481 ();
 FILLCELL_X32 FILLER_82_513 ();
 FILLCELL_X32 FILLER_82_545 ();
 FILLCELL_X32 FILLER_82_577 ();
 FILLCELL_X16 FILLER_82_609 ();
 FILLCELL_X4 FILLER_82_625 ();
 FILLCELL_X2 FILLER_82_629 ();
 FILLCELL_X32 FILLER_82_632 ();
 FILLCELL_X32 FILLER_82_664 ();
 FILLCELL_X32 FILLER_82_696 ();
 FILLCELL_X32 FILLER_82_728 ();
 FILLCELL_X16 FILLER_82_760 ();
 FILLCELL_X8 FILLER_82_776 ();
 FILLCELL_X4 FILLER_82_784 ();
 FILLCELL_X2 FILLER_82_788 ();
 FILLCELL_X32 FILLER_83_1 ();
 FILLCELL_X32 FILLER_83_33 ();
 FILLCELL_X32 FILLER_83_65 ();
 FILLCELL_X32 FILLER_83_97 ();
 FILLCELL_X32 FILLER_83_129 ();
 FILLCELL_X32 FILLER_83_161 ();
 FILLCELL_X32 FILLER_83_193 ();
 FILLCELL_X32 FILLER_83_225 ();
 FILLCELL_X32 FILLER_83_257 ();
 FILLCELL_X32 FILLER_83_289 ();
 FILLCELL_X32 FILLER_83_321 ();
 FILLCELL_X32 FILLER_83_353 ();
 FILLCELL_X32 FILLER_83_385 ();
 FILLCELL_X32 FILLER_83_417 ();
 FILLCELL_X32 FILLER_83_449 ();
 FILLCELL_X32 FILLER_83_481 ();
 FILLCELL_X32 FILLER_83_513 ();
 FILLCELL_X32 FILLER_83_545 ();
 FILLCELL_X32 FILLER_83_577 ();
 FILLCELL_X32 FILLER_83_609 ();
 FILLCELL_X32 FILLER_83_641 ();
 FILLCELL_X32 FILLER_83_673 ();
 FILLCELL_X32 FILLER_83_705 ();
 FILLCELL_X32 FILLER_83_737 ();
 FILLCELL_X16 FILLER_83_769 ();
 FILLCELL_X4 FILLER_83_785 ();
 FILLCELL_X1 FILLER_83_789 ();
 FILLCELL_X32 FILLER_84_1 ();
 FILLCELL_X32 FILLER_84_33 ();
 FILLCELL_X32 FILLER_84_65 ();
 FILLCELL_X32 FILLER_84_97 ();
 FILLCELL_X32 FILLER_84_129 ();
 FILLCELL_X32 FILLER_84_161 ();
 FILLCELL_X32 FILLER_84_193 ();
 FILLCELL_X32 FILLER_84_225 ();
 FILLCELL_X32 FILLER_84_257 ();
 FILLCELL_X32 FILLER_84_289 ();
 FILLCELL_X32 FILLER_84_321 ();
 FILLCELL_X32 FILLER_84_353 ();
 FILLCELL_X32 FILLER_84_385 ();
 FILLCELL_X32 FILLER_84_417 ();
 FILLCELL_X32 FILLER_84_449 ();
 FILLCELL_X32 FILLER_84_481 ();
 FILLCELL_X32 FILLER_84_513 ();
 FILLCELL_X32 FILLER_84_545 ();
 FILLCELL_X32 FILLER_84_577 ();
 FILLCELL_X16 FILLER_84_609 ();
 FILLCELL_X4 FILLER_84_625 ();
 FILLCELL_X2 FILLER_84_629 ();
 FILLCELL_X32 FILLER_84_632 ();
 FILLCELL_X32 FILLER_84_664 ();
 FILLCELL_X32 FILLER_84_696 ();
 FILLCELL_X32 FILLER_84_728 ();
 FILLCELL_X16 FILLER_84_760 ();
 FILLCELL_X8 FILLER_84_776 ();
 FILLCELL_X4 FILLER_84_784 ();
 FILLCELL_X2 FILLER_84_788 ();
 FILLCELL_X32 FILLER_85_1 ();
 FILLCELL_X32 FILLER_85_33 ();
 FILLCELL_X32 FILLER_85_65 ();
 FILLCELL_X32 FILLER_85_97 ();
 FILLCELL_X32 FILLER_85_129 ();
 FILLCELL_X32 FILLER_85_161 ();
 FILLCELL_X32 FILLER_85_193 ();
 FILLCELL_X32 FILLER_85_225 ();
 FILLCELL_X32 FILLER_85_257 ();
 FILLCELL_X32 FILLER_85_289 ();
 FILLCELL_X32 FILLER_85_321 ();
 FILLCELL_X32 FILLER_85_353 ();
 FILLCELL_X32 FILLER_85_385 ();
 FILLCELL_X32 FILLER_85_417 ();
 FILLCELL_X32 FILLER_85_449 ();
 FILLCELL_X32 FILLER_85_481 ();
 FILLCELL_X32 FILLER_85_513 ();
 FILLCELL_X32 FILLER_85_545 ();
 FILLCELL_X32 FILLER_85_577 ();
 FILLCELL_X32 FILLER_85_609 ();
 FILLCELL_X32 FILLER_85_641 ();
 FILLCELL_X32 FILLER_85_673 ();
 FILLCELL_X32 FILLER_85_705 ();
 FILLCELL_X32 FILLER_85_737 ();
 FILLCELL_X16 FILLER_85_769 ();
 FILLCELL_X4 FILLER_85_785 ();
 FILLCELL_X1 FILLER_85_789 ();
 FILLCELL_X32 FILLER_86_1 ();
 FILLCELL_X32 FILLER_86_33 ();
 FILLCELL_X32 FILLER_86_65 ();
 FILLCELL_X32 FILLER_86_97 ();
 FILLCELL_X32 FILLER_86_129 ();
 FILLCELL_X32 FILLER_86_161 ();
 FILLCELL_X32 FILLER_86_193 ();
 FILLCELL_X32 FILLER_86_225 ();
 FILLCELL_X32 FILLER_86_257 ();
 FILLCELL_X32 FILLER_86_289 ();
 FILLCELL_X32 FILLER_86_321 ();
 FILLCELL_X32 FILLER_86_353 ();
 FILLCELL_X32 FILLER_86_385 ();
 FILLCELL_X32 FILLER_86_417 ();
 FILLCELL_X32 FILLER_86_449 ();
 FILLCELL_X32 FILLER_86_481 ();
 FILLCELL_X32 FILLER_86_513 ();
 FILLCELL_X32 FILLER_86_545 ();
 FILLCELL_X32 FILLER_86_577 ();
 FILLCELL_X16 FILLER_86_609 ();
 FILLCELL_X4 FILLER_86_625 ();
 FILLCELL_X2 FILLER_86_629 ();
 FILLCELL_X32 FILLER_86_632 ();
 FILLCELL_X32 FILLER_86_664 ();
 FILLCELL_X32 FILLER_86_696 ();
 FILLCELL_X32 FILLER_86_728 ();
 FILLCELL_X16 FILLER_86_760 ();
 FILLCELL_X8 FILLER_86_776 ();
 FILLCELL_X4 FILLER_86_784 ();
 FILLCELL_X2 FILLER_86_788 ();
 FILLCELL_X32 FILLER_87_1 ();
 FILLCELL_X32 FILLER_87_33 ();
 FILLCELL_X32 FILLER_87_65 ();
 FILLCELL_X32 FILLER_87_97 ();
 FILLCELL_X32 FILLER_87_129 ();
 FILLCELL_X32 FILLER_87_161 ();
 FILLCELL_X32 FILLER_87_193 ();
 FILLCELL_X32 FILLER_87_225 ();
 FILLCELL_X32 FILLER_87_257 ();
 FILLCELL_X32 FILLER_87_289 ();
 FILLCELL_X32 FILLER_87_321 ();
 FILLCELL_X32 FILLER_87_353 ();
 FILLCELL_X32 FILLER_87_385 ();
 FILLCELL_X32 FILLER_87_417 ();
 FILLCELL_X32 FILLER_87_449 ();
 FILLCELL_X32 FILLER_87_481 ();
 FILLCELL_X32 FILLER_87_513 ();
 FILLCELL_X32 FILLER_87_545 ();
 FILLCELL_X32 FILLER_87_577 ();
 FILLCELL_X32 FILLER_87_609 ();
 FILLCELL_X32 FILLER_87_641 ();
 FILLCELL_X32 FILLER_87_673 ();
 FILLCELL_X32 FILLER_87_705 ();
 FILLCELL_X32 FILLER_87_737 ();
 FILLCELL_X16 FILLER_87_769 ();
 FILLCELL_X4 FILLER_87_785 ();
 FILLCELL_X1 FILLER_87_789 ();
 FILLCELL_X32 FILLER_88_1 ();
 FILLCELL_X32 FILLER_88_33 ();
 FILLCELL_X32 FILLER_88_65 ();
 FILLCELL_X32 FILLER_88_97 ();
 FILLCELL_X32 FILLER_88_129 ();
 FILLCELL_X32 FILLER_88_161 ();
 FILLCELL_X32 FILLER_88_193 ();
 FILLCELL_X32 FILLER_88_225 ();
 FILLCELL_X32 FILLER_88_257 ();
 FILLCELL_X32 FILLER_88_289 ();
 FILLCELL_X32 FILLER_88_321 ();
 FILLCELL_X32 FILLER_88_353 ();
 FILLCELL_X32 FILLER_88_385 ();
 FILLCELL_X32 FILLER_88_417 ();
 FILLCELL_X32 FILLER_88_449 ();
 FILLCELL_X32 FILLER_88_481 ();
 FILLCELL_X32 FILLER_88_513 ();
 FILLCELL_X32 FILLER_88_545 ();
 FILLCELL_X32 FILLER_88_577 ();
 FILLCELL_X16 FILLER_88_609 ();
 FILLCELL_X4 FILLER_88_625 ();
 FILLCELL_X2 FILLER_88_629 ();
 FILLCELL_X32 FILLER_88_632 ();
 FILLCELL_X32 FILLER_88_664 ();
 FILLCELL_X32 FILLER_88_696 ();
 FILLCELL_X32 FILLER_88_728 ();
 FILLCELL_X16 FILLER_88_760 ();
 FILLCELL_X8 FILLER_88_776 ();
 FILLCELL_X4 FILLER_88_784 ();
 FILLCELL_X2 FILLER_88_788 ();
 FILLCELL_X32 FILLER_89_1 ();
 FILLCELL_X32 FILLER_89_33 ();
 FILLCELL_X32 FILLER_89_65 ();
 FILLCELL_X32 FILLER_89_97 ();
 FILLCELL_X32 FILLER_89_129 ();
 FILLCELL_X32 FILLER_89_161 ();
 FILLCELL_X32 FILLER_89_193 ();
 FILLCELL_X32 FILLER_89_225 ();
 FILLCELL_X32 FILLER_89_257 ();
 FILLCELL_X32 FILLER_89_289 ();
 FILLCELL_X32 FILLER_89_321 ();
 FILLCELL_X32 FILLER_89_353 ();
 FILLCELL_X32 FILLER_89_385 ();
 FILLCELL_X32 FILLER_89_417 ();
 FILLCELL_X32 FILLER_89_449 ();
 FILLCELL_X32 FILLER_89_481 ();
 FILLCELL_X32 FILLER_89_513 ();
 FILLCELL_X32 FILLER_89_545 ();
 FILLCELL_X32 FILLER_89_577 ();
 FILLCELL_X32 FILLER_89_609 ();
 FILLCELL_X32 FILLER_89_641 ();
 FILLCELL_X32 FILLER_89_673 ();
 FILLCELL_X32 FILLER_89_705 ();
 FILLCELL_X32 FILLER_89_737 ();
 FILLCELL_X16 FILLER_89_769 ();
 FILLCELL_X4 FILLER_89_785 ();
 FILLCELL_X1 FILLER_89_789 ();
 FILLCELL_X32 FILLER_90_1 ();
 FILLCELL_X32 FILLER_90_33 ();
 FILLCELL_X32 FILLER_90_65 ();
 FILLCELL_X32 FILLER_90_97 ();
 FILLCELL_X32 FILLER_90_129 ();
 FILLCELL_X32 FILLER_90_161 ();
 FILLCELL_X32 FILLER_90_193 ();
 FILLCELL_X32 FILLER_90_225 ();
 FILLCELL_X32 FILLER_90_257 ();
 FILLCELL_X32 FILLER_90_289 ();
 FILLCELL_X32 FILLER_90_321 ();
 FILLCELL_X32 FILLER_90_353 ();
 FILLCELL_X32 FILLER_90_385 ();
 FILLCELL_X32 FILLER_90_417 ();
 FILLCELL_X32 FILLER_90_449 ();
 FILLCELL_X32 FILLER_90_481 ();
 FILLCELL_X32 FILLER_90_513 ();
 FILLCELL_X32 FILLER_90_545 ();
 FILLCELL_X32 FILLER_90_577 ();
 FILLCELL_X16 FILLER_90_609 ();
 FILLCELL_X4 FILLER_90_625 ();
 FILLCELL_X2 FILLER_90_629 ();
 FILLCELL_X32 FILLER_90_632 ();
 FILLCELL_X32 FILLER_90_664 ();
 FILLCELL_X32 FILLER_90_696 ();
 FILLCELL_X32 FILLER_90_728 ();
 FILLCELL_X16 FILLER_90_760 ();
 FILLCELL_X8 FILLER_90_776 ();
 FILLCELL_X4 FILLER_90_784 ();
 FILLCELL_X2 FILLER_90_788 ();
 FILLCELL_X32 FILLER_91_1 ();
 FILLCELL_X32 FILLER_91_33 ();
 FILLCELL_X32 FILLER_91_65 ();
 FILLCELL_X32 FILLER_91_97 ();
 FILLCELL_X32 FILLER_91_129 ();
 FILLCELL_X32 FILLER_91_161 ();
 FILLCELL_X32 FILLER_91_193 ();
 FILLCELL_X32 FILLER_91_225 ();
 FILLCELL_X32 FILLER_91_257 ();
 FILLCELL_X32 FILLER_91_289 ();
 FILLCELL_X32 FILLER_91_321 ();
 FILLCELL_X32 FILLER_91_353 ();
 FILLCELL_X32 FILLER_91_385 ();
 FILLCELL_X32 FILLER_91_417 ();
 FILLCELL_X32 FILLER_91_449 ();
 FILLCELL_X32 FILLER_91_481 ();
 FILLCELL_X32 FILLER_91_513 ();
 FILLCELL_X32 FILLER_91_545 ();
 FILLCELL_X32 FILLER_91_577 ();
 FILLCELL_X32 FILLER_91_609 ();
 FILLCELL_X32 FILLER_91_641 ();
 FILLCELL_X32 FILLER_91_673 ();
 FILLCELL_X32 FILLER_91_705 ();
 FILLCELL_X32 FILLER_91_737 ();
 FILLCELL_X16 FILLER_91_769 ();
 FILLCELL_X4 FILLER_91_785 ();
 FILLCELL_X1 FILLER_91_789 ();
 FILLCELL_X32 FILLER_92_1 ();
 FILLCELL_X32 FILLER_92_33 ();
 FILLCELL_X32 FILLER_92_65 ();
 FILLCELL_X32 FILLER_92_97 ();
 FILLCELL_X32 FILLER_92_129 ();
 FILLCELL_X32 FILLER_92_161 ();
 FILLCELL_X32 FILLER_92_193 ();
 FILLCELL_X32 FILLER_92_225 ();
 FILLCELL_X32 FILLER_92_257 ();
 FILLCELL_X32 FILLER_92_289 ();
 FILLCELL_X32 FILLER_92_321 ();
 FILLCELL_X32 FILLER_92_353 ();
 FILLCELL_X32 FILLER_92_385 ();
 FILLCELL_X32 FILLER_92_417 ();
 FILLCELL_X32 FILLER_92_449 ();
 FILLCELL_X32 FILLER_92_481 ();
 FILLCELL_X32 FILLER_92_513 ();
 FILLCELL_X32 FILLER_92_545 ();
 FILLCELL_X32 FILLER_92_577 ();
 FILLCELL_X16 FILLER_92_609 ();
 FILLCELL_X4 FILLER_92_625 ();
 FILLCELL_X2 FILLER_92_629 ();
 FILLCELL_X32 FILLER_92_632 ();
 FILLCELL_X32 FILLER_92_664 ();
 FILLCELL_X32 FILLER_92_696 ();
 FILLCELL_X32 FILLER_92_728 ();
 FILLCELL_X16 FILLER_92_760 ();
 FILLCELL_X8 FILLER_92_776 ();
 FILLCELL_X4 FILLER_92_784 ();
 FILLCELL_X2 FILLER_92_788 ();
 FILLCELL_X32 FILLER_93_1 ();
 FILLCELL_X32 FILLER_93_33 ();
 FILLCELL_X32 FILLER_93_65 ();
 FILLCELL_X32 FILLER_93_97 ();
 FILLCELL_X32 FILLER_93_129 ();
 FILLCELL_X32 FILLER_93_161 ();
 FILLCELL_X32 FILLER_93_193 ();
 FILLCELL_X32 FILLER_93_225 ();
 FILLCELL_X32 FILLER_93_257 ();
 FILLCELL_X32 FILLER_93_289 ();
 FILLCELL_X32 FILLER_93_321 ();
 FILLCELL_X32 FILLER_93_353 ();
 FILLCELL_X32 FILLER_93_385 ();
 FILLCELL_X32 FILLER_93_417 ();
 FILLCELL_X32 FILLER_93_449 ();
 FILLCELL_X32 FILLER_93_481 ();
 FILLCELL_X32 FILLER_93_513 ();
 FILLCELL_X32 FILLER_93_545 ();
 FILLCELL_X32 FILLER_93_577 ();
 FILLCELL_X32 FILLER_93_609 ();
 FILLCELL_X32 FILLER_93_641 ();
 FILLCELL_X32 FILLER_93_673 ();
 FILLCELL_X32 FILLER_93_705 ();
 FILLCELL_X32 FILLER_93_737 ();
 FILLCELL_X16 FILLER_93_769 ();
 FILLCELL_X4 FILLER_93_785 ();
 FILLCELL_X1 FILLER_93_789 ();
 FILLCELL_X32 FILLER_94_1 ();
 FILLCELL_X32 FILLER_94_33 ();
 FILLCELL_X32 FILLER_94_65 ();
 FILLCELL_X32 FILLER_94_97 ();
 FILLCELL_X32 FILLER_94_129 ();
 FILLCELL_X32 FILLER_94_161 ();
 FILLCELL_X32 FILLER_94_193 ();
 FILLCELL_X32 FILLER_94_225 ();
 FILLCELL_X32 FILLER_94_257 ();
 FILLCELL_X32 FILLER_94_289 ();
 FILLCELL_X32 FILLER_94_321 ();
 FILLCELL_X32 FILLER_94_353 ();
 FILLCELL_X32 FILLER_94_385 ();
 FILLCELL_X32 FILLER_94_417 ();
 FILLCELL_X32 FILLER_94_449 ();
 FILLCELL_X32 FILLER_94_481 ();
 FILLCELL_X32 FILLER_94_513 ();
 FILLCELL_X32 FILLER_94_545 ();
 FILLCELL_X32 FILLER_94_577 ();
 FILLCELL_X16 FILLER_94_609 ();
 FILLCELL_X4 FILLER_94_625 ();
 FILLCELL_X2 FILLER_94_629 ();
 FILLCELL_X32 FILLER_94_632 ();
 FILLCELL_X32 FILLER_94_664 ();
 FILLCELL_X32 FILLER_94_696 ();
 FILLCELL_X32 FILLER_94_728 ();
 FILLCELL_X16 FILLER_94_760 ();
 FILLCELL_X8 FILLER_94_776 ();
 FILLCELL_X4 FILLER_94_784 ();
 FILLCELL_X2 FILLER_94_788 ();
 FILLCELL_X32 FILLER_95_1 ();
 FILLCELL_X32 FILLER_95_33 ();
 FILLCELL_X32 FILLER_95_65 ();
 FILLCELL_X32 FILLER_95_97 ();
 FILLCELL_X32 FILLER_95_129 ();
 FILLCELL_X32 FILLER_95_161 ();
 FILLCELL_X32 FILLER_95_193 ();
 FILLCELL_X32 FILLER_95_225 ();
 FILLCELL_X32 FILLER_95_257 ();
 FILLCELL_X32 FILLER_95_289 ();
 FILLCELL_X32 FILLER_95_321 ();
 FILLCELL_X32 FILLER_95_353 ();
 FILLCELL_X32 FILLER_95_385 ();
 FILLCELL_X32 FILLER_95_417 ();
 FILLCELL_X32 FILLER_95_449 ();
 FILLCELL_X32 FILLER_95_481 ();
 FILLCELL_X32 FILLER_95_513 ();
 FILLCELL_X32 FILLER_95_545 ();
 FILLCELL_X32 FILLER_95_577 ();
 FILLCELL_X32 FILLER_95_609 ();
 FILLCELL_X32 FILLER_95_641 ();
 FILLCELL_X32 FILLER_95_673 ();
 FILLCELL_X32 FILLER_95_705 ();
 FILLCELL_X32 FILLER_95_737 ();
 FILLCELL_X16 FILLER_95_769 ();
 FILLCELL_X4 FILLER_95_785 ();
 FILLCELL_X1 FILLER_95_789 ();
 FILLCELL_X32 FILLER_96_1 ();
 FILLCELL_X32 FILLER_96_33 ();
 FILLCELL_X32 FILLER_96_65 ();
 FILLCELL_X32 FILLER_96_97 ();
 FILLCELL_X32 FILLER_96_129 ();
 FILLCELL_X32 FILLER_96_161 ();
 FILLCELL_X32 FILLER_96_193 ();
 FILLCELL_X32 FILLER_96_225 ();
 FILLCELL_X32 FILLER_96_257 ();
 FILLCELL_X32 FILLER_96_289 ();
 FILLCELL_X32 FILLER_96_321 ();
 FILLCELL_X32 FILLER_96_353 ();
 FILLCELL_X32 FILLER_96_385 ();
 FILLCELL_X32 FILLER_96_417 ();
 FILLCELL_X32 FILLER_96_449 ();
 FILLCELL_X32 FILLER_96_481 ();
 FILLCELL_X32 FILLER_96_513 ();
 FILLCELL_X32 FILLER_96_545 ();
 FILLCELL_X32 FILLER_96_577 ();
 FILLCELL_X16 FILLER_96_609 ();
 FILLCELL_X4 FILLER_96_625 ();
 FILLCELL_X2 FILLER_96_629 ();
 FILLCELL_X32 FILLER_96_632 ();
 FILLCELL_X32 FILLER_96_664 ();
 FILLCELL_X32 FILLER_96_696 ();
 FILLCELL_X32 FILLER_96_728 ();
 FILLCELL_X16 FILLER_96_760 ();
 FILLCELL_X8 FILLER_96_776 ();
 FILLCELL_X4 FILLER_96_784 ();
 FILLCELL_X2 FILLER_96_788 ();
 FILLCELL_X32 FILLER_97_1 ();
 FILLCELL_X32 FILLER_97_33 ();
 FILLCELL_X32 FILLER_97_65 ();
 FILLCELL_X32 FILLER_97_97 ();
 FILLCELL_X32 FILLER_97_129 ();
 FILLCELL_X32 FILLER_97_161 ();
 FILLCELL_X32 FILLER_97_193 ();
 FILLCELL_X32 FILLER_97_225 ();
 FILLCELL_X32 FILLER_97_257 ();
 FILLCELL_X32 FILLER_97_289 ();
 FILLCELL_X32 FILLER_97_321 ();
 FILLCELL_X32 FILLER_97_353 ();
 FILLCELL_X32 FILLER_97_385 ();
 FILLCELL_X32 FILLER_97_417 ();
 FILLCELL_X32 FILLER_97_449 ();
 FILLCELL_X32 FILLER_97_481 ();
 FILLCELL_X32 FILLER_97_513 ();
 FILLCELL_X32 FILLER_97_545 ();
 FILLCELL_X32 FILLER_97_577 ();
 FILLCELL_X32 FILLER_97_609 ();
 FILLCELL_X32 FILLER_97_641 ();
 FILLCELL_X32 FILLER_97_673 ();
 FILLCELL_X32 FILLER_97_705 ();
 FILLCELL_X32 FILLER_97_737 ();
 FILLCELL_X16 FILLER_97_769 ();
 FILLCELL_X4 FILLER_97_785 ();
 FILLCELL_X1 FILLER_97_789 ();
 FILLCELL_X32 FILLER_98_1 ();
 FILLCELL_X32 FILLER_98_33 ();
 FILLCELL_X32 FILLER_98_65 ();
 FILLCELL_X32 FILLER_98_97 ();
 FILLCELL_X32 FILLER_98_129 ();
 FILLCELL_X32 FILLER_98_161 ();
 FILLCELL_X32 FILLER_98_193 ();
 FILLCELL_X32 FILLER_98_225 ();
 FILLCELL_X32 FILLER_98_257 ();
 FILLCELL_X32 FILLER_98_289 ();
 FILLCELL_X32 FILLER_98_321 ();
 FILLCELL_X32 FILLER_98_353 ();
 FILLCELL_X32 FILLER_98_385 ();
 FILLCELL_X32 FILLER_98_417 ();
 FILLCELL_X32 FILLER_98_449 ();
 FILLCELL_X32 FILLER_98_481 ();
 FILLCELL_X32 FILLER_98_513 ();
 FILLCELL_X32 FILLER_98_545 ();
 FILLCELL_X32 FILLER_98_577 ();
 FILLCELL_X16 FILLER_98_609 ();
 FILLCELL_X4 FILLER_98_625 ();
 FILLCELL_X2 FILLER_98_629 ();
 FILLCELL_X32 FILLER_98_632 ();
 FILLCELL_X32 FILLER_98_664 ();
 FILLCELL_X32 FILLER_98_696 ();
 FILLCELL_X32 FILLER_98_728 ();
 FILLCELL_X16 FILLER_98_760 ();
 FILLCELL_X8 FILLER_98_776 ();
 FILLCELL_X4 FILLER_98_784 ();
 FILLCELL_X2 FILLER_98_788 ();
 FILLCELL_X32 FILLER_99_1 ();
 FILLCELL_X32 FILLER_99_33 ();
 FILLCELL_X32 FILLER_99_65 ();
 FILLCELL_X32 FILLER_99_97 ();
 FILLCELL_X32 FILLER_99_129 ();
 FILLCELL_X32 FILLER_99_161 ();
 FILLCELL_X32 FILLER_99_193 ();
 FILLCELL_X32 FILLER_99_225 ();
 FILLCELL_X32 FILLER_99_257 ();
 FILLCELL_X32 FILLER_99_289 ();
 FILLCELL_X32 FILLER_99_321 ();
 FILLCELL_X32 FILLER_99_353 ();
 FILLCELL_X32 FILLER_99_385 ();
 FILLCELL_X32 FILLER_99_417 ();
 FILLCELL_X32 FILLER_99_449 ();
 FILLCELL_X32 FILLER_99_481 ();
 FILLCELL_X32 FILLER_99_513 ();
 FILLCELL_X32 FILLER_99_545 ();
 FILLCELL_X32 FILLER_99_577 ();
 FILLCELL_X32 FILLER_99_609 ();
 FILLCELL_X32 FILLER_99_641 ();
 FILLCELL_X32 FILLER_99_673 ();
 FILLCELL_X32 FILLER_99_705 ();
 FILLCELL_X32 FILLER_99_737 ();
 FILLCELL_X16 FILLER_99_769 ();
 FILLCELL_X4 FILLER_99_785 ();
 FILLCELL_X1 FILLER_99_789 ();
 FILLCELL_X32 FILLER_100_1 ();
 FILLCELL_X32 FILLER_100_33 ();
 FILLCELL_X32 FILLER_100_65 ();
 FILLCELL_X32 FILLER_100_97 ();
 FILLCELL_X32 FILLER_100_129 ();
 FILLCELL_X32 FILLER_100_161 ();
 FILLCELL_X32 FILLER_100_193 ();
 FILLCELL_X32 FILLER_100_225 ();
 FILLCELL_X32 FILLER_100_257 ();
 FILLCELL_X32 FILLER_100_289 ();
 FILLCELL_X32 FILLER_100_321 ();
 FILLCELL_X32 FILLER_100_353 ();
 FILLCELL_X32 FILLER_100_385 ();
 FILLCELL_X32 FILLER_100_417 ();
 FILLCELL_X32 FILLER_100_449 ();
 FILLCELL_X32 FILLER_100_481 ();
 FILLCELL_X32 FILLER_100_513 ();
 FILLCELL_X32 FILLER_100_545 ();
 FILLCELL_X32 FILLER_100_577 ();
 FILLCELL_X16 FILLER_100_609 ();
 FILLCELL_X4 FILLER_100_625 ();
 FILLCELL_X2 FILLER_100_629 ();
 FILLCELL_X32 FILLER_100_632 ();
 FILLCELL_X32 FILLER_100_664 ();
 FILLCELL_X32 FILLER_100_696 ();
 FILLCELL_X32 FILLER_100_728 ();
 FILLCELL_X16 FILLER_100_760 ();
 FILLCELL_X8 FILLER_100_776 ();
 FILLCELL_X4 FILLER_100_784 ();
 FILLCELL_X2 FILLER_100_788 ();
 FILLCELL_X32 FILLER_101_1 ();
 FILLCELL_X32 FILLER_101_33 ();
 FILLCELL_X32 FILLER_101_65 ();
 FILLCELL_X32 FILLER_101_97 ();
 FILLCELL_X32 FILLER_101_129 ();
 FILLCELL_X32 FILLER_101_161 ();
 FILLCELL_X32 FILLER_101_193 ();
 FILLCELL_X32 FILLER_101_225 ();
 FILLCELL_X32 FILLER_101_257 ();
 FILLCELL_X32 FILLER_101_289 ();
 FILLCELL_X32 FILLER_101_321 ();
 FILLCELL_X32 FILLER_101_353 ();
 FILLCELL_X32 FILLER_101_385 ();
 FILLCELL_X32 FILLER_101_417 ();
 FILLCELL_X32 FILLER_101_449 ();
 FILLCELL_X32 FILLER_101_481 ();
 FILLCELL_X32 FILLER_101_513 ();
 FILLCELL_X32 FILLER_101_545 ();
 FILLCELL_X32 FILLER_101_577 ();
 FILLCELL_X32 FILLER_101_609 ();
 FILLCELL_X32 FILLER_101_641 ();
 FILLCELL_X32 FILLER_101_673 ();
 FILLCELL_X32 FILLER_101_705 ();
 FILLCELL_X32 FILLER_101_737 ();
 FILLCELL_X16 FILLER_101_769 ();
 FILLCELL_X4 FILLER_101_785 ();
 FILLCELL_X1 FILLER_101_789 ();
 FILLCELL_X32 FILLER_102_1 ();
 FILLCELL_X32 FILLER_102_33 ();
 FILLCELL_X32 FILLER_102_65 ();
 FILLCELL_X32 FILLER_102_97 ();
 FILLCELL_X32 FILLER_102_129 ();
 FILLCELL_X32 FILLER_102_161 ();
 FILLCELL_X32 FILLER_102_193 ();
 FILLCELL_X32 FILLER_102_225 ();
 FILLCELL_X32 FILLER_102_257 ();
 FILLCELL_X32 FILLER_102_289 ();
 FILLCELL_X32 FILLER_102_321 ();
 FILLCELL_X32 FILLER_102_353 ();
 FILLCELL_X32 FILLER_102_385 ();
 FILLCELL_X32 FILLER_102_417 ();
 FILLCELL_X32 FILLER_102_449 ();
 FILLCELL_X32 FILLER_102_481 ();
 FILLCELL_X32 FILLER_102_513 ();
 FILLCELL_X32 FILLER_102_545 ();
 FILLCELL_X32 FILLER_102_577 ();
 FILLCELL_X16 FILLER_102_609 ();
 FILLCELL_X4 FILLER_102_625 ();
 FILLCELL_X2 FILLER_102_629 ();
 FILLCELL_X32 FILLER_102_632 ();
 FILLCELL_X32 FILLER_102_664 ();
 FILLCELL_X32 FILLER_102_696 ();
 FILLCELL_X32 FILLER_102_728 ();
 FILLCELL_X16 FILLER_102_760 ();
 FILLCELL_X8 FILLER_102_776 ();
 FILLCELL_X4 FILLER_102_784 ();
 FILLCELL_X2 FILLER_102_788 ();
 FILLCELL_X32 FILLER_103_1 ();
 FILLCELL_X32 FILLER_103_33 ();
 FILLCELL_X32 FILLER_103_65 ();
 FILLCELL_X32 FILLER_103_97 ();
 FILLCELL_X32 FILLER_103_129 ();
 FILLCELL_X32 FILLER_103_161 ();
 FILLCELL_X32 FILLER_103_193 ();
 FILLCELL_X32 FILLER_103_225 ();
 FILLCELL_X32 FILLER_103_257 ();
 FILLCELL_X32 FILLER_103_289 ();
 FILLCELL_X32 FILLER_103_321 ();
 FILLCELL_X32 FILLER_103_353 ();
 FILLCELL_X32 FILLER_103_385 ();
 FILLCELL_X32 FILLER_103_417 ();
 FILLCELL_X32 FILLER_103_449 ();
 FILLCELL_X32 FILLER_103_481 ();
 FILLCELL_X32 FILLER_103_513 ();
 FILLCELL_X32 FILLER_103_545 ();
 FILLCELL_X32 FILLER_103_577 ();
 FILLCELL_X32 FILLER_103_609 ();
 FILLCELL_X32 FILLER_103_641 ();
 FILLCELL_X32 FILLER_103_673 ();
 FILLCELL_X32 FILLER_103_705 ();
 FILLCELL_X32 FILLER_103_737 ();
 FILLCELL_X16 FILLER_103_769 ();
 FILLCELL_X4 FILLER_103_785 ();
 FILLCELL_X1 FILLER_103_789 ();
 FILLCELL_X32 FILLER_104_1 ();
 FILLCELL_X32 FILLER_104_33 ();
 FILLCELL_X32 FILLER_104_65 ();
 FILLCELL_X32 FILLER_104_97 ();
 FILLCELL_X32 FILLER_104_129 ();
 FILLCELL_X32 FILLER_104_161 ();
 FILLCELL_X32 FILLER_104_193 ();
 FILLCELL_X32 FILLER_104_225 ();
 FILLCELL_X32 FILLER_104_257 ();
 FILLCELL_X32 FILLER_104_289 ();
 FILLCELL_X32 FILLER_104_321 ();
 FILLCELL_X32 FILLER_104_353 ();
 FILLCELL_X16 FILLER_104_385 ();
 FILLCELL_X8 FILLER_104_401 ();
 FILLCELL_X2 FILLER_104_409 ();
 FILLCELL_X32 FILLER_104_416 ();
 FILLCELL_X32 FILLER_104_448 ();
 FILLCELL_X32 FILLER_104_480 ();
 FILLCELL_X32 FILLER_104_512 ();
 FILLCELL_X32 FILLER_104_544 ();
 FILLCELL_X32 FILLER_104_576 ();
 FILLCELL_X16 FILLER_104_608 ();
 FILLCELL_X4 FILLER_104_624 ();
 FILLCELL_X2 FILLER_104_628 ();
 FILLCELL_X1 FILLER_104_630 ();
 FILLCELL_X32 FILLER_104_632 ();
 FILLCELL_X32 FILLER_104_664 ();
 FILLCELL_X32 FILLER_104_696 ();
 FILLCELL_X32 FILLER_104_728 ();
 FILLCELL_X16 FILLER_104_760 ();
 FILLCELL_X8 FILLER_104_776 ();
 FILLCELL_X4 FILLER_104_784 ();
 FILLCELL_X2 FILLER_104_788 ();
 FILLCELL_X32 FILLER_105_1 ();
 FILLCELL_X32 FILLER_105_33 ();
 FILLCELL_X32 FILLER_105_65 ();
 FILLCELL_X32 FILLER_105_97 ();
 FILLCELL_X32 FILLER_105_129 ();
 FILLCELL_X32 FILLER_105_161 ();
 FILLCELL_X32 FILLER_105_193 ();
 FILLCELL_X32 FILLER_105_225 ();
 FILLCELL_X32 FILLER_105_257 ();
 FILLCELL_X32 FILLER_105_289 ();
 FILLCELL_X32 FILLER_105_321 ();
 FILLCELL_X32 FILLER_105_353 ();
 FILLCELL_X16 FILLER_105_385 ();
 FILLCELL_X4 FILLER_105_401 ();
 FILLCELL_X2 FILLER_105_418 ();
 FILLCELL_X4 FILLER_105_427 ();
 FILLCELL_X32 FILLER_105_439 ();
 FILLCELL_X32 FILLER_105_471 ();
 FILLCELL_X32 FILLER_105_503 ();
 FILLCELL_X32 FILLER_105_535 ();
 FILLCELL_X32 FILLER_105_567 ();
 FILLCELL_X32 FILLER_105_599 ();
 FILLCELL_X32 FILLER_105_631 ();
 FILLCELL_X32 FILLER_105_663 ();
 FILLCELL_X32 FILLER_105_695 ();
 FILLCELL_X32 FILLER_105_727 ();
 FILLCELL_X16 FILLER_105_759 ();
 FILLCELL_X8 FILLER_105_775 ();
 FILLCELL_X4 FILLER_105_783 ();
 FILLCELL_X2 FILLER_105_787 ();
 FILLCELL_X1 FILLER_105_789 ();
 FILLCELL_X32 FILLER_106_1 ();
 FILLCELL_X32 FILLER_106_33 ();
 FILLCELL_X32 FILLER_106_65 ();
 FILLCELL_X32 FILLER_106_97 ();
 FILLCELL_X32 FILLER_106_129 ();
 FILLCELL_X32 FILLER_106_161 ();
 FILLCELL_X32 FILLER_106_193 ();
 FILLCELL_X32 FILLER_106_225 ();
 FILLCELL_X32 FILLER_106_257 ();
 FILLCELL_X32 FILLER_106_289 ();
 FILLCELL_X32 FILLER_106_321 ();
 FILLCELL_X32 FILLER_106_353 ();
 FILLCELL_X4 FILLER_106_385 ();
 FILLCELL_X1 FILLER_106_389 ();
 FILLCELL_X16 FILLER_106_396 ();
 FILLCELL_X1 FILLER_106_412 ();
 FILLCELL_X8 FILLER_106_416 ();
 FILLCELL_X4 FILLER_106_437 ();
 FILLCELL_X2 FILLER_106_441 ();
 FILLCELL_X8 FILLER_106_446 ();
 FILLCELL_X1 FILLER_106_454 ();
 FILLCELL_X32 FILLER_106_459 ();
 FILLCELL_X32 FILLER_106_491 ();
 FILLCELL_X32 FILLER_106_523 ();
 FILLCELL_X32 FILLER_106_555 ();
 FILLCELL_X32 FILLER_106_587 ();
 FILLCELL_X8 FILLER_106_619 ();
 FILLCELL_X4 FILLER_106_627 ();
 FILLCELL_X32 FILLER_106_632 ();
 FILLCELL_X32 FILLER_106_664 ();
 FILLCELL_X32 FILLER_106_696 ();
 FILLCELL_X32 FILLER_106_728 ();
 FILLCELL_X16 FILLER_106_760 ();
 FILLCELL_X8 FILLER_106_776 ();
 FILLCELL_X4 FILLER_106_784 ();
 FILLCELL_X2 FILLER_106_788 ();
endmodule
