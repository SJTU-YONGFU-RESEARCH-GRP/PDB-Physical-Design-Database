module floating_point_adder (clk,
    inexact,
    invalid_op,
    overflow,
    rst_n,
    underflow,
    valid_in,
    valid_out,
    a,
    b,
    result);
 input clk;
 output inexact;
 output invalid_op;
 output overflow;
 input rst_n;
 output underflow;
 input valid_in;
 output valid_out;
 input [31:0] a;
 input [31:0] b;
 output [31:0] result;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire a_exp_larger;
 wire a_sign_stage1;
 wire \add_result[10] ;
 wire \add_result[11] ;
 wire \add_result[12] ;
 wire \add_result[13] ;
 wire \add_result[14] ;
 wire \add_result[15] ;
 wire \add_result[16] ;
 wire \add_result[17] ;
 wire \add_result[18] ;
 wire \add_result[19] ;
 wire \add_result[20] ;
 wire \add_result[21] ;
 wire \add_result[22] ;
 wire \add_result[23] ;
 wire \add_result[24] ;
 wire \add_result[25] ;
 wire \add_result[26] ;
 wire \add_result[2] ;
 wire \add_result[3] ;
 wire \add_result[4] ;
 wire \add_result[5] ;
 wire \add_result[6] ;
 wire \add_result[7] ;
 wire \add_result[8] ;
 wire \add_result[9] ;
 wire \aligned_a_mant[0] ;
 wire \aligned_a_mant[10] ;
 wire \aligned_a_mant[11] ;
 wire \aligned_a_mant[12] ;
 wire \aligned_a_mant[13] ;
 wire \aligned_a_mant[14] ;
 wire \aligned_a_mant[15] ;
 wire \aligned_a_mant[16] ;
 wire \aligned_a_mant[17] ;
 wire \aligned_a_mant[18] ;
 wire \aligned_a_mant[19] ;
 wire \aligned_a_mant[1] ;
 wire \aligned_a_mant[20] ;
 wire \aligned_a_mant[21] ;
 wire \aligned_a_mant[22] ;
 wire \aligned_a_mant[23] ;
 wire \aligned_a_mant[24] ;
 wire \aligned_a_mant[25] ;
 wire \aligned_a_mant[2] ;
 wire \aligned_a_mant[3] ;
 wire \aligned_a_mant[4] ;
 wire \aligned_a_mant[5] ;
 wire \aligned_a_mant[6] ;
 wire \aligned_a_mant[7] ;
 wire \aligned_a_mant[8] ;
 wire \aligned_a_mant[9] ;
 wire \aligned_b_mant[0] ;
 wire \aligned_b_mant[10] ;
 wire \aligned_b_mant[11] ;
 wire \aligned_b_mant[12] ;
 wire \aligned_b_mant[13] ;
 wire \aligned_b_mant[14] ;
 wire \aligned_b_mant[15] ;
 wire \aligned_b_mant[16] ;
 wire \aligned_b_mant[17] ;
 wire \aligned_b_mant[18] ;
 wire \aligned_b_mant[19] ;
 wire \aligned_b_mant[1] ;
 wire \aligned_b_mant[20] ;
 wire \aligned_b_mant[21] ;
 wire \aligned_b_mant[22] ;
 wire \aligned_b_mant[23] ;
 wire \aligned_b_mant[24] ;
 wire \aligned_b_mant[25] ;
 wire \aligned_b_mant[2] ;
 wire \aligned_b_mant[3] ;
 wire \aligned_b_mant[4] ;
 wire \aligned_b_mant[5] ;
 wire \aligned_b_mant[6] ;
 wire \aligned_b_mant[7] ;
 wire \aligned_b_mant[8] ;
 wire \aligned_b_mant[9] ;
 wire b_sign_stage1;
 wire \final_exp[0] ;
 wire \final_exp[1] ;
 wire \final_exp[2] ;
 wire \final_exp[3] ;
 wire \final_exp[4] ;
 wire \final_exp[5] ;
 wire \final_exp[6] ;
 wire \final_exp[7] ;
 wire \final_mant[0] ;
 wire \final_mant[10] ;
 wire \final_mant[11] ;
 wire \final_mant[12] ;
 wire \final_mant[13] ;
 wire \final_mant[14] ;
 wire \final_mant[15] ;
 wire \final_mant[16] ;
 wire \final_mant[17] ;
 wire \final_mant[18] ;
 wire \final_mant[19] ;
 wire \final_mant[1] ;
 wire \final_mant[20] ;
 wire \final_mant[21] ;
 wire \final_mant[22] ;
 wire \final_mant[2] ;
 wire \final_mant[3] ;
 wire \final_mant[4] ;
 wire \final_mant[5] ;
 wire \final_mant[6] ;
 wire \final_mant[7] ;
 wire \final_mant[8] ;
 wire \final_mant[9] ;
 wire inexact_stage2;
 wire invalid_op_stage2;
 wire is_a_larger_stage1;
 wire \larger_exp_stage1[0] ;
 wire \larger_exp_stage1[1] ;
 wire \larger_exp_stage1[2] ;
 wire \larger_exp_stage1[3] ;
 wire \larger_exp_stage1[4] ;
 wire \larger_exp_stage1[5] ;
 wire \larger_exp_stage1[6] ;
 wire \larger_exp_stage1[7] ;
 wire \result_exp_stage2[0] ;
 wire \result_exp_stage2[1] ;
 wire \result_exp_stage2[2] ;
 wire \result_exp_stage2[3] ;
 wire \result_exp_stage2[4] ;
 wire \result_exp_stage2[5] ;
 wire \result_exp_stage2[6] ;
 wire \result_exp_stage2[7] ;
 wire result_sign_stage2;
 wire valid_stage1;
 wire valid_stage2;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net105;
 wire net106;
 wire net107;

 sky130_fd_sc_hd__o22ai_2 _1920_ (.A1(_1267_),
    .A2(_1268_),
    .B1(_1354_),
    .B2(_1355_),
    .Y(_1356_));
 sky130_fd_sc_hd__nor2b_1 _1921_ (.A(_1571_),
    .B_N(_1269_),
    .Y(_1357_));
 sky130_fd_sc_hd__nor2b_1 _1922_ (.A(_1269_),
    .B_N(_1571_),
    .Y(_1358_));
 sky130_fd_sc_hd__clkbuf_4 _1923_ (.A(_1233_),
    .X(_1359_));
 sky130_fd_sc_hd__clkbuf_4 _1924_ (.A(_1248_),
    .X(_1360_));
 sky130_fd_sc_hd__o211ai_2 _1925_ (.A1(_1357_),
    .A2(_1358_),
    .B1(_1359_),
    .C1(_1360_),
    .Y(_1361_));
 sky130_fd_sc_hd__and2_0 _1926_ (.A(_1356_),
    .B(_1361_),
    .X(_1362_));
 sky130_fd_sc_hd__clkbuf_4 _1927_ (.A(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__buf_4 _1928_ (.A(_1299_),
    .X(_1364_));
 sky130_fd_sc_hd__mux4_1 _1929_ (.A0(_1331_),
    .A1(_1335_),
    .A2(_1347_),
    .A3(_1353_),
    .S0(_1363_),
    .S1(_1364_),
    .X(_1365_));
 sky130_fd_sc_hd__and2_0 _1930_ (.A(_1274_),
    .B(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__nand2_1 _1931_ (.A(_1269_),
    .B(_1571_),
    .Y(_1367_));
 sky130_fd_sc_hd__or2_0 _1932_ (.A(_1269_),
    .B(_1571_),
    .X(_1368_));
 sky130_fd_sc_hd__a22o_1 _1933_ (.A1(_1299_),
    .A2(_1572_),
    .B1(_1367_),
    .B2(_1368_),
    .X(_1369_));
 sky130_fd_sc_hd__nand2_2 _1934_ (.A(_1234_),
    .B(_1235_),
    .Y(_1370_));
 sky130_fd_sc_hd__xnor2_1 _1935_ (.A(_1263_),
    .B(_1370_),
    .Y(_1371_));
 sky130_fd_sc_hd__nor2_1 _1936_ (.A(_1310_),
    .B(_1601_),
    .Y(_1372_));
 sky130_fd_sc_hd__a311o_1 _1937_ (.A1(_1271_),
    .A2(_1369_),
    .A3(_1371_),
    .B1(_1372_),
    .C1(_1238_),
    .X(_1373_));
 sky130_fd_sc_hd__a21oi_1 _1938_ (.A1(_1204_),
    .A2(_1370_),
    .B1(_1607_),
    .Y(_1374_));
 sky130_fd_sc_hd__nand3b_1 _1939_ (.A_N(_1271_),
    .B(_1369_),
    .C(_1371_),
    .Y(_1375_));
 sky130_fd_sc_hd__o211ai_1 _1940_ (.A1(_1239_),
    .A2(_1374_),
    .B1(_1375_),
    .C1(_1238_),
    .Y(_1376_));
 sky130_fd_sc_hd__and2_0 _1941_ (.A(_1374_),
    .B(_1372_),
    .X(_1377_));
 sky130_fd_sc_hd__a221o_2 _1942_ (.A1(_1310_),
    .A2(_1601_),
    .B1(_1373_),
    .B2(_1376_),
    .C1(_1377_),
    .X(_1378_));
 sky130_fd_sc_hd__nand3_4 _1943_ (.A(_1359_),
    .B(_1360_),
    .C(_1328_),
    .Y(_1379_));
 sky130_fd_sc_hd__nor3_4 _1944_ (.A(_1378_),
    .B(_1341_),
    .C(_1379_),
    .Y(_1380_));
 sky130_fd_sc_hd__mux2i_4 _1945_ (.A0(_1370_),
    .A1(_1296_),
    .S(_1249_),
    .Y(_1381_));
 sky130_fd_sc_hd__xnor2_4 _1946_ (.A(_1204_),
    .B(_1381_),
    .Y(_1382_));
 sky130_fd_sc_hd__nor2_4 _1947_ (.A(_1330_),
    .B(_1293_),
    .Y(_1383_));
 sky130_fd_sc_hd__a2111oi_1 _1948_ (.A1(_1367_),
    .A2(_1368_),
    .B1(_1318_),
    .C1(_1267_),
    .D1(_1268_),
    .Y(_1384_));
 sky130_fd_sc_hd__a221oi_1 _1949_ (.A1(_1359_),
    .A2(_1360_),
    .B1(_1300_),
    .B2(_1301_),
    .C1(_1344_),
    .Y(_1385_));
 sky130_fd_sc_hd__nor2_2 _1950_ (.A(_1384_),
    .B(_1385_),
    .Y(_1386_));
 sky130_fd_sc_hd__mux2_1 _1951_ (.A0(net16),
    .A1(_1180_),
    .S(_1299_),
    .X(_1387_));
 sky130_fd_sc_hd__nand2_1 _1952_ (.A(net48),
    .B(_1298_),
    .Y(_1388_));
 sky130_fd_sc_hd__o21ai_1 _1953_ (.A1(_1298_),
    .A2(_1192_),
    .B1(_1388_),
    .Y(_1389_));
 sky130_fd_sc_hd__a2111o_1 _1954_ (.A1(_1233_),
    .A2(_1248_),
    .B1(_1341_),
    .C1(_1292_),
    .D1(_1342_),
    .X(_1390_));
 sky130_fd_sc_hd__buf_6 _1955_ (.A(_1390_),
    .X(_1391_));
 sky130_fd_sc_hd__mux2i_4 _1956_ (.A0(_1387_),
    .A1(_1389_),
    .S(_1391_),
    .Y(_1392_));
 sky130_fd_sc_hd__nor3_4 _1957_ (.A(_1383_),
    .B(_1386_),
    .C(_1392_),
    .Y(_1393_));
 sky130_fd_sc_hd__xnor2_2 _1958_ (.A(_1308_),
    .B(_1273_),
    .Y(_1394_));
 sky130_fd_sc_hd__nand2b_1 _1959_ (.A_N(_1393_),
    .B(_1394_),
    .Y(_1395_));
 sky130_fd_sc_hd__nand3_1 _1960_ (.A(_1380_),
    .B(_1382_),
    .C(_1395_),
    .Y(_1396_));
 sky130_fd_sc_hd__xnor2_4 _1961_ (.A(_1263_),
    .B(_1381_),
    .Y(_1397_));
 sky130_fd_sc_hd__nand2_2 _1962_ (.A(_1380_),
    .B(_1397_),
    .Y(_1398_));
 sky130_fd_sc_hd__buf_4 _1963_ (.A(_1394_),
    .X(_1399_));
 sky130_fd_sc_hd__buf_4 _1964_ (.A(_1364_),
    .X(_1400_));
 sky130_fd_sc_hd__buf_4 _1965_ (.A(_1363_),
    .X(_1401_));
 sky130_fd_sc_hd__clkbuf_4 _1966_ (.A(_1401_),
    .X(_1402_));
 sky130_fd_sc_hd__nor2_2 _1967_ (.A(_1341_),
    .B(_1342_),
    .Y(_1403_));
 sky130_fd_sc_hd__nand2_4 _1968_ (.A(_1293_),
    .B(_1403_),
    .Y(_1404_));
 sky130_fd_sc_hd__clkbuf_4 _1969_ (.A(_1344_),
    .X(_1405_));
 sky130_fd_sc_hd__mux2i_2 _1970_ (.A0(net12),
    .A1(net15),
    .S(_1405_),
    .Y(_1406_));
 sky130_fd_sc_hd__clkbuf_4 _1971_ (.A(_1318_),
    .X(_1407_));
 sky130_fd_sc_hd__mux2i_2 _1972_ (.A0(net44),
    .A1(net47),
    .S(_1407_),
    .Y(_1408_));
 sky130_fd_sc_hd__mux2i_1 _1973_ (.A0(net44),
    .A1(net47),
    .S(_1344_),
    .Y(_1409_));
 sky130_fd_sc_hd__or4_1 _1974_ (.A(a_exp_larger),
    .B(_1292_),
    .C(_1343_),
    .D(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__o221ai_4 _1975_ (.A1(_1404_),
    .A2(_1406_),
    .B1(_1408_),
    .B2(_1379_),
    .C1(_1410_),
    .Y(_1411_));
 sky130_fd_sc_hd__buf_4 _1976_ (.A(_1293_),
    .X(_1412_));
 sky130_fd_sc_hd__buf_4 _1977_ (.A(_1294_),
    .X(_1413_));
 sky130_fd_sc_hd__mux2i_1 _1978_ (.A0(net8),
    .A1(net10),
    .S(_1413_),
    .Y(_1414_));
 sky130_fd_sc_hd__nand3_1 _1979_ (.A(_1295_),
    .B(_1315_),
    .C(_1414_),
    .Y(_1415_));
 sky130_fd_sc_hd__nand2_1 _1980_ (.A(net42),
    .B(_1413_),
    .Y(_1416_));
 sky130_fd_sc_hd__o221ai_4 _1981_ (.A1(_1643_),
    .A2(_1413_),
    .B1(_1341_),
    .B2(_1342_),
    .C1(_1416_),
    .Y(_1417_));
 sky130_fd_sc_hd__nand2_1 _1982_ (.A(net42),
    .B(_1319_),
    .Y(_1418_));
 sky130_fd_sc_hd__o21ai_1 _1983_ (.A1(_1643_),
    .A2(_1407_),
    .B1(_1418_),
    .Y(_1419_));
 sky130_fd_sc_hd__a32oi_4 _1984_ (.A1(_1412_),
    .A2(_1415_),
    .A3(_1417_),
    .B1(_1419_),
    .B2(_1330_),
    .Y(_1420_));
 sky130_fd_sc_hd__nand2_1 _1985_ (.A(_1363_),
    .B(_1420_),
    .Y(_1421_));
 sky130_fd_sc_hd__o21a_1 _1986_ (.A1(_1402_),
    .A2(_1411_),
    .B1(_1421_),
    .X(_1422_));
 sky130_fd_sc_hd__nand4_1 _1987_ (.A(_1319_),
    .B(_1359_),
    .C(_1360_),
    .D(_1328_),
    .Y(_1423_));
 sky130_fd_sc_hd__inv_1 _1988_ (.A(_1294_),
    .Y(_1424_));
 sky130_fd_sc_hd__a211o_1 _1989_ (.A1(_1359_),
    .A2(_1360_),
    .B1(_1292_),
    .C1(_1424_),
    .X(_1425_));
 sky130_fd_sc_hd__inv_1 _1990_ (.A(net14),
    .Y(_1426_));
 sky130_fd_sc_hd__a21oi_1 _1991_ (.A1(_1423_),
    .A2(_1425_),
    .B1(_1426_),
    .Y(_1427_));
 sky130_fd_sc_hd__inv_1 _1992_ (.A(_1318_),
    .Y(_1428_));
 sky130_fd_sc_hd__nand4_2 _1993_ (.A(_1428_),
    .B(_1359_),
    .C(_1360_),
    .D(_1328_),
    .Y(_1429_));
 sky130_fd_sc_hd__a211o_1 _1994_ (.A1(_1359_),
    .A2(_1360_),
    .B1(_1292_),
    .C1(_1344_),
    .X(_1430_));
 sky130_fd_sc_hd__inv_1 _1995_ (.A(net11),
    .Y(_1431_));
 sky130_fd_sc_hd__a21oi_1 _1996_ (.A1(_1429_),
    .A2(_1430_),
    .B1(_1431_),
    .Y(_1432_));
 sky130_fd_sc_hd__o21ai_2 _1997_ (.A1(_1427_),
    .A2(_1432_),
    .B1(_1337_),
    .Y(_1433_));
 sky130_fd_sc_hd__a21oi_1 _1998_ (.A1(_1429_),
    .A2(_1430_),
    .B1(_1670_),
    .Y(_1434_));
 sky130_fd_sc_hd__a21oi_1 _1999_ (.A1(_1423_),
    .A2(_1425_),
    .B1(_1685_),
    .Y(_1435_));
 sky130_fd_sc_hd__o21ai_2 _2000_ (.A1(_1434_),
    .A2(_1435_),
    .B1(_1404_),
    .Y(_1436_));
 sky130_fd_sc_hd__nand2_4 _2001_ (.A(_1356_),
    .B(_1361_),
    .Y(_1437_));
 sky130_fd_sc_hd__clkbuf_4 _2002_ (.A(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__nand2_1 _2003_ (.A(net41),
    .B(_1413_),
    .Y(_1439_));
 sky130_fd_sc_hd__o221ai_4 _2004_ (.A1(_1646_),
    .A2(_1413_),
    .B1(_1336_),
    .B2(_1316_),
    .C1(_1439_),
    .Y(_1440_));
 sky130_fd_sc_hd__mux2i_1 _2005_ (.A0(net7),
    .A1(net9),
    .S(_1413_),
    .Y(_1441_));
 sky130_fd_sc_hd__nand3_1 _2006_ (.A(_1293_),
    .B(_1403_),
    .C(_1441_),
    .Y(_1442_));
 sky130_fd_sc_hd__mux2i_1 _2007_ (.A0(net39),
    .A1(net41),
    .S(_1319_),
    .Y(_1443_));
 sky130_fd_sc_hd__nor2_1 _2008_ (.A(_1379_),
    .B(_1443_),
    .Y(_1444_));
 sky130_fd_sc_hd__a311oi_2 _2009_ (.A1(_1412_),
    .A2(_1440_),
    .A3(_1442_),
    .B1(_1444_),
    .C1(_1437_),
    .Y(_1445_));
 sky130_fd_sc_hd__a311oi_2 _2010_ (.A1(_1433_),
    .A2(_1436_),
    .A3(_1438_),
    .B1(_1445_),
    .C1(_1400_),
    .Y(_1446_));
 sky130_fd_sc_hd__a21oi_4 _2011_ (.A1(_1400_),
    .A2(_1422_),
    .B1(_1446_),
    .Y(_1447_));
 sky130_fd_sc_hd__buf_4 _2012_ (.A(_1391_),
    .X(_1448_));
 sky130_fd_sc_hd__nand2_1 _2013_ (.A(net60),
    .B(_1448_),
    .Y(_1449_));
 sky130_fd_sc_hd__buf_4 _2014_ (.A(_1343_),
    .X(_1450_));
 sky130_fd_sc_hd__nand2_1 _2015_ (.A(net28),
    .B(_1450_),
    .Y(_1451_));
 sky130_fd_sc_hd__nand3_2 _2016_ (.A(_1318_),
    .B(_1359_),
    .C(_1360_),
    .Y(_1452_));
 sky130_fd_sc_hd__o21ai_2 _2017_ (.A1(_1267_),
    .A2(_1268_),
    .B1(_1344_),
    .Y(_1453_));
 sky130_fd_sc_hd__and2_0 _2018_ (.A(_1452_),
    .B(_1453_),
    .X(_1454_));
 sky130_fd_sc_hd__buf_2 _2019_ (.A(_1454_),
    .X(_1455_));
 sky130_fd_sc_hd__a21oi_1 _2020_ (.A1(_1449_),
    .A2(_1451_),
    .B1(_1455_),
    .Y(_1456_));
 sky130_fd_sc_hd__nand2_1 _2021_ (.A(net56),
    .B(_1448_),
    .Y(_1457_));
 sky130_fd_sc_hd__nand2_1 _2022_ (.A(net24),
    .B(_1450_),
    .Y(_1458_));
 sky130_fd_sc_hd__nand2_8 _2023_ (.A(_1452_),
    .B(_1453_),
    .Y(_1459_));
 sky130_fd_sc_hd__a21oi_1 _2024_ (.A1(_1457_),
    .A2(_1458_),
    .B1(_1459_),
    .Y(_1460_));
 sky130_fd_sc_hd__nor2_1 _2025_ (.A(_1456_),
    .B(_1460_),
    .Y(_1461_));
 sky130_fd_sc_hd__nand2_4 _2026_ (.A(_1429_),
    .B(_1430_),
    .Y(_1462_));
 sky130_fd_sc_hd__mux2_1 _2027_ (.A0(net27),
    .A1(net59),
    .S(_1391_),
    .X(_1463_));
 sky130_fd_sc_hd__mux2_1 _2028_ (.A0(net29),
    .A1(net61),
    .S(_1391_),
    .X(_1464_));
 sky130_fd_sc_hd__nand2_2 _2029_ (.A(_1423_),
    .B(_1425_),
    .Y(_1465_));
 sky130_fd_sc_hd__a22oi_2 _2030_ (.A1(_1462_),
    .A2(_1463_),
    .B1(_1464_),
    .B2(_1465_),
    .Y(_1466_));
 sky130_fd_sc_hd__nor2_1 _2031_ (.A(_1298_),
    .B(_1363_),
    .Y(_1467_));
 sky130_fd_sc_hd__nand2b_1 _2032_ (.A_N(_1466_),
    .B(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__o41ai_1 _2033_ (.A1(_1400_),
    .A2(_1383_),
    .A3(_1402_),
    .A4(_1461_),
    .B1(_1468_),
    .Y(_1469_));
 sky130_fd_sc_hd__clkbuf_4 _2034_ (.A(_1274_),
    .X(_1470_));
 sky130_fd_sc_hd__mux4_1 _2035_ (.A0(net13),
    .A1(net2),
    .A2(net45),
    .A3(net34),
    .S0(_1298_),
    .S1(_1404_),
    .X(_1471_));
 sky130_fd_sc_hd__nand3_1 _2036_ (.A(_1465_),
    .B(_1402_),
    .C(_1471_),
    .Y(_1472_));
 sky130_fd_sc_hd__nand2_1 _2037_ (.A(_1470_),
    .B(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hd__o2bb2ai_1 _2038_ (.A1_N(_1399_),
    .A2_N(_1447_),
    .B1(_1469_),
    .B2(_1473_),
    .Y(_1474_));
 sky130_fd_sc_hd__o22ai_1 _2039_ (.A1(_1366_),
    .A2(_1396_),
    .B1(_1398_),
    .B2(_1474_),
    .Y(_0051_));
 sky130_fd_sc_hd__nand2_4 _2040_ (.A(_1379_),
    .B(_1336_),
    .Y(_1475_));
 sky130_fd_sc_hd__nand2_1 _2041_ (.A(net41),
    .B(_1424_),
    .Y(_1476_));
 sky130_fd_sc_hd__nand2_1 _2042_ (.A(net43),
    .B(_1294_),
    .Y(_1477_));
 sky130_fd_sc_hd__a22oi_1 _2043_ (.A1(_1359_),
    .A2(_1360_),
    .B1(_1476_),
    .B2(_1477_),
    .Y(_1478_));
 sky130_fd_sc_hd__nor4_1 _2044_ (.A(_1676_),
    .B(_1318_),
    .C(_1267_),
    .D(_1268_),
    .Y(_1479_));
 sky130_fd_sc_hd__a311o_1 _2045_ (.A1(net43),
    .A2(_1318_),
    .A3(a_exp_larger),
    .B1(_1478_),
    .C1(_1479_),
    .X(_1480_));
 sky130_fd_sc_hd__nand2_1 _2046_ (.A(net9),
    .B(_1424_),
    .Y(_1481_));
 sky130_fd_sc_hd__nand2_1 _2047_ (.A(net11),
    .B(_1344_),
    .Y(_1482_));
 sky130_fd_sc_hd__a22oi_1 _2048_ (.A1(_1359_),
    .A2(_1360_),
    .B1(_1481_),
    .B2(_1482_),
    .Y(_1483_));
 sky130_fd_sc_hd__nand2_1 _2049_ (.A(net9),
    .B(_1428_),
    .Y(_1484_));
 sky130_fd_sc_hd__nand2_1 _2050_ (.A(net11),
    .B(_1318_),
    .Y(_1485_));
 sky130_fd_sc_hd__a211oi_1 _2051_ (.A1(_1484_),
    .A2(_1485_),
    .B1(_1267_),
    .C1(_1268_),
    .Y(_1486_));
 sky130_fd_sc_hd__o21a_1 _2052_ (.A1(_1483_),
    .A2(_1486_),
    .B1(_1450_),
    .X(_1487_));
 sky130_fd_sc_hd__a31oi_4 _2053_ (.A1(_1475_),
    .A2(_1391_),
    .A3(_1480_),
    .B1(_1487_),
    .Y(_1488_));
 sky130_fd_sc_hd__clkbuf_4 _2054_ (.A(_1298_),
    .X(_1489_));
 sky130_fd_sc_hd__nor2_1 _2055_ (.A(_1489_),
    .B(_1437_),
    .Y(_1490_));
 sky130_fd_sc_hd__nand2_1 _2056_ (.A(_1298_),
    .B(_1437_),
    .Y(_1491_));
 sky130_fd_sc_hd__o22ai_2 _2057_ (.A1(_1491_),
    .A2(_1411_),
    .B1(_1421_),
    .B2(_1364_),
    .Y(_1492_));
 sky130_fd_sc_hd__mux2i_1 _2058_ (.A0(net14),
    .A1(net16),
    .S(_1459_),
    .Y(_1493_));
 sky130_fd_sc_hd__mux2i_1 _2059_ (.A0(net46),
    .A1(net48),
    .S(_1459_),
    .Y(_1494_));
 sky130_fd_sc_hd__nand2_1 _2060_ (.A(_1475_),
    .B(_1448_),
    .Y(_1495_));
 sky130_fd_sc_hd__o221a_1 _2061_ (.A1(_1448_),
    .A2(_1493_),
    .B1(_1494_),
    .B2(_1495_),
    .C1(_1467_),
    .X(_1496_));
 sky130_fd_sc_hd__a211oi_4 _2062_ (.A1(_1488_),
    .A2(_1490_),
    .B1(_1492_),
    .C1(_1496_),
    .Y(_1497_));
 sky130_fd_sc_hd__mux2i_1 _2063_ (.A0(net28),
    .A1(net30),
    .S(_1405_),
    .Y(_1498_));
 sky130_fd_sc_hd__nand3_1 _2064_ (.A(_1412_),
    .B(_1403_),
    .C(_1498_),
    .Y(_1499_));
 sky130_fd_sc_hd__nand2_1 _2065_ (.A(net62),
    .B(_1405_),
    .Y(_1500_));
 sky130_fd_sc_hd__o221ai_1 _2066_ (.A1(_1640_),
    .A2(_1405_),
    .B1(_1336_),
    .B2(_1316_),
    .C1(_1500_),
    .Y(_1501_));
 sky130_fd_sc_hd__mux2i_1 _2067_ (.A0(net60),
    .A1(net62),
    .S(_1407_),
    .Y(_1502_));
 sky130_fd_sc_hd__nor2_1 _2068_ (.A(_1379_),
    .B(_1502_),
    .Y(_1503_));
 sky130_fd_sc_hd__a31oi_2 _2069_ (.A1(_1412_),
    .A2(_1499_),
    .A3(_1501_),
    .B1(_1503_),
    .Y(_1504_));
 sky130_fd_sc_hd__mux2_1 _2070_ (.A0(_1466_),
    .A1(_1504_),
    .S(_1364_),
    .X(_1505_));
 sky130_fd_sc_hd__mux4_1 _2071_ (.A0(net13),
    .A1(net24),
    .A2(net45),
    .A3(net56),
    .S0(_1364_),
    .S1(_1404_),
    .X(_1506_));
 sky130_fd_sc_hd__nand2_1 _2072_ (.A(_1475_),
    .B(_1506_),
    .Y(_1507_));
 sky130_fd_sc_hd__nor2_1 _2073_ (.A(_1455_),
    .B(_1437_),
    .Y(_1508_));
 sky130_fd_sc_hd__mux2i_1 _2074_ (.A0(net2),
    .A1(net34),
    .S(_1448_),
    .Y(_1509_));
 sky130_fd_sc_hd__nor3_1 _2075_ (.A(_1489_),
    .B(_1383_),
    .C(_1509_),
    .Y(_1510_));
 sky130_fd_sc_hd__o211ai_1 _2076_ (.A1(_1386_),
    .A2(_1510_),
    .B1(_1274_),
    .C1(_1397_),
    .Y(_1511_));
 sky130_fd_sc_hd__a221oi_1 _2077_ (.A1(_1438_),
    .A2(_1505_),
    .B1(_1507_),
    .B2(_1508_),
    .C1(_1511_),
    .Y(_1512_));
 sky130_fd_sc_hd__nand2_1 _2078_ (.A(_1489_),
    .B(_1363_),
    .Y(_1513_));
 sky130_fd_sc_hd__o22ai_1 _2079_ (.A1(_1491_),
    .A2(_1347_),
    .B1(_1353_),
    .B2(_1513_),
    .Y(_1514_));
 sky130_fd_sc_hd__nand2_1 _2080_ (.A(net35),
    .B(_1405_),
    .Y(_1515_));
 sky130_fd_sc_hd__o221ai_2 _2081_ (.A1(_1664_),
    .A2(_1405_),
    .B1(_1336_),
    .B2(_1316_),
    .C1(_1515_),
    .Y(_1516_));
 sky130_fd_sc_hd__inv_1 _2082_ (.A(net32),
    .Y(_1517_));
 sky130_fd_sc_hd__nand2_1 _2083_ (.A(net3),
    .B(_1405_),
    .Y(_1518_));
 sky130_fd_sc_hd__o2111ai_2 _2084_ (.A1(_1517_),
    .A2(_1405_),
    .B1(_1412_),
    .C1(_1403_),
    .D1(_1518_),
    .Y(_1519_));
 sky130_fd_sc_hd__mux2i_1 _2085_ (.A0(net64),
    .A1(net35),
    .S(_1407_),
    .Y(_1520_));
 sky130_fd_sc_hd__nor2_1 _2086_ (.A(_1379_),
    .B(_1520_),
    .Y(_1521_));
 sky130_fd_sc_hd__a31oi_4 _2087_ (.A1(_1412_),
    .A2(_1516_),
    .A3(_1519_),
    .B1(_1521_),
    .Y(_1522_));
 sky130_fd_sc_hd__mux2i_1 _2088_ (.A0(net5),
    .A1(net7),
    .S(_1344_),
    .Y(_1523_));
 sky130_fd_sc_hd__nand3_1 _2089_ (.A(_1295_),
    .B(_1315_),
    .C(_1523_),
    .Y(_1524_));
 sky130_fd_sc_hd__nand2_1 _2090_ (.A(net39),
    .B(_1413_),
    .Y(_1525_));
 sky130_fd_sc_hd__o221ai_4 _2091_ (.A1(_1652_),
    .A2(_1413_),
    .B1(_1341_),
    .B2(_1342_),
    .C1(_1525_),
    .Y(_1526_));
 sky130_fd_sc_hd__nand2_1 _2092_ (.A(net39),
    .B(_1319_),
    .Y(_1527_));
 sky130_fd_sc_hd__o21ai_1 _2093_ (.A1(_1652_),
    .A2(_1407_),
    .B1(_1527_),
    .Y(_1528_));
 sky130_fd_sc_hd__a32oi_4 _2094_ (.A1(_1293_),
    .A2(_1524_),
    .A3(_1526_),
    .B1(_1528_),
    .B2(_1330_),
    .Y(_1529_));
 sky130_fd_sc_hd__and2_0 _2095_ (.A(_1437_),
    .B(_1529_),
    .X(_1530_));
 sky130_fd_sc_hd__a211oi_1 _2096_ (.A1(_1363_),
    .A2(_1522_),
    .B1(_1530_),
    .C1(_1489_),
    .Y(_1531_));
 sky130_fd_sc_hd__and2_0 _2097_ (.A(_1178_),
    .B(_1179_),
    .X(_1532_));
 sky130_fd_sc_hd__mux2i_2 _2098_ (.A0(_1532_),
    .A1(_1192_),
    .S(_1391_),
    .Y(_1533_));
 sky130_fd_sc_hd__or4b_1 _2099_ (.A(_1299_),
    .B(_1383_),
    .C(_1386_),
    .D_N(_1533_),
    .X(_1534_));
 sky130_fd_sc_hd__buf_2 _2100_ (.A(_1534_),
    .X(_1535_));
 sky130_fd_sc_hd__nand2_1 _2101_ (.A(_1399_),
    .B(_1535_),
    .Y(_1536_));
 sky130_fd_sc_hd__o311a_1 _2102_ (.A1(_1399_),
    .A2(_1514_),
    .A3(_1531_),
    .B1(_1536_),
    .C1(_1382_),
    .X(_1537_));
 sky130_fd_sc_hd__a311o_1 _2103_ (.A1(_1399_),
    .A2(_1397_),
    .A3(_1497_),
    .B1(_1512_),
    .C1(_1537_),
    .X(_1538_));
 sky130_fd_sc_hd__and2_0 _2104_ (.A(_1380_),
    .B(_1538_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _2105_ (.A0(net33),
    .A1(net4),
    .S(_1405_),
    .X(_1539_));
 sky130_fd_sc_hd__nand2_1 _2106_ (.A(net36),
    .B(_1407_),
    .Y(_1540_));
 sky130_fd_sc_hd__o21ai_1 _2107_ (.A1(_1661_),
    .A2(_1407_),
    .B1(_1540_),
    .Y(_1541_));
 sky130_fd_sc_hd__mux2i_1 _2108_ (.A0(net65),
    .A1(net36),
    .S(_1405_),
    .Y(_1542_));
 sky130_fd_sc_hd__nor4_1 _2109_ (.A(a_exp_larger),
    .B(_1292_),
    .C(_1450_),
    .D(_1542_),
    .Y(_1543_));
 sky130_fd_sc_hd__a221oi_4 _2110_ (.A1(_1337_),
    .A2(_1539_),
    .B1(_1541_),
    .B2(_1330_),
    .C1(_1543_),
    .Y(_1544_));
 sky130_fd_sc_hd__mux4_1 _2111_ (.A0(net6),
    .A1(net8),
    .A2(net38),
    .A3(net40),
    .S0(_1413_),
    .S1(_1316_),
    .X(_1545_));
 sky130_fd_sc_hd__mux2i_1 _2112_ (.A0(net38),
    .A1(net40),
    .S(_1407_),
    .Y(_1546_));
 sky130_fd_sc_hd__nor2_1 _2113_ (.A(_1379_),
    .B(_1546_),
    .Y(_1547_));
 sky130_fd_sc_hd__a211oi_1 _2114_ (.A1(_1412_),
    .A2(_1545_),
    .B1(_1547_),
    .C1(_1401_),
    .Y(_1548_));
 sky130_fd_sc_hd__a21oi_2 _2115_ (.A1(_1401_),
    .A2(_1544_),
    .B1(_1548_),
    .Y(_1549_));
 sky130_fd_sc_hd__a211oi_2 _2116_ (.A1(_1401_),
    .A2(_1522_),
    .B1(_1530_),
    .C1(_1400_),
    .Y(_1550_));
 sky130_fd_sc_hd__a21oi_4 _2117_ (.A1(_1400_),
    .A2(_1549_),
    .B1(_1550_),
    .Y(_1551_));
 sky130_fd_sc_hd__nand3_4 _2118_ (.A(_1380_),
    .B(_1470_),
    .C(_1382_),
    .Y(_1552_));
 sky130_fd_sc_hd__or2_0 _2119_ (.A(_1189_),
    .B(_1250_),
    .X(_1553_));
 sky130_fd_sc_hd__buf_2 _2120_ (.A(_1553_),
    .X(_1554_));
 sky130_fd_sc_hd__nor2_4 _2121_ (.A(_1399_),
    .B(_1398_),
    .Y(_1555_));
 sky130_fd_sc_hd__nand2_2 _2122_ (.A(_1475_),
    .B(_1401_),
    .Y(_1556_));
 sky130_fd_sc_hd__mux4_1 _2123_ (.A0(net27),
    .A1(net24),
    .A2(net59),
    .A3(net56),
    .S0(_1298_),
    .S1(_1404_),
    .X(_1557_));
 sky130_fd_sc_hd__mux2i_1 _2124_ (.A0(_1471_),
    .A1(_1557_),
    .S(_1459_),
    .Y(_1558_));
 sky130_fd_sc_hd__mux4_1 _2125_ (.A0(net29),
    .A1(net31),
    .A2(net61),
    .A3(net63),
    .S0(_1413_),
    .S1(_1316_),
    .X(_1559_));
 sky130_fd_sc_hd__nand2_1 _2126_ (.A(net63),
    .B(_1407_),
    .Y(_1560_));
 sky130_fd_sc_hd__o21ai_1 _2127_ (.A1(_1637_),
    .A2(_1407_),
    .B1(_1560_),
    .Y(_1561_));
 sky130_fd_sc_hd__a22oi_4 _2128_ (.A1(_1412_),
    .A2(_1559_),
    .B1(_1561_),
    .B2(_1330_),
    .Y(_1562_));
 sky130_fd_sc_hd__mux2_1 _2129_ (.A0(_1504_),
    .A1(_1562_),
    .S(_1364_),
    .X(_1563_));
 sky130_fd_sc_hd__o22ai_1 _2130_ (.A1(_1556_),
    .A2(_1558_),
    .B1(_1563_),
    .B2(_1402_),
    .Y(_1564_));
 sky130_fd_sc_hd__a22oi_1 _2131_ (.A1(net34),
    .A2(_1554_),
    .B1(_1555_),
    .B2(_1564_),
    .Y(_0122_));
 sky130_fd_sc_hd__nand2_1 _2132_ (.A(net44),
    .B(_1391_),
    .Y(_0123_));
 sky130_fd_sc_hd__nand2_1 _2133_ (.A(net12),
    .B(_1450_),
    .Y(_0124_));
 sky130_fd_sc_hd__a21oi_1 _2134_ (.A1(_0123_),
    .A2(_0124_),
    .B1(_1455_),
    .Y(_0125_));
 sky130_fd_sc_hd__nand2_1 _2135_ (.A(net42),
    .B(_1448_),
    .Y(_0126_));
 sky130_fd_sc_hd__nand2_1 _2136_ (.A(net10),
    .B(_1450_),
    .Y(_0127_));
 sky130_fd_sc_hd__a21oi_1 _2137_ (.A1(_0126_),
    .A2(_0127_),
    .B1(_1459_),
    .Y(_0128_));
 sky130_fd_sc_hd__o211ai_2 _2138_ (.A1(_0125_),
    .A2(_0128_),
    .B1(_1364_),
    .C1(_1475_),
    .Y(_0129_));
 sky130_fd_sc_hd__or2_0 _2139_ (.A(_1364_),
    .B(_1488_),
    .X(_0130_));
 sky130_fd_sc_hd__nor2_2 _2140_ (.A(_1383_),
    .B(_1392_),
    .Y(_0131_));
 sky130_fd_sc_hd__mux4_2 _2141_ (.A0(net15),
    .A1(net14),
    .A2(net47),
    .A3(net46),
    .S0(_1298_),
    .S1(_1391_),
    .X(_0132_));
 sky130_fd_sc_hd__a221oi_4 _2142_ (.A1(_1459_),
    .A2(_0131_),
    .B1(_0132_),
    .B2(_1462_),
    .C1(_1363_),
    .Y(_0133_));
 sky130_fd_sc_hd__a31oi_4 _2143_ (.A1(_1401_),
    .A2(_0129_),
    .A3(_0130_),
    .B1(_0133_),
    .Y(_0134_));
 sky130_fd_sc_hd__nor2_2 _2144_ (.A(_1470_),
    .B(_1398_),
    .Y(_0135_));
 sky130_fd_sc_hd__nand2_1 _2145_ (.A(_0134_),
    .B(_0135_),
    .Y(_0136_));
 sky130_fd_sc_hd__o211ai_1 _2146_ (.A1(_1551_),
    .A2(_1552_),
    .B1(_0122_),
    .C1(_0136_),
    .Y(_0069_));
 sky130_fd_sc_hd__nor2_1 _2147_ (.A(_0125_),
    .B(_0128_),
    .Y(_0137_));
 sky130_fd_sc_hd__or2_0 _2148_ (.A(_1455_),
    .B(_1533_),
    .X(_0138_));
 sky130_fd_sc_hd__nand2_1 _2149_ (.A(net15),
    .B(_1450_),
    .Y(_0139_));
 sky130_fd_sc_hd__o211ai_2 _2150_ (.A1(_1682_),
    .A2(_1337_),
    .B1(_1455_),
    .C1(_0139_),
    .Y(_0140_));
 sky130_fd_sc_hd__mux2i_1 _2151_ (.A0(net16),
    .A1(net48),
    .S(_1448_),
    .Y(_0141_));
 sky130_fd_sc_hd__nor3_1 _2152_ (.A(_1489_),
    .B(_1459_),
    .C(_0141_),
    .Y(_0142_));
 sky130_fd_sc_hd__a31oi_4 _2153_ (.A1(_1489_),
    .A2(_0138_),
    .A3(_0140_),
    .B1(_0142_),
    .Y(_0143_));
 sky130_fd_sc_hd__o22ai_2 _2154_ (.A1(_1513_),
    .A2(_0137_),
    .B1(_0143_),
    .B2(_1402_),
    .Y(_0144_));
 sky130_fd_sc_hd__clkbuf_4 _2155_ (.A(_1489_),
    .X(_0145_));
 sky130_fd_sc_hd__and2_0 _2156_ (.A(_1433_),
    .B(_1436_),
    .X(_0146_));
 sky130_fd_sc_hd__nor3_1 _2157_ (.A(_0145_),
    .B(_0146_),
    .C(_1438_),
    .Y(_0147_));
 sky130_fd_sc_hd__a21oi_4 _2158_ (.A1(_1475_),
    .A2(_0144_),
    .B1(_0147_),
    .Y(_0148_));
 sky130_fd_sc_hd__a31oi_2 _2159_ (.A1(_1412_),
    .A2(_1440_),
    .A3(_1442_),
    .B1(_1444_),
    .Y(_0149_));
 sky130_fd_sc_hd__nor3_1 _2160_ (.A(_0145_),
    .B(_1401_),
    .C(_0149_),
    .Y(_0150_));
 sky130_fd_sc_hd__nor3_1 _2161_ (.A(_0145_),
    .B(_1438_),
    .C(_1331_),
    .Y(_0151_));
 sky130_fd_sc_hd__a211oi_4 _2162_ (.A1(_0145_),
    .A2(_1549_),
    .B1(_0150_),
    .C1(_0151_),
    .Y(_0152_));
 sky130_fd_sc_hd__mux4_1 _2163_ (.A0(net27),
    .A1(net28),
    .A2(net59),
    .A3(net60),
    .S0(_1364_),
    .S1(_1404_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2i_1 _2164_ (.A0(_1506_),
    .A1(_0153_),
    .S(_1459_),
    .Y(_0154_));
 sky130_fd_sc_hd__mux2i_1 _2165_ (.A0(_1335_),
    .A1(_1562_),
    .S(_0145_),
    .Y(_0155_));
 sky130_fd_sc_hd__a2bb2oi_1 _2166_ (.A1_N(_1556_),
    .A2_N(_0154_),
    .B1(_0155_),
    .B2(_1438_),
    .Y(_0156_));
 sky130_fd_sc_hd__nand3_1 _2167_ (.A(_1380_),
    .B(_1274_),
    .C(_1397_),
    .Y(_0157_));
 sky130_fd_sc_hd__clkbuf_4 _2168_ (.A(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__nand2_1 _2169_ (.A(net45),
    .B(_1554_),
    .Y(_0159_));
 sky130_fd_sc_hd__o221a_1 _2170_ (.A1(_1552_),
    .A2(_0152_),
    .B1(_0156_),
    .B2(_0158_),
    .C1(_0159_),
    .X(_0160_));
 sky130_fd_sc_hd__o31ai_1 _2171_ (.A1(_1470_),
    .A2(_1398_),
    .A3(_0148_),
    .B1(_0160_),
    .Y(_0070_));
 sky130_fd_sc_hd__nor2_1 _2172_ (.A(_1438_),
    .B(_1466_),
    .Y(_0161_));
 sky130_fd_sc_hd__o21ai_0 _2173_ (.A1(_1402_),
    .A2(_1353_),
    .B1(_1400_),
    .Y(_0162_));
 sky130_fd_sc_hd__o22ai_1 _2174_ (.A1(_1461_),
    .A2(_1556_),
    .B1(_1335_),
    .B2(_1402_),
    .Y(_0163_));
 sky130_fd_sc_hd__o22ai_2 _2175_ (.A1(_0161_),
    .A2(_0162_),
    .B1(_0163_),
    .B2(_1400_),
    .Y(_0164_));
 sky130_fd_sc_hd__clkbuf_4 _2176_ (.A(_1554_),
    .X(_0165_));
 sky130_fd_sc_hd__mux4_2 _2177_ (.A0(_1420_),
    .A1(_0149_),
    .A2(_1347_),
    .A3(_1331_),
    .S0(_1298_),
    .S1(_1363_),
    .X(_0166_));
 sky130_fd_sc_hd__nor2_1 _2178_ (.A(_1552_),
    .B(_0166_),
    .Y(_0167_));
 sky130_fd_sc_hd__a21oi_1 _2179_ (.A1(net56),
    .A2(_0165_),
    .B1(_0167_),
    .Y(_0168_));
 sky130_fd_sc_hd__and3_1 _2180_ (.A(_1489_),
    .B(_1433_),
    .C(_1436_),
    .X(_0169_));
 sky130_fd_sc_hd__nor2_1 _2181_ (.A(_1489_),
    .B(_1411_),
    .Y(_0170_));
 sky130_fd_sc_hd__nand3_1 _2182_ (.A(_1455_),
    .B(_1438_),
    .C(_0131_),
    .Y(_0171_));
 sky130_fd_sc_hd__o31a_2 _2183_ (.A1(_1437_),
    .A2(_0169_),
    .A3(_0170_),
    .B1(_0171_),
    .X(_0172_));
 sky130_fd_sc_hd__nand2b_1 _2184_ (.A_N(_0172_),
    .B(_0135_),
    .Y(_0173_));
 sky130_fd_sc_hd__o211ai_2 _2185_ (.A1(_0158_),
    .A2(_0164_),
    .B1(_0168_),
    .C1(_0173_),
    .Y(_0071_));
 sky130_fd_sc_hd__nand4_1 _2186_ (.A(_0145_),
    .B(_1475_),
    .C(_1455_),
    .D(_1533_),
    .Y(_0174_));
 sky130_fd_sc_hd__o22ai_1 _2187_ (.A1(_1448_),
    .A2(_1493_),
    .B1(_1494_),
    .B2(_1495_),
    .Y(_0175_));
 sky130_fd_sc_hd__a21o_1 _2188_ (.A1(_1489_),
    .A2(_1411_),
    .B1(_1437_),
    .X(_0176_));
 sky130_fd_sc_hd__a21oi_1 _2189_ (.A1(_1400_),
    .A2(_0175_),
    .B1(_0176_),
    .Y(_0177_));
 sky130_fd_sc_hd__a21oi_4 _2190_ (.A1(_1438_),
    .A2(_0174_),
    .B1(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__mux2i_1 _2191_ (.A0(_1504_),
    .A1(_1522_),
    .S(_1437_),
    .Y(_0179_));
 sky130_fd_sc_hd__o21ai_0 _2192_ (.A1(_1402_),
    .A2(_1353_),
    .B1(_0145_),
    .Y(_0180_));
 sky130_fd_sc_hd__o22ai_1 _2193_ (.A1(_0145_),
    .A2(_0179_),
    .B1(_0180_),
    .B2(_0161_),
    .Y(_0181_));
 sky130_fd_sc_hd__nor2_1 _2194_ (.A(_0158_),
    .B(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__and3_1 _2195_ (.A(_1380_),
    .B(_1274_),
    .C(_1382_),
    .X(_0183_));
 sky130_fd_sc_hd__clkbuf_2 _2196_ (.A(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2i_1 _2197_ (.A0(_1420_),
    .A1(_1347_),
    .S(_1401_),
    .Y(_0185_));
 sky130_fd_sc_hd__mux2i_2 _2198_ (.A0(_1488_),
    .A1(_1529_),
    .S(_1401_),
    .Y(_0186_));
 sky130_fd_sc_hd__mux2_1 _2199_ (.A0(_0185_),
    .A1(_0186_),
    .S(_1364_),
    .X(_0187_));
 sky130_fd_sc_hd__a22o_1 _2200_ (.A1(net59),
    .A2(_1554_),
    .B1(_0184_),
    .B2(_0187_),
    .X(_0188_));
 sky130_fd_sc_hd__a211o_1 _2201_ (.A1(_0135_),
    .A2(_0178_),
    .B1(_0182_),
    .C1(_0188_),
    .X(_0072_));
 sky130_fd_sc_hd__o21ai_0 _2202_ (.A1(_0125_),
    .A2(_0128_),
    .B1(_1475_),
    .Y(_0189_));
 sky130_fd_sc_hd__a211oi_1 _2203_ (.A1(_1412_),
    .A2(_1545_),
    .B1(_1547_),
    .C1(_1437_),
    .Y(_0190_));
 sky130_fd_sc_hd__a21oi_1 _2204_ (.A1(_1438_),
    .A2(_0189_),
    .B1(_0190_),
    .Y(_0191_));
 sky130_fd_sc_hd__mux2i_4 _2205_ (.A0(_0186_),
    .A1(_0191_),
    .S(_1400_),
    .Y(_0192_));
 sky130_fd_sc_hd__mux2i_2 _2206_ (.A0(_1544_),
    .A1(_1562_),
    .S(_1401_),
    .Y(_0193_));
 sky130_fd_sc_hd__mux2_1 _2207_ (.A0(_0179_),
    .A1(_0193_),
    .S(_1400_),
    .X(_0194_));
 sky130_fd_sc_hd__a32o_4 _2208_ (.A1(_1462_),
    .A2(_1402_),
    .A3(_0132_),
    .B1(_1508_),
    .B2(_0131_),
    .X(_0195_));
 sky130_fd_sc_hd__a222oi_1 _2209_ (.A1(net60),
    .A2(_1554_),
    .B1(_1555_),
    .B2(_0194_),
    .C1(_0195_),
    .C2(_0135_),
    .Y(_0196_));
 sky130_fd_sc_hd__o21ai_0 _2210_ (.A1(_1552_),
    .A2(_0192_),
    .B1(_0196_),
    .Y(_0073_));
 sky130_fd_sc_hd__a21oi_1 _2211_ (.A1(_0146_),
    .A2(_1438_),
    .B1(_1445_),
    .Y(_0197_));
 sky130_fd_sc_hd__mux2_2 _2212_ (.A0(_0197_),
    .A1(_0191_),
    .S(_0145_),
    .X(_0198_));
 sky130_fd_sc_hd__nor2_2 _2213_ (.A(_1556_),
    .B(_0143_),
    .Y(_0199_));
 sky130_fd_sc_hd__a22o_1 _2214_ (.A1(net61),
    .A2(_1554_),
    .B1(_0135_),
    .B2(_0199_),
    .X(_0200_));
 sky130_fd_sc_hd__mux2i_1 _2215_ (.A0(_1331_),
    .A1(_1335_),
    .S(_1402_),
    .Y(_0201_));
 sky130_fd_sc_hd__mux2i_2 _2216_ (.A0(_0201_),
    .A1(_0193_),
    .S(_0145_),
    .Y(_0202_));
 sky130_fd_sc_hd__nor2_1 _2217_ (.A(_0158_),
    .B(_0202_),
    .Y(_0203_));
 sky130_fd_sc_hd__a211o_1 _2218_ (.A1(_0184_),
    .A2(_0198_),
    .B1(_0200_),
    .C1(_0203_),
    .X(_0074_));
 sky130_fd_sc_hd__nand2b_1 _2219_ (.A_N(_1366_),
    .B(_1395_),
    .Y(_0204_));
 sky130_fd_sc_hd__nand2_1 _2220_ (.A(net62),
    .B(_0165_),
    .Y(_0205_));
 sky130_fd_sc_hd__o221ai_2 _2221_ (.A1(_0204_),
    .A2(_1398_),
    .B1(_1552_),
    .B2(_1447_),
    .C1(_0205_),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_1 _2222_ (.A(_1497_),
    .Y(_0206_));
 sky130_fd_sc_hd__nor2_1 _2223_ (.A(_1514_),
    .B(_1531_),
    .Y(_0207_));
 sky130_fd_sc_hd__or3_1 _2224_ (.A(_1274_),
    .B(_1398_),
    .C(_1535_),
    .X(_0208_));
 sky130_fd_sc_hd__o221a_1 _2225_ (.A1(_1631_),
    .A2(_1251_),
    .B1(_0207_),
    .B2(_0157_),
    .C1(_0208_),
    .X(_0209_));
 sky130_fd_sc_hd__o21ai_0 _2226_ (.A1(_0206_),
    .A2(_1552_),
    .B1(_0209_),
    .Y(_0076_));
 sky130_fd_sc_hd__nand2_1 _2227_ (.A(_0134_),
    .B(_0184_),
    .Y(_0210_));
 sky130_fd_sc_hd__o221ai_2 _2228_ (.A1(_1664_),
    .A2(_1260_),
    .B1(_1551_),
    .B2(_0158_),
    .C1(_0210_),
    .Y(_0052_));
 sky130_fd_sc_hd__nand2_1 _2229_ (.A(net65),
    .B(_0165_),
    .Y(_0211_));
 sky130_fd_sc_hd__o221ai_1 _2230_ (.A1(_0158_),
    .A2(_0152_),
    .B1(_0148_),
    .B2(_1552_),
    .C1(_0211_),
    .Y(_0053_));
 sky130_fd_sc_hd__nand2_1 _2231_ (.A(_1192_),
    .B(_1201_),
    .Y(_0212_));
 sky130_fd_sc_hd__nor2_1 _2232_ (.A(_1189_),
    .B(_1249_),
    .Y(_0213_));
 sky130_fd_sc_hd__o22ai_1 _2233_ (.A1(_1378_),
    .A2(_1379_),
    .B1(_1336_),
    .B2(_1342_),
    .Y(_0214_));
 sky130_fd_sc_hd__nand2_1 _2234_ (.A(_1274_),
    .B(_0214_),
    .Y(_0215_));
 sky130_fd_sc_hd__and2_0 _2235_ (.A(_1397_),
    .B(_0166_),
    .X(_0216_));
 sky130_fd_sc_hd__a211oi_1 _2236_ (.A1(_1382_),
    .A2(_0172_),
    .B1(_0215_),
    .C1(_0216_),
    .Y(_0217_));
 sky130_fd_sc_hd__a32o_1 _2237_ (.A1(_0212_),
    .A2(_0213_),
    .A3(_0217_),
    .B1(_0165_),
    .B2(net35),
    .X(_0054_));
 sky130_fd_sc_hd__clkbuf_4 _2238_ (.A(_1251_),
    .X(_0218_));
 sky130_fd_sc_hd__nor2_1 _2239_ (.A(_1655_),
    .B(_0218_),
    .Y(_0219_));
 sky130_fd_sc_hd__a221o_1 _2240_ (.A1(_0184_),
    .A2(_0178_),
    .B1(_0187_),
    .B2(_1555_),
    .C1(_0219_),
    .X(_0055_));
 sky130_fd_sc_hd__a22oi_1 _2241_ (.A1(net37),
    .A2(_0165_),
    .B1(_0184_),
    .B2(_0195_),
    .Y(_0220_));
 sky130_fd_sc_hd__o21ai_0 _2242_ (.A1(_0158_),
    .A2(_0192_),
    .B1(_0220_),
    .Y(_0056_));
 sky130_fd_sc_hd__nor3_1 _2243_ (.A(_1556_),
    .B(_1552_),
    .C(_0143_),
    .Y(_0221_));
 sky130_fd_sc_hd__a221o_1 _2244_ (.A1(net38),
    .A2(_1554_),
    .B1(_1555_),
    .B2(_0198_),
    .C1(_0221_),
    .X(_0057_));
 sky130_fd_sc_hd__a22oi_1 _2245_ (.A1(net39),
    .A2(_0165_),
    .B1(_1393_),
    .B2(_0184_),
    .Y(_0222_));
 sky130_fd_sc_hd__o21ai_0 _2246_ (.A1(_1447_),
    .A2(_0158_),
    .B1(_0222_),
    .Y(_0058_));
 sky130_fd_sc_hd__nand2_1 _2247_ (.A(_1497_),
    .B(_1555_),
    .Y(_0223_));
 sky130_fd_sc_hd__o221ai_1 _2248_ (.A1(_1643_),
    .A2(_1260_),
    .B1(_1535_),
    .B2(_1552_),
    .C1(_0223_),
    .Y(_0059_));
 sky130_fd_sc_hd__nand2_1 _2249_ (.A(_0134_),
    .B(_1555_),
    .Y(_0224_));
 sky130_fd_sc_hd__o21ai_0 _2250_ (.A1(_1676_),
    .A2(_1253_),
    .B1(_0224_),
    .Y(_0060_));
 sky130_fd_sc_hd__o22ai_1 _2251_ (.A1(_1673_),
    .A2(_1252_),
    .B1(_0158_),
    .B2(_0148_),
    .Y(_0061_));
 sky130_fd_sc_hd__o22ai_1 _2252_ (.A1(_1670_),
    .A2(_1252_),
    .B1(_0158_),
    .B2(_0172_),
    .Y(_0063_));
 sky130_fd_sc_hd__a22o_1 _2253_ (.A1(net44),
    .A2(_0165_),
    .B1(_1555_),
    .B2(_0178_),
    .X(_0064_));
 sky130_fd_sc_hd__nand2_1 _2254_ (.A(_1555_),
    .B(_0195_),
    .Y(_0225_));
 sky130_fd_sc_hd__o21ai_0 _2255_ (.A1(_1685_),
    .A2(_1253_),
    .B1(_0225_),
    .Y(_0065_));
 sky130_fd_sc_hd__nand2_1 _2256_ (.A(_1555_),
    .B(_0199_),
    .Y(_0226_));
 sky130_fd_sc_hd__o21ai_0 _2257_ (.A1(_1682_),
    .A2(_1253_),
    .B1(_0226_),
    .Y(_0066_));
 sky130_fd_sc_hd__nand2_1 _2258_ (.A(_1393_),
    .B(_1555_),
    .Y(_0227_));
 sky130_fd_sc_hd__o21ai_0 _2259_ (.A1(_1679_),
    .A2(_1253_),
    .B1(_0227_),
    .Y(_0067_));
 sky130_fd_sc_hd__o21ai_0 _2260_ (.A1(_1197_),
    .A2(_1200_),
    .B1(_0213_),
    .Y(_0228_));
 sky130_fd_sc_hd__o31a_1 _2261_ (.A1(_1382_),
    .A2(_1535_),
    .A3(_0215_),
    .B1(_0213_),
    .X(_0229_));
 sky130_fd_sc_hd__a21oi_1 _2262_ (.A1(_1192_),
    .A2(_0228_),
    .B1(_0229_),
    .Y(_0068_));
 sky130_fd_sc_hd__nand3_1 _2263_ (.A(_1450_),
    .B(_1382_),
    .C(_1395_),
    .Y(_0230_));
 sky130_fd_sc_hd__nand2_1 _2264_ (.A(_1450_),
    .B(_1397_),
    .Y(_0231_));
 sky130_fd_sc_hd__o22ai_1 _2265_ (.A1(_1366_),
    .A2(_0230_),
    .B1(_0231_),
    .B2(_1474_),
    .Y(_0025_));
 sky130_fd_sc_hd__and2_0 _2266_ (.A(_1337_),
    .B(_1538_),
    .X(_0036_));
 sky130_fd_sc_hd__nor2_1 _2267_ (.A(_1470_),
    .B(_0231_),
    .Y(_0232_));
 sky130_fd_sc_hd__nor2_4 _2268_ (.A(_1399_),
    .B(_0231_),
    .Y(_0233_));
 sky130_fd_sc_hd__nand3_2 _2269_ (.A(_1470_),
    .B(_1450_),
    .C(_1382_),
    .Y(_0234_));
 sky130_fd_sc_hd__o2bb2ai_1 _2270_ (.A1_N(_0233_),
    .A2_N(_1564_),
    .B1(_1551_),
    .B2(_0234_),
    .Y(_0235_));
 sky130_fd_sc_hd__a221o_1 _2271_ (.A1(net2),
    .A2(_0218_),
    .B1(_0134_),
    .B2(_0232_),
    .C1(_0235_),
    .X(_0043_));
 sky130_fd_sc_hd__nor2_1 _2272_ (.A(_1448_),
    .B(_1382_),
    .Y(_0236_));
 sky130_fd_sc_hd__nand2_1 _2273_ (.A(_1399_),
    .B(_0236_),
    .Y(_0237_));
 sky130_fd_sc_hd__nand2_1 _2274_ (.A(net13),
    .B(_1260_),
    .Y(_0238_));
 sky130_fd_sc_hd__nand2_1 _2275_ (.A(_1337_),
    .B(_1397_),
    .Y(_0239_));
 sky130_fd_sc_hd__nand3_1 _2276_ (.A(_1470_),
    .B(_1337_),
    .C(_1382_),
    .Y(_0240_));
 sky130_fd_sc_hd__o32a_1 _2277_ (.A1(_1399_),
    .A2(_0156_),
    .A3(_0239_),
    .B1(_0240_),
    .B2(_0152_),
    .X(_0241_));
 sky130_fd_sc_hd__o211ai_1 _2278_ (.A1(_0148_),
    .A2(_0237_),
    .B1(_0238_),
    .C1(_0241_),
    .Y(_0044_));
 sky130_fd_sc_hd__nand2_1 _2279_ (.A(_1470_),
    .B(_0236_),
    .Y(_0242_));
 sky130_fd_sc_hd__clkbuf_4 _2280_ (.A(_0242_),
    .X(_0243_));
 sky130_fd_sc_hd__nand2_1 _2281_ (.A(net24),
    .B(_1260_),
    .Y(_0244_));
 sky130_fd_sc_hd__o32a_1 _2282_ (.A1(_1470_),
    .A2(_0172_),
    .A3(_0239_),
    .B1(_0240_),
    .B2(_0166_),
    .X(_0245_));
 sky130_fd_sc_hd__o211ai_2 _2283_ (.A1(_0164_),
    .A2(_0243_),
    .B1(_0244_),
    .C1(_0245_),
    .Y(_0045_));
 sky130_fd_sc_hd__nor3_4 _2284_ (.A(_1399_),
    .B(_1448_),
    .C(_1397_),
    .Y(_0246_));
 sky130_fd_sc_hd__o2bb2ai_1 _2285_ (.A1_N(_0187_),
    .A2_N(_0246_),
    .B1(_0242_),
    .B2(_0181_),
    .Y(_0247_));
 sky130_fd_sc_hd__a221o_1 _2286_ (.A1(net27),
    .A2(_1251_),
    .B1(_0178_),
    .B2(_0232_),
    .C1(_0247_),
    .X(_0046_));
 sky130_fd_sc_hd__nand2_1 _2287_ (.A(net28),
    .B(_1260_),
    .Y(_0248_));
 sky130_fd_sc_hd__o21a_1 _2288_ (.A1(_1470_),
    .A2(_0195_),
    .B1(_0236_),
    .X(_0249_));
 sky130_fd_sc_hd__o21ai_0 _2289_ (.A1(_1399_),
    .A2(_0194_),
    .B1(_0249_),
    .Y(_0250_));
 sky130_fd_sc_hd__o211ai_1 _2290_ (.A1(_0192_),
    .A2(_0234_),
    .B1(_0248_),
    .C1(_0250_),
    .Y(_0047_));
 sky130_fd_sc_hd__o2bb2ai_1 _2291_ (.A1_N(_0199_),
    .A2_N(_0232_),
    .B1(_0242_),
    .B2(_0202_),
    .Y(_0251_));
 sky130_fd_sc_hd__a221o_1 _2292_ (.A1(net29),
    .A2(_1251_),
    .B1(_0198_),
    .B2(_0246_),
    .C1(_0251_),
    .X(_0048_));
 sky130_fd_sc_hd__nand2_1 _2293_ (.A(net30),
    .B(_1260_),
    .Y(_0252_));
 sky130_fd_sc_hd__o221ai_2 _2294_ (.A1(_0204_),
    .A2(_0239_),
    .B1(_0240_),
    .B2(_1447_),
    .C1(_0252_),
    .Y(_0049_));
 sky130_fd_sc_hd__nand2_1 _2295_ (.A(net31),
    .B(_1251_),
    .Y(_0253_));
 sky130_fd_sc_hd__o221ai_1 _2296_ (.A1(_0207_),
    .A2(_0243_),
    .B1(_0237_),
    .B2(_1535_),
    .C1(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hd__a21o_1 _2297_ (.A1(_1497_),
    .A2(_0246_),
    .B1(_0254_),
    .X(_0050_));
 sky130_fd_sc_hd__nor2_1 _2298_ (.A(a_exp_larger),
    .B(_1341_),
    .Y(_0255_));
 sky130_fd_sc_hd__nand4bb_1 _2299_ (.A_N(_1397_),
    .B_N(_0215_),
    .C(_0255_),
    .D(_0134_),
    .Y(_0256_));
 sky130_fd_sc_hd__o221ai_2 _2300_ (.A1(_1517_),
    .A2(_0165_),
    .B1(_1551_),
    .B2(_0243_),
    .C1(_0256_),
    .Y(_0026_));
 sky130_fd_sc_hd__a2bb2oi_1 _2301_ (.A1_N(_0152_),
    .A2_N(_0243_),
    .B1(net33),
    .B2(_0218_),
    .Y(_0257_));
 sky130_fd_sc_hd__o21ai_1 _2302_ (.A1(_0148_),
    .A2(_0234_),
    .B1(_0257_),
    .Y(_0027_));
 sky130_fd_sc_hd__a22o_1 _2303_ (.A1(net3),
    .A2(_0218_),
    .B1(_0217_),
    .B2(_0255_),
    .X(_0028_));
 sky130_fd_sc_hd__and2_0 _2304_ (.A(net4),
    .B(_1251_),
    .X(_0258_));
 sky130_fd_sc_hd__and2_0 _2305_ (.A(_0187_),
    .B(_0233_),
    .X(_0259_));
 sky130_fd_sc_hd__a211o_1 _2306_ (.A1(_0178_),
    .A2(_0246_),
    .B1(_0258_),
    .C1(_0259_),
    .X(_0029_));
 sky130_fd_sc_hd__a22oi_1 _2307_ (.A1(net5),
    .A2(_0218_),
    .B1(_0195_),
    .B2(_0246_),
    .Y(_0260_));
 sky130_fd_sc_hd__o21ai_0 _2308_ (.A1(_0192_),
    .A2(_0243_),
    .B1(_0260_),
    .Y(_0030_));
 sky130_fd_sc_hd__and2_0 _2309_ (.A(net6),
    .B(_1251_),
    .X(_0261_));
 sky130_fd_sc_hd__a221o_1 _2310_ (.A1(_0199_),
    .A2(_0246_),
    .B1(_0233_),
    .B2(_0198_),
    .C1(_0261_),
    .X(_0031_));
 sky130_fd_sc_hd__a22oi_1 _2311_ (.A1(net7),
    .A2(_0218_),
    .B1(_1393_),
    .B2(_0246_),
    .Y(_0262_));
 sky130_fd_sc_hd__o21ai_0 _2312_ (.A1(_1447_),
    .A2(_0243_),
    .B1(_0262_),
    .Y(_0032_));
 sky130_fd_sc_hd__nand2_1 _2313_ (.A(net8),
    .B(_1260_),
    .Y(_0263_));
 sky130_fd_sc_hd__o221ai_1 _2314_ (.A1(_1535_),
    .A2(_0234_),
    .B1(_0243_),
    .B2(_0206_),
    .C1(_0263_),
    .Y(_0033_));
 sky130_fd_sc_hd__a22o_1 _2315_ (.A1(net9),
    .A2(_0218_),
    .B1(_0134_),
    .B2(_0233_),
    .X(_0034_));
 sky130_fd_sc_hd__nand2_1 _2316_ (.A(net10),
    .B(_1260_),
    .Y(_0264_));
 sky130_fd_sc_hd__o21ai_0 _2317_ (.A1(_0148_),
    .A2(_0243_),
    .B1(_0264_),
    .Y(_0035_));
 sky130_fd_sc_hd__o22ai_1 _2318_ (.A1(_1431_),
    .A2(_0165_),
    .B1(_0172_),
    .B2(_0243_),
    .Y(_0037_));
 sky130_fd_sc_hd__a22o_1 _2319_ (.A1(net12),
    .A2(_0218_),
    .B1(_0178_),
    .B2(_0233_),
    .X(_0038_));
 sky130_fd_sc_hd__nand2_1 _2320_ (.A(_0195_),
    .B(_0233_),
    .Y(_0265_));
 sky130_fd_sc_hd__o21ai_0 _2321_ (.A1(_1426_),
    .A2(_0165_),
    .B1(_0265_),
    .Y(_0039_));
 sky130_fd_sc_hd__a22o_1 _2322_ (.A1(net15),
    .A2(_0218_),
    .B1(_0199_),
    .B2(_0233_),
    .X(_0040_));
 sky130_fd_sc_hd__a22o_1 _2323_ (.A1(net16),
    .A2(_0218_),
    .B1(_1393_),
    .B2(_0233_),
    .X(_0041_));
 sky130_fd_sc_hd__o22ai_1 _2324_ (.A1(_1532_),
    .A2(_1250_),
    .B1(_1535_),
    .B2(_0243_),
    .Y(_0042_));
 sky130_fd_sc_hd__buf_4 _2325_ (.A(\add_result[26] ),
    .X(_0266_));
 sky130_fd_sc_hd__buf_2 _2326_ (.A(\add_result[22] ),
    .X(_0267_));
 sky130_fd_sc_hd__buf_2 _2327_ (.A(\add_result[24] ),
    .X(_0268_));
 sky130_fd_sc_hd__buf_2 _2328_ (.A(\add_result[23] ),
    .X(_0269_));
 sky130_fd_sc_hd__nor3_1 _2329_ (.A(_0267_),
    .B(_0268_),
    .C(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__buf_4 _2330_ (.A(\add_result[4] ),
    .X(_0271_));
 sky130_fd_sc_hd__nor4_1 _2331_ (.A(_0271_),
    .B(\add_result[17] ),
    .C(\add_result[19] ),
    .D(\add_result[25] ),
    .Y(_0272_));
 sky130_fd_sc_hd__buf_4 _2332_ (.A(\add_result[3] ),
    .X(_0273_));
 sky130_fd_sc_hd__buf_4 _2333_ (.A(\add_result[9] ),
    .X(_0274_));
 sky130_fd_sc_hd__clkbuf_4 _2334_ (.A(\add_result[12] ),
    .X(_0275_));
 sky130_fd_sc_hd__nor4_1 _2335_ (.A(_0273_),
    .B(_0274_),
    .C(_0275_),
    .D(\add_result[11] ),
    .Y(_0276_));
 sky130_fd_sc_hd__clkbuf_4 _2336_ (.A(\add_result[13] ),
    .X(_0277_));
 sky130_fd_sc_hd__clkbuf_4 _2337_ (.A(\add_result[16] ),
    .X(_0278_));
 sky130_fd_sc_hd__clkbuf_4 _2338_ (.A(\add_result[15] ),
    .X(_0279_));
 sky130_fd_sc_hd__nor4_1 _2339_ (.A(_0277_),
    .B(_0278_),
    .C(_0279_),
    .D(\add_result[18] ),
    .Y(_0280_));
 sky130_fd_sc_hd__nand4_2 _2340_ (.A(_0270_),
    .B(_0272_),
    .C(_0276_),
    .D(_0280_),
    .Y(_0281_));
 sky130_fd_sc_hd__buf_4 _2341_ (.A(\add_result[5] ),
    .X(_0282_));
 sky130_fd_sc_hd__buf_4 _2342_ (.A(\add_result[8] ),
    .X(_0283_));
 sky130_fd_sc_hd__buf_4 _2343_ (.A(\add_result[7] ),
    .X(_0284_));
 sky130_fd_sc_hd__nor4_1 _2344_ (.A(_0282_),
    .B(_0283_),
    .C(_0284_),
    .D(\add_result[10] ),
    .Y(_0285_));
 sky130_fd_sc_hd__buf_2 _2345_ (.A(\add_result[20] ),
    .X(_0286_));
 sky130_fd_sc_hd__buf_2 _2346_ (.A(\add_result[21] ),
    .X(_0287_));
 sky130_fd_sc_hd__nor2_2 _2347_ (.A(_0286_),
    .B(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__buf_4 _2348_ (.A(\add_result[6] ),
    .X(_0289_));
 sky130_fd_sc_hd__clkbuf_4 _2349_ (.A(\add_result[14] ),
    .X(_0290_));
 sky130_fd_sc_hd__nor2_1 _2350_ (.A(_0289_),
    .B(_0290_),
    .Y(_0291_));
 sky130_fd_sc_hd__nand3_1 _2351_ (.A(_0285_),
    .B(_0288_),
    .C(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__o31a_1 _2352_ (.A1(_0266_),
    .A2(_0281_),
    .A3(_0292_),
    .B1(inexact_stage2),
    .X(_0108_));
 sky130_fd_sc_hd__nor2_2 _2353_ (.A(\add_result[25] ),
    .B(\add_result[26] ),
    .Y(_0293_));
 sky130_fd_sc_hd__nand2_1 _2354_ (.A(_0270_),
    .B(_0293_),
    .Y(_0294_));
 sky130_fd_sc_hd__inv_2 _2355_ (.A(_0294_),
    .Y(_0295_));
 sky130_fd_sc_hd__clkbuf_4 _2356_ (.A(_0295_),
    .X(_1695_));
 sky130_fd_sc_hd__or2_0 _2357_ (.A(\add_result[25] ),
    .B(\add_result[26] ),
    .X(_0296_));
 sky130_fd_sc_hd__nor2_2 _2358_ (.A(_0268_),
    .B(_0296_),
    .Y(_0297_));
 sky130_fd_sc_hd__o31ai_4 _2359_ (.A1(_0267_),
    .A2(_0269_),
    .A3(_0288_),
    .B1(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__buf_4 _2360_ (.A(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__clkinvlp_4 _2361_ (.A(_0299_),
    .Y(_1702_));
 sky130_fd_sc_hd__inv_1 _2362_ (.A(_0267_),
    .Y(_0300_));
 sky130_fd_sc_hd__nand2b_1 _2363_ (.A_N(_0287_),
    .B(_0286_),
    .Y(_0301_));
 sky130_fd_sc_hd__a21oi_1 _2364_ (.A1(_0300_),
    .A2(_0301_),
    .B1(_0269_),
    .Y(_0302_));
 sky130_fd_sc_hd__o21ai_4 _2365_ (.A1(\add_result[24] ),
    .A2(_0302_),
    .B1(_0293_),
    .Y(_0303_));
 sky130_fd_sc_hd__buf_4 _2366_ (.A(_0303_),
    .X(_1711_));
 sky130_fd_sc_hd__inv_1 _2367_ (.A(_1711_),
    .Y(_1708_));
 sky130_fd_sc_hd__buf_4 _2368_ (.A(\add_result[25] ),
    .X(_0304_));
 sky130_fd_sc_hd__clkbuf_4 _2369_ (.A(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__inv_2 _2370_ (.A(\add_result[26] ),
    .Y(_0306_));
 sky130_fd_sc_hd__o21ai_4 _2371_ (.A1(_0281_),
    .A2(_0292_),
    .B1(_0306_),
    .Y(_0307_));
 sky130_fd_sc_hd__buf_2 _2372_ (.A(_0307_),
    .X(_0308_));
 sky130_fd_sc_hd__buf_2 _2373_ (.A(\result_exp_stage2[7] ),
    .X(_0309_));
 sky130_fd_sc_hd__nand2b_1 _2374_ (.A_N(_1710_),
    .B(_1712_),
    .Y(_0310_));
 sky130_fd_sc_hd__a21o_1 _2375_ (.A1(_1704_),
    .A2(_0310_),
    .B1(_1703_),
    .X(_0311_));
 sky130_fd_sc_hd__a21oi_1 _2376_ (.A1(_1697_),
    .A2(_0311_),
    .B1(_1696_),
    .Y(_0312_));
 sky130_fd_sc_hd__clkbuf_4 _2377_ (.A(\result_exp_stage2[4] ),
    .X(_0313_));
 sky130_fd_sc_hd__nor3_1 _2378_ (.A(\result_exp_stage2[5] ),
    .B(_0313_),
    .C(\result_exp_stage2[3] ),
    .Y(_0314_));
 sky130_fd_sc_hd__nand2b_1 _2379_ (.A_N(\result_exp_stage2[6] ),
    .B(_0314_),
    .Y(_0315_));
 sky130_fd_sc_hd__or3_1 _2380_ (.A(_0309_),
    .B(_0312_),
    .C(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__clkbuf_4 _2381_ (.A(_0316_),
    .X(_0317_));
 sky130_fd_sc_hd__clkbuf_4 _2382_ (.A(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__nor3_1 _2383_ (.A(_0305_),
    .B(_0308_),
    .C(_0318_),
    .Y(_0120_));
 sky130_fd_sc_hd__clkbuf_4 _2384_ (.A(\result_exp_stage2[0] ),
    .X(_0319_));
 sky130_fd_sc_hd__inv_1 _2385_ (.A(_0319_),
    .Y(_1707_));
 sky130_fd_sc_hd__clkbuf_4 _2386_ (.A(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__buf_4 _2387_ (.A(\result_exp_stage2[5] ),
    .X(_0321_));
 sky130_fd_sc_hd__buf_4 _2388_ (.A(\result_exp_stage2[3] ),
    .X(_0322_));
 sky130_fd_sc_hd__nand4_2 _2389_ (.A(\result_exp_stage2[6] ),
    .B(_0321_),
    .C(_0313_),
    .D(_0322_),
    .Y(_0323_));
 sky130_fd_sc_hd__buf_6 _2390_ (.A(\result_exp_stage2[2] ),
    .X(_0324_));
 sky130_fd_sc_hd__nand3_1 _2391_ (.A(_0309_),
    .B(_0324_),
    .C(_1716_),
    .Y(_0325_));
 sky130_fd_sc_hd__nor2_2 _2392_ (.A(_0323_),
    .B(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__buf_4 _2393_ (.A(_0304_),
    .X(_0327_));
 sky130_fd_sc_hd__nor2_1 _2394_ (.A(_0327_),
    .B(_1710_),
    .Y(_0328_));
 sky130_fd_sc_hd__a21oi_1 _2395_ (.A1(_0305_),
    .A2(_0320_),
    .B1(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__nor2_1 _2396_ (.A(_0304_),
    .B(_0317_),
    .Y(_0330_));
 sky130_fd_sc_hd__or2_0 _2397_ (.A(_0307_),
    .B(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__buf_2 _2398_ (.A(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__o32ai_1 _2399_ (.A1(_0306_),
    .A2(_0320_),
    .A3(_0326_),
    .B1(_0329_),
    .B2(_0332_),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_1 _2400_ (.A(\result_exp_stage2[1] ),
    .Y(_1701_));
 sky130_fd_sc_hd__inv_1 _2401_ (.A(_1715_),
    .Y(_0333_));
 sky130_fd_sc_hd__buf_2 _2402_ (.A(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__mux2i_1 _2403_ (.A0(_1576_),
    .A1(\result_exp_stage2[1] ),
    .S(_0327_),
    .Y(_0335_));
 sky130_fd_sc_hd__o22ai_1 _2404_ (.A1(_0306_),
    .A2(_0334_),
    .B1(_0332_),
    .B2(_0335_),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_1 _2405_ (.A(_0324_),
    .Y(_1694_));
 sky130_fd_sc_hd__xnor2_1 _2406_ (.A(_1697_),
    .B(_1575_),
    .Y(_0336_));
 sky130_fd_sc_hd__nor2_1 _2407_ (.A(_0327_),
    .B(_0336_),
    .Y(_0337_));
 sky130_fd_sc_hd__a21oi_1 _2408_ (.A1(_0305_),
    .A2(_0324_),
    .B1(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__xor2_1 _2409_ (.A(_0324_),
    .B(_1718_),
    .X(_0339_));
 sky130_fd_sc_hd__clkbuf_4 _2410_ (.A(_0266_),
    .X(_0340_));
 sky130_fd_sc_hd__o21ai_0 _2411_ (.A1(_0326_),
    .A2(_0339_),
    .B1(_0340_),
    .Y(_0341_));
 sky130_fd_sc_hd__o21ai_0 _2412_ (.A1(_0332_),
    .A2(_0338_),
    .B1(_0341_),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_1 _2413_ (.A(_1709_),
    .Y(_1573_));
 sky130_fd_sc_hd__nor2_1 _2414_ (.A(_0304_),
    .B(_1699_),
    .Y(_0342_));
 sky130_fd_sc_hd__nor2b_1 _2415_ (.A(_1709_),
    .B_N(_1704_),
    .Y(_0343_));
 sky130_fd_sc_hd__o21ai_1 _2416_ (.A1(_1705_),
    .A2(_0343_),
    .B1(_1697_),
    .Y(_0344_));
 sky130_fd_sc_hd__nand2_1 _2417_ (.A(_0342_),
    .B(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__nand3_1 _2418_ (.A(_0324_),
    .B(\result_exp_stage2[1] ),
    .C(_0320_),
    .Y(_0346_));
 sky130_fd_sc_hd__inv_1 _2419_ (.A(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__nor2_1 _2420_ (.A(_0307_),
    .B(_0330_),
    .Y(_0348_));
 sky130_fd_sc_hd__nand2_1 _2421_ (.A(_0348_),
    .B(_0345_),
    .Y(_0349_));
 sky130_fd_sc_hd__o21ai_0 _2422_ (.A1(_0306_),
    .A2(_0347_),
    .B1(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__nand2_1 _2423_ (.A(_0322_),
    .B(_0350_),
    .Y(_0351_));
 sky130_fd_sc_hd__nor2_1 _2424_ (.A(_0322_),
    .B(_0346_),
    .Y(_0352_));
 sky130_fd_sc_hd__o21ai_0 _2425_ (.A1(_0326_),
    .A2(_0352_),
    .B1(_0340_),
    .Y(_0353_));
 sky130_fd_sc_hd__o311ai_0 _2426_ (.A1(_0322_),
    .A2(_0332_),
    .A3(_0345_),
    .B1(_0351_),
    .C1(_0353_),
    .Y(_0080_));
 sky130_fd_sc_hd__nand3_1 _2427_ (.A(_0322_),
    .B(_0324_),
    .C(_1718_),
    .Y(_0354_));
 sky130_fd_sc_hd__o22ai_1 _2428_ (.A1(_0323_),
    .A2(_0325_),
    .B1(_0354_),
    .B2(_0313_),
    .Y(_0355_));
 sky130_fd_sc_hd__a211oi_1 _2429_ (.A1(_1697_),
    .A2(_1575_),
    .B1(_1699_),
    .C1(_0304_),
    .Y(_0356_));
 sky130_fd_sc_hd__nor2b_1 _2430_ (.A(_0322_),
    .B_N(_0356_),
    .Y(_0357_));
 sky130_fd_sc_hd__nand2_1 _2431_ (.A(_0266_),
    .B(_0354_),
    .Y(_0358_));
 sky130_fd_sc_hd__o21ai_0 _2432_ (.A1(_0332_),
    .A2(_0357_),
    .B1(_0358_),
    .Y(_0359_));
 sky130_fd_sc_hd__nor3b_1 _2433_ (.A(_0313_),
    .B(_0332_),
    .C_N(_0357_),
    .Y(_0360_));
 sky130_fd_sc_hd__a221o_1 _2434_ (.A1(_0266_),
    .A2(_0355_),
    .B1(_0359_),
    .B2(_0313_),
    .C1(_0360_),
    .X(_0081_));
 sky130_fd_sc_hd__nor2_1 _2435_ (.A(_0313_),
    .B(\result_exp_stage2[3] ),
    .Y(_0361_));
 sky130_fd_sc_hd__nand3_1 _2436_ (.A(_0361_),
    .B(_0342_),
    .C(_0344_),
    .Y(_0362_));
 sky130_fd_sc_hd__nand3_1 _2437_ (.A(_0313_),
    .B(_0322_),
    .C(_0347_),
    .Y(_0363_));
 sky130_fd_sc_hd__a22o_1 _2438_ (.A1(_0266_),
    .A2(_0363_),
    .B1(_0362_),
    .B2(_0348_),
    .X(_0364_));
 sky130_fd_sc_hd__nand2_1 _2439_ (.A(_0321_),
    .B(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__nor2_1 _2440_ (.A(_0321_),
    .B(_0363_),
    .Y(_0366_));
 sky130_fd_sc_hd__o21ai_0 _2441_ (.A1(_0326_),
    .A2(_0366_),
    .B1(_0340_),
    .Y(_0367_));
 sky130_fd_sc_hd__o311ai_1 _2442_ (.A1(_0321_),
    .A2(_0332_),
    .A3(_0362_),
    .B1(_0365_),
    .C1(_0367_),
    .Y(_0082_));
 sky130_fd_sc_hd__nand2_1 _2443_ (.A(_0314_),
    .B(_0356_),
    .Y(_0368_));
 sky130_fd_sc_hd__nand2_1 _2444_ (.A(_0321_),
    .B(_0313_),
    .Y(_0369_));
 sky130_fd_sc_hd__or2_0 _2445_ (.A(_0369_),
    .B(_0354_),
    .X(_0370_));
 sky130_fd_sc_hd__a22o_1 _2446_ (.A1(_0266_),
    .A2(_0370_),
    .B1(_0368_),
    .B2(_0348_),
    .X(_0371_));
 sky130_fd_sc_hd__nand2_1 _2447_ (.A(\result_exp_stage2[6] ),
    .B(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__nor2_1 _2448_ (.A(\result_exp_stage2[6] ),
    .B(_0370_),
    .Y(_0373_));
 sky130_fd_sc_hd__o21ai_0 _2449_ (.A1(_0326_),
    .A2(_0373_),
    .B1(_0266_),
    .Y(_0374_));
 sky130_fd_sc_hd__o311ai_2 _2450_ (.A1(\result_exp_stage2[6] ),
    .A2(_0332_),
    .A3(_0368_),
    .B1(_0372_),
    .C1(_0374_),
    .Y(_0083_));
 sky130_fd_sc_hd__nor2_1 _2451_ (.A(_0315_),
    .B(_0345_),
    .Y(_0375_));
 sky130_fd_sc_hd__xnor2_1 _2452_ (.A(_0309_),
    .B(_0375_),
    .Y(_0376_));
 sky130_fd_sc_hd__nor2_1 _2453_ (.A(_0323_),
    .B(_0346_),
    .Y(_0377_));
 sky130_fd_sc_hd__xor2_1 _2454_ (.A(_0309_),
    .B(_0377_),
    .X(_0378_));
 sky130_fd_sc_hd__o21ai_0 _2455_ (.A1(_0326_),
    .A2(_0378_),
    .B1(_0340_),
    .Y(_0379_));
 sky130_fd_sc_hd__o21ai_0 _2456_ (.A1(_0332_),
    .A2(_0376_),
    .B1(_0379_),
    .Y(_0084_));
 sky130_fd_sc_hd__nor3_2 _2457_ (.A(_0309_),
    .B(_0312_),
    .C(_0315_),
    .Y(_0380_));
 sky130_fd_sc_hd__nor2_1 _2458_ (.A(_0309_),
    .B(\result_exp_stage2[6] ),
    .Y(_0381_));
 sky130_fd_sc_hd__clkinvlp_4 _2459_ (.A(_0381_),
    .Y(_0382_));
 sky130_fd_sc_hd__or4b_2 _2460_ (.A(_0313_),
    .B(\result_exp_stage2[3] ),
    .C(\result_exp_stage2[2] ),
    .D_N(_1714_),
    .X(_0383_));
 sky130_fd_sc_hd__nor3_4 _2461_ (.A(_0321_),
    .B(_0382_),
    .C(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__a21o_1 _2462_ (.A1(_0380_),
    .A2(_0384_),
    .B1(_0304_),
    .X(_0385_));
 sky130_fd_sc_hd__clkbuf_4 _2463_ (.A(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__buf_2 _2464_ (.A(_0317_),
    .X(_0387_));
 sky130_fd_sc_hd__clkbuf_4 _2465_ (.A(_1715_),
    .X(_0388_));
 sky130_fd_sc_hd__clkbuf_4 _2466_ (.A(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__buf_4 _2467_ (.A(_0319_),
    .X(_0390_));
 sky130_fd_sc_hd__and2_2 _2468_ (.A(_0390_),
    .B(\add_result[2] ),
    .X(_0391_));
 sky130_fd_sc_hd__nor3_4 _2469_ (.A(_0324_),
    .B(\result_exp_stage2[1] ),
    .C(\result_exp_stage2[0] ),
    .Y(_0392_));
 sky130_fd_sc_hd__nand2_1 _2470_ (.A(_0361_),
    .B(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__a21oi_2 _2471_ (.A1(_0383_),
    .A2(_0393_),
    .B1(\result_exp_stage2[5] ),
    .Y(_0394_));
 sky130_fd_sc_hd__nor2b_1 _2472_ (.A(\result_exp_stage2[6] ),
    .B_N(_0309_),
    .Y(_0395_));
 sky130_fd_sc_hd__nand4_1 _2473_ (.A(_0361_),
    .B(_0383_),
    .C(_0392_),
    .D(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__or3b_1 _2474_ (.A(_0383_),
    .B(_0309_),
    .C_N(\result_exp_stage2[6] ),
    .X(_0397_));
 sky130_fd_sc_hd__a21oi_1 _2475_ (.A1(_0396_),
    .A2(_0397_),
    .B1(_0321_),
    .Y(_0398_));
 sky130_fd_sc_hd__o21bai_4 _2476_ (.A1(_0382_),
    .A2(_0394_),
    .B1_N(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__clkbuf_4 _2477_ (.A(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__xnor2_4 _2478_ (.A(_0324_),
    .B(_1714_),
    .Y(_0401_));
 sky130_fd_sc_hd__buf_4 _2479_ (.A(_0401_),
    .X(_0402_));
 sky130_fd_sc_hd__clkbuf_4 _2480_ (.A(_0402_),
    .X(_0403_));
 sky130_fd_sc_hd__nand4_2 _2481_ (.A(_0389_),
    .B(_0391_),
    .C(_0400_),
    .D(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__xnor2_2 _2482_ (.A(_0322_),
    .B(_0392_),
    .Y(_0405_));
 sky130_fd_sc_hd__buf_2 _2483_ (.A(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__nor3b_2 _2484_ (.A(_0322_),
    .B(_0324_),
    .C_N(_1714_),
    .Y(_0407_));
 sky130_fd_sc_hd__xnor2_4 _2485_ (.A(_0313_),
    .B(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__xor2_2 _2486_ (.A(_0321_),
    .B(_0393_),
    .X(_0409_));
 sky130_fd_sc_hd__and2_0 _2487_ (.A(_0408_),
    .B(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__buf_2 _2488_ (.A(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__nand2_1 _2489_ (.A(_0406_),
    .B(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__nor4_1 _2490_ (.A(_0304_),
    .B(_0387_),
    .C(_0404_),
    .D(_0412_),
    .Y(_0413_));
 sky130_fd_sc_hd__a21oi_1 _2491_ (.A1(\add_result[2] ),
    .A2(_0386_),
    .B1(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__clkbuf_4 _2492_ (.A(_0266_),
    .X(_0415_));
 sky130_fd_sc_hd__nand2_1 _2493_ (.A(_0273_),
    .B(_0415_),
    .Y(_0416_));
 sky130_fd_sc_hd__o21ai_0 _2494_ (.A1(_0308_),
    .A2(_0414_),
    .B1(_0416_),
    .Y(_0085_));
 sky130_fd_sc_hd__clkbuf_4 _2495_ (.A(_0304_),
    .X(_0417_));
 sky130_fd_sc_hd__buf_2 _2496_ (.A(_0380_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_1 _2497_ (.A0(\add_result[2] ),
    .A1(_0273_),
    .S(_0390_),
    .X(_0419_));
 sky130_fd_sc_hd__nand4_2 _2498_ (.A(_0389_),
    .B(_0400_),
    .C(_0403_),
    .D(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__buf_2 _2499_ (.A(_0384_),
    .X(_0421_));
 sky130_fd_sc_hd__nand2_1 _2500_ (.A(_0273_),
    .B(_0421_),
    .Y(_0422_));
 sky130_fd_sc_hd__o21ai_0 _2501_ (.A1(_0412_),
    .A2(_0420_),
    .B1(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__clkbuf_4 _2502_ (.A(_0380_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2i_2 _2503_ (.A0(\add_result[2] ),
    .A1(_0273_),
    .S(_1711_),
    .Y(_0425_));
 sky130_fd_sc_hd__nor3_1 _2504_ (.A(_0297_),
    .B(_0424_),
    .C(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__a21oi_1 _2505_ (.A1(_0418_),
    .A2(_0423_),
    .B1(_0426_),
    .Y(_0427_));
 sky130_fd_sc_hd__nor2_1 _2506_ (.A(_0417_),
    .B(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__a21oi_1 _2507_ (.A1(_0273_),
    .A2(_0305_),
    .B1(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__nand2_1 _2508_ (.A(_0271_),
    .B(_0415_),
    .Y(_0430_));
 sky130_fd_sc_hd__o21ai_0 _2509_ (.A1(_0308_),
    .A2(_0429_),
    .B1(_0430_),
    .Y(_0096_));
 sky130_fd_sc_hd__clkbuf_4 _2510_ (.A(_0304_),
    .X(_0431_));
 sky130_fd_sc_hd__buf_2 _2511_ (.A(_0388_),
    .X(_0432_));
 sky130_fd_sc_hd__mux2i_2 _2512_ (.A0(_0273_),
    .A1(_0271_),
    .S(_0390_),
    .Y(_0433_));
 sky130_fd_sc_hd__nand2_1 _2513_ (.A(_0432_),
    .B(_0433_),
    .Y(_0434_));
 sky130_fd_sc_hd__o2111ai_4 _2514_ (.A1(_0389_),
    .A2(_0391_),
    .B1(_0399_),
    .C1(_0402_),
    .D1(_0434_),
    .Y(_0435_));
 sky130_fd_sc_hd__nor2_1 _2515_ (.A(_0412_),
    .B(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__a211oi_1 _2516_ (.A1(_0271_),
    .A2(_0421_),
    .B1(_0436_),
    .C1(_0387_),
    .Y(_0437_));
 sky130_fd_sc_hd__buf_4 _2517_ (.A(_0294_),
    .X(_1698_));
 sky130_fd_sc_hd__buf_4 _2518_ (.A(_0298_),
    .X(_1574_));
 sky130_fd_sc_hd__mux2i_2 _2519_ (.A0(_0273_),
    .A1(_0271_),
    .S(_1711_),
    .Y(_0438_));
 sky130_fd_sc_hd__a21oi_1 _2520_ (.A1(\add_result[2] ),
    .A2(_1711_),
    .B1(_1574_),
    .Y(_0439_));
 sky130_fd_sc_hd__a21oi_1 _2521_ (.A1(_1574_),
    .A2(_0438_),
    .B1(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__a21oi_1 _2522_ (.A1(_1698_),
    .A2(_0440_),
    .B1(_0418_),
    .Y(_0441_));
 sky130_fd_sc_hd__nor3_1 _2523_ (.A(_0431_),
    .B(_0437_),
    .C(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__a21oi_1 _2524_ (.A1(_0271_),
    .A2(_0305_),
    .B1(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__nand2_1 _2525_ (.A(_0282_),
    .B(_0415_),
    .Y(_0444_));
 sky130_fd_sc_hd__o21ai_0 _2526_ (.A1(_0308_),
    .A2(_0443_),
    .B1(_0444_),
    .Y(_0100_));
 sky130_fd_sc_hd__xor2_4 _2527_ (.A(_0322_),
    .B(_0392_),
    .X(_0445_));
 sky130_fd_sc_hd__nand2_2 _2528_ (.A(_0408_),
    .B(_0409_),
    .Y(_0446_));
 sky130_fd_sc_hd__nor2_1 _2529_ (.A(_0445_),
    .B(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__o21ba_2 _2530_ (.A1(_0382_),
    .A2(_0394_),
    .B1_N(_0398_),
    .X(_0448_));
 sky130_fd_sc_hd__xor2_4 _2531_ (.A(_0324_),
    .B(_1714_),
    .X(_0449_));
 sky130_fd_sc_hd__buf_2 _2532_ (.A(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__buf_2 _2533_ (.A(_0388_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2i_2 _2534_ (.A0(_0271_),
    .A1(_0282_),
    .S(_0390_),
    .Y(_0452_));
 sky130_fd_sc_hd__nand2_1 _2535_ (.A(_0451_),
    .B(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__o21ai_0 _2536_ (.A1(_0451_),
    .A2(_0419_),
    .B1(_0453_),
    .Y(_0454_));
 sky130_fd_sc_hd__nor3_1 _2537_ (.A(_0448_),
    .B(_0450_),
    .C(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__a221oi_1 _2538_ (.A1(_0282_),
    .A2(_0421_),
    .B1(_0447_),
    .B2(_0455_),
    .C1(_0387_),
    .Y(_0456_));
 sky130_fd_sc_hd__mux2i_1 _2539_ (.A0(_0271_),
    .A1(_0282_),
    .S(_1711_),
    .Y(_0457_));
 sky130_fd_sc_hd__mux2i_1 _2540_ (.A0(_0425_),
    .A1(_0457_),
    .S(_1574_),
    .Y(_0458_));
 sky130_fd_sc_hd__a21oi_1 _2541_ (.A1(_1698_),
    .A2(_0458_),
    .B1(_0424_),
    .Y(_0459_));
 sky130_fd_sc_hd__nor3_1 _2542_ (.A(_0431_),
    .B(_0456_),
    .C(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__a21oi_1 _2543_ (.A1(_0282_),
    .A2(_0305_),
    .B1(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__nand2_1 _2544_ (.A(_0289_),
    .B(_0415_),
    .Y(_0462_));
 sky130_fd_sc_hd__o21ai_0 _2545_ (.A1(_0308_),
    .A2(_0461_),
    .B1(_0462_),
    .Y(_0101_));
 sky130_fd_sc_hd__mux2i_1 _2546_ (.A0(_0282_),
    .A1(_0289_),
    .S(_1711_),
    .Y(_0463_));
 sky130_fd_sc_hd__mux2i_2 _2547_ (.A0(_0438_),
    .A1(_0463_),
    .S(_0299_),
    .Y(_0464_));
 sky130_fd_sc_hd__nand2_1 _2548_ (.A(_1698_),
    .B(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__nand4_1 _2549_ (.A(\add_result[2] ),
    .B(_1695_),
    .C(_1574_),
    .D(_1711_),
    .Y(_0466_));
 sky130_fd_sc_hd__nor2_1 _2550_ (.A(_0391_),
    .B(_0401_),
    .Y(_0467_));
 sky130_fd_sc_hd__mux2_1 _2551_ (.A0(_0282_),
    .A1(_0289_),
    .S(_0319_),
    .X(_0468_));
 sky130_fd_sc_hd__nor2_1 _2552_ (.A(_0449_),
    .B(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__nor3_1 _2553_ (.A(_0334_),
    .B(_0467_),
    .C(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__nor3_1 _2554_ (.A(_0432_),
    .B(_0449_),
    .C(_0433_),
    .Y(_0471_));
 sky130_fd_sc_hd__o21ai_2 _2555_ (.A1(_0470_),
    .A2(_0471_),
    .B1(_0399_),
    .Y(_0472_));
 sky130_fd_sc_hd__nor2_1 _2556_ (.A(_0412_),
    .B(_0472_),
    .Y(_0473_));
 sky130_fd_sc_hd__a211oi_1 _2557_ (.A1(_0289_),
    .A2(_0421_),
    .B1(_0473_),
    .C1(_0387_),
    .Y(_0474_));
 sky130_fd_sc_hd__a311oi_1 _2558_ (.A1(_0318_),
    .A2(_0465_),
    .A3(_0466_),
    .B1(_0474_),
    .C1(_0431_),
    .Y(_0475_));
 sky130_fd_sc_hd__a21oi_1 _2559_ (.A1(_0289_),
    .A2(_0305_),
    .B1(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__nand2_1 _2560_ (.A(_0284_),
    .B(_0415_),
    .Y(_0477_));
 sky130_fd_sc_hd__o21ai_0 _2561_ (.A1(_0308_),
    .A2(_0476_),
    .B1(_0477_),
    .Y(_0102_));
 sky130_fd_sc_hd__buf_2 _2562_ (.A(_0294_),
    .X(_0478_));
 sky130_fd_sc_hd__buf_4 _2563_ (.A(_0303_),
    .X(_0479_));
 sky130_fd_sc_hd__mux2i_1 _2564_ (.A0(_0289_),
    .A1(_0284_),
    .S(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__mux2i_1 _2565_ (.A0(_0457_),
    .A1(_0480_),
    .S(_0299_),
    .Y(_0481_));
 sky130_fd_sc_hd__nor3_1 _2566_ (.A(_0478_),
    .B(_1702_),
    .C(_0425_),
    .Y(_0482_));
 sky130_fd_sc_hd__a211oi_1 _2567_ (.A1(_0478_),
    .A2(_0481_),
    .B1(_0482_),
    .C1(_0424_),
    .Y(_0483_));
 sky130_fd_sc_hd__mux4_1 _2568_ (.A0(_0273_),
    .A1(_0284_),
    .A2(\add_result[2] ),
    .A3(_0289_),
    .S0(_0401_),
    .S1(_1707_),
    .X(_0484_));
 sky130_fd_sc_hd__nor3_1 _2569_ (.A(_0388_),
    .B(_0449_),
    .C(_0452_),
    .Y(_0485_));
 sky130_fd_sc_hd__a21oi_1 _2570_ (.A1(_0432_),
    .A2(_0484_),
    .B1(_0485_),
    .Y(_0486_));
 sky130_fd_sc_hd__nor2_1 _2571_ (.A(_0448_),
    .B(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__a221oi_1 _2572_ (.A1(_0284_),
    .A2(_0421_),
    .B1(_0447_),
    .B2(_0487_),
    .C1(_0387_),
    .Y(_0488_));
 sky130_fd_sc_hd__nor3_1 _2573_ (.A(_0431_),
    .B(_0483_),
    .C(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__a21oi_1 _2574_ (.A1(_0284_),
    .A2(_0305_),
    .B1(_0489_),
    .Y(_0490_));
 sky130_fd_sc_hd__nand2_1 _2575_ (.A(_0283_),
    .B(_0415_),
    .Y(_0491_));
 sky130_fd_sc_hd__o21ai_0 _2576_ (.A1(_0308_),
    .A2(_0490_),
    .B1(_0491_),
    .Y(_0103_));
 sky130_fd_sc_hd__nand2_1 _2577_ (.A(_1695_),
    .B(_0440_),
    .Y(_0492_));
 sky130_fd_sc_hd__mux2i_1 _2578_ (.A0(_0284_),
    .A1(_0283_),
    .S(_0479_),
    .Y(_0493_));
 sky130_fd_sc_hd__mux2i_1 _2579_ (.A0(_0463_),
    .A1(_0493_),
    .S(_1574_),
    .Y(_0494_));
 sky130_fd_sc_hd__nand2_1 _2580_ (.A(_1698_),
    .B(_0494_),
    .Y(_0495_));
 sky130_fd_sc_hd__mux2i_1 _2581_ (.A0(_0284_),
    .A1(_0283_),
    .S(_0319_),
    .Y(_0496_));
 sky130_fd_sc_hd__nand2_1 _2582_ (.A(_0388_),
    .B(_0496_),
    .Y(_0497_));
 sky130_fd_sc_hd__o211ai_2 _2583_ (.A1(_0388_),
    .A2(_0468_),
    .B1(_0497_),
    .C1(_0399_),
    .Y(_0498_));
 sky130_fd_sc_hd__o2111ai_1 _2584_ (.A1(_0432_),
    .A2(_0391_),
    .B1(_0399_),
    .C1(_0449_),
    .D1(_0434_),
    .Y(_0499_));
 sky130_fd_sc_hd__o21ai_2 _2585_ (.A1(_0449_),
    .A2(_0498_),
    .B1(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__a221oi_1 _2586_ (.A1(_0283_),
    .A2(_0421_),
    .B1(_0447_),
    .B2(_0500_),
    .C1(_0317_),
    .Y(_0501_));
 sky130_fd_sc_hd__a311oi_1 _2587_ (.A1(_0318_),
    .A2(_0492_),
    .A3(_0495_),
    .B1(_0501_),
    .C1(_0431_),
    .Y(_0502_));
 sky130_fd_sc_hd__a21oi_1 _2588_ (.A1(_0283_),
    .A2(_0305_),
    .B1(_0502_),
    .Y(_0503_));
 sky130_fd_sc_hd__nand2_1 _2589_ (.A(_0274_),
    .B(_0415_),
    .Y(_0504_));
 sky130_fd_sc_hd__o21ai_0 _2590_ (.A1(_0308_),
    .A2(_0503_),
    .B1(_0504_),
    .Y(_0104_));
 sky130_fd_sc_hd__nand2_1 _2591_ (.A(_1695_),
    .B(_0458_),
    .Y(_0505_));
 sky130_fd_sc_hd__mux2i_1 _2592_ (.A0(_0283_),
    .A1(_0274_),
    .S(_0479_),
    .Y(_0506_));
 sky130_fd_sc_hd__mux2i_1 _2593_ (.A0(_0480_),
    .A1(_0506_),
    .S(_0299_),
    .Y(_0507_));
 sky130_fd_sc_hd__nand2_1 _2594_ (.A(_1698_),
    .B(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__and2_0 _2595_ (.A(_0284_),
    .B(_0390_),
    .X(_0509_));
 sky130_fd_sc_hd__nor2b_1 _2596_ (.A(_0319_),
    .B_N(_0289_),
    .Y(_0510_));
 sky130_fd_sc_hd__mux2i_1 _2597_ (.A0(_0283_),
    .A1(_0274_),
    .S(_0319_),
    .Y(_0511_));
 sky130_fd_sc_hd__nand2_1 _2598_ (.A(_0432_),
    .B(_0511_),
    .Y(_0512_));
 sky130_fd_sc_hd__o31a_1 _2599_ (.A1(_0388_),
    .A2(_0509_),
    .A3(_0510_),
    .B1(_0512_),
    .X(_0513_));
 sky130_fd_sc_hd__nand2_1 _2600_ (.A(_0402_),
    .B(_0513_),
    .Y(_0514_));
 sky130_fd_sc_hd__o21ai_0 _2601_ (.A1(_0402_),
    .A2(_0454_),
    .B1(_0514_),
    .Y(_0515_));
 sky130_fd_sc_hd__nand2_1 _2602_ (.A(_0400_),
    .B(_0515_),
    .Y(_0516_));
 sky130_fd_sc_hd__nand2_1 _2603_ (.A(_0274_),
    .B(_0384_),
    .Y(_0517_));
 sky130_fd_sc_hd__o21ai_0 _2604_ (.A1(_0412_),
    .A2(_0516_),
    .B1(_0517_),
    .Y(_0518_));
 sky130_fd_sc_hd__nor2_1 _2605_ (.A(_0387_),
    .B(_0518_),
    .Y(_0519_));
 sky130_fd_sc_hd__a311oi_1 _2606_ (.A1(_0318_),
    .A2(_0505_),
    .A3(_0508_),
    .B1(_0519_),
    .C1(_0431_),
    .Y(_0520_));
 sky130_fd_sc_hd__a21oi_1 _2607_ (.A1(_0274_),
    .A2(_0327_),
    .B1(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__nand2_1 _2608_ (.A(\add_result[10] ),
    .B(_0415_),
    .Y(_0522_));
 sky130_fd_sc_hd__o21ai_0 _2609_ (.A1(_0308_),
    .A2(_0521_),
    .B1(_0522_),
    .Y(_0105_));
 sky130_fd_sc_hd__clkbuf_2 _2610_ (.A(\add_result[26] ),
    .X(_0523_));
 sky130_fd_sc_hd__clkbuf_2 _2611_ (.A(_0406_),
    .X(_0524_));
 sky130_fd_sc_hd__nand2_1 _2612_ (.A(_0334_),
    .B(_0496_),
    .Y(_0525_));
 sky130_fd_sc_hd__mux2i_1 _2613_ (.A0(_0274_),
    .A1(\add_result[10] ),
    .S(_0319_),
    .Y(_0526_));
 sky130_fd_sc_hd__nand2_1 _2614_ (.A(_0451_),
    .B(_0526_),
    .Y(_0527_));
 sky130_fd_sc_hd__nand3_1 _2615_ (.A(_0399_),
    .B(_0525_),
    .C(_0527_),
    .Y(_0528_));
 sky130_fd_sc_hd__nand2_1 _2616_ (.A(_0451_),
    .B(_0468_),
    .Y(_0529_));
 sky130_fd_sc_hd__o21ai_1 _2617_ (.A1(_0451_),
    .A2(_0433_),
    .B1(_0529_),
    .Y(_0530_));
 sky130_fd_sc_hd__a21oi_1 _2618_ (.A1(_0400_),
    .A2(_0530_),
    .B1(_0402_),
    .Y(_0531_));
 sky130_fd_sc_hd__a21oi_1 _2619_ (.A1(_0403_),
    .A2(_0528_),
    .B1(_0531_),
    .Y(_0532_));
 sky130_fd_sc_hd__nand2_1 _2620_ (.A(_0524_),
    .B(_0532_),
    .Y(_0533_));
 sky130_fd_sc_hd__o21ai_0 _2621_ (.A1(_0404_),
    .A2(_0524_),
    .B1(_0533_),
    .Y(_0534_));
 sky130_fd_sc_hd__nand2_1 _2622_ (.A(_0295_),
    .B(_0464_),
    .Y(_0535_));
 sky130_fd_sc_hd__mux2i_1 _2623_ (.A0(_0274_),
    .A1(\add_result[10] ),
    .S(_0479_),
    .Y(_0536_));
 sky130_fd_sc_hd__mux2i_1 _2624_ (.A0(_0493_),
    .A1(_0536_),
    .S(_0299_),
    .Y(_0537_));
 sky130_fd_sc_hd__nand2_1 _2625_ (.A(_0478_),
    .B(_0537_),
    .Y(_0538_));
 sky130_fd_sc_hd__a21oi_1 _2626_ (.A1(_0535_),
    .A2(_0538_),
    .B1(_0424_),
    .Y(_0539_));
 sky130_fd_sc_hd__a31oi_1 _2627_ (.A1(_0418_),
    .A2(_0411_),
    .A3(_0534_),
    .B1(_0539_),
    .Y(_0540_));
 sky130_fd_sc_hd__a2bb2oi_1 _2628_ (.A1_N(_0417_),
    .A2_N(_0540_),
    .B1(_0386_),
    .B2(\add_result[10] ),
    .Y(_0541_));
 sky130_fd_sc_hd__nand2_1 _2629_ (.A(\add_result[11] ),
    .B(_0415_),
    .Y(_0542_));
 sky130_fd_sc_hd__o21ai_0 _2630_ (.A1(_0523_),
    .A2(_0541_),
    .B1(_0542_),
    .Y(_0106_));
 sky130_fd_sc_hd__nand2_1 _2631_ (.A(_1695_),
    .B(_0481_),
    .Y(_0543_));
 sky130_fd_sc_hd__mux2i_1 _2632_ (.A0(\add_result[10] ),
    .A1(\add_result[11] ),
    .S(_0479_),
    .Y(_0544_));
 sky130_fd_sc_hd__mux2i_1 _2633_ (.A0(_0506_),
    .A1(_0544_),
    .S(_0299_),
    .Y(_0545_));
 sky130_fd_sc_hd__nand2_1 _2634_ (.A(_0478_),
    .B(_0545_),
    .Y(_0546_));
 sky130_fd_sc_hd__nand2_1 _2635_ (.A(_0543_),
    .B(_0546_),
    .Y(_0547_));
 sky130_fd_sc_hd__mux2_1 _2636_ (.A0(\add_result[10] ),
    .A1(\add_result[11] ),
    .S(\result_exp_stage2[0] ),
    .X(_0548_));
 sky130_fd_sc_hd__nor2_1 _2637_ (.A(_0333_),
    .B(_0548_),
    .Y(_0549_));
 sky130_fd_sc_hd__a21oi_1 _2638_ (.A1(_0334_),
    .A2(_0511_),
    .B1(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__nor3_1 _2639_ (.A(_0334_),
    .B(_0509_),
    .C(_0510_),
    .Y(_0551_));
 sky130_fd_sc_hd__a211oi_1 _2640_ (.A1(_0334_),
    .A2(_0452_),
    .B1(_0551_),
    .C1(_0402_),
    .Y(_0552_));
 sky130_fd_sc_hd__a21oi_1 _2641_ (.A1(_0402_),
    .A2(_0550_),
    .B1(_0552_),
    .Y(_0553_));
 sky130_fd_sc_hd__nor2_1 _2642_ (.A(_0448_),
    .B(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__nor2_1 _2643_ (.A(_0406_),
    .B(_0420_),
    .Y(_0555_));
 sky130_fd_sc_hd__a21oi_1 _2644_ (.A1(_0524_),
    .A2(_0554_),
    .B1(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__nor3_1 _2645_ (.A(_0387_),
    .B(_0446_),
    .C(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__a21oi_1 _2646_ (.A1(_0387_),
    .A2(_0547_),
    .B1(_0557_),
    .Y(_0558_));
 sky130_fd_sc_hd__a2bb2oi_1 _2647_ (.A1_N(_0417_),
    .A2_N(_0558_),
    .B1(_0386_),
    .B2(\add_result[11] ),
    .Y(_0559_));
 sky130_fd_sc_hd__buf_2 _2648_ (.A(_0266_),
    .X(_0560_));
 sky130_fd_sc_hd__nand2_1 _2649_ (.A(_0275_),
    .B(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__o21ai_0 _2650_ (.A1(_0523_),
    .A2(_0559_),
    .B1(_0561_),
    .Y(_0107_));
 sky130_fd_sc_hd__nand2_1 _2651_ (.A(_1695_),
    .B(_0494_),
    .Y(_0562_));
 sky130_fd_sc_hd__mux2i_1 _2652_ (.A0(\add_result[11] ),
    .A1(_0275_),
    .S(_0479_),
    .Y(_0563_));
 sky130_fd_sc_hd__mux2i_1 _2653_ (.A0(_0536_),
    .A1(_0563_),
    .S(_0299_),
    .Y(_0564_));
 sky130_fd_sc_hd__nand2_1 _2654_ (.A(_1698_),
    .B(_0564_),
    .Y(_0565_));
 sky130_fd_sc_hd__mux2_1 _2655_ (.A0(\add_result[11] ),
    .A1(_0275_),
    .S(\result_exp_stage2[0] ),
    .X(_0566_));
 sky130_fd_sc_hd__nand2_1 _2656_ (.A(_0334_),
    .B(_0526_),
    .Y(_0567_));
 sky130_fd_sc_hd__o211ai_1 _2657_ (.A1(_0334_),
    .A2(_0566_),
    .B1(_0567_),
    .C1(_0399_),
    .Y(_0568_));
 sky130_fd_sc_hd__mux2_1 _2658_ (.A0(_0498_),
    .A1(_0568_),
    .S(_0401_),
    .X(_0569_));
 sky130_fd_sc_hd__mux2i_1 _2659_ (.A0(_0435_),
    .A1(_0569_),
    .S(_0406_),
    .Y(_0570_));
 sky130_fd_sc_hd__a221oi_2 _2660_ (.A1(_0275_),
    .A2(_0384_),
    .B1(_0411_),
    .B2(_0570_),
    .C1(_0317_),
    .Y(_0571_));
 sky130_fd_sc_hd__a311oi_2 _2661_ (.A1(_0318_),
    .A2(_0562_),
    .A3(_0565_),
    .B1(_0571_),
    .C1(_0431_),
    .Y(_0572_));
 sky130_fd_sc_hd__a21oi_1 _2662_ (.A1(_0275_),
    .A2(_0327_),
    .B1(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__nand2_1 _2663_ (.A(_0277_),
    .B(_0560_),
    .Y(_0574_));
 sky130_fd_sc_hd__o21ai_0 _2664_ (.A1(_0523_),
    .A2(_0573_),
    .B1(_0574_),
    .Y(_0086_));
 sky130_fd_sc_hd__mux2i_1 _2665_ (.A0(_0275_),
    .A1(_0277_),
    .S(_0390_),
    .Y(_0575_));
 sky130_fd_sc_hd__nand2_1 _2666_ (.A(_0451_),
    .B(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__o21ai_0 _2667_ (.A1(_0451_),
    .A2(_0548_),
    .B1(_0576_),
    .Y(_0577_));
 sky130_fd_sc_hd__nand2_1 _2668_ (.A(_0450_),
    .B(_0513_),
    .Y(_0578_));
 sky130_fd_sc_hd__o21ai_0 _2669_ (.A1(_0450_),
    .A2(_0577_),
    .B1(_0578_),
    .Y(_0579_));
 sky130_fd_sc_hd__nand2_1 _2670_ (.A(_0400_),
    .B(_0579_),
    .Y(_0580_));
 sky130_fd_sc_hd__nand2_1 _2671_ (.A(_0445_),
    .B(_0455_),
    .Y(_0581_));
 sky130_fd_sc_hd__o21ai_0 _2672_ (.A1(_0445_),
    .A2(_0580_),
    .B1(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__a22oi_1 _2673_ (.A1(_0277_),
    .A2(_0421_),
    .B1(_0411_),
    .B2(_0582_),
    .Y(_0583_));
 sky130_fd_sc_hd__nand2_1 _2674_ (.A(_0295_),
    .B(_0507_),
    .Y(_0584_));
 sky130_fd_sc_hd__mux2i_1 _2675_ (.A0(_0275_),
    .A1(_0277_),
    .S(_0303_),
    .Y(_0585_));
 sky130_fd_sc_hd__mux2i_1 _2676_ (.A0(_0544_),
    .A1(_0585_),
    .S(_0298_),
    .Y(_0586_));
 sky130_fd_sc_hd__nand2_1 _2677_ (.A(_0478_),
    .B(_0586_),
    .Y(_0587_));
 sky130_fd_sc_hd__and3_1 _2678_ (.A(_0317_),
    .B(_0584_),
    .C(_0587_),
    .X(_0588_));
 sky130_fd_sc_hd__a211oi_2 _2679_ (.A1(_0418_),
    .A2(_0583_),
    .B1(_0588_),
    .C1(_0417_),
    .Y(_0589_));
 sky130_fd_sc_hd__a21oi_1 _2680_ (.A1(_0277_),
    .A2(_0327_),
    .B1(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__nand2_1 _2681_ (.A(_0290_),
    .B(_0560_),
    .Y(_0591_));
 sky130_fd_sc_hd__o21ai_1 _2682_ (.A1(_0523_),
    .A2(_0590_),
    .B1(_0591_),
    .Y(_0087_));
 sky130_fd_sc_hd__nor2_1 _2683_ (.A(_0388_),
    .B(_0566_),
    .Y(_0592_));
 sky130_fd_sc_hd__mux2_1 _2684_ (.A0(_0277_),
    .A1(_0290_),
    .S(_0319_),
    .X(_0593_));
 sky130_fd_sc_hd__nor2_1 _2685_ (.A(_0333_),
    .B(_0593_),
    .Y(_0594_));
 sky130_fd_sc_hd__or3_1 _2686_ (.A(_0448_),
    .B(_0592_),
    .C(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__mux2i_1 _2687_ (.A0(_0528_),
    .A1(_0595_),
    .S(_0402_),
    .Y(_0596_));
 sky130_fd_sc_hd__nor2_1 _2688_ (.A(_0406_),
    .B(_0472_),
    .Y(_0597_));
 sky130_fd_sc_hd__a21oi_1 _2689_ (.A1(_0406_),
    .A2(_0596_),
    .B1(_0597_),
    .Y(_0598_));
 sky130_fd_sc_hd__a2bb2oi_1 _2690_ (.A1_N(_0446_),
    .A2_N(_0598_),
    .B1(_0290_),
    .B2(_0421_),
    .Y(_0599_));
 sky130_fd_sc_hd__nand2_1 _2691_ (.A(_0295_),
    .B(_0537_),
    .Y(_0600_));
 sky130_fd_sc_hd__mux2i_1 _2692_ (.A0(_0277_),
    .A1(_0290_),
    .S(_0303_),
    .Y(_0601_));
 sky130_fd_sc_hd__mux2i_1 _2693_ (.A0(_0563_),
    .A1(_0601_),
    .S(_0298_),
    .Y(_0602_));
 sky130_fd_sc_hd__nand2_1 _2694_ (.A(_0478_),
    .B(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__and3_1 _2695_ (.A(_0317_),
    .B(_0600_),
    .C(_0603_),
    .X(_0604_));
 sky130_fd_sc_hd__a211oi_1 _2696_ (.A1(_0418_),
    .A2(_0599_),
    .B1(_0604_),
    .C1(_0417_),
    .Y(_0605_));
 sky130_fd_sc_hd__a21oi_1 _2697_ (.A1(_0290_),
    .A2(_0327_),
    .B1(_0605_),
    .Y(_0606_));
 sky130_fd_sc_hd__nand2_1 _2698_ (.A(_0279_),
    .B(_0560_),
    .Y(_0607_));
 sky130_fd_sc_hd__o21ai_0 _2699_ (.A1(_0523_),
    .A2(_0606_),
    .B1(_0607_),
    .Y(_0088_));
 sky130_fd_sc_hd__nand2_1 _2700_ (.A(_1695_),
    .B(_0545_),
    .Y(_0608_));
 sky130_fd_sc_hd__mux2i_1 _2701_ (.A0(_0290_),
    .A1(_0279_),
    .S(_1711_),
    .Y(_0609_));
 sky130_fd_sc_hd__mux2i_1 _2702_ (.A0(_0585_),
    .A1(_0609_),
    .S(_1574_),
    .Y(_0610_));
 sky130_fd_sc_hd__nand2_1 _2703_ (.A(_1698_),
    .B(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__mux2i_1 _2704_ (.A0(_0290_),
    .A1(_0279_),
    .S(_0390_),
    .Y(_0612_));
 sky130_fd_sc_hd__mux2i_1 _2705_ (.A0(_0575_),
    .A1(_0612_),
    .S(_0388_),
    .Y(_0613_));
 sky130_fd_sc_hd__nand2_1 _2706_ (.A(_0401_),
    .B(_0613_),
    .Y(_0614_));
 sky130_fd_sc_hd__nand2_1 _2707_ (.A(_0449_),
    .B(_0550_),
    .Y(_0615_));
 sky130_fd_sc_hd__a21oi_1 _2708_ (.A1(_0614_),
    .A2(_0615_),
    .B1(_0448_),
    .Y(_0616_));
 sky130_fd_sc_hd__mux2_1 _2709_ (.A0(_0487_),
    .A1(_0616_),
    .S(_0405_),
    .X(_0617_));
 sky130_fd_sc_hd__a221oi_2 _2710_ (.A1(_0279_),
    .A2(_0384_),
    .B1(_0411_),
    .B2(_0617_),
    .C1(_0317_),
    .Y(_0618_));
 sky130_fd_sc_hd__a311oi_2 _2711_ (.A1(_0318_),
    .A2(_0608_),
    .A3(_0611_),
    .B1(_0618_),
    .C1(_0431_),
    .Y(_0619_));
 sky130_fd_sc_hd__a21oi_1 _2712_ (.A1(_0279_),
    .A2(_0327_),
    .B1(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__nand2_1 _2713_ (.A(_0278_),
    .B(_0560_),
    .Y(_0621_));
 sky130_fd_sc_hd__o21ai_0 _2714_ (.A1(_0523_),
    .A2(_0620_),
    .B1(_0621_),
    .Y(_0089_));
 sky130_fd_sc_hd__mux2i_1 _2715_ (.A0(_0279_),
    .A1(_0278_),
    .S(_0390_),
    .Y(_0622_));
 sky130_fd_sc_hd__nand2_1 _2716_ (.A(_0432_),
    .B(_0622_),
    .Y(_0623_));
 sky130_fd_sc_hd__o211ai_1 _2717_ (.A1(_0432_),
    .A2(_0593_),
    .B1(_0623_),
    .C1(_0399_),
    .Y(_0624_));
 sky130_fd_sc_hd__mux2i_2 _2718_ (.A0(_0568_),
    .A1(_0624_),
    .S(_0402_),
    .Y(_0625_));
 sky130_fd_sc_hd__mux2_1 _2719_ (.A0(_0500_),
    .A1(_0625_),
    .S(_0405_),
    .X(_0626_));
 sky130_fd_sc_hd__a22oi_1 _2720_ (.A1(_0278_),
    .A2(_0421_),
    .B1(_0411_),
    .B2(_0626_),
    .Y(_0627_));
 sky130_fd_sc_hd__nand2_1 _2721_ (.A(_0295_),
    .B(_0564_),
    .Y(_0628_));
 sky130_fd_sc_hd__mux2i_2 _2722_ (.A0(_0279_),
    .A1(_0278_),
    .S(_0303_),
    .Y(_0629_));
 sky130_fd_sc_hd__mux2i_1 _2723_ (.A0(_0601_),
    .A1(_0629_),
    .S(_0298_),
    .Y(_0630_));
 sky130_fd_sc_hd__nand2_1 _2724_ (.A(_0478_),
    .B(_0630_),
    .Y(_0631_));
 sky130_fd_sc_hd__and3_1 _2725_ (.A(_0317_),
    .B(_0628_),
    .C(_0631_),
    .X(_0632_));
 sky130_fd_sc_hd__a211oi_1 _2726_ (.A1(_0418_),
    .A2(_0627_),
    .B1(_0632_),
    .C1(_0431_),
    .Y(_0633_));
 sky130_fd_sc_hd__a21oi_1 _2727_ (.A1(_0278_),
    .A2(_0327_),
    .B1(_0633_),
    .Y(_0634_));
 sky130_fd_sc_hd__nand2_1 _2728_ (.A(\add_result[17] ),
    .B(_0560_),
    .Y(_0635_));
 sky130_fd_sc_hd__o21ai_0 _2729_ (.A1(_0523_),
    .A2(_0634_),
    .B1(_0635_),
    .Y(_0090_));
 sky130_fd_sc_hd__nand2_1 _2730_ (.A(_1695_),
    .B(_0586_),
    .Y(_0636_));
 sky130_fd_sc_hd__mux2i_1 _2731_ (.A0(_0278_),
    .A1(\add_result[17] ),
    .S(_0479_),
    .Y(_0637_));
 sky130_fd_sc_hd__mux2i_1 _2732_ (.A0(_0609_),
    .A1(_0637_),
    .S(_0299_),
    .Y(_0638_));
 sky130_fd_sc_hd__nand2_1 _2733_ (.A(_1698_),
    .B(_0638_),
    .Y(_0639_));
 sky130_fd_sc_hd__mux2_1 _2734_ (.A0(_0278_),
    .A1(\add_result[17] ),
    .S(_0319_),
    .X(_0640_));
 sky130_fd_sc_hd__nor2_1 _2735_ (.A(_0334_),
    .B(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__a21oi_1 _2736_ (.A1(_0334_),
    .A2(_0612_),
    .B1(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__nand2_1 _2737_ (.A(_0402_),
    .B(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__o21ai_0 _2738_ (.A1(_0403_),
    .A2(_0577_),
    .B1(_0643_),
    .Y(_0644_));
 sky130_fd_sc_hd__nand3_1 _2739_ (.A(_0400_),
    .B(_0406_),
    .C(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__o21ai_0 _2740_ (.A1(_0524_),
    .A2(_0516_),
    .B1(_0645_),
    .Y(_0646_));
 sky130_fd_sc_hd__a21oi_1 _2741_ (.A1(_0411_),
    .A2(_0646_),
    .B1(_0387_),
    .Y(_0647_));
 sky130_fd_sc_hd__a311oi_2 _2742_ (.A1(_0318_),
    .A2(_0636_),
    .A3(_0639_),
    .B1(_0647_),
    .C1(_0431_),
    .Y(_0648_));
 sky130_fd_sc_hd__a21oi_1 _2743_ (.A1(\add_result[17] ),
    .A2(_0386_),
    .B1(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__nand2_1 _2744_ (.A(\add_result[18] ),
    .B(_0560_),
    .Y(_0650_));
 sky130_fd_sc_hd__o21ai_1 _2745_ (.A1(_0523_),
    .A2(_0649_),
    .B1(_0650_),
    .Y(_0091_));
 sky130_fd_sc_hd__and2_0 _2746_ (.A(\add_result[18] ),
    .B(_0390_),
    .X(_0651_));
 sky130_fd_sc_hd__nor2b_1 _2747_ (.A(_0390_),
    .B_N(\add_result[17] ),
    .Y(_0652_));
 sky130_fd_sc_hd__o21ai_0 _2748_ (.A1(_0651_),
    .A2(_0652_),
    .B1(_0451_),
    .Y(_0653_));
 sky130_fd_sc_hd__o21ai_1 _2749_ (.A1(_0451_),
    .A2(_0622_),
    .B1(_0653_),
    .Y(_0654_));
 sky130_fd_sc_hd__nand3_1 _2750_ (.A(_0400_),
    .B(_0403_),
    .C(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__o211ai_1 _2751_ (.A1(_0403_),
    .A2(_0595_),
    .B1(_0655_),
    .C1(_0406_),
    .Y(_0656_));
 sky130_fd_sc_hd__o21ai_0 _2752_ (.A1(_0524_),
    .A2(_0532_),
    .B1(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__nand2_1 _2753_ (.A(_0408_),
    .B(_0657_),
    .Y(_0658_));
 sky130_fd_sc_hd__or3_1 _2754_ (.A(_0321_),
    .B(_0384_),
    .C(_0445_),
    .X(_0659_));
 sky130_fd_sc_hd__o21ai_0 _2755_ (.A1(_0404_),
    .A2(_0659_),
    .B1(_0446_),
    .Y(_0660_));
 sky130_fd_sc_hd__nand2_1 _2756_ (.A(_0295_),
    .B(_0602_),
    .Y(_0661_));
 sky130_fd_sc_hd__mux2i_2 _2757_ (.A0(\add_result[17] ),
    .A1(\add_result[18] ),
    .S(_0303_),
    .Y(_0662_));
 sky130_fd_sc_hd__mux2i_2 _2758_ (.A0(_0629_),
    .A1(_0662_),
    .S(_0298_),
    .Y(_0663_));
 sky130_fd_sc_hd__nand2_1 _2759_ (.A(_0478_),
    .B(_0663_),
    .Y(_0664_));
 sky130_fd_sc_hd__a21oi_1 _2760_ (.A1(_0661_),
    .A2(_0664_),
    .B1(_0424_),
    .Y(_0665_));
 sky130_fd_sc_hd__a31oi_1 _2761_ (.A1(_0418_),
    .A2(_0658_),
    .A3(_0660_),
    .B1(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__a2bb2oi_1 _2762_ (.A1_N(_0417_),
    .A2_N(_0666_),
    .B1(_0386_),
    .B2(\add_result[18] ),
    .Y(_0667_));
 sky130_fd_sc_hd__nand2_1 _2763_ (.A(\add_result[19] ),
    .B(_0560_),
    .Y(_0668_));
 sky130_fd_sc_hd__o21ai_0 _2764_ (.A1(_0340_),
    .A2(_0667_),
    .B1(_0668_),
    .Y(_0092_));
 sky130_fd_sc_hd__nand2_1 _2765_ (.A(_1695_),
    .B(_0610_),
    .Y(_0669_));
 sky130_fd_sc_hd__mux2i_1 _2766_ (.A0(\add_result[18] ),
    .A1(\add_result[19] ),
    .S(_0479_),
    .Y(_0670_));
 sky130_fd_sc_hd__mux2i_1 _2767_ (.A0(_0637_),
    .A1(_0670_),
    .S(_0299_),
    .Y(_0671_));
 sky130_fd_sc_hd__nand2_1 _2768_ (.A(_1698_),
    .B(_0671_),
    .Y(_0672_));
 sky130_fd_sc_hd__mux2i_1 _2769_ (.A0(\add_result[18] ),
    .A1(\add_result[19] ),
    .S(_0320_),
    .Y(_0673_));
 sky130_fd_sc_hd__nand2_1 _2770_ (.A(_0432_),
    .B(_0673_),
    .Y(_0674_));
 sky130_fd_sc_hd__o21ai_1 _2771_ (.A1(_0432_),
    .A2(_0640_),
    .B1(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__nor2_1 _2772_ (.A(_0449_),
    .B(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__a21oi_1 _2773_ (.A1(_0450_),
    .A2(_0613_),
    .B1(_0676_),
    .Y(_0677_));
 sky130_fd_sc_hd__nand2_1 _2774_ (.A(_0445_),
    .B(_0554_),
    .Y(_0678_));
 sky130_fd_sc_hd__o311ai_1 _2775_ (.A1(_0448_),
    .A2(_0445_),
    .A3(_0677_),
    .B1(_0678_),
    .C1(_0408_),
    .Y(_0679_));
 sky130_fd_sc_hd__o21ai_0 _2776_ (.A1(_0420_),
    .A2(_0659_),
    .B1(_0446_),
    .Y(_0680_));
 sky130_fd_sc_hd__a21oi_1 _2777_ (.A1(_0679_),
    .A2(_0680_),
    .B1(_0387_),
    .Y(_0681_));
 sky130_fd_sc_hd__a311oi_2 _2778_ (.A1(_0318_),
    .A2(_0669_),
    .A3(_0672_),
    .B1(_0681_),
    .C1(_0304_),
    .Y(_0682_));
 sky130_fd_sc_hd__a21oi_1 _2779_ (.A1(\add_result[19] ),
    .A2(_0386_),
    .B1(_0682_),
    .Y(_0683_));
 sky130_fd_sc_hd__nand2_1 _2780_ (.A(_0286_),
    .B(_0560_),
    .Y(_0684_));
 sky130_fd_sc_hd__o21ai_0 _2781_ (.A1(_0340_),
    .A2(_0683_),
    .B1(_0684_),
    .Y(_0093_));
 sky130_fd_sc_hd__and2_0 _2782_ (.A(_0445_),
    .B(_0569_),
    .X(_0685_));
 sky130_fd_sc_hd__mux2i_1 _2783_ (.A0(\add_result[19] ),
    .A1(_0286_),
    .S(_0320_),
    .Y(_0686_));
 sky130_fd_sc_hd__nand2_1 _2784_ (.A(_0432_),
    .B(_0686_),
    .Y(_0687_));
 sky130_fd_sc_hd__o311a_1 _2785_ (.A1(_0388_),
    .A2(_0651_),
    .A3(_0652_),
    .B1(_0687_),
    .C1(_0399_),
    .X(_0688_));
 sky130_fd_sc_hd__nor2_1 _2786_ (.A(_0403_),
    .B(_0624_),
    .Y(_0689_));
 sky130_fd_sc_hd__a211oi_1 _2787_ (.A1(_0403_),
    .A2(_0688_),
    .B1(_0689_),
    .C1(_0445_),
    .Y(_0690_));
 sky130_fd_sc_hd__o21ai_0 _2788_ (.A1(_0685_),
    .A2(_0690_),
    .B1(_0408_),
    .Y(_0691_));
 sky130_fd_sc_hd__o21ai_0 _2789_ (.A1(_0435_),
    .A2(_0659_),
    .B1(_0446_),
    .Y(_0692_));
 sky130_fd_sc_hd__nand2_1 _2790_ (.A(_0295_),
    .B(_0630_),
    .Y(_0693_));
 sky130_fd_sc_hd__mux2i_2 _2791_ (.A0(\add_result[19] ),
    .A1(_0286_),
    .S(_0479_),
    .Y(_0694_));
 sky130_fd_sc_hd__mux2i_2 _2792_ (.A0(_0662_),
    .A1(_0694_),
    .S(_0299_),
    .Y(_0695_));
 sky130_fd_sc_hd__nand2_1 _2793_ (.A(_0478_),
    .B(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__a21oi_1 _2794_ (.A1(_0693_),
    .A2(_0696_),
    .B1(_0424_),
    .Y(_0697_));
 sky130_fd_sc_hd__a31oi_1 _2795_ (.A1(_0418_),
    .A2(_0691_),
    .A3(_0692_),
    .B1(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__a2bb2oi_1 _2796_ (.A1_N(_0417_),
    .A2_N(_0698_),
    .B1(_0386_),
    .B2(_0286_),
    .Y(_0699_));
 sky130_fd_sc_hd__nand2_1 _2797_ (.A(_0287_),
    .B(_0560_),
    .Y(_0700_));
 sky130_fd_sc_hd__o21ai_0 _2798_ (.A1(_0340_),
    .A2(_0699_),
    .B1(_0700_),
    .Y(_0094_));
 sky130_fd_sc_hd__nor3_1 _2799_ (.A(_0321_),
    .B(_0384_),
    .C(_0445_),
    .Y(_0701_));
 sky130_fd_sc_hd__nand2_1 _2800_ (.A(_0455_),
    .B(_0701_),
    .Y(_0702_));
 sky130_fd_sc_hd__nand2_1 _2801_ (.A(_0446_),
    .B(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__mux2_1 _2802_ (.A0(_0286_),
    .A1(_0287_),
    .S(_0320_),
    .X(_0704_));
 sky130_fd_sc_hd__nor2_1 _2803_ (.A(_0389_),
    .B(_0673_),
    .Y(_0705_));
 sky130_fd_sc_hd__a21oi_1 _2804_ (.A1(_0389_),
    .A2(_0704_),
    .B1(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hd__nand2_1 _2805_ (.A(_0450_),
    .B(_0642_),
    .Y(_0707_));
 sky130_fd_sc_hd__o21ai_0 _2806_ (.A1(_0450_),
    .A2(_0706_),
    .B1(_0707_),
    .Y(_0708_));
 sky130_fd_sc_hd__nand3_1 _2807_ (.A(_0400_),
    .B(_0524_),
    .C(_0708_),
    .Y(_0709_));
 sky130_fd_sc_hd__o211ai_1 _2808_ (.A1(_0524_),
    .A2(_0580_),
    .B1(_0709_),
    .C1(_0408_),
    .Y(_0710_));
 sky130_fd_sc_hd__nand2_1 _2809_ (.A(_0295_),
    .B(_0638_),
    .Y(_0711_));
 sky130_fd_sc_hd__nand2_1 _2810_ (.A(_1702_),
    .B(_0670_),
    .Y(_0712_));
 sky130_fd_sc_hd__mux2i_1 _2811_ (.A0(_0286_),
    .A1(_0287_),
    .S(_1711_),
    .Y(_0713_));
 sky130_fd_sc_hd__nand2_1 _2812_ (.A(_1574_),
    .B(_0713_),
    .Y(_0714_));
 sky130_fd_sc_hd__nand3_1 _2813_ (.A(_0478_),
    .B(_0712_),
    .C(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__a21oi_1 _2814_ (.A1(_0711_),
    .A2(_0715_),
    .B1(_0424_),
    .Y(_0716_));
 sky130_fd_sc_hd__a31oi_1 _2815_ (.A1(_0424_),
    .A2(_0703_),
    .A3(_0710_),
    .B1(_0716_),
    .Y(_0717_));
 sky130_fd_sc_hd__nor2_1 _2816_ (.A(_0417_),
    .B(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__a211oi_1 _2817_ (.A1(_0287_),
    .A2(_0386_),
    .B1(_0718_),
    .C1(_0266_),
    .Y(_0719_));
 sky130_fd_sc_hd__a21oi_1 _2818_ (.A1(_0300_),
    .A2(_0415_),
    .B1(_0719_),
    .Y(_0095_));
 sky130_fd_sc_hd__mux2_1 _2819_ (.A0(_0287_),
    .A1(_0267_),
    .S(_0320_),
    .X(_0720_));
 sky130_fd_sc_hd__nor2_1 _2820_ (.A(_0451_),
    .B(_0686_),
    .Y(_0721_));
 sky130_fd_sc_hd__a21oi_1 _2821_ (.A1(_0389_),
    .A2(_0720_),
    .B1(_0721_),
    .Y(_0722_));
 sky130_fd_sc_hd__nand3_1 _2822_ (.A(_0400_),
    .B(_0450_),
    .C(_0654_),
    .Y(_0723_));
 sky130_fd_sc_hd__o311ai_0 _2823_ (.A1(_0448_),
    .A2(_0450_),
    .A3(_0722_),
    .B1(_0723_),
    .C1(_0406_),
    .Y(_0724_));
 sky130_fd_sc_hd__o21ai_0 _2824_ (.A1(_0524_),
    .A2(_0596_),
    .B1(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__nand2_1 _2825_ (.A(_0408_),
    .B(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__o21ai_0 _2826_ (.A1(_0472_),
    .A2(_0659_),
    .B1(_0446_),
    .Y(_0727_));
 sky130_fd_sc_hd__mux2_1 _2827_ (.A0(_0287_),
    .A1(_0267_),
    .S(_0479_),
    .X(_0728_));
 sky130_fd_sc_hd__nor2_1 _2828_ (.A(_1574_),
    .B(_0694_),
    .Y(_0729_));
 sky130_fd_sc_hd__a221oi_2 _2829_ (.A1(_0295_),
    .A2(_0663_),
    .B1(_0728_),
    .B2(_1574_),
    .C1(_0729_),
    .Y(_0730_));
 sky130_fd_sc_hd__nor2_1 _2830_ (.A(_0424_),
    .B(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__a31oi_1 _2831_ (.A1(_0418_),
    .A2(_0726_),
    .A3(_0727_),
    .B1(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__a2bb2oi_1 _2832_ (.A1_N(_0417_),
    .A2_N(_0732_),
    .B1(_0386_),
    .B2(_0267_),
    .Y(_0733_));
 sky130_fd_sc_hd__nand2_1 _2833_ (.A(_0269_),
    .B(_0523_),
    .Y(_0734_));
 sky130_fd_sc_hd__o21ai_0 _2834_ (.A1(_0340_),
    .A2(_0733_),
    .B1(_0734_),
    .Y(_0097_));
 sky130_fd_sc_hd__nand2_1 _2835_ (.A(_0445_),
    .B(_0616_),
    .Y(_0735_));
 sky130_fd_sc_hd__nand2_1 _2836_ (.A(_0269_),
    .B(_0320_),
    .Y(_0736_));
 sky130_fd_sc_hd__o211ai_1 _2837_ (.A1(_0300_),
    .A2(_0320_),
    .B1(_0736_),
    .C1(_0389_),
    .Y(_0737_));
 sky130_fd_sc_hd__o211ai_1 _2838_ (.A1(_0389_),
    .A2(_0704_),
    .B1(_0737_),
    .C1(_0403_),
    .Y(_0738_));
 sky130_fd_sc_hd__o21ai_0 _2839_ (.A1(_0403_),
    .A2(_0675_),
    .B1(_0738_),
    .Y(_0739_));
 sky130_fd_sc_hd__nand3_1 _2840_ (.A(_0400_),
    .B(_0524_),
    .C(_0739_),
    .Y(_0740_));
 sky130_fd_sc_hd__a21oi_1 _2841_ (.A1(_0487_),
    .A2(_0701_),
    .B1(_0411_),
    .Y(_0741_));
 sky130_fd_sc_hd__a31oi_1 _2842_ (.A1(_0408_),
    .A2(_0735_),
    .A3(_0740_),
    .B1(_0741_),
    .Y(_0742_));
 sky130_fd_sc_hd__nor2b_1 _2843_ (.A(_0268_),
    .B_N(_0287_),
    .Y(_0743_));
 sky130_fd_sc_hd__o21ai_0 _2844_ (.A1(_0296_),
    .A2(_0743_),
    .B1(_0269_),
    .Y(_0744_));
 sky130_fd_sc_hd__nor2b_1 _2845_ (.A(_0269_),
    .B_N(_0286_),
    .Y(_0745_));
 sky130_fd_sc_hd__o211ai_1 _2846_ (.A1(_0268_),
    .A2(_0745_),
    .B1(_0293_),
    .C1(_0267_),
    .Y(_0746_));
 sky130_fd_sc_hd__nand2_1 _2847_ (.A(_0295_),
    .B(_0671_),
    .Y(_0747_));
 sky130_fd_sc_hd__a31oi_1 _2848_ (.A1(_0744_),
    .A2(_0746_),
    .A3(_0747_),
    .B1(_0424_),
    .Y(_0748_));
 sky130_fd_sc_hd__a21oi_1 _2849_ (.A1(_0418_),
    .A2(_0742_),
    .B1(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__nor2_1 _2850_ (.A(_0417_),
    .B(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__a21oi_1 _2851_ (.A1(_0269_),
    .A2(_0386_),
    .B1(_0750_),
    .Y(_0751_));
 sky130_fd_sc_hd__nand2_1 _2852_ (.A(_0268_),
    .B(_0523_),
    .Y(_0752_));
 sky130_fd_sc_hd__o21ai_0 _2853_ (.A1(_0340_),
    .A2(_0751_),
    .B1(_0752_),
    .Y(_0098_));
 sky130_fd_sc_hd__mux2i_1 _2854_ (.A0(_0269_),
    .A1(_0268_),
    .S(_0320_),
    .Y(_0753_));
 sky130_fd_sc_hd__nand2_1 _2855_ (.A(_0389_),
    .B(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__o21ai_0 _2856_ (.A1(_0389_),
    .A2(_0720_),
    .B1(_0754_),
    .Y(_0755_));
 sky130_fd_sc_hd__nand2_1 _2857_ (.A(_0450_),
    .B(_0688_),
    .Y(_0756_));
 sky130_fd_sc_hd__o311ai_1 _2858_ (.A1(_0448_),
    .A2(_0450_),
    .A3(_0755_),
    .B1(_0756_),
    .C1(_0406_),
    .Y(_0757_));
 sky130_fd_sc_hd__o21ai_0 _2859_ (.A1(_0524_),
    .A2(_0625_),
    .B1(_0757_),
    .Y(_0758_));
 sky130_fd_sc_hd__a21oi_1 _2860_ (.A1(_0500_),
    .A2(_0701_),
    .B1(_0411_),
    .Y(_0759_));
 sky130_fd_sc_hd__a21oi_1 _2861_ (.A1(_0408_),
    .A2(_0758_),
    .B1(_0759_),
    .Y(_0760_));
 sky130_fd_sc_hd__a211oi_1 _2862_ (.A1(_0268_),
    .A2(_0421_),
    .B1(_0760_),
    .C1(_0318_),
    .Y(_0761_));
 sky130_fd_sc_hd__a211oi_1 _2863_ (.A1(_0268_),
    .A2(_0296_),
    .B1(_0743_),
    .C1(_0269_),
    .Y(_0762_));
 sky130_fd_sc_hd__a21oi_1 _2864_ (.A1(_0267_),
    .A2(_0293_),
    .B1(_0268_),
    .Y(_0763_));
 sky130_fd_sc_hd__o21ai_0 _2865_ (.A1(_0762_),
    .A2(_0763_),
    .B1(_0318_),
    .Y(_0764_));
 sky130_fd_sc_hd__a21oi_1 _2866_ (.A1(_1695_),
    .A2(_0695_),
    .B1(_0764_),
    .Y(_0765_));
 sky130_fd_sc_hd__o21ai_0 _2867_ (.A1(_0268_),
    .A2(_0340_),
    .B1(_0305_),
    .Y(_0766_));
 sky130_fd_sc_hd__o41ai_1 _2868_ (.A1(_0327_),
    .A2(_0308_),
    .A3(_0761_),
    .A4(_0765_),
    .B1(_0766_),
    .Y(_0099_));
 sky130_fd_sc_hd__nand4_4 _2869_ (.A(net22),
    .B(net21),
    .C(net25),
    .D(net23),
    .Y(_0767_));
 sky130_fd_sc_hd__nand4_2 _2870_ (.A(net18),
    .B(net17),
    .C(net20),
    .D(net19),
    .Y(_0768_));
 sky130_fd_sc_hd__nand4_1 _2871_ (.A(net54),
    .B(net53),
    .C(net57),
    .D(net55),
    .Y(_0769_));
 sky130_fd_sc_hd__nand2_1 _2872_ (.A(net50),
    .B(net49),
    .Y(_0770_));
 sky130_fd_sc_hd__or4_1 _2873_ (.A(_1606_),
    .B(_1612_),
    .C(_0769_),
    .D(_0770_),
    .X(_0771_));
 sky130_fd_sc_hd__clkbuf_2 _2874_ (.A(_0771_),
    .X(_0772_));
 sky130_fd_sc_hd__o21ai_4 _2875_ (.A1(_0767_),
    .A2(_0768_),
    .B1(_0772_),
    .Y(_0773_));
 sky130_fd_sc_hd__buf_2 _2876_ (.A(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__inv_1 _2877_ (.A(_1730_),
    .Y(_0775_));
 sky130_fd_sc_hd__a31oi_2 _2878_ (.A1(\aligned_a_mant[0] ),
    .A2(\aligned_b_mant[0] ),
    .A3(_0775_),
    .B1(_1734_),
    .Y(_0776_));
 sky130_fd_sc_hd__xnor2_4 _2879_ (.A(a_sign_stage1),
    .B(b_sign_stage1),
    .Y(_0777_));
 sky130_fd_sc_hd__buf_4 _2880_ (.A(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__buf_4 _2881_ (.A(_0778_),
    .X(_0779_));
 sky130_fd_sc_hd__clkbuf_4 _2882_ (.A(is_a_larger_stage1),
    .X(_0780_));
 sky130_fd_sc_hd__clkbuf_4 _2883_ (.A(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__clkbuf_4 _2884_ (.A(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__nand2b_1 _2885_ (.A_N(_1732_),
    .B(_0781_),
    .Y(_0783_));
 sky130_fd_sc_hd__o21ai_0 _2886_ (.A1(_1729_),
    .A2(_0782_),
    .B1(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__nand2b_1 _2887_ (.A_N(\aligned_b_mant[0] ),
    .B(\aligned_a_mant[0] ),
    .Y(_0785_));
 sky130_fd_sc_hd__nor3_1 _2888_ (.A(_1729_),
    .B(_0782_),
    .C(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__nand2b_1 _2889_ (.A_N(\aligned_a_mant[0] ),
    .B(\aligned_b_mant[0] ),
    .Y(_0787_));
 sky130_fd_sc_hd__nor2_1 _2890_ (.A(_0783_),
    .B(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__a2111oi_0 _2891_ (.A1(_0775_),
    .A2(_0784_),
    .B1(_0786_),
    .C1(_0788_),
    .D1(_0778_),
    .Y(_0789_));
 sky130_fd_sc_hd__a21oi_1 _2892_ (.A1(_0776_),
    .A2(_0779_),
    .B1(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__xor2_2 _2893_ (.A(_1722_),
    .B(_0790_),
    .X(_0791_));
 sky130_fd_sc_hd__nor2_1 _2894_ (.A(_0774_),
    .B(_0791_),
    .Y(_0017_));
 sky130_fd_sc_hd__clkbuf_4 _2895_ (.A(_0777_),
    .X(_0792_));
 sky130_fd_sc_hd__clkinv_4 _2896_ (.A(is_a_larger_stage1),
    .Y(_0793_));
 sky130_fd_sc_hd__a21o_1 _2897_ (.A1(_1730_),
    .A2(_0787_),
    .B1(_1732_),
    .X(_0794_));
 sky130_fd_sc_hd__a21o_1 _2898_ (.A1(_1722_),
    .A2(_0794_),
    .B1(_1724_),
    .X(_0795_));
 sky130_fd_sc_hd__nor2_1 _2899_ (.A(_0793_),
    .B(_0795_),
    .Y(_0796_));
 sky130_fd_sc_hd__buf_4 _2900_ (.A(_0782_),
    .X(_0797_));
 sky130_fd_sc_hd__a21o_1 _2901_ (.A1(_1730_),
    .A2(_0785_),
    .B1(_1729_),
    .X(_0798_));
 sky130_fd_sc_hd__a21o_1 _2902_ (.A1(_1722_),
    .A2(_0798_),
    .B1(_1721_),
    .X(_0799_));
 sky130_fd_sc_hd__nor2_1 _2903_ (.A(_0797_),
    .B(_0799_),
    .Y(_0800_));
 sky130_fd_sc_hd__nor2_1 _2904_ (.A(_0796_),
    .B(_0800_),
    .Y(_0801_));
 sky130_fd_sc_hd__o21bai_2 _2905_ (.A1(_1722_),
    .A2(_0776_),
    .B1_N(_1726_),
    .Y(_0802_));
 sky130_fd_sc_hd__nand2_1 _2906_ (.A(_0792_),
    .B(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__o21ai_1 _2907_ (.A1(_0792_),
    .A2(_0801_),
    .B1(_0803_),
    .Y(_0804_));
 sky130_fd_sc_hd__xor2_2 _2908_ (.A(_1738_),
    .B(_0804_),
    .X(_0805_));
 sky130_fd_sc_hd__nor2_1 _2909_ (.A(_0774_),
    .B(_0805_),
    .Y(_0018_));
 sky130_fd_sc_hd__clkbuf_2 _2910_ (.A(_1746_),
    .X(_0806_));
 sky130_fd_sc_hd__xor2_4 _2911_ (.A(a_sign_stage1),
    .B(b_sign_stage1),
    .X(_0807_));
 sky130_fd_sc_hd__buf_4 _2912_ (.A(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__nor2b_1 _2913_ (.A(_1738_),
    .B_N(_0802_),
    .Y(_0809_));
 sky130_fd_sc_hd__a21o_1 _2914_ (.A1(_1738_),
    .A2(_0799_),
    .B1(_1737_),
    .X(_0810_));
 sky130_fd_sc_hd__a21oi_2 _2915_ (.A1(_1738_),
    .A2(_0795_),
    .B1(_1740_),
    .Y(_0811_));
 sky130_fd_sc_hd__nand2_1 _2916_ (.A(_0797_),
    .B(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__o211ai_1 _2917_ (.A1(_0797_),
    .A2(_0810_),
    .B1(_0812_),
    .C1(_0808_),
    .Y(_0813_));
 sky130_fd_sc_hd__o31ai_1 _2918_ (.A1(_1742_),
    .A2(_0808_),
    .A3(_0809_),
    .B1(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__xnor2_1 _2919_ (.A(_0806_),
    .B(_0814_),
    .Y(_0815_));
 sky130_fd_sc_hd__nor2_1 _2920_ (.A(_0774_),
    .B(_0815_),
    .Y(_0019_));
 sky130_fd_sc_hd__buf_2 _2921_ (.A(_1754_),
    .X(_0816_));
 sky130_fd_sc_hd__inv_1 _2922_ (.A(_0806_),
    .Y(_0817_));
 sky130_fd_sc_hd__o21bai_1 _2923_ (.A1(_0817_),
    .A2(_0811_),
    .B1_N(_1748_),
    .Y(_0818_));
 sky130_fd_sc_hd__a21oi_1 _2924_ (.A1(_0806_),
    .A2(_0810_),
    .B1(_1745_),
    .Y(_0819_));
 sky130_fd_sc_hd__nor2_1 _2925_ (.A(_0797_),
    .B(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hd__a21oi_1 _2926_ (.A1(_0797_),
    .A2(_0818_),
    .B1(_0820_),
    .Y(_0821_));
 sky130_fd_sc_hd__nor2_1 _2927_ (.A(_1738_),
    .B(_0806_),
    .Y(_0822_));
 sky130_fd_sc_hd__a21o_1 _2928_ (.A1(_1742_),
    .A2(_0817_),
    .B1(_1750_),
    .X(_0823_));
 sky130_fd_sc_hd__a21oi_1 _2929_ (.A1(_0802_),
    .A2(_0822_),
    .B1(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__nand2_1 _2930_ (.A(_0779_),
    .B(_0824_),
    .Y(_0825_));
 sky130_fd_sc_hd__o21ai_1 _2931_ (.A1(_0792_),
    .A2(_0821_),
    .B1(_0825_),
    .Y(_0826_));
 sky130_fd_sc_hd__xnor2_1 _2932_ (.A(_0816_),
    .B(_0826_),
    .Y(_0827_));
 sky130_fd_sc_hd__nor2_1 _2933_ (.A(_0774_),
    .B(_0827_),
    .Y(_0020_));
 sky130_fd_sc_hd__buf_2 _2934_ (.A(_1762_),
    .X(_0828_));
 sky130_fd_sc_hd__nor2_1 _2935_ (.A(_0816_),
    .B(_0824_),
    .Y(_0829_));
 sky130_fd_sc_hd__nor2_1 _2936_ (.A(_1758_),
    .B(_0829_),
    .Y(_0830_));
 sky130_fd_sc_hd__clkbuf_4 _2937_ (.A(_0782_),
    .X(_0831_));
 sky130_fd_sc_hd__and3_1 _2938_ (.A(_1738_),
    .B(_0806_),
    .C(_0816_),
    .X(_0832_));
 sky130_fd_sc_hd__a21oi_1 _2939_ (.A1(_0806_),
    .A2(_1737_),
    .B1(_1745_),
    .Y(_0833_));
 sky130_fd_sc_hd__nor2b_1 _2940_ (.A(_0833_),
    .B_N(_0816_),
    .Y(_0834_));
 sky130_fd_sc_hd__a211o_1 _2941_ (.A1(_0799_),
    .A2(_0832_),
    .B1(_0834_),
    .C1(_1753_),
    .X(_0835_));
 sky130_fd_sc_hd__nor2_1 _2942_ (.A(_0831_),
    .B(_0835_),
    .Y(_0836_));
 sky130_fd_sc_hd__a211oi_1 _2943_ (.A1(_0816_),
    .A2(_0818_),
    .B1(_1756_),
    .C1(_0793_),
    .Y(_0837_));
 sky130_fd_sc_hd__nor3_1 _2944_ (.A(_0778_),
    .B(_0836_),
    .C(_0837_),
    .Y(_0838_));
 sky130_fd_sc_hd__a21oi_1 _2945_ (.A1(_0779_),
    .A2(_0830_),
    .B1(_0838_),
    .Y(_0839_));
 sky130_fd_sc_hd__xor2_1 _2946_ (.A(_0828_),
    .B(_0839_),
    .X(_0840_));
 sky130_fd_sc_hd__nor2_1 _2947_ (.A(_0774_),
    .B(_0840_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_1 _2948_ (.A(_1770_),
    .Y(_0841_));
 sky130_fd_sc_hd__inv_1 _2949_ (.A(_1766_),
    .Y(_0842_));
 sky130_fd_sc_hd__o21ai_0 _2950_ (.A1(_0828_),
    .A2(_0830_),
    .B1(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hd__nor2_1 _2951_ (.A(_0808_),
    .B(_0843_),
    .Y(_0844_));
 sky130_fd_sc_hd__nand3_1 _2952_ (.A(_0806_),
    .B(_0816_),
    .C(_0828_),
    .Y(_0845_));
 sky130_fd_sc_hd__nand3_1 _2953_ (.A(_0816_),
    .B(_1748_),
    .C(_0828_),
    .Y(_0846_));
 sky130_fd_sc_hd__nand2_1 _2954_ (.A(_0828_),
    .B(_1756_),
    .Y(_0847_));
 sky130_fd_sc_hd__and2_0 _2955_ (.A(_0846_),
    .B(_0847_),
    .X(_0848_));
 sky130_fd_sc_hd__inv_1 _2956_ (.A(_1764_),
    .Y(_0849_));
 sky130_fd_sc_hd__o2111a_1 _2957_ (.A1(_0811_),
    .A2(_0845_),
    .B1(_0848_),
    .C1(_0849_),
    .D1(_0780_),
    .X(_0850_));
 sky130_fd_sc_hd__a211oi_2 _2958_ (.A1(_0828_),
    .A2(_0835_),
    .B1(_1761_),
    .C1(_0780_),
    .Y(_0851_));
 sky130_fd_sc_hd__nor3_1 _2959_ (.A(_0778_),
    .B(_0850_),
    .C(_0851_),
    .Y(_0852_));
 sky130_fd_sc_hd__nor2_1 _2960_ (.A(_0844_),
    .B(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__xnor2_1 _2961_ (.A(_0841_),
    .B(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__nor2_1 _2962_ (.A(_0774_),
    .B(_0854_),
    .Y(_0022_));
 sky130_fd_sc_hd__clkbuf_4 _2963_ (.A(_1778_),
    .X(_0855_));
 sky130_fd_sc_hd__a21oi_1 _2964_ (.A1(_0841_),
    .A2(_0843_),
    .B1(_1774_),
    .Y(_0856_));
 sky130_fd_sc_hd__nand4_1 _2965_ (.A(_0806_),
    .B(_0816_),
    .C(_0828_),
    .D(_1770_),
    .Y(_0857_));
 sky130_fd_sc_hd__a31oi_1 _2966_ (.A1(_0849_),
    .A2(_0846_),
    .A3(_0847_),
    .B1(_0841_),
    .Y(_0858_));
 sky130_fd_sc_hd__nor2_1 _2967_ (.A(_1772_),
    .B(_0858_),
    .Y(_0859_));
 sky130_fd_sc_hd__o21ai_2 _2968_ (.A1(_0811_),
    .A2(_0857_),
    .B1(_0859_),
    .Y(_0860_));
 sky130_fd_sc_hd__a21oi_2 _2969_ (.A1(_0828_),
    .A2(_0835_),
    .B1(_1761_),
    .Y(_0861_));
 sky130_fd_sc_hd__nor2_1 _2970_ (.A(_0831_),
    .B(_1769_),
    .Y(_0862_));
 sky130_fd_sc_hd__o21ai_0 _2971_ (.A1(_0841_),
    .A2(_0861_),
    .B1(_0862_),
    .Y(_0863_));
 sky130_fd_sc_hd__o211ai_1 _2972_ (.A1(_0793_),
    .A2(_0860_),
    .B1(_0863_),
    .C1(_0808_),
    .Y(_0864_));
 sky130_fd_sc_hd__a21boi_0 _2973_ (.A1(_0792_),
    .A2(_0856_),
    .B1_N(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__xor2_1 _2974_ (.A(_0855_),
    .B(_0865_),
    .X(_0866_));
 sky130_fd_sc_hd__nor2_1 _2975_ (.A(_0774_),
    .B(_0866_),
    .Y(_0023_));
 sky130_fd_sc_hd__buf_2 _2976_ (.A(_1786_),
    .X(_0867_));
 sky130_fd_sc_hd__inv_1 _2977_ (.A(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__a21oi_2 _2978_ (.A1(_0855_),
    .A2(_0860_),
    .B1(_1780_),
    .Y(_0869_));
 sky130_fd_sc_hd__nand2_1 _2979_ (.A(_1770_),
    .B(_0855_),
    .Y(_0870_));
 sky130_fd_sc_hd__a21oi_2 _2980_ (.A1(_0855_),
    .A2(_1769_),
    .B1(_1777_),
    .Y(_0871_));
 sky130_fd_sc_hd__o21ai_0 _2981_ (.A1(_0861_),
    .A2(_0870_),
    .B1(_0871_),
    .Y(_0872_));
 sky130_fd_sc_hd__nor2_1 _2982_ (.A(_0797_),
    .B(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__a21oi_1 _2983_ (.A1(_0797_),
    .A2(_0869_),
    .B1(_0873_),
    .Y(_0874_));
 sky130_fd_sc_hd__nor4_1 _2984_ (.A(_1758_),
    .B(_1766_),
    .C(_1774_),
    .D(_1782_),
    .Y(_0875_));
 sky130_fd_sc_hd__a21oi_1 _2985_ (.A1(_0828_),
    .A2(_0842_),
    .B1(_1770_),
    .Y(_0876_));
 sky130_fd_sc_hd__nor3_1 _2986_ (.A(_1758_),
    .B(_1766_),
    .C(_1774_),
    .Y(_0877_));
 sky130_fd_sc_hd__a21oi_1 _2987_ (.A1(_0816_),
    .A2(_0877_),
    .B1(_0855_),
    .Y(_0878_));
 sky130_fd_sc_hd__o21ai_0 _2988_ (.A1(_1774_),
    .A2(_0876_),
    .B1(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__nor2b_1 _2989_ (.A(_1782_),
    .B_N(_0879_),
    .Y(_0880_));
 sky130_fd_sc_hd__a21oi_1 _2990_ (.A1(_0824_),
    .A2(_0875_),
    .B1(_0880_),
    .Y(_0881_));
 sky130_fd_sc_hd__nand2_1 _2991_ (.A(_0779_),
    .B(_0881_),
    .Y(_0882_));
 sky130_fd_sc_hd__o21ai_0 _2992_ (.A1(_0792_),
    .A2(_0874_),
    .B1(_0882_),
    .Y(_0883_));
 sky130_fd_sc_hd__xnor2_1 _2993_ (.A(_0868_),
    .B(_0883_),
    .Y(_0884_));
 sky130_fd_sc_hd__nor2_1 _2994_ (.A(_0774_),
    .B(_0884_),
    .Y(_0024_));
 sky130_fd_sc_hd__clkbuf_4 _2995_ (.A(_1794_),
    .X(_0885_));
 sky130_fd_sc_hd__a21oi_1 _2996_ (.A1(_0868_),
    .A2(_0881_),
    .B1(_1790_),
    .Y(_0886_));
 sky130_fd_sc_hd__a211oi_1 _2997_ (.A1(_0867_),
    .A2(_0872_),
    .B1(_1785_),
    .C1(_0831_),
    .Y(_0887_));
 sky130_fd_sc_hd__inv_1 _2998_ (.A(_1788_),
    .Y(_0888_));
 sky130_fd_sc_hd__o211a_1 _2999_ (.A1(_0868_),
    .A2(_0869_),
    .B1(_0888_),
    .C1(_0831_),
    .X(_0889_));
 sky130_fd_sc_hd__nor3_1 _3000_ (.A(_0778_),
    .B(_0887_),
    .C(_0889_),
    .Y(_0890_));
 sky130_fd_sc_hd__a21oi_1 _3001_ (.A1(_0779_),
    .A2(_0886_),
    .B1(_0890_),
    .Y(_0891_));
 sky130_fd_sc_hd__xor2_1 _3002_ (.A(_0885_),
    .B(_0891_),
    .X(_0892_));
 sky130_fd_sc_hd__nor2_1 _3003_ (.A(_0774_),
    .B(_0892_),
    .Y(_0000_));
 sky130_fd_sc_hd__buf_2 _3004_ (.A(_1802_),
    .X(_0893_));
 sky130_fd_sc_hd__nand4_2 _3005_ (.A(_1770_),
    .B(_0855_),
    .C(_0867_),
    .D(_0885_),
    .Y(_0894_));
 sky130_fd_sc_hd__o21bai_1 _3006_ (.A1(_0868_),
    .A2(_0871_),
    .B1_N(_1785_),
    .Y(_0895_));
 sky130_fd_sc_hd__a211o_1 _3007_ (.A1(_0885_),
    .A2(_0895_),
    .B1(_1793_),
    .C1(_0780_),
    .X(_0896_));
 sky130_fd_sc_hd__a21oi_1 _3008_ (.A1(_0855_),
    .A2(_1772_),
    .B1(_1780_),
    .Y(_0897_));
 sky130_fd_sc_hd__o21ai_0 _3009_ (.A1(_0868_),
    .A2(_0897_),
    .B1(_0888_),
    .Y(_0898_));
 sky130_fd_sc_hd__a211o_1 _3010_ (.A1(_0885_),
    .A2(_0898_),
    .B1(_1796_),
    .C1(_0793_),
    .X(_0899_));
 sky130_fd_sc_hd__nand2_1 _3011_ (.A(_0896_),
    .B(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__o31ai_4 _3012_ (.A1(_0850_),
    .A2(_0851_),
    .A3(_0894_),
    .B1(_0900_),
    .Y(_0901_));
 sky130_fd_sc_hd__nor2_1 _3013_ (.A(_0885_),
    .B(_0886_),
    .Y(_0902_));
 sky130_fd_sc_hd__o21ai_0 _3014_ (.A1(_1798_),
    .A2(_0902_),
    .B1(_0778_),
    .Y(_0903_));
 sky130_fd_sc_hd__o21ai_0 _3015_ (.A1(_0792_),
    .A2(_0901_),
    .B1(_0903_),
    .Y(_0904_));
 sky130_fd_sc_hd__xor2_1 _3016_ (.A(_0893_),
    .B(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__nor2_1 _3017_ (.A(_0774_),
    .B(_0905_),
    .Y(_0001_));
 sky130_fd_sc_hd__buf_2 _3018_ (.A(_0773_),
    .X(_0906_));
 sky130_fd_sc_hd__buf_2 _3019_ (.A(_1810_),
    .X(_0907_));
 sky130_fd_sc_hd__inv_1 _3020_ (.A(_1798_),
    .Y(_0908_));
 sky130_fd_sc_hd__nand2b_1 _3021_ (.A_N(_1794_),
    .B(_1790_),
    .Y(_0909_));
 sky130_fd_sc_hd__a21oi_1 _3022_ (.A1(_0908_),
    .A2(_0909_),
    .B1(_0893_),
    .Y(_0910_));
 sky130_fd_sc_hd__or3b_1 _3023_ (.A(_1806_),
    .B(_0910_),
    .C_N(_0875_),
    .X(_0911_));
 sky130_fd_sc_hd__a211oi_2 _3024_ (.A1(_0802_),
    .A2(_0822_),
    .B1(_0823_),
    .C1(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__nor2_1 _3025_ (.A(_1806_),
    .B(_0910_),
    .Y(_0913_));
 sky130_fd_sc_hd__or3_1 _3026_ (.A(_0867_),
    .B(_1794_),
    .C(_0893_),
    .X(_0914_));
 sky130_fd_sc_hd__nor3_1 _3027_ (.A(_1782_),
    .B(_1806_),
    .C(_0910_),
    .Y(_0915_));
 sky130_fd_sc_hd__a22o_1 _3028_ (.A1(_0913_),
    .A2(_0914_),
    .B1(_0915_),
    .B2(_0879_),
    .X(_0916_));
 sky130_fd_sc_hd__nor2_1 _3029_ (.A(_0912_),
    .B(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__a21o_1 _3030_ (.A1(_0893_),
    .A2(_1796_),
    .B1(_1804_),
    .X(_0918_));
 sky130_fd_sc_hd__nor3_1 _3031_ (.A(_0793_),
    .B(_1788_),
    .C(_0918_),
    .Y(_0919_));
 sky130_fd_sc_hd__nand2_1 _3032_ (.A(_0885_),
    .B(_0893_),
    .Y(_0920_));
 sky130_fd_sc_hd__a21o_1 _3033_ (.A1(_0893_),
    .A2(_1793_),
    .B1(_1801_),
    .X(_0921_));
 sky130_fd_sc_hd__mux2i_1 _3034_ (.A0(_0921_),
    .A1(_0918_),
    .S(is_a_larger_stage1),
    .Y(_0922_));
 sky130_fd_sc_hd__nor3_1 _3035_ (.A(is_a_larger_stage1),
    .B(_1785_),
    .C(_0921_),
    .Y(_0923_));
 sky130_fd_sc_hd__nor2_1 _3036_ (.A(_0923_),
    .B(_0919_),
    .Y(_0924_));
 sky130_fd_sc_hd__o2bb2ai_1 _3037_ (.A1_N(_0920_),
    .A2_N(_0922_),
    .B1(_0924_),
    .B2(_0867_),
    .Y(_0925_));
 sky130_fd_sc_hd__o211a_1 _3038_ (.A1(_0861_),
    .A2(_0870_),
    .B1(_0923_),
    .C1(_0871_),
    .X(_0926_));
 sky130_fd_sc_hd__a2111o_1 _3039_ (.A1(_0869_),
    .A2(_0919_),
    .B1(_0925_),
    .C1(_0926_),
    .D1(_0778_),
    .X(_0927_));
 sky130_fd_sc_hd__o21ai_0 _3040_ (.A1(_0808_),
    .A2(_0917_),
    .B1(_0927_),
    .Y(_0928_));
 sky130_fd_sc_hd__xnor2_1 _3041_ (.A(_0907_),
    .B(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__nor2_1 _3042_ (.A(_0906_),
    .B(_0929_),
    .Y(_0002_));
 sky130_fd_sc_hd__buf_2 _3043_ (.A(_1818_),
    .X(_0930_));
 sky130_fd_sc_hd__inv_1 _3044_ (.A(_0930_),
    .Y(_0931_));
 sky130_fd_sc_hd__inv_1 _3045_ (.A(_0907_),
    .Y(_0932_));
 sky130_fd_sc_hd__a21oi_1 _3046_ (.A1(_0932_),
    .A2(_0917_),
    .B1(_1814_),
    .Y(_0933_));
 sky130_fd_sc_hd__o21bai_2 _3047_ (.A1(_0861_),
    .A2(_0894_),
    .B1_N(_0896_),
    .Y(_0934_));
 sky130_fd_sc_hd__nand3_1 _3048_ (.A(_0867_),
    .B(_1780_),
    .C(_0885_),
    .Y(_0935_));
 sky130_fd_sc_hd__nand2_1 _3049_ (.A(_0780_),
    .B(_0935_),
    .Y(_0936_));
 sky130_fd_sc_hd__a41o_1 _3050_ (.A1(_0855_),
    .A2(_0867_),
    .A3(_0885_),
    .A4(_0860_),
    .B1(_0936_),
    .X(_0937_));
 sky130_fd_sc_hd__nand4_1 _3051_ (.A(_0893_),
    .B(_0907_),
    .C(_0934_),
    .D(_0937_),
    .Y(_0938_));
 sky130_fd_sc_hd__a21o_1 _3052_ (.A1(_0885_),
    .A2(_1788_),
    .B1(_1796_),
    .X(_0939_));
 sky130_fd_sc_hd__a21oi_1 _3053_ (.A1(_0893_),
    .A2(_0939_),
    .B1(_1804_),
    .Y(_0940_));
 sky130_fd_sc_hd__o21bai_1 _3054_ (.A1(_0932_),
    .A2(_0940_),
    .B1_N(_1812_),
    .Y(_0941_));
 sky130_fd_sc_hd__a21oi_1 _3055_ (.A1(_0907_),
    .A2(_1801_),
    .B1(_1809_),
    .Y(_0942_));
 sky130_fd_sc_hd__nor2_1 _3056_ (.A(_0780_),
    .B(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__a21oi_1 _3057_ (.A1(_0780_),
    .A2(_0941_),
    .B1(_0943_),
    .Y(_0944_));
 sky130_fd_sc_hd__a21oi_1 _3058_ (.A1(_0938_),
    .A2(_0944_),
    .B1(_0792_),
    .Y(_0945_));
 sky130_fd_sc_hd__a21oi_1 _3059_ (.A1(_0779_),
    .A2(_0933_),
    .B1(_0945_),
    .Y(_0946_));
 sky130_fd_sc_hd__xnor2_1 _3060_ (.A(_0931_),
    .B(_0946_),
    .Y(_0947_));
 sky130_fd_sc_hd__nor2_1 _3061_ (.A(_0906_),
    .B(_0947_),
    .Y(_0003_));
 sky130_fd_sc_hd__buf_2 _3062_ (.A(_1826_),
    .X(_0948_));
 sky130_fd_sc_hd__nor2_1 _3063_ (.A(_0930_),
    .B(_0933_),
    .Y(_0949_));
 sky130_fd_sc_hd__a21oi_1 _3064_ (.A1(_0907_),
    .A2(_0918_),
    .B1(_1812_),
    .Y(_0950_));
 sky130_fd_sc_hd__nand2_1 _3065_ (.A(_0893_),
    .B(_0907_),
    .Y(_0951_));
 sky130_fd_sc_hd__nand2_1 _3066_ (.A(_0885_),
    .B(_0930_),
    .Y(_0952_));
 sky130_fd_sc_hd__nor2_1 _3067_ (.A(_0951_),
    .B(_0952_),
    .Y(_0953_));
 sky130_fd_sc_hd__a211oi_1 _3068_ (.A1(_1788_),
    .A2(_0953_),
    .B1(_1820_),
    .C1(_0793_),
    .Y(_0954_));
 sky130_fd_sc_hd__o21ai_1 _3069_ (.A1(_0931_),
    .A2(_0950_),
    .B1(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__a211oi_2 _3070_ (.A1(_0855_),
    .A2(_0860_),
    .B1(_0955_),
    .C1(_1780_),
    .Y(_0956_));
 sky130_fd_sc_hd__a21oi_1 _3071_ (.A1(_0907_),
    .A2(_0921_),
    .B1(_1809_),
    .Y(_0957_));
 sky130_fd_sc_hd__a211oi_1 _3072_ (.A1(_1785_),
    .A2(_0953_),
    .B1(_1817_),
    .C1(_0780_),
    .Y(_0958_));
 sky130_fd_sc_hd__o21ai_1 _3073_ (.A1(_0931_),
    .A2(_0957_),
    .B1(_0958_),
    .Y(_0959_));
 sky130_fd_sc_hd__inv_1 _3074_ (.A(_0959_),
    .Y(_0960_));
 sky130_fd_sc_hd__o211a_1 _3075_ (.A1(_0861_),
    .A2(_0870_),
    .B1(_0960_),
    .C1(_0871_),
    .X(_0961_));
 sky130_fd_sc_hd__a22oi_2 _3076_ (.A1(_0867_),
    .A2(_0953_),
    .B1(_0955_),
    .B2(_0959_),
    .Y(_0962_));
 sky130_fd_sc_hd__or4_1 _3077_ (.A(_0777_),
    .B(_0956_),
    .C(_0961_),
    .D(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__o31ai_1 _3078_ (.A1(_1822_),
    .A2(_0808_),
    .A3(_0949_),
    .B1(_0963_),
    .Y(_0964_));
 sky130_fd_sc_hd__xnor2_1 _3079_ (.A(_0948_),
    .B(_0964_),
    .Y(_0965_));
 sky130_fd_sc_hd__nor2_1 _3080_ (.A(_0906_),
    .B(_0965_),
    .Y(_0004_));
 sky130_fd_sc_hd__buf_2 _3081_ (.A(_1834_),
    .X(_0966_));
 sky130_fd_sc_hd__or3_1 _3082_ (.A(_0907_),
    .B(_0930_),
    .C(_0948_),
    .X(_0967_));
 sky130_fd_sc_hd__nor2b_1 _3083_ (.A(_0930_),
    .B_N(_1814_),
    .Y(_0968_));
 sky130_fd_sc_hd__o21bai_1 _3084_ (.A1(_1822_),
    .A2(_0968_),
    .B1_N(_0948_),
    .Y(_0969_));
 sky130_fd_sc_hd__o31ai_1 _3085_ (.A1(_0912_),
    .A2(_0916_),
    .A3(_0967_),
    .B1(_0969_),
    .Y(_0970_));
 sky130_fd_sc_hd__nor2_1 _3086_ (.A(_1830_),
    .B(_0970_),
    .Y(_0971_));
 sky130_fd_sc_hd__nand2_1 _3087_ (.A(_0930_),
    .B(_0948_),
    .Y(_0972_));
 sky130_fd_sc_hd__a21oi_1 _3088_ (.A1(_0907_),
    .A2(_1804_),
    .B1(_1812_),
    .Y(_0973_));
 sky130_fd_sc_hd__a21oi_1 _3089_ (.A1(_0948_),
    .A2(_1820_),
    .B1(_1828_),
    .Y(_0974_));
 sky130_fd_sc_hd__o211ai_2 _3090_ (.A1(_0972_),
    .A2(_0973_),
    .B1(_0781_),
    .C1(_0974_),
    .Y(_0975_));
 sky130_fd_sc_hd__a21oi_1 _3091_ (.A1(_0948_),
    .A2(_1817_),
    .B1(_1825_),
    .Y(_0976_));
 sky130_fd_sc_hd__o211ai_2 _3092_ (.A1(_0942_),
    .A2(_0972_),
    .B1(_0976_),
    .C1(_0793_),
    .Y(_0977_));
 sky130_fd_sc_hd__nor2_1 _3093_ (.A(_0951_),
    .B(_0972_),
    .Y(_0978_));
 sky130_fd_sc_hd__a22oi_4 _3094_ (.A1(_0975_),
    .A2(_0977_),
    .B1(_0978_),
    .B2(_0901_),
    .Y(_0979_));
 sky130_fd_sc_hd__nor2_1 _3095_ (.A(_0778_),
    .B(_0979_),
    .Y(_0980_));
 sky130_fd_sc_hd__a21oi_1 _3096_ (.A1(_0779_),
    .A2(_0971_),
    .B1(_0980_),
    .Y(_0981_));
 sky130_fd_sc_hd__xor2_1 _3097_ (.A(_0966_),
    .B(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__nor2_1 _3098_ (.A(_0906_),
    .B(_0982_),
    .Y(_0005_));
 sky130_fd_sc_hd__buf_2 _3099_ (.A(_1842_),
    .X(_0983_));
 sky130_fd_sc_hd__nand2_1 _3100_ (.A(_0948_),
    .B(_0966_),
    .Y(_0984_));
 sky130_fd_sc_hd__a21oi_1 _3101_ (.A1(_0930_),
    .A2(_1809_),
    .B1(_1817_),
    .Y(_0985_));
 sky130_fd_sc_hd__a21oi_1 _3102_ (.A1(_0966_),
    .A2(_1825_),
    .B1(_1833_),
    .Y(_0986_));
 sky130_fd_sc_hd__o21ai_0 _3103_ (.A1(_0984_),
    .A2(_0985_),
    .B1(_0986_),
    .Y(_0987_));
 sky130_fd_sc_hd__a21oi_1 _3104_ (.A1(_0930_),
    .A2(_1812_),
    .B1(_1820_),
    .Y(_0988_));
 sky130_fd_sc_hd__a21oi_1 _3105_ (.A1(_0966_),
    .A2(_1828_),
    .B1(_1836_),
    .Y(_0989_));
 sky130_fd_sc_hd__o211ai_1 _3106_ (.A1(_0984_),
    .A2(_0988_),
    .B1(_0781_),
    .C1(_0989_),
    .Y(_0990_));
 sky130_fd_sc_hd__o21ai_1 _3107_ (.A1(_0781_),
    .A2(_0987_),
    .B1(_0990_),
    .Y(_0991_));
 sky130_fd_sc_hd__nand4_1 _3108_ (.A(_0907_),
    .B(_0930_),
    .C(_0948_),
    .D(_0966_),
    .Y(_0992_));
 sky130_fd_sc_hd__a2111o_1 _3109_ (.A1(_0869_),
    .A2(_0919_),
    .B1(_0925_),
    .C1(_0992_),
    .D1(_0926_),
    .X(_0993_));
 sky130_fd_sc_hd__a21oi_1 _3110_ (.A1(_0991_),
    .A2(_0993_),
    .B1(_0792_),
    .Y(_0994_));
 sky130_fd_sc_hd__nor2_1 _3111_ (.A(_0966_),
    .B(_0971_),
    .Y(_0995_));
 sky130_fd_sc_hd__nor3_1 _3112_ (.A(_1838_),
    .B(_0808_),
    .C(_0995_),
    .Y(_0996_));
 sky130_fd_sc_hd__nor3_1 _3113_ (.A(_0983_),
    .B(_0994_),
    .C(_0996_),
    .Y(_0997_));
 sky130_fd_sc_hd__o21a_1 _3114_ (.A1(_0994_),
    .A2(_0996_),
    .B1(_0983_),
    .X(_0998_));
 sky130_fd_sc_hd__nor3_1 _3115_ (.A(_0773_),
    .B(_0997_),
    .C(_0998_),
    .Y(_0006_));
 sky130_fd_sc_hd__buf_2 _3116_ (.A(_1850_),
    .X(_0999_));
 sky130_fd_sc_hd__or3_1 _3117_ (.A(_1830_),
    .B(_1838_),
    .C(_1846_),
    .X(_1000_));
 sky130_fd_sc_hd__inv_1 _3118_ (.A(_1838_),
    .Y(_1001_));
 sky130_fd_sc_hd__a21oi_1 _3119_ (.A1(_0966_),
    .A2(_1001_),
    .B1(_0983_),
    .Y(_1002_));
 sky130_fd_sc_hd__o22a_2 _3120_ (.A1(_0970_),
    .A2(_1000_),
    .B1(_1002_),
    .B2(_1846_),
    .X(_1003_));
 sky130_fd_sc_hd__nand4_1 _3121_ (.A(_0930_),
    .B(_0948_),
    .C(_0966_),
    .D(_0983_),
    .Y(_1004_));
 sky130_fd_sc_hd__nor2_1 _3122_ (.A(_0951_),
    .B(_1004_),
    .Y(_1005_));
 sky130_fd_sc_hd__nand2_1 _3123_ (.A(_0966_),
    .B(_0983_),
    .Y(_1006_));
 sky130_fd_sc_hd__a21oi_1 _3124_ (.A1(_0983_),
    .A2(_1833_),
    .B1(_1841_),
    .Y(_1007_));
 sky130_fd_sc_hd__o21ai_0 _3125_ (.A1(_0976_),
    .A2(_1006_),
    .B1(_1007_),
    .Y(_1008_));
 sky130_fd_sc_hd__a21oi_1 _3126_ (.A1(_0983_),
    .A2(_1836_),
    .B1(_1844_),
    .Y(_1009_));
 sky130_fd_sc_hd__o211ai_1 _3127_ (.A1(_0974_),
    .A2(_1006_),
    .B1(_1009_),
    .C1(_0780_),
    .Y(_1010_));
 sky130_fd_sc_hd__o21ai_0 _3128_ (.A1(_0780_),
    .A2(_1008_),
    .B1(_1010_),
    .Y(_1011_));
 sky130_fd_sc_hd__o21ai_1 _3129_ (.A1(_0944_),
    .A2(_1004_),
    .B1(_1011_),
    .Y(_1012_));
 sky130_fd_sc_hd__a31oi_4 _3130_ (.A1(_0934_),
    .A2(_0937_),
    .A3(_1005_),
    .B1(_1012_),
    .Y(_1013_));
 sky130_fd_sc_hd__mux2i_1 _3131_ (.A0(_1003_),
    .A1(_1013_),
    .S(_0808_),
    .Y(_1014_));
 sky130_fd_sc_hd__xnor2_1 _3132_ (.A(_0999_),
    .B(_1014_),
    .Y(_1015_));
 sky130_fd_sc_hd__nor2_1 _3133_ (.A(_0906_),
    .B(_1015_),
    .Y(_0007_));
 sky130_fd_sc_hd__buf_2 _3134_ (.A(_1858_),
    .X(_1016_));
 sky130_fd_sc_hd__inv_1 _3135_ (.A(_1016_),
    .Y(_1017_));
 sky130_fd_sc_hd__nand4_1 _3136_ (.A(_0948_),
    .B(_0966_),
    .C(_0983_),
    .D(_0999_),
    .Y(_1018_));
 sky130_fd_sc_hd__nand2_1 _3137_ (.A(_0983_),
    .B(_0999_),
    .Y(_1019_));
 sky130_fd_sc_hd__a21oi_1 _3138_ (.A1(_1850_),
    .A2(_1841_),
    .B1(_1849_),
    .Y(_1020_));
 sky130_fd_sc_hd__o21ai_0 _3139_ (.A1(_0986_),
    .A2(_1019_),
    .B1(_1020_),
    .Y(_1021_));
 sky130_fd_sc_hd__a21oi_1 _3140_ (.A1(_0999_),
    .A2(_1844_),
    .B1(_1852_),
    .Y(_1022_));
 sky130_fd_sc_hd__o211ai_1 _3141_ (.A1(_0989_),
    .A2(_1019_),
    .B1(_1022_),
    .C1(_0782_),
    .Y(_1023_));
 sky130_fd_sc_hd__o21ai_1 _3142_ (.A1(_0782_),
    .A2(_1021_),
    .B1(_1023_),
    .Y(_1024_));
 sky130_fd_sc_hd__o41ai_4 _3143_ (.A1(_0956_),
    .A2(_0961_),
    .A3(_0962_),
    .A4(_1018_),
    .B1(_1024_),
    .Y(_1025_));
 sky130_fd_sc_hd__inv_1 _3144_ (.A(_0999_),
    .Y(_1026_));
 sky130_fd_sc_hd__a21oi_1 _3145_ (.A1(_1026_),
    .A2(_1003_),
    .B1(_1854_),
    .Y(_1027_));
 sky130_fd_sc_hd__mux2i_1 _3146_ (.A0(_1025_),
    .A1(_1027_),
    .S(_0792_),
    .Y(_1028_));
 sky130_fd_sc_hd__xnor2_1 _3147_ (.A(_1017_),
    .B(_1028_),
    .Y(_1029_));
 sky130_fd_sc_hd__nor2_1 _3148_ (.A(_0906_),
    .B(_1029_),
    .Y(_0008_));
 sky130_fd_sc_hd__buf_2 _3149_ (.A(_1866_),
    .X(_1030_));
 sky130_fd_sc_hd__o21bai_1 _3150_ (.A1(_1026_),
    .A2(_1009_),
    .B1_N(_1852_),
    .Y(_1031_));
 sky130_fd_sc_hd__a21oi_1 _3151_ (.A1(_1016_),
    .A2(_1031_),
    .B1(_1860_),
    .Y(_1032_));
 sky130_fd_sc_hd__nor2b_1 _3152_ (.A(_1007_),
    .B_N(_0999_),
    .Y(_1033_));
 sky130_fd_sc_hd__o21ai_0 _3153_ (.A1(_1849_),
    .A2(_1033_),
    .B1(_1016_),
    .Y(_1034_));
 sky130_fd_sc_hd__nand2b_1 _3154_ (.A_N(_1857_),
    .B(_1034_),
    .Y(_1035_));
 sky130_fd_sc_hd__nor2_1 _3155_ (.A(_0831_),
    .B(_1035_),
    .Y(_1036_));
 sky130_fd_sc_hd__a211oi_1 _3156_ (.A1(_0831_),
    .A2(_1032_),
    .B1(_1036_),
    .C1(_0777_),
    .Y(_1037_));
 sky130_fd_sc_hd__inv_1 _3157_ (.A(_1854_),
    .Y(_1038_));
 sky130_fd_sc_hd__a21oi_1 _3158_ (.A1(_0999_),
    .A2(_1038_),
    .B1(_1016_),
    .Y(_1039_));
 sky130_fd_sc_hd__nor3_1 _3159_ (.A(_1862_),
    .B(_0807_),
    .C(_1039_),
    .Y(_1040_));
 sky130_fd_sc_hd__nand3_1 _3160_ (.A(_0999_),
    .B(_1016_),
    .C(_0807_),
    .Y(_1041_));
 sky130_fd_sc_hd__nor3_1 _3161_ (.A(_0979_),
    .B(_1006_),
    .C(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__nor4_1 _3162_ (.A(_1854_),
    .B(_1862_),
    .C(_0807_),
    .D(_1003_),
    .Y(_1043_));
 sky130_fd_sc_hd__nor4_1 _3163_ (.A(_1037_),
    .B(_1040_),
    .C(_1042_),
    .D(_1043_),
    .Y(_1044_));
 sky130_fd_sc_hd__xor2_1 _3164_ (.A(_1030_),
    .B(_1044_),
    .X(_1045_));
 sky130_fd_sc_hd__nor2_1 _3165_ (.A(_0906_),
    .B(_1045_),
    .Y(_0009_));
 sky130_fd_sc_hd__clkinvlp_4 _3166_ (.A(_1874_),
    .Y(_1046_));
 sky130_fd_sc_hd__nand2_1 _3167_ (.A(_1016_),
    .B(_1030_),
    .Y(_1047_));
 sky130_fd_sc_hd__a2111oi_2 _3168_ (.A1(_0991_),
    .A2(_0993_),
    .B1(_1019_),
    .C1(_1047_),
    .D1(_0777_),
    .Y(_1048_));
 sky130_fd_sc_hd__a21oi_1 _3169_ (.A1(_1030_),
    .A2(_1860_),
    .B1(_1868_),
    .Y(_1049_));
 sky130_fd_sc_hd__o21ai_1 _3170_ (.A1(_1022_),
    .A2(_1047_),
    .B1(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__nor2_1 _3171_ (.A(_0793_),
    .B(_1050_),
    .Y(_1051_));
 sky130_fd_sc_hd__o21bai_1 _3172_ (.A1(_1017_),
    .A2(_1020_),
    .B1_N(_1857_),
    .Y(_1052_));
 sky130_fd_sc_hd__a21o_1 _3173_ (.A1(_1030_),
    .A2(_1052_),
    .B1(_1865_),
    .X(_1053_));
 sky130_fd_sc_hd__nor2_1 _3174_ (.A(_0831_),
    .B(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__o21ai_0 _3175_ (.A1(_1051_),
    .A2(_1054_),
    .B1(_0808_),
    .Y(_1055_));
 sky130_fd_sc_hd__nor3_1 _3176_ (.A(_0999_),
    .B(_1016_),
    .C(_1866_),
    .Y(_1056_));
 sky130_fd_sc_hd__a21oi_1 _3177_ (.A1(_1854_),
    .A2(_1017_),
    .B1(_1862_),
    .Y(_1057_));
 sky130_fd_sc_hd__nor2_1 _3178_ (.A(_1866_),
    .B(_1057_),
    .Y(_1058_));
 sky130_fd_sc_hd__a211o_1 _3179_ (.A1(_1003_),
    .A2(_1056_),
    .B1(_1058_),
    .C1(_1870_),
    .X(_1059_));
 sky130_fd_sc_hd__nand2_1 _3180_ (.A(_0792_),
    .B(_1059_),
    .Y(_1060_));
 sky130_fd_sc_hd__o21ai_0 _3181_ (.A1(_1048_),
    .A2(_1055_),
    .B1(_1060_),
    .Y(_1061_));
 sky130_fd_sc_hd__xnor2_1 _3182_ (.A(_1046_),
    .B(_1061_),
    .Y(_1062_));
 sky130_fd_sc_hd__nor2_1 _3183_ (.A(_0906_),
    .B(_1062_),
    .Y(_0010_));
 sky130_fd_sc_hd__buf_2 _3184_ (.A(_1882_),
    .X(_1063_));
 sky130_fd_sc_hd__a21o_1 _3185_ (.A1(_1016_),
    .A2(_1852_),
    .B1(_1860_),
    .X(_1064_));
 sky130_fd_sc_hd__a21oi_1 _3186_ (.A1(_1030_),
    .A2(_1064_),
    .B1(_1868_),
    .Y(_1065_));
 sky130_fd_sc_hd__nor2_1 _3187_ (.A(_1046_),
    .B(_1065_),
    .Y(_1066_));
 sky130_fd_sc_hd__nor2_1 _3188_ (.A(_1876_),
    .B(_1066_),
    .Y(_1067_));
 sky130_fd_sc_hd__a21o_1 _3189_ (.A1(_1016_),
    .A2(_1849_),
    .B1(_1857_),
    .X(_1068_));
 sky130_fd_sc_hd__a21oi_1 _3190_ (.A1(_1030_),
    .A2(_1068_),
    .B1(_1865_),
    .Y(_1069_));
 sky130_fd_sc_hd__nor2_1 _3191_ (.A(_1046_),
    .B(_1069_),
    .Y(_1070_));
 sky130_fd_sc_hd__nor3_1 _3192_ (.A(_0781_),
    .B(_1873_),
    .C(_1070_),
    .Y(_1071_));
 sky130_fd_sc_hd__a21oi_1 _3193_ (.A1(_0781_),
    .A2(_1067_),
    .B1(_1071_),
    .Y(_1072_));
 sky130_fd_sc_hd__nand4_1 _3194_ (.A(_0999_),
    .B(_1016_),
    .C(_1030_),
    .D(_1874_),
    .Y(_1073_));
 sky130_fd_sc_hd__nor2_1 _3195_ (.A(_1013_),
    .B(_1073_),
    .Y(_1074_));
 sky130_fd_sc_hd__nor2_1 _3196_ (.A(_1046_),
    .B(_1878_),
    .Y(_1075_));
 sky130_fd_sc_hd__a2111oi_4 _3197_ (.A1(_1003_),
    .A2(_1056_),
    .B1(_1058_),
    .C1(_1870_),
    .D1(_1878_),
    .Y(_1076_));
 sky130_fd_sc_hd__or3_1 _3198_ (.A(_0807_),
    .B(_1075_),
    .C(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__o31ai_1 _3199_ (.A1(_0778_),
    .A2(_1072_),
    .A3(_1074_),
    .B1(_1077_),
    .Y(_1078_));
 sky130_fd_sc_hd__xor2_1 _3200_ (.A(_1063_),
    .B(_1078_),
    .X(_1079_));
 sky130_fd_sc_hd__nor2_1 _3201_ (.A(_0906_),
    .B(_1079_),
    .Y(_0011_));
 sky130_fd_sc_hd__buf_2 _3202_ (.A(_1890_),
    .X(_1080_));
 sky130_fd_sc_hd__inv_1 _3203_ (.A(_1886_),
    .Y(_1081_));
 sky130_fd_sc_hd__o31ai_1 _3204_ (.A1(_1063_),
    .A2(_1075_),
    .A3(_1076_),
    .B1(_1081_),
    .Y(_1082_));
 sky130_fd_sc_hd__nand2_1 _3205_ (.A(_1874_),
    .B(_1063_),
    .Y(_1083_));
 sky130_fd_sc_hd__nor2_1 _3206_ (.A(_1047_),
    .B(_1083_),
    .Y(_1084_));
 sky130_fd_sc_hd__o21bai_1 _3207_ (.A1(_1046_),
    .A2(_1049_),
    .B1_N(_1876_),
    .Y(_1085_));
 sky130_fd_sc_hd__a21oi_1 _3208_ (.A1(_1063_),
    .A2(_1085_),
    .B1(_1884_),
    .Y(_1086_));
 sky130_fd_sc_hd__nor2_1 _3209_ (.A(_0793_),
    .B(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__a21oi_1 _3210_ (.A1(_1030_),
    .A2(_1857_),
    .B1(_1865_),
    .Y(_1088_));
 sky130_fd_sc_hd__o21bai_1 _3211_ (.A1(_1046_),
    .A2(_1088_),
    .B1_N(_1873_),
    .Y(_1089_));
 sky130_fd_sc_hd__a21oi_1 _3212_ (.A1(_1063_),
    .A2(_1089_),
    .B1(_1881_),
    .Y(_1090_));
 sky130_fd_sc_hd__nor2_1 _3213_ (.A(_0831_),
    .B(_1090_),
    .Y(_1091_));
 sky130_fd_sc_hd__a2111oi_0 _3214_ (.A1(_1025_),
    .A2(_1084_),
    .B1(_1087_),
    .C1(_1091_),
    .D1(_0778_),
    .Y(_1092_));
 sky130_fd_sc_hd__a21oi_1 _3215_ (.A1(_0779_),
    .A2(_1082_),
    .B1(_1092_),
    .Y(_1093_));
 sky130_fd_sc_hd__xnor2_1 _3216_ (.A(_1080_),
    .B(_1093_),
    .Y(_1094_));
 sky130_fd_sc_hd__nor2_1 _3217_ (.A(_0906_),
    .B(_1094_),
    .Y(_0012_));
 sky130_fd_sc_hd__clkbuf_2 _3218_ (.A(_1898_),
    .X(_1095_));
 sky130_fd_sc_hd__inv_1 _3219_ (.A(_1080_),
    .Y(_1096_));
 sky130_fd_sc_hd__a21oi_1 _3220_ (.A1(_1886_),
    .A2(_1096_),
    .B1(_1894_),
    .Y(_1097_));
 sky130_fd_sc_hd__o41ai_4 _3221_ (.A1(_1882_),
    .A2(_1080_),
    .A3(_1075_),
    .A4(_1076_),
    .B1(_1097_),
    .Y(_1098_));
 sky130_fd_sc_hd__inv_1 _3222_ (.A(_1073_),
    .Y(_1099_));
 sky130_fd_sc_hd__nand3_1 _3223_ (.A(_1063_),
    .B(_1080_),
    .C(_1099_),
    .Y(_1100_));
 sky130_fd_sc_hd__or3_1 _3224_ (.A(_0979_),
    .B(_1006_),
    .C(_1100_),
    .X(_1101_));
 sky130_fd_sc_hd__a21oi_1 _3225_ (.A1(_1080_),
    .A2(_1884_),
    .B1(_1892_),
    .Y(_1102_));
 sky130_fd_sc_hd__a21o_1 _3226_ (.A1(_1080_),
    .A2(_1881_),
    .B1(_1889_),
    .X(_1103_));
 sky130_fd_sc_hd__nor2_1 _3227_ (.A(_0781_),
    .B(_1103_),
    .Y(_1104_));
 sky130_fd_sc_hd__a21oi_1 _3228_ (.A1(_0782_),
    .A2(_1102_),
    .B1(_1104_),
    .Y(_1105_));
 sky130_fd_sc_hd__a211oi_1 _3229_ (.A1(_1874_),
    .A2(_1868_),
    .B1(_1876_),
    .C1(_1892_),
    .Y(_1106_));
 sky130_fd_sc_hd__nand2_1 _3230_ (.A(_0782_),
    .B(_1106_),
    .Y(_1107_));
 sky130_fd_sc_hd__o22ai_1 _3231_ (.A1(_1063_),
    .A2(_1105_),
    .B1(_1107_),
    .B2(_1884_),
    .Y(_1108_));
 sky130_fd_sc_hd__a21oi_1 _3232_ (.A1(_1105_),
    .A2(_1107_),
    .B1(_1080_),
    .Y(_1109_));
 sky130_fd_sc_hd__nor2_1 _3233_ (.A(_1108_),
    .B(_1109_),
    .Y(_1110_));
 sky130_fd_sc_hd__a21oi_1 _3234_ (.A1(_1030_),
    .A2(_1035_),
    .B1(_1865_),
    .Y(_1111_));
 sky130_fd_sc_hd__nor3_1 _3235_ (.A(_0831_),
    .B(_1873_),
    .C(_1103_),
    .Y(_1112_));
 sky130_fd_sc_hd__o21ai_0 _3236_ (.A1(_1046_),
    .A2(_1111_),
    .B1(_1112_),
    .Y(_1113_));
 sky130_fd_sc_hd__nand3_1 _3237_ (.A(_0831_),
    .B(_1030_),
    .C(_1080_),
    .Y(_1114_));
 sky130_fd_sc_hd__o31ai_1 _3238_ (.A1(_1032_),
    .A2(_1083_),
    .A3(_1114_),
    .B1(_0807_),
    .Y(_1115_));
 sky130_fd_sc_hd__a21oi_1 _3239_ (.A1(_1110_),
    .A2(_1113_),
    .B1(_1115_),
    .Y(_1116_));
 sky130_fd_sc_hd__a22oi_1 _3240_ (.A1(_0779_),
    .A2(_1098_),
    .B1(_1101_),
    .B2(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__xnor2_1 _3241_ (.A(_1095_),
    .B(_1117_),
    .Y(_1118_));
 sky130_fd_sc_hd__nor2_1 _3242_ (.A(_0773_),
    .B(_1118_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_1 _3243_ (.A(_1906_),
    .Y(_1119_));
 sky130_fd_sc_hd__nor2_1 _3244_ (.A(_1119_),
    .B(_0773_),
    .Y(_1120_));
 sky130_fd_sc_hd__nor2_1 _3245_ (.A(_1906_),
    .B(_0773_),
    .Y(_1121_));
 sky130_fd_sc_hd__inv_1 _3246_ (.A(_1095_),
    .Y(_1122_));
 sky130_fd_sc_hd__a21oi_1 _3247_ (.A1(_1122_),
    .A2(_1098_),
    .B1(_1902_),
    .Y(_1123_));
 sky130_fd_sc_hd__nor3_1 _3248_ (.A(_1096_),
    .B(_1122_),
    .C(_1083_),
    .Y(_1124_));
 sky130_fd_sc_hd__inv_1 _3249_ (.A(_1900_),
    .Y(_1125_));
 sky130_fd_sc_hd__a21o_1 _3250_ (.A1(_1874_),
    .A2(_1050_),
    .B1(_1876_),
    .X(_1126_));
 sky130_fd_sc_hd__a21oi_1 _3251_ (.A1(_1063_),
    .A2(_1126_),
    .B1(_1884_),
    .Y(_1127_));
 sky130_fd_sc_hd__nor2_1 _3252_ (.A(_1096_),
    .B(_1127_),
    .Y(_1128_));
 sky130_fd_sc_hd__o21ai_0 _3253_ (.A1(_1892_),
    .A2(_1128_),
    .B1(_1095_),
    .Y(_1129_));
 sky130_fd_sc_hd__a21o_1 _3254_ (.A1(_1874_),
    .A2(_1053_),
    .B1(_1873_),
    .X(_1130_));
 sky130_fd_sc_hd__a21oi_1 _3255_ (.A1(_1882_),
    .A2(_1130_),
    .B1(_1881_),
    .Y(_1131_));
 sky130_fd_sc_hd__o21bai_1 _3256_ (.A1(_1096_),
    .A2(_1131_),
    .B1_N(_1889_),
    .Y(_1132_));
 sky130_fd_sc_hd__a211oi_1 _3257_ (.A1(_1095_),
    .A2(_1132_),
    .B1(_1897_),
    .C1(_0782_),
    .Y(_1133_));
 sky130_fd_sc_hd__a311oi_1 _3258_ (.A1(_0782_),
    .A2(_1125_),
    .A3(_1129_),
    .B1(_1133_),
    .C1(_0777_),
    .Y(_1134_));
 sky130_fd_sc_hd__a221o_1 _3259_ (.A1(_0777_),
    .A2(_1123_),
    .B1(_1124_),
    .B2(_1048_),
    .C1(_1134_),
    .X(_1135_));
 sky130_fd_sc_hd__mux2_1 _3260_ (.A0(_1120_),
    .A1(_1121_),
    .S(_1135_),
    .X(_0014_));
 sky130_fd_sc_hd__a2111oi_1 _3261_ (.A1(_1122_),
    .A2(_1098_),
    .B1(_0807_),
    .C1(_1910_),
    .D1(_1902_),
    .Y(_1136_));
 sky130_fd_sc_hd__nor3_1 _3262_ (.A(_1096_),
    .B(_1122_),
    .C(_1119_),
    .Y(_1137_));
 sky130_fd_sc_hd__nand3_1 _3263_ (.A(_1063_),
    .B(_1099_),
    .C(_1137_),
    .Y(_1138_));
 sky130_fd_sc_hd__inv_1 _3264_ (.A(_1908_),
    .Y(_1139_));
 sky130_fd_sc_hd__o21ai_0 _3265_ (.A1(_1122_),
    .A2(_1102_),
    .B1(_1125_),
    .Y(_1140_));
 sky130_fd_sc_hd__nand2_1 _3266_ (.A(_1906_),
    .B(_1140_),
    .Y(_1141_));
 sky130_fd_sc_hd__a21oi_1 _3267_ (.A1(_1095_),
    .A2(_1103_),
    .B1(_1897_),
    .Y(_1142_));
 sky130_fd_sc_hd__nor2_1 _3268_ (.A(_1119_),
    .B(_1142_),
    .Y(_1143_));
 sky130_fd_sc_hd__nor3_1 _3269_ (.A(_0781_),
    .B(_1905_),
    .C(_1143_),
    .Y(_1144_));
 sky130_fd_sc_hd__a31oi_1 _3270_ (.A1(_0781_),
    .A2(_1139_),
    .A3(_1141_),
    .B1(_1144_),
    .Y(_1145_));
 sky130_fd_sc_hd__a31oi_1 _3271_ (.A1(_1063_),
    .A2(_1072_),
    .A3(_1137_),
    .B1(_1145_),
    .Y(_1146_));
 sky130_fd_sc_hd__o21ai_0 _3272_ (.A1(_1013_),
    .A2(_1138_),
    .B1(_1146_),
    .Y(_1147_));
 sky130_fd_sc_hd__o21ai_0 _3273_ (.A1(_1119_),
    .A2(_1910_),
    .B1(_0777_),
    .Y(_1148_));
 sky130_fd_sc_hd__o21a_1 _3274_ (.A1(_0777_),
    .A2(_1147_),
    .B1(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__o21ai_0 _3275_ (.A1(_1136_),
    .A2(_1149_),
    .B1(_1914_),
    .Y(_1150_));
 sky130_fd_sc_hd__or3_1 _3276_ (.A(_1914_),
    .B(_1136_),
    .C(_1149_),
    .X(_1151_));
 sky130_fd_sc_hd__a21o_1 _3277_ (.A1(_1150_),
    .A2(_1151_),
    .B1(_0773_),
    .X(_0015_));
 sky130_fd_sc_hd__a21oi_1 _3278_ (.A1(_1025_),
    .A2(_1084_),
    .B1(_1091_),
    .Y(_1152_));
 sky130_fd_sc_hd__nand2_1 _3279_ (.A(_1914_),
    .B(_1137_),
    .Y(_1153_));
 sky130_fd_sc_hd__a21oi_1 _3280_ (.A1(_1095_),
    .A2(_1889_),
    .B1(_1897_),
    .Y(_1154_));
 sky130_fd_sc_hd__o21bai_1 _3281_ (.A1(_1119_),
    .A2(_1154_),
    .B1_N(_1905_),
    .Y(_1155_));
 sky130_fd_sc_hd__a21oi_1 _3282_ (.A1(_1914_),
    .A2(_1155_),
    .B1(_1913_),
    .Y(_1156_));
 sky130_fd_sc_hd__inv_1 _3283_ (.A(_1914_),
    .Y(_1157_));
 sky130_fd_sc_hd__o21bai_1 _3284_ (.A1(_1096_),
    .A2(_1086_),
    .B1_N(_1892_),
    .Y(_1158_));
 sky130_fd_sc_hd__a21oi_1 _3285_ (.A1(_1095_),
    .A2(_1158_),
    .B1(_1900_),
    .Y(_1159_));
 sky130_fd_sc_hd__nor2_1 _3286_ (.A(_1119_),
    .B(_1159_),
    .Y(_1160_));
 sky130_fd_sc_hd__nor2_1 _3287_ (.A(_1908_),
    .B(_1160_),
    .Y(_1161_));
 sky130_fd_sc_hd__nor2_1 _3288_ (.A(_1157_),
    .B(_1161_),
    .Y(_1162_));
 sky130_fd_sc_hd__o21ai_0 _3289_ (.A1(_1916_),
    .A2(_1162_),
    .B1(_0797_),
    .Y(_1163_));
 sky130_fd_sc_hd__o221ai_1 _3290_ (.A1(_1152_),
    .A2(_1153_),
    .B1(_1156_),
    .B2(_0797_),
    .C1(_1163_),
    .Y(_1164_));
 sky130_fd_sc_hd__a21oi_1 _3291_ (.A1(_1910_),
    .A2(_1157_),
    .B1(_1918_),
    .Y(_1165_));
 sky130_fd_sc_hd__o311a_1 _3292_ (.A1(_1906_),
    .A2(_1914_),
    .A3(_1123_),
    .B1(_1165_),
    .C1(_0779_),
    .X(_1166_));
 sky130_fd_sc_hd__a211oi_1 _3293_ (.A1(_0808_),
    .A2(_1164_),
    .B1(_1166_),
    .C1(_0773_),
    .Y(_0016_));
 sky130_fd_sc_hd__nor2_1 _3294_ (.A(_1185_),
    .B(_1188_),
    .Y(_1167_));
 sky130_fd_sc_hd__nor2_1 _3295_ (.A(_0767_),
    .B(_0768_),
    .Y(_1168_));
 sky130_fd_sc_hd__nand2_1 _3296_ (.A(_1577_),
    .B(_1201_),
    .Y(_1169_));
 sky130_fd_sc_hd__nand2_1 _3297_ (.A(net26),
    .B(_0772_),
    .Y(_1170_));
 sky130_fd_sc_hd__o21ai_0 _3298_ (.A1(_0772_),
    .A2(_1169_),
    .B1(_1170_),
    .Y(_1171_));
 sky130_fd_sc_hd__mux2i_1 _3299_ (.A0(b_sign_stage1),
    .A1(a_sign_stage1),
    .S(_0797_),
    .Y(_1172_));
 sky130_fd_sc_hd__a21oi_1 _3300_ (.A1(net58),
    .A2(_1201_),
    .B1(_0772_),
    .Y(_1173_));
 sky130_fd_sc_hd__a211oi_1 _3301_ (.A1(_0772_),
    .A2(_1172_),
    .B1(_1173_),
    .C1(_1168_),
    .Y(_1174_));
 sky130_fd_sc_hd__a31o_1 _3302_ (.A1(_1167_),
    .A2(_1168_),
    .A3(_1171_),
    .B1(_1174_),
    .X(_0119_));
 sky130_fd_sc_hd__nor3_1 _3303_ (.A(_0306_),
    .B(_0323_),
    .C(_0325_),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_1 _3304_ (.A(net25),
    .Y(_1579_));
 sky130_fd_sc_hd__inv_1 _3305_ (.A(net23),
    .Y(_1585_));
 sky130_fd_sc_hd__inv_1 _3306_ (.A(net22),
    .Y(_1591_));
 sky130_fd_sc_hd__inv_1 _3307_ (.A(net21),
    .Y(_1597_));
 sky130_fd_sc_hd__inv_1 _3308_ (.A(net20),
    .Y(_1603_));
 sky130_fd_sc_hd__inv_1 _3309_ (.A(net19),
    .Y(_1609_));
 sky130_fd_sc_hd__inv_1 _3310_ (.A(net18),
    .Y(_1565_));
 sky130_fd_sc_hd__inv_1 _3311_ (.A(_1692_),
    .Y(_1566_));
 sky130_fd_sc_hd__inv_1 _3312_ (.A(_1689_),
    .Y(_1570_));
 sky130_fd_sc_hd__inv_1 _3313_ (.A(net17),
    .Y(_1688_));
 sky130_fd_sc_hd__inv_1 _3314_ (.A(\aligned_a_mant[2] ),
    .Y(_1720_));
 sky130_fd_sc_hd__inv_1 _3315_ (.A(\aligned_a_mant[1] ),
    .Y(_1728_));
 sky130_fd_sc_hd__inv_1 _3316_ (.A(\aligned_a_mant[3] ),
    .Y(_1736_));
 sky130_fd_sc_hd__inv_1 _3317_ (.A(\aligned_a_mant[4] ),
    .Y(_1744_));
 sky130_fd_sc_hd__inv_1 _3318_ (.A(\aligned_a_mant[5] ),
    .Y(_1752_));
 sky130_fd_sc_hd__inv_1 _3319_ (.A(\aligned_a_mant[6] ),
    .Y(_1760_));
 sky130_fd_sc_hd__inv_1 _3320_ (.A(\aligned_a_mant[7] ),
    .Y(_1768_));
 sky130_fd_sc_hd__inv_1 _3321_ (.A(\aligned_a_mant[8] ),
    .Y(_1776_));
 sky130_fd_sc_hd__inv_1 _3322_ (.A(\aligned_a_mant[9] ),
    .Y(_1784_));
 sky130_fd_sc_hd__inv_1 _3323_ (.A(\aligned_a_mant[10] ),
    .Y(_1792_));
 sky130_fd_sc_hd__inv_1 _3324_ (.A(\aligned_a_mant[11] ),
    .Y(_1800_));
 sky130_fd_sc_hd__inv_1 _3325_ (.A(\aligned_a_mant[12] ),
    .Y(_1808_));
 sky130_fd_sc_hd__inv_1 _3326_ (.A(\aligned_a_mant[13] ),
    .Y(_1816_));
 sky130_fd_sc_hd__inv_1 _3327_ (.A(\aligned_a_mant[14] ),
    .Y(_1824_));
 sky130_fd_sc_hd__inv_1 _3328_ (.A(\aligned_a_mant[15] ),
    .Y(_1832_));
 sky130_fd_sc_hd__inv_1 _3329_ (.A(\aligned_a_mant[16] ),
    .Y(_1840_));
 sky130_fd_sc_hd__inv_1 _3330_ (.A(\aligned_a_mant[17] ),
    .Y(_1848_));
 sky130_fd_sc_hd__inv_1 _3331_ (.A(\aligned_a_mant[18] ),
    .Y(_1856_));
 sky130_fd_sc_hd__inv_1 _3332_ (.A(\aligned_a_mant[19] ),
    .Y(_1864_));
 sky130_fd_sc_hd__inv_1 _3333_ (.A(\aligned_a_mant[20] ),
    .Y(_1872_));
 sky130_fd_sc_hd__inv_1 _3334_ (.A(\aligned_a_mant[21] ),
    .Y(_1880_));
 sky130_fd_sc_hd__inv_1 _3335_ (.A(\aligned_a_mant[22] ),
    .Y(_1888_));
 sky130_fd_sc_hd__inv_1 _3336_ (.A(\aligned_a_mant[23] ),
    .Y(_1896_));
 sky130_fd_sc_hd__inv_1 _3337_ (.A(\aligned_a_mant[24] ),
    .Y(_1904_));
 sky130_fd_sc_hd__inv_1 _3338_ (.A(\aligned_a_mant[25] ),
    .Y(_1912_));
 sky130_fd_sc_hd__inv_1 _3339_ (.A(\aligned_b_mant[2] ),
    .Y(_1723_));
 sky130_fd_sc_hd__inv_1 _3340_ (.A(\aligned_b_mant[1] ),
    .Y(_1731_));
 sky130_fd_sc_hd__inv_1 _3341_ (.A(\aligned_b_mant[3] ),
    .Y(_1739_));
 sky130_fd_sc_hd__inv_1 _3342_ (.A(\aligned_b_mant[4] ),
    .Y(_1747_));
 sky130_fd_sc_hd__inv_1 _3343_ (.A(\aligned_b_mant[5] ),
    .Y(_1755_));
 sky130_fd_sc_hd__inv_1 _3344_ (.A(\aligned_b_mant[6] ),
    .Y(_1763_));
 sky130_fd_sc_hd__inv_1 _3345_ (.A(\aligned_b_mant[7] ),
    .Y(_1771_));
 sky130_fd_sc_hd__inv_1 _3346_ (.A(\aligned_b_mant[8] ),
    .Y(_1779_));
 sky130_fd_sc_hd__inv_1 _3347_ (.A(\aligned_b_mant[9] ),
    .Y(_1787_));
 sky130_fd_sc_hd__inv_1 _3348_ (.A(\aligned_b_mant[10] ),
    .Y(_1795_));
 sky130_fd_sc_hd__inv_1 _3349_ (.A(\aligned_b_mant[11] ),
    .Y(_1803_));
 sky130_fd_sc_hd__inv_1 _3350_ (.A(\aligned_b_mant[12] ),
    .Y(_1811_));
 sky130_fd_sc_hd__inv_1 _3351_ (.A(\aligned_b_mant[13] ),
    .Y(_1819_));
 sky130_fd_sc_hd__inv_1 _3352_ (.A(\aligned_b_mant[14] ),
    .Y(_1827_));
 sky130_fd_sc_hd__inv_1 _3353_ (.A(\aligned_b_mant[15] ),
    .Y(_1835_));
 sky130_fd_sc_hd__inv_1 _3354_ (.A(\aligned_b_mant[16] ),
    .Y(_1843_));
 sky130_fd_sc_hd__inv_1 _3355_ (.A(\aligned_b_mant[17] ),
    .Y(_1851_));
 sky130_fd_sc_hd__inv_1 _3356_ (.A(\aligned_b_mant[18] ),
    .Y(_1859_));
 sky130_fd_sc_hd__inv_1 _3357_ (.A(\aligned_b_mant[19] ),
    .Y(_1867_));
 sky130_fd_sc_hd__inv_1 _3358_ (.A(\aligned_b_mant[20] ),
    .Y(_1875_));
 sky130_fd_sc_hd__inv_1 _3359_ (.A(\aligned_b_mant[21] ),
    .Y(_1883_));
 sky130_fd_sc_hd__inv_1 _3360_ (.A(\aligned_b_mant[22] ),
    .Y(_1891_));
 sky130_fd_sc_hd__inv_1 _3361_ (.A(\aligned_b_mant[23] ),
    .Y(_1899_));
 sky130_fd_sc_hd__inv_1 _3362_ (.A(\aligned_b_mant[24] ),
    .Y(_1907_));
 sky130_fd_sc_hd__inv_1 _3363_ (.A(\aligned_b_mant[25] ),
    .Y(_1915_));
 sky130_fd_sc_hd__nand2_1 _3364_ (.A(_1578_),
    .B(_1168_),
    .Y(_1175_));
 sky130_fd_sc_hd__a21oi_1 _3365_ (.A1(_1201_),
    .A2(_1175_),
    .B1(_0772_),
    .Y(_1176_));
 sky130_fd_sc_hd__nor3_1 _3366_ (.A(_1167_),
    .B(_0767_),
    .C(_0768_),
    .Y(_1177_));
 sky130_fd_sc_hd__or3_1 _3367_ (.A(invalid_op_stage2),
    .B(_1176_),
    .C(_1177_),
    .X(_0121_));
 sky130_fd_sc_hd__or4_2 _3368_ (.A(\aligned_a_mant[1] ),
    .B(\aligned_a_mant[0] ),
    .C(\aligned_b_mant[1] ),
    .D(\aligned_b_mant[0] ),
    .X(_0109_));
 sky130_fd_sc_hd__inv_1 _3369_ (.A(net49),
    .Y(_1691_));
 sky130_fd_sc_hd__nor4_2 _3370_ (.A(net22),
    .B(net21),
    .C(net25),
    .D(net23),
    .Y(_1178_));
 sky130_fd_sc_hd__nor4_1 _3371_ (.A(net18),
    .B(net17),
    .C(net20),
    .D(net19),
    .Y(_1179_));
 sky130_fd_sc_hd__nand2_2 _3372_ (.A(_1178_),
    .B(_1179_),
    .Y(_1180_));
 sky130_fd_sc_hd__nor4_2 _3373_ (.A(net13),
    .B(net2),
    .C(net27),
    .D(net16),
    .Y(_1181_));
 sky130_fd_sc_hd__nor4_1 _3374_ (.A(net9),
    .B(net11),
    .C(net15),
    .D(net14),
    .Y(_1182_));
 sky130_fd_sc_hd__nor4_1 _3375_ (.A(net3),
    .B(net7),
    .C(net10),
    .D(net12),
    .Y(_1183_));
 sky130_fd_sc_hd__nor3_1 _3376_ (.A(net6),
    .B(net5),
    .C(net8),
    .Y(_1184_));
 sky130_fd_sc_hd__nand4_2 _3377_ (.A(_1181_),
    .B(_1182_),
    .C(_1183_),
    .D(_1184_),
    .Y(_1185_));
 sky130_fd_sc_hd__nor4_1 _3378_ (.A(net28),
    .B(net30),
    .C(net33),
    .D(net32),
    .Y(_1186_));
 sky130_fd_sc_hd__nor4_1 _3379_ (.A(net24),
    .B(net29),
    .C(net31),
    .D(net4),
    .Y(_1187_));
 sky130_fd_sc_hd__nand2_2 _3380_ (.A(_1186_),
    .B(_1187_),
    .Y(_1188_));
 sky130_fd_sc_hd__nor3_4 _3381_ (.A(_1180_),
    .B(_1185_),
    .C(_1188_),
    .Y(_1189_));
 sky130_fd_sc_hd__inv_1 _3382_ (.A(net54),
    .Y(_1594_));
 sky130_fd_sc_hd__inv_1 _3383_ (.A(net53),
    .Y(_1600_));
 sky130_fd_sc_hd__inv_1 _3384_ (.A(net57),
    .Y(_1582_));
 sky130_fd_sc_hd__inv_1 _3385_ (.A(net55),
    .Y(_1588_));
 sky130_fd_sc_hd__nand4_2 _3386_ (.A(_1594_),
    .B(_1600_),
    .C(_1582_),
    .D(_1588_),
    .Y(_1190_));
 sky130_fd_sc_hd__inv_1 _3387_ (.A(net50),
    .Y(_1569_));
 sky130_fd_sc_hd__inv_1 _3388_ (.A(net52),
    .Y(_1606_));
 sky130_fd_sc_hd__inv_1 _3389_ (.A(net51),
    .Y(_1612_));
 sky130_fd_sc_hd__nand4_1 _3390_ (.A(_1569_),
    .B(_1691_),
    .C(_1606_),
    .D(_1612_),
    .Y(_1191_));
 sky130_fd_sc_hd__nor2_4 _3391_ (.A(_1190_),
    .B(_1191_),
    .Y(_1192_));
 sky130_fd_sc_hd__nor4_2 _3392_ (.A(net45),
    .B(net34),
    .C(net59),
    .D(net48),
    .Y(_1193_));
 sky130_fd_sc_hd__nor4_1 _3393_ (.A(net41),
    .B(net43),
    .C(net47),
    .D(net46),
    .Y(_1194_));
 sky130_fd_sc_hd__nor4_1 _3394_ (.A(net35),
    .B(net39),
    .C(net42),
    .D(net44),
    .Y(_1195_));
 sky130_fd_sc_hd__nor3_1 _3395_ (.A(net38),
    .B(net37),
    .C(net40),
    .Y(_1196_));
 sky130_fd_sc_hd__nand4_2 _3396_ (.A(_1193_),
    .B(_1194_),
    .C(_1195_),
    .D(_1196_),
    .Y(_1197_));
 sky130_fd_sc_hd__nor4_1 _3397_ (.A(net60),
    .B(net62),
    .C(net65),
    .D(net64),
    .Y(_1198_));
 sky130_fd_sc_hd__nor4_1 _3398_ (.A(net56),
    .B(net61),
    .C(net63),
    .D(net36),
    .Y(_1199_));
 sky130_fd_sc_hd__nand2_2 _3399_ (.A(_1198_),
    .B(_1199_),
    .Y(_1200_));
 sky130_fd_sc_hd__nor2_4 _3400_ (.A(_1197_),
    .B(_1200_),
    .Y(_1201_));
 sky130_fd_sc_hd__a21o_1 _3401_ (.A1(_1687_),
    .A2(_1668_),
    .B1(_1686_),
    .X(_1202_));
 sky130_fd_sc_hd__a21o_1 _3402_ (.A1(_1684_),
    .A2(_1202_),
    .B1(_1683_),
    .X(_1203_));
 sky130_fd_sc_hd__buf_6 _3403_ (.A(_1605_),
    .X(_1204_));
 sky130_fd_sc_hd__nand4_2 _3404_ (.A(_1611_),
    .B(_1204_),
    .C(_1690_),
    .D(_1616_),
    .Y(_1205_));
 sky130_fd_sc_hd__nand4_4 _3405_ (.A(_1587_),
    .B(_1599_),
    .C(_1581_),
    .D(_1593_),
    .Y(_1206_));
 sky130_fd_sc_hd__a2111oi_4 _3406_ (.A1(_1681_),
    .A2(_1203_),
    .B1(_1205_),
    .C1(_1206_),
    .D1(_1680_),
    .Y(_1207_));
 sky130_fd_sc_hd__and4_1 _3407_ (.A(_1645_),
    .B(_1672_),
    .C(_1675_),
    .D(_1678_),
    .X(_1208_));
 sky130_fd_sc_hd__and3_1 _3408_ (.A(_1648_),
    .B(_1651_),
    .C(_1654_),
    .X(_1209_));
 sky130_fd_sc_hd__and4_1 _3409_ (.A(_1633_),
    .B(_1660_),
    .C(_1663_),
    .D(_1666_),
    .X(_1210_));
 sky130_fd_sc_hd__nand4_1 _3410_ (.A(_1657_),
    .B(_1208_),
    .C(_1209_),
    .D(_1210_),
    .Y(_1211_));
 sky130_fd_sc_hd__a21oi_1 _3411_ (.A1(_1626_),
    .A2(_1642_),
    .B1(_1641_),
    .Y(_1212_));
 sky130_fd_sc_hd__nand2_1 _3412_ (.A(_1636_),
    .B(_1639_),
    .Y(_1213_));
 sky130_fd_sc_hd__a21oi_1 _3413_ (.A1(_1636_),
    .A2(_1638_),
    .B1(_1635_),
    .Y(_1214_));
 sky130_fd_sc_hd__o21a_1 _3414_ (.A1(_1212_),
    .A2(_1213_),
    .B1(_1214_),
    .X(_1215_));
 sky130_fd_sc_hd__nand2_1 _3415_ (.A(_1660_),
    .B(_1663_),
    .Y(_1216_));
 sky130_fd_sc_hd__a21oi_1 _3416_ (.A1(_1632_),
    .A2(_1666_),
    .B1(_1665_),
    .Y(_1217_));
 sky130_fd_sc_hd__a21oi_1 _3417_ (.A1(_1662_),
    .A2(_1660_),
    .B1(_1659_),
    .Y(_1218_));
 sky130_fd_sc_hd__o21ai_1 _3418_ (.A1(_1216_),
    .A2(_1217_),
    .B1(_1218_),
    .Y(_1219_));
 sky130_fd_sc_hd__and3_1 _3419_ (.A(_1657_),
    .B(_1208_),
    .C(_1209_),
    .X(_1220_));
 sky130_fd_sc_hd__a2bb2oi_2 _3420_ (.A1_N(_1211_),
    .A2_N(_1215_),
    .B1(_1219_),
    .B2(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hd__a21o_1 _3421_ (.A1(_1644_),
    .A2(_1678_),
    .B1(_1677_),
    .X(_1222_));
 sky130_fd_sc_hd__a21o_1 _3422_ (.A1(_1675_),
    .A2(_1222_),
    .B1(_1674_),
    .X(_1223_));
 sky130_fd_sc_hd__a21oi_1 _3423_ (.A1(_1672_),
    .A2(_1223_),
    .B1(_1671_),
    .Y(_1224_));
 sky130_fd_sc_hd__nand2b_1 _3424_ (.A_N(_1624_),
    .B(_1623_),
    .Y(_1225_));
 sky130_fd_sc_hd__a21o_1 _3425_ (.A1(_1620_),
    .A2(_1630_),
    .B1(_1629_),
    .X(_1226_));
 sky130_fd_sc_hd__a31oi_2 _3426_ (.A1(_1621_),
    .A2(_1630_),
    .A3(_1225_),
    .B1(_1226_),
    .Y(_1227_));
 sky130_fd_sc_hd__nand4_1 _3427_ (.A(_1636_),
    .B(_1627_),
    .C(_1639_),
    .D(_1642_),
    .Y(_1228_));
 sky130_fd_sc_hd__a21o_1 _3428_ (.A1(_1651_),
    .A2(_1653_),
    .B1(_1650_),
    .X(_1229_));
 sky130_fd_sc_hd__a221oi_1 _3429_ (.A1(_1656_),
    .A2(_1209_),
    .B1(_1229_),
    .B2(_1648_),
    .C1(_1647_),
    .Y(_1230_));
 sky130_fd_sc_hd__nand4_1 _3430_ (.A(_1645_),
    .B(_1672_),
    .C(_1675_),
    .D(_1678_),
    .Y(_1231_));
 sky130_fd_sc_hd__o32a_1 _3431_ (.A1(_1211_),
    .A2(_1227_),
    .A3(_1228_),
    .B1(_1230_),
    .B2(_1231_),
    .X(_1232_));
 sky130_fd_sc_hd__nand4_4 _3432_ (.A(_1207_),
    .B(_1221_),
    .C(_1224_),
    .D(_1232_),
    .Y(_1233_));
 sky130_fd_sc_hd__nand3b_1 _3433_ (.A_N(_1689_),
    .B(_1616_),
    .C(_1611_),
    .Y(_1234_));
 sky130_fd_sc_hd__a21oi_1 _3434_ (.A1(_1611_),
    .A2(_1617_),
    .B1(_1613_),
    .Y(_1235_));
 sky130_fd_sc_hd__nand4_1 _3435_ (.A(_1587_),
    .B(_1599_),
    .C(_1204_),
    .D(_1593_),
    .Y(_1236_));
 sky130_fd_sc_hd__a21oi_2 _3436_ (.A1(_1234_),
    .A2(_1235_),
    .B1(_1236_),
    .Y(_1237_));
 sky130_fd_sc_hd__buf_6 _3437_ (.A(_1599_),
    .X(_1238_));
 sky130_fd_sc_hd__buf_6 _3438_ (.A(_1593_),
    .X(_1239_));
 sky130_fd_sc_hd__nand3_1 _3439_ (.A(_1238_),
    .B(_1239_),
    .C(_1607_),
    .Y(_1240_));
 sky130_fd_sc_hd__a21oi_1 _3440_ (.A1(_1239_),
    .A2(_1601_),
    .B1(_1595_),
    .Y(_1241_));
 sky130_fd_sc_hd__inv_1 _3441_ (.A(_1587_),
    .Y(_1242_));
 sky130_fd_sc_hd__a21oi_1 _3442_ (.A1(_1240_),
    .A2(_1241_),
    .B1(_1242_),
    .Y(_1243_));
 sky130_fd_sc_hd__o31ai_4 _3443_ (.A1(_1589_),
    .A2(_1237_),
    .A3(_1243_),
    .B1(_1581_),
    .Y(_1244_));
 sky130_fd_sc_hd__nor2_1 _3444_ (.A(_1206_),
    .B(_1205_),
    .Y(_1245_));
 sky130_fd_sc_hd__nor2_1 _3445_ (.A(_1583_),
    .B(_1245_),
    .Y(_1246_));
 sky130_fd_sc_hd__nand4_2 _3446_ (.A(_1687_),
    .B(_1681_),
    .C(_1669_),
    .D(_1684_),
    .Y(_1247_));
 sky130_fd_sc_hd__a22oi_4 _3447_ (.A1(_1244_),
    .A2(_1246_),
    .B1(_1207_),
    .B2(_1247_),
    .Y(_1248_));
 sky130_fd_sc_hd__nand2_4 _3448_ (.A(_1233_),
    .B(_1248_),
    .Y(_1249_));
 sky130_fd_sc_hd__inv_2 _3449_ (.A(_1249_),
    .Y(a_exp_larger));
 sky130_fd_sc_hd__a21oi_2 _3450_ (.A1(_1192_),
    .A2(_1201_),
    .B1(a_exp_larger),
    .Y(_1250_));
 sky130_fd_sc_hd__nor2_4 _3451_ (.A(_1189_),
    .B(_1250_),
    .Y(_1251_));
 sky130_fd_sc_hd__buf_2 _3452_ (.A(_1251_),
    .X(_1252_));
 sky130_fd_sc_hd__buf_2 _3453_ (.A(_1251_),
    .X(_1253_));
 sky130_fd_sc_hd__nand2_1 _3454_ (.A(net17),
    .B(_1253_),
    .Y(_1254_));
 sky130_fd_sc_hd__o21ai_0 _3455_ (.A1(_1691_),
    .A2(_1252_),
    .B1(_1254_),
    .Y(_0110_));
 sky130_fd_sc_hd__nand2_1 _3456_ (.A(net18),
    .B(_1253_),
    .Y(_1255_));
 sky130_fd_sc_hd__o21ai_0 _3457_ (.A1(_1569_),
    .A2(_1252_),
    .B1(_1255_),
    .Y(_0111_));
 sky130_fd_sc_hd__nand2_1 _3458_ (.A(net19),
    .B(_1253_),
    .Y(_1256_));
 sky130_fd_sc_hd__o21ai_0 _3459_ (.A1(_1612_),
    .A2(_1252_),
    .B1(_1256_),
    .Y(_0112_));
 sky130_fd_sc_hd__nand2_1 _3460_ (.A(net20),
    .B(_1253_),
    .Y(_1257_));
 sky130_fd_sc_hd__o21ai_0 _3461_ (.A1(_1606_),
    .A2(_1252_),
    .B1(_1257_),
    .Y(_0113_));
 sky130_fd_sc_hd__nand2_1 _3462_ (.A(net21),
    .B(_1253_),
    .Y(_1258_));
 sky130_fd_sc_hd__o21ai_0 _3463_ (.A1(_1600_),
    .A2(_1252_),
    .B1(_1258_),
    .Y(_0114_));
 sky130_fd_sc_hd__nand2_1 _3464_ (.A(net22),
    .B(_1253_),
    .Y(_1259_));
 sky130_fd_sc_hd__o21ai_0 _3465_ (.A1(_1594_),
    .A2(_1252_),
    .B1(_1259_),
    .Y(_0115_));
 sky130_fd_sc_hd__buf_4 _3466_ (.A(_1251_),
    .X(_1260_));
 sky130_fd_sc_hd__nand2_1 _3467_ (.A(net23),
    .B(_1260_),
    .Y(_1261_));
 sky130_fd_sc_hd__o21ai_0 _3468_ (.A1(_1588_),
    .A2(_1252_),
    .B1(_1261_),
    .Y(_0116_));
 sky130_fd_sc_hd__nand2_1 _3469_ (.A(net25),
    .B(_1260_),
    .Y(_1262_));
 sky130_fd_sc_hd__o21ai_0 _3470_ (.A1(_1582_),
    .A2(_1252_),
    .B1(_1262_),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_1 _3471_ (.A(net2),
    .Y(_1622_));
 sky130_fd_sc_hd__inv_1 _3472_ (.A(net45),
    .Y(_1619_));
 sky130_fd_sc_hd__inv_1 _3473_ (.A(net56),
    .Y(_1628_));
 sky130_fd_sc_hd__inv_1 _3474_ (.A(net59),
    .Y(_1625_));
 sky130_fd_sc_hd__inv_1 _3475_ (.A(net60),
    .Y(_1640_));
 sky130_fd_sc_hd__inv_1 _3476_ (.A(net61),
    .Y(_1637_));
 sky130_fd_sc_hd__inv_1 _3477_ (.A(net62),
    .Y(_1634_));
 sky130_fd_sc_hd__inv_1 _3478_ (.A(net63),
    .Y(_1631_));
 sky130_fd_sc_hd__clkinvlp_4 _3479_ (.A(net64),
    .Y(_1664_));
 sky130_fd_sc_hd__inv_1 _3480_ (.A(net65),
    .Y(_1661_));
 sky130_fd_sc_hd__inv_1 _3481_ (.A(net35),
    .Y(_1658_));
 sky130_fd_sc_hd__inv_1 _3482_ (.A(net36),
    .Y(_1655_));
 sky130_fd_sc_hd__inv_1 _3483_ (.A(net37),
    .Y(_1652_));
 sky130_fd_sc_hd__inv_1 _3484_ (.A(net38),
    .Y(_1649_));
 sky130_fd_sc_hd__inv_1 _3485_ (.A(net39),
    .Y(_1646_));
 sky130_fd_sc_hd__clkinv_2 _3486_ (.A(net40),
    .Y(_1643_));
 sky130_fd_sc_hd__inv_1 _3487_ (.A(net41),
    .Y(_1676_));
 sky130_fd_sc_hd__inv_1 _3488_ (.A(net42),
    .Y(_1673_));
 sky130_fd_sc_hd__inv_1 _3489_ (.A(net43),
    .Y(_1670_));
 sky130_fd_sc_hd__inv_1 _3490_ (.A(net44),
    .Y(_1667_));
 sky130_fd_sc_hd__inv_1 _3491_ (.A(net46),
    .Y(_1685_));
 sky130_fd_sc_hd__inv_1 _3492_ (.A(net47),
    .Y(_1682_));
 sky130_fd_sc_hd__inv_1 _3493_ (.A(net48),
    .Y(_1679_));
 sky130_fd_sc_hd__inv_2 _3494_ (.A(_1204_),
    .Y(_1263_));
 sky130_fd_sc_hd__a21oi_1 _3495_ (.A1(_1611_),
    .A2(_1567_),
    .B1(_1610_),
    .Y(_1264_));
 sky130_fd_sc_hd__o21ba_2 _3496_ (.A1(_1263_),
    .A2(_1264_),
    .B1_N(_1604_),
    .X(_1265_));
 sky130_fd_sc_hd__and4_1 _3497_ (.A(_1207_),
    .B(_1221_),
    .C(_1224_),
    .D(_1232_),
    .X(_1266_));
 sky130_fd_sc_hd__clkbuf_2 _3498_ (.A(_1266_),
    .X(_1267_));
 sky130_fd_sc_hd__a22o_2 _3499_ (.A1(_1244_),
    .A2(_1246_),
    .B1(_1207_),
    .B2(_1247_),
    .X(_1268_));
 sky130_fd_sc_hd__clkbuf_2 _3500_ (.A(_1611_),
    .X(_1269_));
 sky130_fd_sc_hd__a21oi_1 _3501_ (.A1(_1269_),
    .A2(_1571_),
    .B1(_1613_),
    .Y(_1270_));
 sky130_fd_sc_hd__o21bai_2 _3502_ (.A1(_1263_),
    .A2(_1270_),
    .B1_N(_1607_),
    .Y(_1271_));
 sky130_fd_sc_hd__nor3_1 _3503_ (.A(_1267_),
    .B(_1268_),
    .C(_1271_),
    .Y(_1272_));
 sky130_fd_sc_hd__a21oi_4 _3504_ (.A1(_1249_),
    .A2(_1265_),
    .B1(_1272_),
    .Y(_1273_));
 sky130_fd_sc_hd__xnor2_4 _3505_ (.A(_1238_),
    .B(_1273_),
    .Y(_1274_));
 sky130_fd_sc_hd__nand2b_1 _3506_ (.A_N(_1692_),
    .B(_1616_),
    .Y(_1275_));
 sky130_fd_sc_hd__nor2_1 _3507_ (.A(_1610_),
    .B(_1615_),
    .Y(_1276_));
 sky130_fd_sc_hd__nor2_1 _3508_ (.A(_1611_),
    .B(_1610_),
    .Y(_1277_));
 sky130_fd_sc_hd__a211oi_1 _3509_ (.A1(_1275_),
    .A2(_1276_),
    .B1(_1277_),
    .C1(_1236_),
    .Y(_1278_));
 sky130_fd_sc_hd__a21oi_1 _3510_ (.A1(_1593_),
    .A2(_1598_),
    .B1(_1592_),
    .Y(_1279_));
 sky130_fd_sc_hd__nand3_1 _3511_ (.A(_1238_),
    .B(_1593_),
    .C(_1604_),
    .Y(_1280_));
 sky130_fd_sc_hd__a21oi_1 _3512_ (.A1(_1279_),
    .A2(_1280_),
    .B1(_1242_),
    .Y(_1281_));
 sky130_fd_sc_hd__o31ai_1 _3513_ (.A1(_1586_),
    .A2(_1278_),
    .A3(_1281_),
    .B1(_1581_),
    .Y(_1282_));
 sky130_fd_sc_hd__or4_1 _3514_ (.A(_1581_),
    .B(_1586_),
    .C(_1278_),
    .D(_1281_),
    .X(_1283_));
 sky130_fd_sc_hd__nand3_1 _3515_ (.A(_1238_),
    .B(_1204_),
    .C(_1239_),
    .Y(_1284_));
 sky130_fd_sc_hd__o211ai_1 _3516_ (.A1(_1284_),
    .A2(_1264_),
    .B1(_1279_),
    .C1(_1280_),
    .Y(_1285_));
 sky130_fd_sc_hd__xnor2_1 _3517_ (.A(_1242_),
    .B(_1285_),
    .Y(_1286_));
 sky130_fd_sc_hd__a211o_1 _3518_ (.A1(_1239_),
    .A2(_1598_),
    .B1(_1592_),
    .C1(_1586_),
    .X(_1287_));
 sky130_fd_sc_hd__o21a_1 _3519_ (.A1(_1587_),
    .A2(_1586_),
    .B1(_1581_),
    .X(_1288_));
 sky130_fd_sc_hd__a21oi_1 _3520_ (.A1(_1287_),
    .A2(_1288_),
    .B1(_1580_),
    .Y(_1289_));
 sky130_fd_sc_hd__o21a_1 _3521_ (.A1(_1206_),
    .A2(_1265_),
    .B1(_1289_),
    .X(_1290_));
 sky130_fd_sc_hd__a211o_1 _3522_ (.A1(_1282_),
    .A2(_1283_),
    .B1(_1286_),
    .C1(_1290_),
    .X(_1291_));
 sky130_fd_sc_hd__buf_6 _3523_ (.A(_1291_),
    .X(_1292_));
 sky130_fd_sc_hd__a21oi_4 _3524_ (.A1(_1233_),
    .A2(_1248_),
    .B1(_1292_),
    .Y(_1293_));
 sky130_fd_sc_hd__clkbuf_4 _3525_ (.A(_1568_),
    .X(_1294_));
 sky130_fd_sc_hd__a21oi_4 _3526_ (.A1(_1192_),
    .A2(_1201_),
    .B1(_1189_),
    .Y(_1295_));
 sky130_fd_sc_hd__a21oi_2 _3527_ (.A1(_1275_),
    .A2(_1276_),
    .B1(_1277_),
    .Y(_1296_));
 sky130_fd_sc_hd__nand2_1 _3528_ (.A(_1204_),
    .B(_1296_),
    .Y(_1297_));
 sky130_fd_sc_hd__buf_4 _3529_ (.A(_1690_),
    .X(_1298_));
 sky130_fd_sc_hd__inv_1 _3530_ (.A(_1298_),
    .Y(_1299_));
 sky130_fd_sc_hd__nand2_1 _3531_ (.A(_1269_),
    .B(_1567_),
    .Y(_1300_));
 sky130_fd_sc_hd__or2_0 _3532_ (.A(_1269_),
    .B(_1567_),
    .X(_1301_));
 sky130_fd_sc_hd__a22o_1 _3533_ (.A1(_1299_),
    .A2(_1294_),
    .B1(_1300_),
    .B2(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__nand2b_1 _3534_ (.A_N(_1296_),
    .B(_1263_),
    .Y(_1303_));
 sky130_fd_sc_hd__xnor2_2 _3535_ (.A(_1238_),
    .B(_1265_),
    .Y(_1304_));
 sky130_fd_sc_hd__o21ai_0 _3536_ (.A1(_1269_),
    .A2(_1610_),
    .B1(_1204_),
    .Y(_1305_));
 sky130_fd_sc_hd__a21oi_1 _3537_ (.A1(_1275_),
    .A2(_1276_),
    .B1(_1305_),
    .Y(_1306_));
 sky130_fd_sc_hd__nand2b_1 _3538_ (.A_N(_1598_),
    .B(_1239_),
    .Y(_1307_));
 sky130_fd_sc_hd__inv_1 _3539_ (.A(_1238_),
    .Y(_1308_));
 sky130_fd_sc_hd__a2111o_1 _3540_ (.A1(_1275_),
    .A2(_1276_),
    .B1(_1305_),
    .C1(_1239_),
    .D1(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__inv_2 _3541_ (.A(_1239_),
    .Y(_1310_));
 sky130_fd_sc_hd__nor2b_1 _3542_ (.A(_1239_),
    .B_N(_1238_),
    .Y(_1311_));
 sky130_fd_sc_hd__nor3b_1 _3543_ (.A(_1238_),
    .B(_1598_),
    .C_N(_1239_),
    .Y(_1312_));
 sky130_fd_sc_hd__a221oi_2 _3544_ (.A1(_1310_),
    .A2(_1598_),
    .B1(_1604_),
    .B2(_1311_),
    .C1(_1312_),
    .Y(_1313_));
 sky130_fd_sc_hd__o311ai_4 _3545_ (.A1(_1604_),
    .A2(_1306_),
    .A3(_1307_),
    .B1(_1309_),
    .C1(_1313_),
    .Y(_1314_));
 sky130_fd_sc_hd__a41oi_4 _3546_ (.A1(_1297_),
    .A2(_1302_),
    .A3(_1303_),
    .A4(_1304_),
    .B1(_1314_),
    .Y(_1315_));
 sky130_fd_sc_hd__nand2_8 _3547_ (.A(_1295_),
    .B(_1315_),
    .Y(_1316_));
 sky130_fd_sc_hd__mux4_1 _3548_ (.A0(net3),
    .A1(net5),
    .A2(net35),
    .A3(net37),
    .S0(_1294_),
    .S1(_1316_),
    .X(_1317_));
 sky130_fd_sc_hd__clkbuf_4 _3549_ (.A(_1572_),
    .X(_1318_));
 sky130_fd_sc_hd__clkbuf_4 _3550_ (.A(_1318_),
    .X(_1319_));
 sky130_fd_sc_hd__nand2_1 _3551_ (.A(net37),
    .B(_1319_),
    .Y(_1320_));
 sky130_fd_sc_hd__o21ai_1 _3552_ (.A1(_1658_),
    .A2(_1319_),
    .B1(_1320_),
    .Y(_1321_));
 sky130_fd_sc_hd__or4_1 _3553_ (.A(_1581_),
    .B(_1589_),
    .C(_1237_),
    .D(_1243_),
    .X(_1322_));
 sky130_fd_sc_hd__inv_1 _3554_ (.A(_1206_),
    .Y(_1323_));
 sky130_fd_sc_hd__o21bai_1 _3555_ (.A1(_1242_),
    .A2(_1241_),
    .B1_N(_1589_),
    .Y(_1324_));
 sky130_fd_sc_hd__a221oi_2 _3556_ (.A1(_1323_),
    .A2(_1271_),
    .B1(_1324_),
    .B2(_1581_),
    .C1(_1583_),
    .Y(_1325_));
 sky130_fd_sc_hd__o211ai_1 _3557_ (.A1(_1284_),
    .A2(_1270_),
    .B1(_1241_),
    .C1(_1240_),
    .Y(_1326_));
 sky130_fd_sc_hd__xnor2_1 _3558_ (.A(_1242_),
    .B(_1326_),
    .Y(_1327_));
 sky130_fd_sc_hd__a211oi_4 _3559_ (.A1(_1244_),
    .A2(_1322_),
    .B1(_1325_),
    .C1(_1327_),
    .Y(_1328_));
 sky130_fd_sc_hd__and3_1 _3560_ (.A(_1233_),
    .B(_1248_),
    .C(_1328_),
    .X(_1329_));
 sky130_fd_sc_hd__buf_8 _3561_ (.A(_1329_),
    .X(_1330_));
 sky130_fd_sc_hd__a22oi_4 _3562_ (.A1(_1293_),
    .A2(_1317_),
    .B1(_1321_),
    .B2(_1330_),
    .Y(_1331_));
 sky130_fd_sc_hd__mux4_1 _3563_ (.A0(net30),
    .A1(net32),
    .A2(net62),
    .A3(net64),
    .S0(_1294_),
    .S1(_1316_),
    .X(_1332_));
 sky130_fd_sc_hd__nand2_1 _3564_ (.A(net64),
    .B(_1319_),
    .Y(_1333_));
 sky130_fd_sc_hd__o21ai_1 _3565_ (.A1(_1634_),
    .A2(_1319_),
    .B1(_1333_),
    .Y(_1334_));
 sky130_fd_sc_hd__a22oi_4 _3566_ (.A1(_1293_),
    .A2(_1332_),
    .B1(_1334_),
    .B2(_1330_),
    .Y(_1335_));
 sky130_fd_sc_hd__a21o_4 _3567_ (.A1(_1233_),
    .A2(_1248_),
    .B1(_1292_),
    .X(_1336_));
 sky130_fd_sc_hd__nor2_8 _3568_ (.A(_1336_),
    .B(_1316_),
    .Y(_1337_));
 sky130_fd_sc_hd__mux2_1 _3569_ (.A0(net4),
    .A1(net6),
    .S(_1294_),
    .X(_1338_));
 sky130_fd_sc_hd__nand2_1 _3570_ (.A(net38),
    .B(_1318_),
    .Y(_1339_));
 sky130_fd_sc_hd__o21ai_1 _3571_ (.A1(_1655_),
    .A2(_1319_),
    .B1(_1339_),
    .Y(_1340_));
 sky130_fd_sc_hd__a21o_4 _3572_ (.A1(_1192_),
    .A2(_1201_),
    .B1(_1189_),
    .X(_1341_));
 sky130_fd_sc_hd__a41o_4 _3573_ (.A1(_1297_),
    .A2(_1302_),
    .A3(_1303_),
    .A4(_1304_),
    .B1(_1314_),
    .X(_1342_));
 sky130_fd_sc_hd__a2111oi_4 _3574_ (.A1(_1233_),
    .A2(_1248_),
    .B1(_1341_),
    .C1(_1292_),
    .D1(_1342_),
    .Y(_1343_));
 sky130_fd_sc_hd__clkbuf_4 _3575_ (.A(_1294_),
    .X(_1344_));
 sky130_fd_sc_hd__mux2i_1 _3576_ (.A0(net36),
    .A1(net38),
    .S(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hd__nor4_1 _3577_ (.A(a_exp_larger),
    .B(_1292_),
    .C(_1343_),
    .D(_1345_),
    .Y(_1346_));
 sky130_fd_sc_hd__a221oi_4 _3578_ (.A1(_1337_),
    .A2(_1338_),
    .B1(_1340_),
    .B2(_1330_),
    .C1(_1346_),
    .Y(_1347_));
 sky130_fd_sc_hd__mux2_1 _3579_ (.A0(net31),
    .A1(net33),
    .S(_1344_),
    .X(_1348_));
 sky130_fd_sc_hd__nand2_1 _3580_ (.A(net65),
    .B(_1318_),
    .Y(_1349_));
 sky130_fd_sc_hd__o21ai_1 _3581_ (.A1(_1631_),
    .A2(_1319_),
    .B1(_1349_),
    .Y(_1350_));
 sky130_fd_sc_hd__mux2i_1 _3582_ (.A0(net63),
    .A1(net65),
    .S(_1344_),
    .Y(_1351_));
 sky130_fd_sc_hd__nor4_1 _3583_ (.A(a_exp_larger),
    .B(_1292_),
    .C(_1343_),
    .D(_1351_),
    .Y(_1352_));
 sky130_fd_sc_hd__a221oi_4 _3584_ (.A1(_1337_),
    .A2(_1348_),
    .B1(_1350_),
    .B2(_1330_),
    .C1(_1352_),
    .Y(_1353_));
 sky130_fd_sc_hd__nor2b_1 _3585_ (.A(_1567_),
    .B_N(_1269_),
    .Y(_1354_));
 sky130_fd_sc_hd__nor2b_1 _3586_ (.A(_1269_),
    .B_N(_1567_),
    .Y(_1355_));
 sky130_fd_sc_hd__fa_1 _3587_ (.A(_1565_),
    .B(net50),
    .CIN(_1566_),
    .COUT(_1567_),
    .SUM(_1568_));
 sky130_fd_sc_hd__fa_1 _3588_ (.A(net18),
    .B(_1569_),
    .CIN(_1570_),
    .COUT(_1571_),
    .SUM(_1572_));
 sky130_fd_sc_hd__fa_1 _3589_ (.A(\result_exp_stage2[1] ),
    .B(_1573_),
    .CIN(_1574_),
    .COUT(_1575_),
    .SUM(_1576_));
 sky130_fd_sc_hd__ha_1 _3590_ (.A(net26),
    .B(net58),
    .COUT(_1577_),
    .SUM(_1578_));
 sky130_fd_sc_hd__ha_2 _3591_ (.A(_1579_),
    .B(net57),
    .COUT(_1580_),
    .SUM(_1581_));
 sky130_fd_sc_hd__ha_1 _3592_ (.A(net25),
    .B(_1582_),
    .COUT(_1583_),
    .SUM(_1584_));
 sky130_fd_sc_hd__ha_1 _3593_ (.A(_1585_),
    .B(net55),
    .COUT(_1586_),
    .SUM(_1587_));
 sky130_fd_sc_hd__ha_1 _3594_ (.A(net23),
    .B(_1588_),
    .COUT(_1589_),
    .SUM(_1590_));
 sky130_fd_sc_hd__ha_2 _3595_ (.A(_1591_),
    .B(net54),
    .COUT(_1592_),
    .SUM(_1593_));
 sky130_fd_sc_hd__ha_1 _3596_ (.A(net22),
    .B(_1594_),
    .COUT(_1595_),
    .SUM(_1596_));
 sky130_fd_sc_hd__ha_1 _3597_ (.A(_1597_),
    .B(net53),
    .COUT(_1598_),
    .SUM(_1599_));
 sky130_fd_sc_hd__ha_1 _3598_ (.A(net21),
    .B(_1600_),
    .COUT(_1601_),
    .SUM(_1602_));
 sky130_fd_sc_hd__ha_1 _3599_ (.A(_1603_),
    .B(net52),
    .COUT(_1604_),
    .SUM(_1605_));
 sky130_fd_sc_hd__ha_1 _3600_ (.A(net20),
    .B(_1606_),
    .COUT(_1607_),
    .SUM(_1608_));
 sky130_fd_sc_hd__ha_1 _3601_ (.A(_1609_),
    .B(net51),
    .COUT(_1610_),
    .SUM(_1611_));
 sky130_fd_sc_hd__ha_1 _3602_ (.A(net19),
    .B(_1612_),
    .COUT(_1613_),
    .SUM(_1614_));
 sky130_fd_sc_hd__ha_1 _3603_ (.A(_1565_),
    .B(net50),
    .COUT(_1615_),
    .SUM(_1616_));
 sky130_fd_sc_hd__ha_1 _3604_ (.A(net18),
    .B(_1569_),
    .COUT(_1617_),
    .SUM(_1618_));
 sky130_fd_sc_hd__ha_1 _3605_ (.A(net13),
    .B(_1619_),
    .COUT(_1620_),
    .SUM(_1621_));
 sky130_fd_sc_hd__ha_1 _3606_ (.A(_1622_),
    .B(net34),
    .COUT(_1623_),
    .SUM(_1624_));
 sky130_fd_sc_hd__ha_1 _3607_ (.A(net27),
    .B(_1625_),
    .COUT(_1626_),
    .SUM(_1627_));
 sky130_fd_sc_hd__ha_1 _3608_ (.A(net24),
    .B(_1628_),
    .COUT(_1629_),
    .SUM(_1630_));
 sky130_fd_sc_hd__ha_1 _3609_ (.A(net31),
    .B(_1631_),
    .COUT(_1632_),
    .SUM(_1633_));
 sky130_fd_sc_hd__ha_1 _3610_ (.A(net30),
    .B(_1634_),
    .COUT(_1635_),
    .SUM(_1636_));
 sky130_fd_sc_hd__ha_1 _3611_ (.A(net29),
    .B(_1637_),
    .COUT(_1638_),
    .SUM(_1639_));
 sky130_fd_sc_hd__ha_1 _3612_ (.A(net28),
    .B(_1640_),
    .COUT(_1641_),
    .SUM(_1642_));
 sky130_fd_sc_hd__ha_1 _3613_ (.A(net8),
    .B(_1643_),
    .COUT(_1644_),
    .SUM(_1645_));
 sky130_fd_sc_hd__ha_1 _3614_ (.A(net7),
    .B(_1646_),
    .COUT(_1647_),
    .SUM(_1648_));
 sky130_fd_sc_hd__ha_1 _3615_ (.A(net6),
    .B(_1649_),
    .COUT(_1650_),
    .SUM(_1651_));
 sky130_fd_sc_hd__ha_1 _3616_ (.A(net5),
    .B(_1652_),
    .COUT(_1653_),
    .SUM(_1654_));
 sky130_fd_sc_hd__ha_1 _3617_ (.A(net4),
    .B(_1655_),
    .COUT(_1656_),
    .SUM(_1657_));
 sky130_fd_sc_hd__ha_1 _3618_ (.A(net3),
    .B(_1658_),
    .COUT(_1659_),
    .SUM(_1660_));
 sky130_fd_sc_hd__ha_1 _3619_ (.A(net33),
    .B(_1661_),
    .COUT(_1662_),
    .SUM(_1663_));
 sky130_fd_sc_hd__ha_1 _3620_ (.A(net32),
    .B(_1664_),
    .COUT(_1665_),
    .SUM(_1666_));
 sky130_fd_sc_hd__ha_1 _3621_ (.A(net12),
    .B(_1667_),
    .COUT(_1668_),
    .SUM(_1669_));
 sky130_fd_sc_hd__ha_1 _3622_ (.A(net11),
    .B(_1670_),
    .COUT(_1671_),
    .SUM(_1672_));
 sky130_fd_sc_hd__ha_1 _3623_ (.A(net10),
    .B(_1673_),
    .COUT(_1674_),
    .SUM(_1675_));
 sky130_fd_sc_hd__ha_1 _3624_ (.A(net9),
    .B(_1676_),
    .COUT(_1677_),
    .SUM(_1678_));
 sky130_fd_sc_hd__ha_1 _3625_ (.A(net16),
    .B(_1679_),
    .COUT(_1680_),
    .SUM(_1681_));
 sky130_fd_sc_hd__ha_1 _3626_ (.A(net15),
    .B(_1682_),
    .COUT(_1683_),
    .SUM(_1684_));
 sky130_fd_sc_hd__ha_1 _3627_ (.A(net14),
    .B(_1685_),
    .COUT(_1686_),
    .SUM(_1687_));
 sky130_fd_sc_hd__ha_1 _3628_ (.A(_1688_),
    .B(net49),
    .COUT(_1689_),
    .SUM(_1690_));
 sky130_fd_sc_hd__ha_1 _3629_ (.A(net17),
    .B(_1691_),
    .COUT(_1692_),
    .SUM(_1693_));
 sky130_fd_sc_hd__ha_1 _3630_ (.A(_1694_),
    .B(_1695_),
    .COUT(_1696_),
    .SUM(_1697_));
 sky130_fd_sc_hd__ha_1 _3631_ (.A(\result_exp_stage2[2] ),
    .B(_1698_),
    .COUT(_1699_),
    .SUM(_1700_));
 sky130_fd_sc_hd__ha_1 _3632_ (.A(_1701_),
    .B(_1702_),
    .COUT(_1703_),
    .SUM(_1704_));
 sky130_fd_sc_hd__ha_1 _3633_ (.A(\result_exp_stage2[1] ),
    .B(_1574_),
    .COUT(_1705_),
    .SUM(_1706_));
 sky130_fd_sc_hd__ha_1 _3634_ (.A(_1707_),
    .B(_1708_),
    .COUT(_1709_),
    .SUM(_1710_));
 sky130_fd_sc_hd__ha_1 _3635_ (.A(\result_exp_stage2[0] ),
    .B(_1711_),
    .COUT(_1712_),
    .SUM(_1713_));
 sky130_fd_sc_hd__ha_2 _3636_ (.A(_1707_),
    .B(_1701_),
    .COUT(_1714_),
    .SUM(_1715_));
 sky130_fd_sc_hd__ha_1 _3637_ (.A(_1707_),
    .B(\result_exp_stage2[1] ),
    .COUT(_1716_),
    .SUM(_1717_));
 sky130_fd_sc_hd__ha_1 _3638_ (.A(\result_exp_stage2[0] ),
    .B(\result_exp_stage2[1] ),
    .COUT(_1718_),
    .SUM(_1719_));
 sky130_fd_sc_hd__ha_1 _3639_ (.A(_1720_),
    .B(\aligned_b_mant[2] ),
    .COUT(_1721_),
    .SUM(_1722_));
 sky130_fd_sc_hd__ha_1 _3640_ (.A(\aligned_a_mant[2] ),
    .B(_1723_),
    .COUT(_1724_),
    .SUM(_1725_));
 sky130_fd_sc_hd__ha_1 _3641_ (.A(\aligned_a_mant[2] ),
    .B(\aligned_b_mant[2] ),
    .COUT(_1726_),
    .SUM(_1727_));
 sky130_fd_sc_hd__ha_1 _3642_ (.A(_1728_),
    .B(\aligned_b_mant[1] ),
    .COUT(_1729_),
    .SUM(_1730_));
 sky130_fd_sc_hd__ha_1 _3643_ (.A(\aligned_a_mant[1] ),
    .B(_1731_),
    .COUT(_1732_),
    .SUM(_1733_));
 sky130_fd_sc_hd__ha_1 _3644_ (.A(\aligned_a_mant[1] ),
    .B(\aligned_b_mant[1] ),
    .COUT(_1734_),
    .SUM(_1735_));
 sky130_fd_sc_hd__ha_2 _3645_ (.A(_1736_),
    .B(\aligned_b_mant[3] ),
    .COUT(_1737_),
    .SUM(_1738_));
 sky130_fd_sc_hd__ha_1 _3646_ (.A(\aligned_a_mant[3] ),
    .B(_1739_),
    .COUT(_1740_),
    .SUM(_1741_));
 sky130_fd_sc_hd__ha_1 _3647_ (.A(\aligned_a_mant[3] ),
    .B(\aligned_b_mant[3] ),
    .COUT(_1742_),
    .SUM(_1743_));
 sky130_fd_sc_hd__ha_1 _3648_ (.A(_1744_),
    .B(\aligned_b_mant[4] ),
    .COUT(_1745_),
    .SUM(_1746_));
 sky130_fd_sc_hd__ha_1 _3649_ (.A(\aligned_a_mant[4] ),
    .B(_1747_),
    .COUT(_1748_),
    .SUM(_1749_));
 sky130_fd_sc_hd__ha_1 _3650_ (.A(\aligned_a_mant[4] ),
    .B(\aligned_b_mant[4] ),
    .COUT(_1750_),
    .SUM(_1751_));
 sky130_fd_sc_hd__ha_1 _3651_ (.A(_1752_),
    .B(\aligned_b_mant[5] ),
    .COUT(_1753_),
    .SUM(_1754_));
 sky130_fd_sc_hd__ha_1 _3652_ (.A(\aligned_a_mant[5] ),
    .B(_1755_),
    .COUT(_1756_),
    .SUM(_1757_));
 sky130_fd_sc_hd__ha_1 _3653_ (.A(\aligned_a_mant[5] ),
    .B(\aligned_b_mant[5] ),
    .COUT(_1758_),
    .SUM(_1759_));
 sky130_fd_sc_hd__ha_1 _3654_ (.A(_1760_),
    .B(\aligned_b_mant[6] ),
    .COUT(_1761_),
    .SUM(_1762_));
 sky130_fd_sc_hd__ha_1 _3655_ (.A(\aligned_a_mant[6] ),
    .B(_1763_),
    .COUT(_1764_),
    .SUM(_1765_));
 sky130_fd_sc_hd__ha_1 _3656_ (.A(\aligned_a_mant[6] ),
    .B(\aligned_b_mant[6] ),
    .COUT(_1766_),
    .SUM(_1767_));
 sky130_fd_sc_hd__ha_2 _3657_ (.A(_1768_),
    .B(\aligned_b_mant[7] ),
    .COUT(_1769_),
    .SUM(_1770_));
 sky130_fd_sc_hd__ha_1 _3658_ (.A(\aligned_a_mant[7] ),
    .B(_1771_),
    .COUT(_1772_),
    .SUM(_1773_));
 sky130_fd_sc_hd__ha_1 _3659_ (.A(\aligned_a_mant[7] ),
    .B(\aligned_b_mant[7] ),
    .COUT(_1774_),
    .SUM(_1775_));
 sky130_fd_sc_hd__ha_1 _3660_ (.A(_1776_),
    .B(\aligned_b_mant[8] ),
    .COUT(_1777_),
    .SUM(_1778_));
 sky130_fd_sc_hd__ha_2 _3661_ (.A(\aligned_a_mant[8] ),
    .B(_1779_),
    .COUT(_1780_),
    .SUM(_1781_));
 sky130_fd_sc_hd__ha_1 _3662_ (.A(\aligned_a_mant[8] ),
    .B(\aligned_b_mant[8] ),
    .COUT(_1782_),
    .SUM(_1783_));
 sky130_fd_sc_hd__ha_1 _3663_ (.A(_1784_),
    .B(\aligned_b_mant[9] ),
    .COUT(_1785_),
    .SUM(_1786_));
 sky130_fd_sc_hd__ha_1 _3664_ (.A(\aligned_a_mant[9] ),
    .B(_1787_),
    .COUT(_1788_),
    .SUM(_1789_));
 sky130_fd_sc_hd__ha_1 _3665_ (.A(\aligned_a_mant[9] ),
    .B(\aligned_b_mant[9] ),
    .COUT(_1790_),
    .SUM(_1791_));
 sky130_fd_sc_hd__ha_1 _3666_ (.A(_1792_),
    .B(\aligned_b_mant[10] ),
    .COUT(_1793_),
    .SUM(_1794_));
 sky130_fd_sc_hd__ha_1 _3667_ (.A(\aligned_a_mant[10] ),
    .B(_1795_),
    .COUT(_1796_),
    .SUM(_1797_));
 sky130_fd_sc_hd__ha_1 _3668_ (.A(\aligned_a_mant[10] ),
    .B(\aligned_b_mant[10] ),
    .COUT(_1798_),
    .SUM(_1799_));
 sky130_fd_sc_hd__ha_1 _3669_ (.A(_1800_),
    .B(\aligned_b_mant[11] ),
    .COUT(_1801_),
    .SUM(_1802_));
 sky130_fd_sc_hd__ha_1 _3670_ (.A(\aligned_a_mant[11] ),
    .B(_1803_),
    .COUT(_1804_),
    .SUM(_1805_));
 sky130_fd_sc_hd__ha_1 _3671_ (.A(\aligned_a_mant[11] ),
    .B(\aligned_b_mant[11] ),
    .COUT(_1806_),
    .SUM(_1807_));
 sky130_fd_sc_hd__ha_1 _3672_ (.A(_1808_),
    .B(\aligned_b_mant[12] ),
    .COUT(_1809_),
    .SUM(_1810_));
 sky130_fd_sc_hd__ha_1 _3673_ (.A(\aligned_a_mant[12] ),
    .B(_1811_),
    .COUT(_1812_),
    .SUM(_1813_));
 sky130_fd_sc_hd__ha_1 _3674_ (.A(\aligned_a_mant[12] ),
    .B(\aligned_b_mant[12] ),
    .COUT(_1814_),
    .SUM(_1815_));
 sky130_fd_sc_hd__ha_1 _3675_ (.A(_1816_),
    .B(\aligned_b_mant[13] ),
    .COUT(_1817_),
    .SUM(_1818_));
 sky130_fd_sc_hd__ha_1 _3676_ (.A(\aligned_a_mant[13] ),
    .B(_1819_),
    .COUT(_1820_),
    .SUM(_1821_));
 sky130_fd_sc_hd__ha_1 _3677_ (.A(\aligned_a_mant[13] ),
    .B(\aligned_b_mant[13] ),
    .COUT(_1822_),
    .SUM(_1823_));
 sky130_fd_sc_hd__ha_1 _3678_ (.A(_1824_),
    .B(\aligned_b_mant[14] ),
    .COUT(_1825_),
    .SUM(_1826_));
 sky130_fd_sc_hd__ha_1 _3679_ (.A(\aligned_a_mant[14] ),
    .B(_1827_),
    .COUT(_1828_),
    .SUM(_1829_));
 sky130_fd_sc_hd__ha_1 _3680_ (.A(\aligned_a_mant[14] ),
    .B(\aligned_b_mant[14] ),
    .COUT(_1830_),
    .SUM(_1831_));
 sky130_fd_sc_hd__ha_1 _3681_ (.A(_1832_),
    .B(\aligned_b_mant[15] ),
    .COUT(_1833_),
    .SUM(_1834_));
 sky130_fd_sc_hd__ha_1 _3682_ (.A(\aligned_a_mant[15] ),
    .B(_1835_),
    .COUT(_1836_),
    .SUM(_1837_));
 sky130_fd_sc_hd__ha_1 _3683_ (.A(\aligned_a_mant[15] ),
    .B(\aligned_b_mant[15] ),
    .COUT(_1838_),
    .SUM(_1839_));
 sky130_fd_sc_hd__ha_1 _3684_ (.A(_1840_),
    .B(\aligned_b_mant[16] ),
    .COUT(_1841_),
    .SUM(_1842_));
 sky130_fd_sc_hd__ha_1 _3685_ (.A(\aligned_a_mant[16] ),
    .B(_1843_),
    .COUT(_1844_),
    .SUM(_1845_));
 sky130_fd_sc_hd__ha_1 _3686_ (.A(\aligned_a_mant[16] ),
    .B(\aligned_b_mant[16] ),
    .COUT(_1846_),
    .SUM(_1847_));
 sky130_fd_sc_hd__ha_1 _3687_ (.A(_1848_),
    .B(\aligned_b_mant[17] ),
    .COUT(_1849_),
    .SUM(_1850_));
 sky130_fd_sc_hd__ha_1 _3688_ (.A(\aligned_a_mant[17] ),
    .B(_1851_),
    .COUT(_1852_),
    .SUM(_1853_));
 sky130_fd_sc_hd__ha_1 _3689_ (.A(\aligned_a_mant[17] ),
    .B(\aligned_b_mant[17] ),
    .COUT(_1854_),
    .SUM(_1855_));
 sky130_fd_sc_hd__ha_1 _3690_ (.A(_1856_),
    .B(\aligned_b_mant[18] ),
    .COUT(_1857_),
    .SUM(_1858_));
 sky130_fd_sc_hd__ha_1 _3691_ (.A(\aligned_a_mant[18] ),
    .B(_1859_),
    .COUT(_1860_),
    .SUM(_1861_));
 sky130_fd_sc_hd__ha_1 _3692_ (.A(\aligned_a_mant[18] ),
    .B(\aligned_b_mant[18] ),
    .COUT(_1862_),
    .SUM(_1863_));
 sky130_fd_sc_hd__ha_1 _3693_ (.A(_1864_),
    .B(\aligned_b_mant[19] ),
    .COUT(_1865_),
    .SUM(_1866_));
 sky130_fd_sc_hd__ha_1 _3694_ (.A(\aligned_a_mant[19] ),
    .B(_1867_),
    .COUT(_1868_),
    .SUM(_1869_));
 sky130_fd_sc_hd__ha_1 _3695_ (.A(\aligned_a_mant[19] ),
    .B(\aligned_b_mant[19] ),
    .COUT(_1870_),
    .SUM(_1871_));
 sky130_fd_sc_hd__ha_2 _3696_ (.A(_1872_),
    .B(\aligned_b_mant[20] ),
    .COUT(_1873_),
    .SUM(_1874_));
 sky130_fd_sc_hd__ha_1 _3697_ (.A(\aligned_a_mant[20] ),
    .B(_1875_),
    .COUT(_1876_),
    .SUM(_1877_));
 sky130_fd_sc_hd__ha_1 _3698_ (.A(\aligned_a_mant[20] ),
    .B(\aligned_b_mant[20] ),
    .COUT(_1878_),
    .SUM(_1879_));
 sky130_fd_sc_hd__ha_1 _3699_ (.A(_1880_),
    .B(\aligned_b_mant[21] ),
    .COUT(_1881_),
    .SUM(_1882_));
 sky130_fd_sc_hd__ha_1 _3700_ (.A(\aligned_a_mant[21] ),
    .B(_1883_),
    .COUT(_1884_),
    .SUM(_1885_));
 sky130_fd_sc_hd__ha_1 _3701_ (.A(\aligned_a_mant[21] ),
    .B(\aligned_b_mant[21] ),
    .COUT(_1886_),
    .SUM(_1887_));
 sky130_fd_sc_hd__ha_1 _3702_ (.A(_1888_),
    .B(\aligned_b_mant[22] ),
    .COUT(_1889_),
    .SUM(_1890_));
 sky130_fd_sc_hd__ha_1 _3703_ (.A(\aligned_a_mant[22] ),
    .B(_1891_),
    .COUT(_1892_),
    .SUM(_1893_));
 sky130_fd_sc_hd__ha_1 _3704_ (.A(\aligned_a_mant[22] ),
    .B(\aligned_b_mant[22] ),
    .COUT(_1894_),
    .SUM(_1895_));
 sky130_fd_sc_hd__ha_1 _3705_ (.A(_1896_),
    .B(\aligned_b_mant[23] ),
    .COUT(_1897_),
    .SUM(_1898_));
 sky130_fd_sc_hd__ha_1 _3706_ (.A(\aligned_a_mant[23] ),
    .B(_1899_),
    .COUT(_1900_),
    .SUM(_1901_));
 sky130_fd_sc_hd__ha_1 _3707_ (.A(\aligned_a_mant[23] ),
    .B(\aligned_b_mant[23] ),
    .COUT(_1902_),
    .SUM(_1903_));
 sky130_fd_sc_hd__ha_1 _3708_ (.A(_1904_),
    .B(\aligned_b_mant[24] ),
    .COUT(_1905_),
    .SUM(_1906_));
 sky130_fd_sc_hd__ha_1 _3709_ (.A(\aligned_a_mant[24] ),
    .B(_1907_),
    .COUT(_1908_),
    .SUM(_1909_));
 sky130_fd_sc_hd__ha_1 _3710_ (.A(\aligned_a_mant[24] ),
    .B(\aligned_b_mant[24] ),
    .COUT(_1910_),
    .SUM(_1911_));
 sky130_fd_sc_hd__ha_1 _3711_ (.A(_1912_),
    .B(\aligned_b_mant[25] ),
    .COUT(_1913_),
    .SUM(_1914_));
 sky130_fd_sc_hd__ha_1 _3712_ (.A(\aligned_a_mant[25] ),
    .B(_1915_),
    .COUT(_1916_),
    .SUM(_1917_));
 sky130_fd_sc_hd__ha_1 _3713_ (.A(\aligned_a_mant[25] ),
    .B(\aligned_b_mant[25] ),
    .COUT(_1918_),
    .SUM(_1919_));
 sky130_fd_sc_hd__dfrtp_4 \a_sign_stage1$_DFF_PN0_  (.D(net26),
    .Q(a_sign_stage1),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \add_result[10]$_DFF_PN0_  (.D(_0000_),
    .Q(\add_result[10] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \add_result[11]$_DFF_PN0_  (.D(_0001_),
    .Q(\add_result[11] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \add_result[12]$_DFF_PN0_  (.D(_0002_),
    .Q(\add_result[12] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \add_result[13]$_DFF_PN0_  (.D(_0003_),
    .Q(\add_result[13] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \add_result[14]$_DFF_PN0_  (.D(_0004_),
    .Q(\add_result[14] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \add_result[15]$_DFF_PN0_  (.D(_0005_),
    .Q(\add_result[15] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \add_result[16]$_DFF_PN0_  (.D(_0006_),
    .Q(\add_result[16] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \add_result[17]$_DFF_PN0_  (.D(_0007_),
    .Q(\add_result[17] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \add_result[18]$_DFF_PN0_  (.D(_0008_),
    .Q(\add_result[18] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \add_result[19]$_DFF_PN0_  (.D(_0009_),
    .Q(\add_result[19] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \add_result[20]$_DFF_PN0_  (.D(_0010_),
    .Q(\add_result[20] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \add_result[21]$_DFF_PN0_  (.D(_0011_),
    .Q(\add_result[21] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \add_result[22]$_DFF_PN0_  (.D(_0012_),
    .Q(\add_result[22] ),
    .RESET_B(net1),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \add_result[23]$_DFF_PN0_  (.D(_0013_),
    .Q(\add_result[23] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \add_result[24]$_DFF_PN0_  (.D(_0014_),
    .Q(\add_result[24] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \add_result[25]$_DFF_PN0_  (.D(_0015_),
    .Q(\add_result[25] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \add_result[26]$_DFF_PN0_  (.D(_0016_),
    .Q(\add_result[26] ),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \add_result[2]$_DFF_PN0_  (.D(_0017_),
    .Q(\add_result[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \add_result[3]$_DFF_PN0_  (.D(_0018_),
    .Q(\add_result[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \add_result[4]$_DFF_PN0_  (.D(_0019_),
    .Q(\add_result[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \add_result[5]$_DFF_PN0_  (.D(_0020_),
    .Q(\add_result[5] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \add_result[6]$_DFF_PN0_  (.D(_0021_),
    .Q(\add_result[6] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \add_result[7]$_DFF_PN0_  (.D(_0022_),
    .Q(\add_result[7] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \add_result[8]$_DFF_PN0_  (.D(_0023_),
    .Q(\add_result[8] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \add_result[9]$_DFF_PN0_  (.D(_0024_),
    .Q(\add_result[9] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[0]$_DFF_PN0_  (.D(_0025_),
    .Q(\aligned_a_mant[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[10]$_DFF_PN0_  (.D(_0026_),
    .Q(\aligned_a_mant[10] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[11]$_DFF_PN0_  (.D(_0027_),
    .Q(\aligned_a_mant[11] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[12]$_DFF_PN0_  (.D(_0028_),
    .Q(\aligned_a_mant[12] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[13]$_DFF_PN0_  (.D(_0029_),
    .Q(\aligned_a_mant[13] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[14]$_DFF_PN0_  (.D(_0030_),
    .Q(\aligned_a_mant[14] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[15]$_DFF_PN0_  (.D(_0031_),
    .Q(\aligned_a_mant[15] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[16]$_DFF_PN0_  (.D(_0032_),
    .Q(\aligned_a_mant[16] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[17]$_DFF_PN0_  (.D(_0033_),
    .Q(\aligned_a_mant[17] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[18]$_DFF_PN0_  (.D(_0034_),
    .Q(\aligned_a_mant[18] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[19]$_DFF_PN0_  (.D(_0035_),
    .Q(\aligned_a_mant[19] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[1]$_DFF_PN0_  (.D(_0036_),
    .Q(\aligned_a_mant[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[20]$_DFF_PN0_  (.D(_0037_),
    .Q(\aligned_a_mant[20] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[21]$_DFF_PN0_  (.D(_0038_),
    .Q(\aligned_a_mant[21] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[22]$_DFF_PN0_  (.D(_0039_),
    .Q(\aligned_a_mant[22] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[23]$_DFF_PN0_  (.D(_0040_),
    .Q(\aligned_a_mant[23] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[24]$_DFF_PN0_  (.D(_0041_),
    .Q(\aligned_a_mant[24] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[25]$_DFF_PN0_  (.D(_0042_),
    .Q(\aligned_a_mant[25] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[2]$_DFF_PN0_  (.D(_0043_),
    .Q(\aligned_a_mant[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[3]$_DFF_PN0_  (.D(_0044_),
    .Q(\aligned_a_mant[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[4]$_DFF_PN0_  (.D(_0045_),
    .Q(\aligned_a_mant[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[5]$_DFF_PN0_  (.D(_0046_),
    .Q(\aligned_a_mant[5] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[6]$_DFF_PN0_  (.D(_0047_),
    .Q(\aligned_a_mant[6] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[7]$_DFF_PN0_  (.D(_0048_),
    .Q(\aligned_a_mant[7] ),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[8]$_DFF_PN0_  (.D(_0049_),
    .Q(\aligned_a_mant[8] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_a_mant[9]$_DFF_PN0_  (.D(_0050_),
    .Q(\aligned_a_mant[9] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[0]$_DFF_PN0_  (.D(_0051_),
    .Q(\aligned_b_mant[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[10]$_DFF_PN0_  (.D(_0052_),
    .Q(\aligned_b_mant[10] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[11]$_DFF_PN0_  (.D(_0053_),
    .Q(\aligned_b_mant[11] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[12]$_DFF_PN0_  (.D(_0054_),
    .Q(\aligned_b_mant[12] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[13]$_DFF_PN0_  (.D(_0055_),
    .Q(\aligned_b_mant[13] ),
    .RESET_B(net1),
    .CLK(clknet_4_9_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[14]$_DFF_PN0_  (.D(_0056_),
    .Q(\aligned_b_mant[14] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[15]$_DFF_PN0_  (.D(_0057_),
    .Q(\aligned_b_mant[15] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[16]$_DFF_PN0_  (.D(_0058_),
    .Q(\aligned_b_mant[16] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[17]$_DFF_PN0_  (.D(_0059_),
    .Q(\aligned_b_mant[17] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[18]$_DFF_PN0_  (.D(_0060_),
    .Q(\aligned_b_mant[18] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[19]$_DFF_PN0_  (.D(_0061_),
    .Q(\aligned_b_mant[19] ),
    .RESET_B(net1),
    .CLK(clknet_4_8_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[1]$_DFF_PN0_  (.D(_0062_),
    .Q(\aligned_b_mant[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[20]$_DFF_PN0_  (.D(_0063_),
    .Q(\aligned_b_mant[20] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[21]$_DFF_PN0_  (.D(_0064_),
    .Q(\aligned_b_mant[21] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[22]$_DFF_PN0_  (.D(_0065_),
    .Q(\aligned_b_mant[22] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[23]$_DFF_PN0_  (.D(_0066_),
    .Q(\aligned_b_mant[23] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[24]$_DFF_PN0_  (.D(_0067_),
    .Q(\aligned_b_mant[24] ),
    .RESET_B(net1),
    .CLK(clknet_4_2_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[25]$_DFF_PN0_  (.D(_0068_),
    .Q(\aligned_b_mant[25] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[2]$_DFF_PN0_  (.D(_0069_),
    .Q(\aligned_b_mant[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[3]$_DFF_PN0_  (.D(_0070_),
    .Q(\aligned_b_mant[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[4]$_DFF_PN0_  (.D(_0071_),
    .Q(\aligned_b_mant[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[5]$_DFF_PN0_  (.D(_0072_),
    .Q(\aligned_b_mant[5] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[6]$_DFF_PN0_  (.D(_0073_),
    .Q(\aligned_b_mant[6] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[7]$_DFF_PN0_  (.D(_0074_),
    .Q(\aligned_b_mant[7] ),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[8]$_DFF_PN0_  (.D(_0075_),
    .Q(\aligned_b_mant[8] ),
    .RESET_B(net1),
    .CLK(clknet_4_11_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \aligned_b_mant[9]$_DFF_PN0_  (.D(_0076_),
    .Q(\aligned_b_mant[9] ),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \b_sign_stage1$_DFF_PN0_  (.D(net58),
    .Q(b_sign_stage1),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_exp[0]$_DFFE_PP_  (.D(_0077_),
    .DE(net66),
    .Q(\final_exp[0] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_exp[1]$_DFFE_PP_  (.D(_0078_),
    .DE(net66),
    .Q(\final_exp[1] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_exp[2]$_DFFE_PP_  (.D(_0079_),
    .DE(net66),
    .Q(\final_exp[2] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_exp[3]$_DFFE_PP_  (.D(_0080_),
    .DE(net66),
    .Q(\final_exp[3] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_exp[4]$_DFFE_PP_  (.D(_0081_),
    .DE(net66),
    .Q(\final_exp[4] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_exp[5]$_DFFE_PP_  (.D(_0082_),
    .DE(net66),
    .Q(\final_exp[5] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_exp[6]$_DFFE_PP_  (.D(_0083_),
    .DE(net66),
    .Q(\final_exp[6] ),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_exp[7]$_DFFE_PP_  (.D(_0084_),
    .DE(net66),
    .Q(\final_exp[7] ),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[0]$_DFFE_PP_  (.D(_0085_),
    .DE(net66),
    .Q(\final_mant[0] ),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[10]$_DFFE_PP_  (.D(_0086_),
    .DE(net66),
    .Q(\final_mant[10] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[11]$_DFFE_PP_  (.D(_0087_),
    .DE(net66),
    .Q(\final_mant[11] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[12]$_DFFE_PP_  (.D(_0088_),
    .DE(net66),
    .Q(\final_mant[12] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[13]$_DFFE_PP_  (.D(_0089_),
    .DE(net66),
    .Q(\final_mant[13] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[14]$_DFFE_PP_  (.D(_0090_),
    .DE(net66),
    .Q(\final_mant[14] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[15]$_DFFE_PP_  (.D(_0091_),
    .DE(net66),
    .Q(\final_mant[15] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[16]$_DFFE_PP_  (.D(_0092_),
    .DE(net66),
    .Q(\final_mant[16] ),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[17]$_DFFE_PP_  (.D(_0093_),
    .DE(net66),
    .Q(\final_mant[17] ),
    .CLK(clknet_4_12_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[18]$_DFFE_PP_  (.D(_0094_),
    .DE(net66),
    .Q(\final_mant[18] ),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[19]$_DFFE_PP_  (.D(_0095_),
    .DE(net66),
    .Q(\final_mant[19] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[1]$_DFFE_PP_  (.D(_0096_),
    .DE(net66),
    .Q(\final_mant[1] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[20]$_DFFE_PP_  (.D(_0097_),
    .DE(net66),
    .Q(\final_mant[20] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[21]$_DFFE_PP_  (.D(_0098_),
    .DE(net66),
    .Q(\final_mant[21] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[22]$_DFFE_PP_  (.D(_0099_),
    .DE(net66),
    .Q(\final_mant[22] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[2]$_DFFE_PP_  (.D(_0100_),
    .DE(net66),
    .Q(\final_mant[2] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[3]$_DFFE_PP_  (.D(_0101_),
    .DE(net66),
    .Q(\final_mant[3] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[4]$_DFFE_PP_  (.D(_0102_),
    .DE(net66),
    .Q(\final_mant[4] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[5]$_DFFE_PP_  (.D(_0103_),
    .DE(net66),
    .Q(\final_mant[5] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[6]$_DFFE_PP_  (.D(_0104_),
    .DE(net66),
    .Q(\final_mant[6] ),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[7]$_DFFE_PP_  (.D(_0105_),
    .DE(net66),
    .Q(\final_mant[7] ),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[8]$_DFFE_PP_  (.D(_0106_),
    .DE(net66),
    .Q(\final_mant[8] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \final_mant[9]$_DFFE_PP_  (.D(_0107_),
    .DE(net66),
    .Q(\final_mant[9] ),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \inexact$_DFF_PN0_  (.D(_0108_),
    .Q(net68),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \inexact_stage2$_DFF_PN0_  (.D(_0109_),
    .Q(inexact_stage2),
    .RESET_B(net1),
    .CLK(clknet_4_6_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \invalid_op$_DFF_PN0_  (.D(invalid_op_stage2),
    .Q(net69),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \invalid_op_stage2$_DFFE_PN0P_  (.D(_0121_),
    .Q(invalid_op_stage2),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \is_a_larger_stage1$_DFF_PN0_  (.D(a_exp_larger),
    .Q(is_a_larger_stage1),
    .RESET_B(net1),
    .CLK(clknet_4_10_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \larger_exp_stage1[0]$_DFF_PN0_  (.D(_0110_),
    .Q(\larger_exp_stage1[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \larger_exp_stage1[1]$_DFF_PN0_  (.D(_0111_),
    .Q(\larger_exp_stage1[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \larger_exp_stage1[2]$_DFF_PN0_  (.D(_0112_),
    .Q(\larger_exp_stage1[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \larger_exp_stage1[3]$_DFF_PN0_  (.D(_0113_),
    .Q(\larger_exp_stage1[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \larger_exp_stage1[4]$_DFF_PN0_  (.D(_0114_),
    .Q(\larger_exp_stage1[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \larger_exp_stage1[5]$_DFF_PN0_  (.D(_0115_),
    .Q(\larger_exp_stage1[5] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \larger_exp_stage1[6]$_DFF_PN0_  (.D(_0116_),
    .Q(\larger_exp_stage1[6] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \larger_exp_stage1[7]$_DFF_PN0_  (.D(_0117_),
    .Q(\larger_exp_stage1[7] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \overflow$_DFF_PN0_  (.D(_0118_),
    .Q(net70),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[0]$_DFF_PN0_  (.D(\final_mant[0] ),
    .Q(net71),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[10]$_DFF_PN0_  (.D(\final_mant[10] ),
    .Q(net72),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[11]$_DFF_PN0_  (.D(\final_mant[11] ),
    .Q(net73),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[12]$_DFF_PN0_  (.D(\final_mant[12] ),
    .Q(net74),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[13]$_DFF_PN0_  (.D(\final_mant[13] ),
    .Q(net75),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[14]$_DFF_PN0_  (.D(\final_mant[14] ),
    .Q(net76),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[15]$_DFF_PN0_  (.D(\final_mant[15] ),
    .Q(net77),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[16]$_DFF_PN0_  (.D(\final_mant[16] ),
    .Q(net78),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[17]$_DFF_PN0_  (.D(\final_mant[17] ),
    .Q(net79),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[18]$_DFF_PN0_  (.D(\final_mant[18] ),
    .Q(net80),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[19]$_DFF_PN0_  (.D(\final_mant[19] ),
    .Q(net81),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[1]$_DFF_PN0_  (.D(\final_mant[1] ),
    .Q(net82),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[20]$_DFF_PN0_  (.D(\final_mant[20] ),
    .Q(net83),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[21]$_DFF_PN0_  (.D(\final_mant[21] ),
    .Q(net84),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[22]$_DFF_PN0_  (.D(\final_mant[22] ),
    .Q(net85),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[23]$_DFF_PN0_  (.D(\final_exp[0] ),
    .Q(net86),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[24]$_DFF_PN0_  (.D(\final_exp[1] ),
    .Q(net87),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[25]$_DFF_PN0_  (.D(\final_exp[2] ),
    .Q(net88),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[26]$_DFF_PN0_  (.D(\final_exp[3] ),
    .Q(net89),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[27]$_DFF_PN0_  (.D(\final_exp[4] ),
    .Q(net90),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[28]$_DFF_PN0_  (.D(\final_exp[5] ),
    .Q(net91),
    .RESET_B(net1),
    .CLK(clknet_4_7_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[29]$_DFF_PN0_  (.D(\final_exp[6] ),
    .Q(net92),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[2]$_DFF_PN0_  (.D(\final_mant[2] ),
    .Q(net93),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[30]$_DFF_PN0_  (.D(\final_exp[7] ),
    .Q(net94),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[31]$_DFF_PN0_  (.D(result_sign_stage2),
    .Q(net95),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[3]$_DFF_PN0_  (.D(\final_mant[3] ),
    .Q(net96),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[4]$_DFF_PN0_  (.D(\final_mant[4] ),
    .Q(net97),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[5]$_DFF_PN0_  (.D(\final_mant[5] ),
    .Q(net98),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[6]$_DFF_PN0_  (.D(\final_mant[6] ),
    .Q(net99),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[7]$_DFF_PN0_  (.D(\final_mant[7] ),
    .Q(net100),
    .RESET_B(net1),
    .CLK(clknet_4_5_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[8]$_DFF_PN0_  (.D(\final_mant[8] ),
    .Q(net101),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[9]$_DFF_PN0_  (.D(\final_mant[9] ),
    .Q(net102),
    .RESET_B(net1),
    .CLK(clknet_4_13_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \result_exp_stage2[0]$_DFF_PN0_  (.D(\larger_exp_stage1[0] ),
    .Q(\result_exp_stage2[0] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \result_exp_stage2[1]$_DFF_PN0_  (.D(\larger_exp_stage1[1] ),
    .Q(\result_exp_stage2[1] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result_exp_stage2[2]$_DFF_PN0_  (.D(\larger_exp_stage1[2] ),
    .Q(\result_exp_stage2[2] ),
    .RESET_B(net1),
    .CLK(clknet_4_3_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result_exp_stage2[3]$_DFF_PN0_  (.D(\larger_exp_stage1[3] ),
    .Q(\result_exp_stage2[3] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result_exp_stage2[4]$_DFF_PN0_  (.D(\larger_exp_stage1[4] ),
    .Q(\result_exp_stage2[4] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result_exp_stage2[5]$_DFF_PN0_  (.D(\larger_exp_stage1[5] ),
    .Q(\result_exp_stage2[5] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_2 \result_exp_stage2[6]$_DFF_PN0_  (.D(\larger_exp_stage1[6] ),
    .Q(\result_exp_stage2[6] ),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result_exp_stage2[7]$_DFF_PN0_  (.D(\larger_exp_stage1[7] ),
    .Q(\result_exp_stage2[7] ),
    .RESET_B(net1),
    .CLK(clknet_4_0_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \result_sign_stage2$_DFF_PN0_  (.D(_0119_),
    .Q(result_sign_stage2),
    .RESET_B(net1),
    .CLK(clknet_4_1_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \underflow$_DFF_PN0_  (.D(_0120_),
    .Q(net103),
    .RESET_B(net1),
    .CLK(clknet_4_4_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_out$_DFF_PN0_  (.D(valid_stage2),
    .Q(net104),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_stage1$_DFF_PN0_  (.D(net67),
    .Q(valid_stage1),
    .RESET_B(net1),
    .CLK(clknet_4_15_0_clk));
 sky130_fd_sc_hd__dfrtp_1 \valid_stage2$_DFF_PN0_  (.D(valid_stage1),
    .Q(valid_stage2),
    .RESET_B(net1),
    .CLK(clknet_4_14_0_clk));
 sky130_fd_sc_hd__buf_16 hold1 (.A(net66),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_377 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(a[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(a[10]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(a[11]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(a[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(a[13]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(a[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(a[15]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 input8 (.A(a[16]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(a[17]),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input10 (.A(a[18]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input11 (.A(a[19]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(a[1]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(a[20]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input14 (.A(a[21]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(a[22]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(a[23]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(a[24]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(a[25]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(a[26]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(a[27]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(a[28]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(a[29]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(a[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(a[30]),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(net107),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(a[3]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(a[4]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input28 (.A(a[5]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(a[6]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(a[7]),
    .X(net31));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(a[8]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(a[9]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(b[0]),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input34 (.A(b[10]),
    .X(net35));
 sky130_fd_sc_hd__dlymetal6s2s_1 input35 (.A(b[11]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(b[12]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(b[13]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(b[14]),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 input39 (.A(b[15]),
    .X(net40));
 sky130_fd_sc_hd__dlymetal6s2s_1 input40 (.A(b[16]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(b[17]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(b[18]),
    .X(net43));
 sky130_fd_sc_hd__buf_2 input43 (.A(b[19]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(b[1]),
    .X(net45));
 sky130_fd_sc_hd__dlymetal6s2s_1 input45 (.A(b[20]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(b[21]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 input47 (.A(b[22]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(b[23]),
    .X(net49));
 sky130_fd_sc_hd__dlymetal6s2s_1 input49 (.A(b[24]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(b[25]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(b[26]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(b[27]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(b[28]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(b[29]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(b[2]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(b[30]),
    .X(net57));
 sky130_fd_sc_hd__dlymetal6s2s_1 input57 (.A(net106),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(b[3]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(b[4]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(b[5]),
    .X(net61));
 sky130_fd_sc_hd__buf_2 input61 (.A(b[6]),
    .X(net62));
 sky130_fd_sc_hd__dlymetal6s2s_1 input62 (.A(b[7]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(b[8]),
    .X(net64));
 sky130_fd_sc_hd__buf_2 input64 (.A(b[9]),
    .X(net65));
 sky130_fd_sc_hd__buf_12 input65 (.A(rst_n),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(net105),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net68),
    .X(inexact));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net69),
    .X(invalid_op));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net70),
    .X(overflow));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net71),
    .X(result[0]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net72),
    .X(result[10]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net73),
    .X(result[11]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net74),
    .X(result[12]));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net75),
    .X(result[13]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net76),
    .X(result[14]));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net77),
    .X(result[15]));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net78),
    .X(result[16]));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net79),
    .X(result[17]));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net80),
    .X(result[18]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net81),
    .X(result[19]));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net82),
    .X(result[1]));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net83),
    .X(result[20]));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net84),
    .X(result[21]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net85),
    .X(result[22]));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(net86),
    .X(result[23]));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(net87),
    .X(result[24]));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(net88),
    .X(result[25]));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(net89),
    .X(result[26]));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net90),
    .X(result[27]));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(net91),
    .X(result[28]));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(net92),
    .X(result[29]));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(net93),
    .X(result[2]));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(net94),
    .X(result[30]));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net95),
    .X(result[31]));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(net96),
    .X(result[3]));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(net97),
    .X(result[4]));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(net98),
    .X(result[5]));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(net99),
    .X(result[6]));
 sky130_fd_sc_hd__clkbuf_1 output99 (.A(net100),
    .X(result[7]));
 sky130_fd_sc_hd__clkbuf_1 output100 (.A(net101),
    .X(result[8]));
 sky130_fd_sc_hd__clkbuf_1 output101 (.A(net102),
    .X(result[9]));
 sky130_fd_sc_hd__clkbuf_1 output102 (.A(net103),
    .X(underflow));
 sky130_fd_sc_hd__clkbuf_1 output103 (.A(net104),
    .X(valid_out));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload1 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__inv_6 clkload2 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__inv_6 clkload3 (.A(clknet_4_3_0_clk));
 sky130_fd_sc_hd__inv_6 clkload4 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__inv_4 clkload5 (.A(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkinv_8 clkload6 (.A(clknet_4_6_0_clk));
 sky130_fd_sc_hd__inv_8 clkload7 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload8 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__inv_8 clkload9 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload10 (.A(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload11 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload12 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload13 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__inv_4 clkload14 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(valid_in),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(b[31]),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(a[31]),
    .X(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0074_));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_207 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_19 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_330 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_5 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_212 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_284 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_354 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_280 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_87 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_140 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_92 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_70 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_150 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_62 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_106 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_182 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_66 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_60 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_272 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_272 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_34 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_353 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_23 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_367 ();
endmodule
