module barrel_rotator (direction,
    data_in,
    data_out,
    rotate_amount);
 input direction;
 input [7:0] data_in;
 output [7:0] data_out;
 input [2:0] rotate_amount;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;

 sky130_fd_sc_hd__buf_2 _119_ (.A(net8),
    .X(_044_));
 sky130_fd_sc_hd__inv_2 _120_ (.A(_044_),
    .Y(_045_));
 sky130_fd_sc_hd__clkbuf_4 _121_ (.A(data_in[1]),
    .X(_046_));
 sky130_fd_sc_hd__buf_6 _122_ (.A(rotate_amount[2]),
    .X(_047_));
 sky130_fd_sc_hd__mux2i_4 _123_ (.A0(net4),
    .A1(_046_),
    .S(_047_),
    .Y(_048_));
 sky130_fd_sc_hd__mux2i_4 _124_ (.A0(net5),
    .A1(net2),
    .S(_047_),
    .Y(_049_));
 sky130_fd_sc_hd__buf_6 _125_ (.A(rotate_amount[0]),
    .X(_050_));
 sky130_fd_sc_hd__inv_2 _126_ (.A(_050_),
    .Y(_051_));
 sky130_fd_sc_hd__mux2_1 _127_ (.A0(_048_),
    .A1(_049_),
    .S(_051_),
    .X(_052_));
 sky130_fd_sc_hd__mux2i_4 _128_ (.A0(net6),
    .A1(net3),
    .S(_047_),
    .Y(_053_));
 sky130_fd_sc_hd__or3_1 _129_ (.A(net8),
    .B(_051_),
    .C(_053_),
    .X(_054_));
 sky130_fd_sc_hd__buf_6 _130_ (.A(_047_),
    .X(_055_));
 sky130_fd_sc_hd__buf_2 _131_ (.A(_055_),
    .X(_056_));
 sky130_fd_sc_hd__clkbuf_4 _132_ (.A(data_in[4]),
    .X(_057_));
 sky130_fd_sc_hd__buf_6 _133_ (.A(_050_),
    .X(_058_));
 sky130_fd_sc_hd__nor2_2 _134_ (.A(_044_),
    .B(_058_),
    .Y(_059_));
 sky130_fd_sc_hd__inv_2 _135_ (.A(net7),
    .Y(_060_));
 sky130_fd_sc_hd__a31oi_1 _136_ (.A1(_056_),
    .A2(_057_),
    .A3(_059_),
    .B1(_060_),
    .Y(_061_));
 sky130_fd_sc_hd__o211a_1 _137_ (.A1(_045_),
    .A2(_052_),
    .B1(_054_),
    .C1(_061_),
    .X(_062_));
 sky130_fd_sc_hd__buf_2 _138_ (.A(_044_),
    .X(_063_));
 sky130_fd_sc_hd__buf_6 _139_ (.A(_050_),
    .X(_064_));
 sky130_fd_sc_hd__mux2i_1 _140_ (.A0(net5),
    .A1(net6),
    .S(_064_),
    .Y(_065_));
 sky130_fd_sc_hd__nand2_1 _141_ (.A(_056_),
    .B(_065_),
    .Y(_066_));
 sky130_fd_sc_hd__nor2_1 _142_ (.A(_064_),
    .B(net2),
    .Y(_067_));
 sky130_fd_sc_hd__clkbuf_4 _143_ (.A(net3),
    .X(_068_));
 sky130_fd_sc_hd__nor2b_1 _144_ (.A(_068_),
    .B_N(_058_),
    .Y(_069_));
 sky130_fd_sc_hd__inv_1 _145_ (.A(_056_),
    .Y(_070_));
 sky130_fd_sc_hd__o21ai_0 _146_ (.A1(_067_),
    .A2(_069_),
    .B1(_070_),
    .Y(_071_));
 sky130_fd_sc_hd__buf_2 _147_ (.A(_064_),
    .X(_072_));
 sky130_fd_sc_hd__buf_6 _148_ (.A(_055_),
    .X(_073_));
 sky130_fd_sc_hd__mux2i_2 _149_ (.A0(_046_),
    .A1(net4),
    .S(_073_),
    .Y(_074_));
 sky130_fd_sc_hd__nand3_1 _150_ (.A(_072_),
    .B(_060_),
    .C(_074_),
    .Y(_075_));
 sky130_fd_sc_hd__clkbuf_4 _151_ (.A(net7),
    .X(_076_));
 sky130_fd_sc_hd__o22ai_1 _152_ (.A1(_044_),
    .A2(_056_),
    .B1(_057_),
    .B2(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__a22oi_1 _153_ (.A1(_063_),
    .A2(_060_),
    .B1(_077_),
    .B2(_051_),
    .Y(_078_));
 sky130_fd_sc_hd__a32oi_1 _154_ (.A1(_063_),
    .A2(_066_),
    .A3(_071_),
    .B1(_075_),
    .B2(_078_),
    .Y(_079_));
 sky130_fd_sc_hd__nand2_2 _155_ (.A(_070_),
    .B(_059_),
    .Y(_080_));
 sky130_fd_sc_hd__inv_1 _156_ (.A(net1),
    .Y(_081_));
 sky130_fd_sc_hd__o22ai_1 _157_ (.A1(_062_),
    .A2(_079_),
    .B1(_080_),
    .B2(_081_),
    .Y(net9));
 sky130_fd_sc_hd__inv_1 _158_ (.A(_068_),
    .Y(_082_));
 sky130_fd_sc_hd__a21oi_1 _159_ (.A1(_056_),
    .A2(net6),
    .B1(_072_),
    .Y(_083_));
 sky130_fd_sc_hd__o21ai_0 _160_ (.A1(_056_),
    .A2(_082_),
    .B1(_083_),
    .Y(_084_));
 sky130_fd_sc_hd__mux2i_2 _161_ (.A0(_057_),
    .A1(net1),
    .S(_055_),
    .Y(_085_));
 sky130_fd_sc_hd__nand2_1 _162_ (.A(_072_),
    .B(_085_),
    .Y(_086_));
 sky130_fd_sc_hd__or2_1 _163_ (.A(net8),
    .B(_058_),
    .X(_087_));
 sky130_fd_sc_hd__nor2b_1 _164_ (.A(net4),
    .B_N(_055_),
    .Y(_088_));
 sky130_fd_sc_hd__mux2i_1 _165_ (.A0(net2),
    .A1(net5),
    .S(_056_),
    .Y(_089_));
 sky130_fd_sc_hd__nand2b_1 _166_ (.A_N(net8),
    .B(_064_),
    .Y(_090_));
 sky130_fd_sc_hd__o221ai_1 _167_ (.A1(_087_),
    .A2(_088_),
    .B1(_089_),
    .B2(_090_),
    .C1(_060_),
    .Y(_091_));
 sky130_fd_sc_hd__a31oi_1 _168_ (.A1(_063_),
    .A2(_084_),
    .A3(_086_),
    .B1(_091_),
    .Y(_092_));
 sky130_fd_sc_hd__mux2i_4 _169_ (.A0(net1),
    .A1(_057_),
    .S(_047_),
    .Y(_093_));
 sky130_fd_sc_hd__mux4_1 _170_ (.A0(_049_),
    .A1(_053_),
    .A2(_093_),
    .A3(_088_),
    .S0(_051_),
    .S1(_045_),
    .X(_094_));
 sky130_fd_sc_hd__o2bb2ai_1 _171_ (.A1_N(_076_),
    .A2_N(_094_),
    .B1(_080_),
    .B2(_046_),
    .Y(_095_));
 sky130_fd_sc_hd__nor2_1 _172_ (.A(_092_),
    .B(_095_),
    .Y(net10));
 sky130_fd_sc_hd__nand2_1 _173_ (.A(_058_),
    .B(_048_),
    .Y(_096_));
 sky130_fd_sc_hd__nand2_1 _174_ (.A(_051_),
    .B(_085_),
    .Y(_097_));
 sky130_fd_sc_hd__nor3b_1 _175_ (.A(_055_),
    .B(_068_),
    .C_N(_064_),
    .Y(_098_));
 sky130_fd_sc_hd__a211oi_1 _176_ (.A1(_073_),
    .A2(_065_),
    .B1(_098_),
    .C1(_044_),
    .Y(_099_));
 sky130_fd_sc_hd__a311o_1 _177_ (.A1(_063_),
    .A2(_096_),
    .A3(_097_),
    .B1(_099_),
    .C1(_076_),
    .X(_100_));
 sky130_fd_sc_hd__nand2_1 _178_ (.A(_072_),
    .B(_053_),
    .Y(_101_));
 sky130_fd_sc_hd__a21oi_1 _179_ (.A1(_051_),
    .A2(_093_),
    .B1(_045_),
    .Y(_102_));
 sky130_fd_sc_hd__mux2i_1 _180_ (.A0(net5),
    .A1(net4),
    .S(_064_),
    .Y(_103_));
 sky130_fd_sc_hd__nor3b_1 _181_ (.A(_055_),
    .B(_046_),
    .C_N(_064_),
    .Y(_104_));
 sky130_fd_sc_hd__a211oi_1 _182_ (.A1(_073_),
    .A2(_103_),
    .B1(_104_),
    .C1(_044_),
    .Y(_105_));
 sky130_fd_sc_hd__a211o_1 _183_ (.A1(_101_),
    .A2(_102_),
    .B1(_105_),
    .C1(_060_),
    .X(_106_));
 sky130_fd_sc_hd__o211a_1 _184_ (.A1(net2),
    .A2(_080_),
    .B1(_100_),
    .C1(_106_),
    .X(net11));
 sky130_fd_sc_hd__nand2_1 _185_ (.A(_072_),
    .B(_049_),
    .Y(_107_));
 sky130_fd_sc_hd__nand2_1 _186_ (.A(_051_),
    .B(_048_),
    .Y(_108_));
 sky130_fd_sc_hd__nor2_1 _187_ (.A(_063_),
    .B(_083_),
    .Y(_109_));
 sky130_fd_sc_hd__a32oi_1 _188_ (.A1(_063_),
    .A2(_107_),
    .A3(_108_),
    .B1(_086_),
    .B2(_109_),
    .Y(_110_));
 sky130_fd_sc_hd__nor2_1 _189_ (.A(_056_),
    .B(_087_),
    .Y(_111_));
 sky130_fd_sc_hd__a21oi_1 _190_ (.A1(_068_),
    .A2(_111_),
    .B1(_076_),
    .Y(_112_));
 sky130_fd_sc_hd__a21oi_1 _191_ (.A1(_068_),
    .A2(_111_),
    .B1(_060_),
    .Y(_113_));
 sky130_fd_sc_hd__mux2i_1 _192_ (.A0(_074_),
    .A1(_093_),
    .S(_072_),
    .Y(_114_));
 sky130_fd_sc_hd__mux2i_1 _193_ (.A0(net6),
    .A1(net5),
    .S(_058_),
    .Y(_115_));
 sky130_fd_sc_hd__nand3b_1 _194_ (.A_N(_056_),
    .B(_072_),
    .C(net2),
    .Y(_116_));
 sky130_fd_sc_hd__o211ai_1 _195_ (.A1(_070_),
    .A2(_115_),
    .B1(_116_),
    .C1(_045_),
    .Y(_117_));
 sky130_fd_sc_hd__o21ai_1 _196_ (.A1(_045_),
    .A2(_114_),
    .B1(_117_),
    .Y(_118_));
 sky130_fd_sc_hd__a22oi_2 _197_ (.A1(_110_),
    .A2(_112_),
    .B1(_113_),
    .B2(_118_),
    .Y(net12));
 sky130_fd_sc_hd__o21ai_0 _198_ (.A1(_070_),
    .A2(net1),
    .B1(_059_),
    .Y(_000_));
 sky130_fd_sc_hd__nor2_1 _199_ (.A(_072_),
    .B(_049_),
    .Y(_001_));
 sky130_fd_sc_hd__nor2_1 _200_ (.A(_051_),
    .B(_053_),
    .Y(_002_));
 sky130_fd_sc_hd__o21ai_0 _201_ (.A1(_051_),
    .A2(_048_),
    .B1(_045_),
    .Y(_003_));
 sky130_fd_sc_hd__o31ai_1 _202_ (.A1(_045_),
    .A2(_001_),
    .A3(_002_),
    .B1(_003_),
    .Y(_004_));
 sky130_fd_sc_hd__nor2b_1 _203_ (.A(net2),
    .B_N(net8),
    .Y(_005_));
 sky130_fd_sc_hd__nand3_1 _204_ (.A(_044_),
    .B(_058_),
    .C(_046_),
    .Y(_006_));
 sky130_fd_sc_hd__o21ai_0 _205_ (.A1(_058_),
    .A2(_005_),
    .B1(_006_),
    .Y(_007_));
 sky130_fd_sc_hd__nand2_1 _206_ (.A(_072_),
    .B(_068_),
    .Y(_008_));
 sky130_fd_sc_hd__mux2i_1 _207_ (.A0(net1),
    .A1(net6),
    .S(_058_),
    .Y(_009_));
 sky130_fd_sc_hd__mux2i_1 _208_ (.A0(_008_),
    .A1(_009_),
    .S(_073_),
    .Y(_010_));
 sky130_fd_sc_hd__nand2_1 _209_ (.A(_044_),
    .B(_073_),
    .Y(_011_));
 sky130_fd_sc_hd__o21ai_1 _210_ (.A1(_103_),
    .A2(_011_),
    .B1(_076_),
    .Y(_012_));
 sky130_fd_sc_hd__a221oi_2 _211_ (.A1(_070_),
    .A2(_007_),
    .B1(_010_),
    .B2(_045_),
    .C1(_012_),
    .Y(_013_));
 sky130_fd_sc_hd__nor2_1 _212_ (.A(_057_),
    .B(_080_),
    .Y(_014_));
 sky130_fd_sc_hd__a311oi_2 _213_ (.A1(_060_),
    .A2(_000_),
    .A3(_004_),
    .B1(_013_),
    .C1(_014_),
    .Y(net13));
 sky130_fd_sc_hd__nor2b_1 _214_ (.A(_055_),
    .B_N(_064_),
    .Y(_015_));
 sky130_fd_sc_hd__mux2_1 _215_ (.A0(_046_),
    .A1(net1),
    .S(_050_),
    .X(_016_));
 sky130_fd_sc_hd__a22oi_1 _216_ (.A1(_057_),
    .A2(_015_),
    .B1(_016_),
    .B2(_073_),
    .Y(_017_));
 sky130_fd_sc_hd__nand2_1 _217_ (.A(net8),
    .B(net2),
    .Y(_018_));
 sky130_fd_sc_hd__nor2_1 _218_ (.A(_064_),
    .B(_068_),
    .Y(_019_));
 sky130_fd_sc_hd__a221o_1 _219_ (.A1(_058_),
    .A2(_018_),
    .B1(_019_),
    .B2(net8),
    .C1(_073_),
    .X(_020_));
 sky130_fd_sc_hd__o221a_1 _220_ (.A1(_115_),
    .A2(_011_),
    .B1(_017_),
    .B2(_044_),
    .C1(_020_),
    .X(_021_));
 sky130_fd_sc_hd__nand2_1 _221_ (.A(_072_),
    .B(_093_),
    .Y(_022_));
 sky130_fd_sc_hd__nand2_1 _222_ (.A(_051_),
    .B(_053_),
    .Y(_023_));
 sky130_fd_sc_hd__nor2b_1 _223_ (.A(_046_),
    .B_N(_055_),
    .Y(_024_));
 sky130_fd_sc_hd__o221ai_1 _224_ (.A1(_049_),
    .A2(_090_),
    .B1(_024_),
    .B2(_087_),
    .C1(_060_),
    .Y(_025_));
 sky130_fd_sc_hd__a31oi_1 _225_ (.A1(_063_),
    .A2(_022_),
    .A3(_023_),
    .B1(_025_),
    .Y(_026_));
 sky130_fd_sc_hd__nor2_1 _226_ (.A(net4),
    .B(_080_),
    .Y(_027_));
 sky130_fd_sc_hd__a211oi_2 _227_ (.A1(_076_),
    .A2(_021_),
    .B1(_026_),
    .C1(_027_),
    .Y(net14));
 sky130_fd_sc_hd__nand2_1 _228_ (.A(_076_),
    .B(_048_),
    .Y(_028_));
 sky130_fd_sc_hd__nand2_1 _229_ (.A(_060_),
    .B(_053_),
    .Y(_029_));
 sky130_fd_sc_hd__a21oi_1 _230_ (.A1(_028_),
    .A2(_029_),
    .B1(_090_),
    .Y(_030_));
 sky130_fd_sc_hd__a21oi_1 _231_ (.A1(_073_),
    .A2(_067_),
    .B1(_044_),
    .Y(_031_));
 sky130_fd_sc_hd__mux4_1 _232_ (.A0(_057_),
    .A1(_068_),
    .A2(net1),
    .A3(net6),
    .S0(_050_),
    .S1(_055_),
    .X(_032_));
 sky130_fd_sc_hd__a211oi_1 _233_ (.A1(_096_),
    .A2(_031_),
    .B1(_032_),
    .C1(_060_),
    .Y(_033_));
 sky130_fd_sc_hd__mux4_1 _234_ (.A0(net1),
    .A1(_046_),
    .A2(_057_),
    .A3(net4),
    .S0(_050_),
    .S1(_055_),
    .X(_034_));
 sky130_fd_sc_hd__a211oi_1 _235_ (.A1(_101_),
    .A2(_031_),
    .B1(_034_),
    .C1(_076_),
    .Y(_035_));
 sky130_fd_sc_hd__a2111oi_2 _236_ (.A1(_059_),
    .A2(_049_),
    .B1(_030_),
    .C1(_033_),
    .D1(_035_),
    .Y(net15));
 sky130_fd_sc_hd__nor2_1 _237_ (.A(net6),
    .B(_080_),
    .Y(_036_));
 sky130_fd_sc_hd__nor2b_1 _238_ (.A(_068_),
    .B_N(_073_),
    .Y(_037_));
 sky130_fd_sc_hd__o221ai_1 _239_ (.A1(_049_),
    .A2(_090_),
    .B1(_037_),
    .B2(_087_),
    .C1(_076_),
    .Y(_038_));
 sky130_fd_sc_hd__a31oi_1 _240_ (.A1(_063_),
    .A2(_086_),
    .A3(_108_),
    .B1(_038_),
    .Y(_039_));
 sky130_fd_sc_hd__mux4_1 _241_ (.A0(_046_),
    .A1(net2),
    .A2(net4),
    .A3(net5),
    .S0(_064_),
    .S1(_073_),
    .X(_040_));
 sky130_fd_sc_hd__mux2i_1 _242_ (.A0(_068_),
    .A1(_057_),
    .S(_058_),
    .Y(_041_));
 sky130_fd_sc_hd__a221oi_1 _243_ (.A1(_081_),
    .A2(_015_),
    .B1(_041_),
    .B2(_056_),
    .C1(_063_),
    .Y(_042_));
 sky130_fd_sc_hd__a211oi_1 _244_ (.A1(_063_),
    .A2(_040_),
    .B1(_042_),
    .C1(_076_),
    .Y(_043_));
 sky130_fd_sc_hd__nor3_1 _245_ (.A(_036_),
    .B(_039_),
    .C(_043_),
    .Y(net16));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_107 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(data_in[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input2 (.A(data_in[2]),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(data_in[3]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input4 (.A(data_in[5]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(data_in[6]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(data_in[7]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(direction),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(rotate_amount[1]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 output9 (.A(net9),
    .X(data_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output10 (.A(net10),
    .X(data_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output11 (.A(net11),
    .X(data_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output12 (.A(net12),
    .X(data_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net13),
    .X(data_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net14),
    .X(data_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net15),
    .X(data_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net16),
    .X(data_out[7]));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_11 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_64 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_152 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_114 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_205 ();
endmodule
