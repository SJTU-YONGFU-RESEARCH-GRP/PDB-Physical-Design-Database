module parameterized_clock_gating (clk_in,
    clk_out,
    enable,
    test_mode);
 input clk_in;
 output clk_out;
 input enable;
 input test_mode;

 wire _0_;
 wire _1_;
 wire _2_;
 wire enable_final;
 wire enable_latch;
 wire \gen_sync.enable_sync_reg[0] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;

 OR2_X1 _3_ (.A1(net3),
    .A2(enable_final),
    .ZN(_0_));
 AND2_X1 _4_ (.A1(enable_latch),
    .A2(net1),
    .ZN(net4));
 DLL_X1 \enable_latch$_DLATCH_N_  (.D(_0_),
    .GN(net1),
    .Q(enable_latch));
 DFF_X1 \gen_sync.enable_sync_reg[0]$_DFF_P_  (.D(net2),
    .CK(net1),
    .Q(\gen_sync.enable_sync_reg[0] ),
    .QN(_2_));
 DFF_X1 \gen_sync.enable_sync_reg[1]$_DFF_P_  (.D(\gen_sync.enable_sync_reg[0] ),
    .CK(net1),
    .Q(enable_final),
    .QN(_1_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_69 ();
 BUF_X1 input1 (.A(clk_in),
    .Z(net1));
 BUF_X1 input2 (.A(enable),
    .Z(net2));
 BUF_X1 input3 (.A(test_mode),
    .Z(net3));
 BUF_X1 output4 (.A(net4),
    .Z(clk_out));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X4 FILLER_0_257 ();
 FILLCELL_X2 FILLER_0_261 ();
 FILLCELL_X1 FILLER_0_263 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X4 FILLER_1_257 ();
 FILLCELL_X2 FILLER_1_261 ();
 FILLCELL_X1 FILLER_1_263 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X4 FILLER_2_257 ();
 FILLCELL_X2 FILLER_2_261 ();
 FILLCELL_X1 FILLER_2_263 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X4 FILLER_3_257 ();
 FILLCELL_X2 FILLER_3_261 ();
 FILLCELL_X1 FILLER_3_263 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X4 FILLER_4_257 ();
 FILLCELL_X2 FILLER_4_261 ();
 FILLCELL_X1 FILLER_4_263 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X4 FILLER_5_257 ();
 FILLCELL_X2 FILLER_5_261 ();
 FILLCELL_X1 FILLER_5_263 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X4 FILLER_6_257 ();
 FILLCELL_X2 FILLER_6_261 ();
 FILLCELL_X1 FILLER_6_263 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X4 FILLER_7_257 ();
 FILLCELL_X2 FILLER_7_261 ();
 FILLCELL_X1 FILLER_7_263 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X4 FILLER_8_257 ();
 FILLCELL_X2 FILLER_8_261 ();
 FILLCELL_X1 FILLER_8_263 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X4 FILLER_9_257 ();
 FILLCELL_X2 FILLER_9_261 ();
 FILLCELL_X1 FILLER_9_263 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X32 FILLER_10_193 ();
 FILLCELL_X32 FILLER_10_225 ();
 FILLCELL_X4 FILLER_10_257 ();
 FILLCELL_X2 FILLER_10_261 ();
 FILLCELL_X1 FILLER_10_263 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X32 FILLER_11_193 ();
 FILLCELL_X32 FILLER_11_225 ();
 FILLCELL_X4 FILLER_11_257 ();
 FILLCELL_X2 FILLER_11_261 ();
 FILLCELL_X1 FILLER_11_263 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X32 FILLER_12_129 ();
 FILLCELL_X32 FILLER_12_161 ();
 FILLCELL_X32 FILLER_12_193 ();
 FILLCELL_X32 FILLER_12_225 ();
 FILLCELL_X4 FILLER_12_257 ();
 FILLCELL_X2 FILLER_12_261 ();
 FILLCELL_X1 FILLER_12_263 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X32 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_193 ();
 FILLCELL_X32 FILLER_13_225 ();
 FILLCELL_X4 FILLER_13_257 ();
 FILLCELL_X2 FILLER_13_261 ();
 FILLCELL_X1 FILLER_13_263 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X32 FILLER_14_193 ();
 FILLCELL_X32 FILLER_14_225 ();
 FILLCELL_X4 FILLER_14_257 ();
 FILLCELL_X2 FILLER_14_261 ();
 FILLCELL_X1 FILLER_14_263 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X32 FILLER_15_193 ();
 FILLCELL_X32 FILLER_15_225 ();
 FILLCELL_X4 FILLER_15_257 ();
 FILLCELL_X2 FILLER_15_261 ();
 FILLCELL_X1 FILLER_15_263 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X32 FILLER_16_193 ();
 FILLCELL_X32 FILLER_16_225 ();
 FILLCELL_X1 FILLER_16_257 ();
 FILLCELL_X2 FILLER_16_261 ();
 FILLCELL_X1 FILLER_16_263 ();
 FILLCELL_X16 FILLER_17_1 ();
 FILLCELL_X2 FILLER_17_17 ();
 FILLCELL_X1 FILLER_17_19 ();
 FILLCELL_X32 FILLER_17_23 ();
 FILLCELL_X32 FILLER_17_55 ();
 FILLCELL_X32 FILLER_17_87 ();
 FILLCELL_X32 FILLER_17_119 ();
 FILLCELL_X32 FILLER_17_151 ();
 FILLCELL_X32 FILLER_17_183 ();
 FILLCELL_X8 FILLER_17_215 ();
 FILLCELL_X4 FILLER_17_223 ();
 FILLCELL_X2 FILLER_17_244 ();
 FILLCELL_X1 FILLER_17_260 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X32 FILLER_18_193 ();
 FILLCELL_X8 FILLER_18_225 ();
 FILLCELL_X4 FILLER_18_233 ();
 FILLCELL_X1 FILLER_18_237 ();
 FILLCELL_X2 FILLER_18_262 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X32 FILLER_19_193 ();
 FILLCELL_X32 FILLER_19_225 ();
 FILLCELL_X4 FILLER_19_257 ();
 FILLCELL_X2 FILLER_19_261 ();
 FILLCELL_X1 FILLER_19_263 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X32 FILLER_20_193 ();
 FILLCELL_X32 FILLER_20_225 ();
 FILLCELL_X4 FILLER_20_257 ();
 FILLCELL_X2 FILLER_20_261 ();
 FILLCELL_X1 FILLER_20_263 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X32 FILLER_21_193 ();
 FILLCELL_X32 FILLER_21_225 ();
 FILLCELL_X4 FILLER_21_257 ();
 FILLCELL_X2 FILLER_21_261 ();
 FILLCELL_X1 FILLER_21_263 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X32 FILLER_22_193 ();
 FILLCELL_X32 FILLER_22_225 ();
 FILLCELL_X4 FILLER_22_257 ();
 FILLCELL_X2 FILLER_22_261 ();
 FILLCELL_X1 FILLER_22_263 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X32 FILLER_23_225 ();
 FILLCELL_X4 FILLER_23_257 ();
 FILLCELL_X2 FILLER_23_261 ();
 FILLCELL_X1 FILLER_23_263 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X32 FILLER_24_193 ();
 FILLCELL_X32 FILLER_24_225 ();
 FILLCELL_X4 FILLER_24_257 ();
 FILLCELL_X2 FILLER_24_261 ();
 FILLCELL_X1 FILLER_24_263 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X32 FILLER_25_193 ();
 FILLCELL_X32 FILLER_25_225 ();
 FILLCELL_X4 FILLER_25_257 ();
 FILLCELL_X2 FILLER_25_261 ();
 FILLCELL_X1 FILLER_25_263 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X32 FILLER_26_225 ();
 FILLCELL_X4 FILLER_26_257 ();
 FILLCELL_X2 FILLER_26_261 ();
 FILLCELL_X1 FILLER_26_263 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X32 FILLER_27_225 ();
 FILLCELL_X4 FILLER_27_257 ();
 FILLCELL_X2 FILLER_27_261 ();
 FILLCELL_X1 FILLER_27_263 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X4 FILLER_28_257 ();
 FILLCELL_X2 FILLER_28_261 ();
 FILLCELL_X1 FILLER_28_263 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X4 FILLER_29_257 ();
 FILLCELL_X2 FILLER_29_261 ();
 FILLCELL_X1 FILLER_29_263 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X4 FILLER_30_257 ();
 FILLCELL_X2 FILLER_30_261 ();
 FILLCELL_X1 FILLER_30_263 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X4 FILLER_31_257 ();
 FILLCELL_X2 FILLER_31_261 ();
 FILLCELL_X1 FILLER_31_263 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X4 FILLER_32_257 ();
 FILLCELL_X2 FILLER_32_261 ();
 FILLCELL_X1 FILLER_32_263 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X4 FILLER_33_257 ();
 FILLCELL_X2 FILLER_33_261 ();
 FILLCELL_X1 FILLER_33_263 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X32 FILLER_34_161 ();
 FILLCELL_X32 FILLER_34_193 ();
 FILLCELL_X32 FILLER_34_225 ();
 FILLCELL_X4 FILLER_34_257 ();
 FILLCELL_X2 FILLER_34_261 ();
 FILLCELL_X1 FILLER_34_263 ();
endmodule
