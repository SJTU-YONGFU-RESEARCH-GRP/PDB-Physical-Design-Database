module parameterized_onehot_counter (clk,
    enable,
    rst_n,
    count);
 input clk;
 input enable;
 input rst_n;
 output [7:0] count;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire _34_;
 wire _35_;
 wire _36_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 BUF_X4 _37_ (.A(rst_n),
    .Z(_08_));
 BUF_X4 _38_ (.A(enable),
    .Z(_09_));
 INV_X4 _39_ (.A(_09_),
    .ZN(_10_));
 NOR2_X1 _40_ (.A1(net8),
    .A2(_10_),
    .ZN(_11_));
 NOR2_X1 _41_ (.A1(net1),
    .A2(_09_),
    .ZN(_12_));
 OAI21_X1 _42_ (.A(_08_),
    .B1(_11_),
    .B2(_12_),
    .ZN(_00_));
 NAND3_X1 _43_ (.A1(net2),
    .A2(_10_),
    .A3(_08_),
    .ZN(_13_));
 NAND2_X2 _44_ (.A1(_09_),
    .A2(_08_),
    .ZN(_14_));
 INV_X2 _45_ (.A(net8),
    .ZN(_15_));
 NAND2_X1 _46_ (.A1(net1),
    .A2(_15_),
    .ZN(_16_));
 OAI21_X1 _47_ (.A(_13_),
    .B1(_14_),
    .B2(_16_),
    .ZN(_01_));
 NAND3_X1 _48_ (.A1(net3),
    .A2(_10_),
    .A3(_08_),
    .ZN(_17_));
 NAND2_X1 _49_ (.A1(_15_),
    .A2(net2),
    .ZN(_18_));
 OAI21_X1 _50_ (.A(_17_),
    .B1(_18_),
    .B2(_14_),
    .ZN(_02_));
 NAND3_X1 _51_ (.A1(net4),
    .A2(_10_),
    .A3(_08_),
    .ZN(_19_));
 NAND2_X1 _52_ (.A1(_15_),
    .A2(net3),
    .ZN(_20_));
 OAI21_X1 _53_ (.A(_19_),
    .B1(_20_),
    .B2(_14_),
    .ZN(_03_));
 NAND3_X1 _54_ (.A1(net5),
    .A2(_10_),
    .A3(_08_),
    .ZN(_21_));
 NAND2_X1 _55_ (.A1(_15_),
    .A2(net4),
    .ZN(_22_));
 OAI21_X1 _56_ (.A(_21_),
    .B1(_22_),
    .B2(_14_),
    .ZN(_04_));
 NAND3_X1 _57_ (.A1(net6),
    .A2(_10_),
    .A3(_08_),
    .ZN(_23_));
 NAND2_X1 _58_ (.A1(_15_),
    .A2(net5),
    .ZN(_24_));
 OAI21_X1 _59_ (.A(_23_),
    .B1(_24_),
    .B2(_14_),
    .ZN(_05_));
 NAND3_X1 _60_ (.A1(net7),
    .A2(_10_),
    .A3(_08_),
    .ZN(_25_));
 NAND2_X1 _61_ (.A1(_15_),
    .A2(net6),
    .ZN(_26_));
 OAI21_X1 _62_ (.A(_25_),
    .B1(_26_),
    .B2(_14_),
    .ZN(_06_));
 NAND3_X1 _63_ (.A1(net8),
    .A2(_10_),
    .A3(_08_),
    .ZN(_27_));
 NAND2_X1 _64_ (.A1(_15_),
    .A2(net7),
    .ZN(_28_));
 OAI21_X1 _65_ (.A(_27_),
    .B1(_28_),
    .B2(_14_),
    .ZN(_07_));
 DFF_X1 \counter_reg[0]$_SDFFE_PN1P_  (.D(_00_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net1),
    .QN(_36_));
 DFF_X1 \counter_reg[1]$_SDFFE_PN0P_  (.D(_01_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net2),
    .QN(_35_));
 DFF_X1 \counter_reg[2]$_SDFFE_PN0P_  (.D(_02_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net3),
    .QN(_34_));
 DFF_X1 \counter_reg[3]$_SDFFE_PN0P_  (.D(_03_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net4),
    .QN(_33_));
 DFF_X1 \counter_reg[4]$_SDFFE_PN0P_  (.D(_04_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net5),
    .QN(_32_));
 DFF_X1 \counter_reg[5]$_SDFFE_PN0P_  (.D(_05_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net6),
    .QN(_31_));
 DFF_X1 \counter_reg[6]$_SDFFE_PN0P_  (.D(_06_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net7),
    .QN(_30_));
 DFF_X2 \counter_reg[7]$_SDFFE_PN0P_  (.D(_07_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net8),
    .QN(_29_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_53 ();
 BUF_X1 output1 (.A(net1),
    .Z(count[0]));
 BUF_X1 output2 (.A(net2),
    .Z(count[1]));
 BUF_X1 output3 (.A(net3),
    .Z(count[2]));
 BUF_X1 output4 (.A(net4),
    .Z(count[3]));
 BUF_X1 output5 (.A(net5),
    .Z(count[4]));
 BUF_X1 output6 (.A(net6),
    .Z(count[5]));
 BUF_X1 output7 (.A(net7),
    .Z(count[6]));
 BUF_X1 output8 (.A(net8),
    .Z(count[7]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 CLKBUF_X1 clkload0 (.A(clknet_1_0__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X16 FILLER_0_65 ();
 FILLCELL_X2 FILLER_0_81 ();
 FILLCELL_X4 FILLER_0_86 ();
 FILLCELL_X2 FILLER_0_90 ();
 FILLCELL_X1 FILLER_0_92 ();
 FILLCELL_X32 FILLER_0_96 ();
 FILLCELL_X32 FILLER_0_128 ();
 FILLCELL_X32 FILLER_0_160 ();
 FILLCELL_X4 FILLER_0_192 ();
 FILLCELL_X2 FILLER_0_196 ();
 FILLCELL_X1 FILLER_0_198 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_104 ();
 FILLCELL_X32 FILLER_1_136 ();
 FILLCELL_X16 FILLER_1_168 ();
 FILLCELL_X8 FILLER_1_184 ();
 FILLCELL_X4 FILLER_1_192 ();
 FILLCELL_X2 FILLER_1_196 ();
 FILLCELL_X1 FILLER_1_198 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X8 FILLER_2_65 ();
 FILLCELL_X4 FILLER_2_73 ();
 FILLCELL_X1 FILLER_2_77 ();
 FILLCELL_X2 FILLER_2_85 ();
 FILLCELL_X32 FILLER_2_104 ();
 FILLCELL_X32 FILLER_2_136 ();
 FILLCELL_X16 FILLER_2_168 ();
 FILLCELL_X8 FILLER_2_184 ();
 FILLCELL_X4 FILLER_2_192 ();
 FILLCELL_X2 FILLER_2_196 ();
 FILLCELL_X1 FILLER_2_198 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X8 FILLER_3_65 ();
 FILLCELL_X2 FILLER_3_73 ();
 FILLCELL_X1 FILLER_3_75 ();
 FILLCELL_X2 FILLER_3_96 ();
 FILLCELL_X2 FILLER_3_103 ();
 FILLCELL_X32 FILLER_3_110 ();
 FILLCELL_X32 FILLER_3_142 ();
 FILLCELL_X16 FILLER_3_174 ();
 FILLCELL_X8 FILLER_3_190 ();
 FILLCELL_X1 FILLER_3_198 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X16 FILLER_4_65 ();
 FILLCELL_X2 FILLER_4_81 ();
 FILLCELL_X1 FILLER_4_96 ();
 FILLCELL_X1 FILLER_4_104 ();
 FILLCELL_X32 FILLER_4_108 ();
 FILLCELL_X32 FILLER_4_140 ();
 FILLCELL_X16 FILLER_4_172 ();
 FILLCELL_X8 FILLER_4_188 ();
 FILLCELL_X2 FILLER_4_196 ();
 FILLCELL_X1 FILLER_4_198 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X16 FILLER_5_65 ();
 FILLCELL_X8 FILLER_5_81 ();
 FILLCELL_X2 FILLER_5_89 ();
 FILLCELL_X8 FILLER_5_94 ();
 FILLCELL_X4 FILLER_5_102 ();
 FILLCELL_X2 FILLER_5_114 ();
 FILLCELL_X1 FILLER_5_116 ();
 FILLCELL_X32 FILLER_5_136 ();
 FILLCELL_X16 FILLER_5_168 ();
 FILLCELL_X8 FILLER_5_184 ();
 FILLCELL_X4 FILLER_5_192 ();
 FILLCELL_X2 FILLER_5_196 ();
 FILLCELL_X1 FILLER_5_198 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X4 FILLER_6_193 ();
 FILLCELL_X2 FILLER_6_197 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X16 FILLER_7_65 ();
 FILLCELL_X4 FILLER_7_81 ();
 FILLCELL_X2 FILLER_7_85 ();
 FILLCELL_X8 FILLER_7_90 ();
 FILLCELL_X4 FILLER_7_98 ();
 FILLCELL_X1 FILLER_7_102 ();
 FILLCELL_X2 FILLER_7_108 ();
 FILLCELL_X32 FILLER_7_113 ();
 FILLCELL_X32 FILLER_7_145 ();
 FILLCELL_X16 FILLER_7_177 ();
 FILLCELL_X4 FILLER_7_193 ();
 FILLCELL_X2 FILLER_7_197 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X2 FILLER_8_65 ();
 FILLCELL_X1 FILLER_8_67 ();
 FILLCELL_X8 FILLER_8_93 ();
 FILLCELL_X4 FILLER_8_101 ();
 FILLCELL_X1 FILLER_8_105 ();
 FILLCELL_X32 FILLER_8_113 ();
 FILLCELL_X16 FILLER_8_145 ();
 FILLCELL_X32 FILLER_8_164 ();
 FILLCELL_X2 FILLER_8_196 ();
 FILLCELL_X1 FILLER_8_198 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X16 FILLER_9_65 ();
 FILLCELL_X4 FILLER_9_81 ();
 FILLCELL_X1 FILLER_9_85 ();
 FILLCELL_X8 FILLER_9_93 ();
 FILLCELL_X4 FILLER_9_101 ();
 FILLCELL_X2 FILLER_9_105 ();
 FILLCELL_X2 FILLER_9_115 ();
 FILLCELL_X32 FILLER_9_134 ();
 FILLCELL_X32 FILLER_9_166 ();
 FILLCELL_X1 FILLER_9_198 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X4 FILLER_10_65 ();
 FILLCELL_X1 FILLER_10_69 ();
 FILLCELL_X2 FILLER_10_91 ();
 FILLCELL_X2 FILLER_10_96 ();
 FILLCELL_X2 FILLER_10_106 ();
 FILLCELL_X1 FILLER_10_111 ();
 FILLCELL_X32 FILLER_10_124 ();
 FILLCELL_X4 FILLER_10_156 ();
 FILLCELL_X32 FILLER_10_163 ();
 FILLCELL_X4 FILLER_10_195 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X4 FILLER_11_97 ();
 FILLCELL_X2 FILLER_11_101 ();
 FILLCELL_X1 FILLER_11_103 ();
 FILLCELL_X32 FILLER_11_138 ();
 FILLCELL_X16 FILLER_11_170 ();
 FILLCELL_X8 FILLER_11_186 ();
 FILLCELL_X4 FILLER_11_194 ();
 FILLCELL_X1 FILLER_11_198 ();
 FILLCELL_X4 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_8 ();
 FILLCELL_X32 FILLER_12_40 ();
 FILLCELL_X32 FILLER_12_72 ();
 FILLCELL_X32 FILLER_12_104 ();
 FILLCELL_X32 FILLER_12_136 ();
 FILLCELL_X4 FILLER_12_168 ();
 FILLCELL_X1 FILLER_12_172 ();
 FILLCELL_X16 FILLER_12_176 ();
 FILLCELL_X4 FILLER_12_192 ();
 FILLCELL_X2 FILLER_12_196 ();
 FILLCELL_X1 FILLER_12_198 ();
 FILLCELL_X16 FILLER_13_1 ();
 FILLCELL_X2 FILLER_13_17 ();
 FILLCELL_X1 FILLER_13_19 ();
 FILLCELL_X32 FILLER_13_23 ();
 FILLCELL_X32 FILLER_13_55 ();
 FILLCELL_X32 FILLER_13_87 ();
 FILLCELL_X32 FILLER_13_119 ();
 FILLCELL_X8 FILLER_13_151 ();
 FILLCELL_X2 FILLER_13_159 ();
 FILLCELL_X1 FILLER_13_161 ();
 FILLCELL_X32 FILLER_13_165 ();
 FILLCELL_X2 FILLER_13_197 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X32 FILLER_14_161 ();
 FILLCELL_X4 FILLER_14_193 ();
 FILLCELL_X2 FILLER_14_197 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X32 FILLER_15_161 ();
 FILLCELL_X4 FILLER_15_193 ();
 FILLCELL_X2 FILLER_15_197 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X32 FILLER_16_161 ();
 FILLCELL_X4 FILLER_16_193 ();
 FILLCELL_X2 FILLER_16_197 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X32 FILLER_17_161 ();
 FILLCELL_X4 FILLER_17_193 ();
 FILLCELL_X2 FILLER_17_197 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X32 FILLER_18_161 ();
 FILLCELL_X4 FILLER_18_193 ();
 FILLCELL_X2 FILLER_18_197 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X4 FILLER_19_193 ();
 FILLCELL_X2 FILLER_19_197 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X4 FILLER_20_193 ();
 FILLCELL_X2 FILLER_20_197 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X4 FILLER_21_193 ();
 FILLCELL_X2 FILLER_21_197 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X4 FILLER_22_193 ();
 FILLCELL_X2 FILLER_22_197 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X4 FILLER_23_193 ();
 FILLCELL_X2 FILLER_23_197 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X4 FILLER_24_193 ();
 FILLCELL_X2 FILLER_24_197 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X4 FILLER_25_193 ();
 FILLCELL_X2 FILLER_25_197 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X4 FILLER_26_193 ();
 FILLCELL_X2 FILLER_26_197 ();
endmodule
