module parameterized_cam (clk,
    compare_enable,
    match,
    rst_n,
    valid,
    write_enable,
    compare_data,
    match_addr,
    write_addr,
    write_data);
 input clk;
 input compare_enable;
 output match;
 input rst_n;
 output valid;
 input write_enable;
 input [7:0] compare_data;
 output [3:0] match_addr;
 input [3:0] write_addr;
 input [7:0] write_data;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire \cam_memory[0][0] ;
 wire \cam_memory[0][1] ;
 wire \cam_memory[0][2] ;
 wire \cam_memory[0][3] ;
 wire \cam_memory[0][4] ;
 wire \cam_memory[0][5] ;
 wire \cam_memory[0][6] ;
 wire \cam_memory[0][7] ;
 wire \cam_memory[10][0] ;
 wire \cam_memory[10][1] ;
 wire \cam_memory[10][2] ;
 wire \cam_memory[10][3] ;
 wire \cam_memory[10][4] ;
 wire \cam_memory[10][5] ;
 wire \cam_memory[10][6] ;
 wire \cam_memory[10][7] ;
 wire \cam_memory[11][0] ;
 wire \cam_memory[11][1] ;
 wire \cam_memory[11][2] ;
 wire \cam_memory[11][3] ;
 wire \cam_memory[11][4] ;
 wire \cam_memory[11][5] ;
 wire \cam_memory[11][6] ;
 wire \cam_memory[11][7] ;
 wire \cam_memory[12][0] ;
 wire \cam_memory[12][1] ;
 wire \cam_memory[12][2] ;
 wire \cam_memory[12][3] ;
 wire \cam_memory[12][4] ;
 wire \cam_memory[12][5] ;
 wire \cam_memory[12][6] ;
 wire \cam_memory[12][7] ;
 wire \cam_memory[13][0] ;
 wire \cam_memory[13][1] ;
 wire \cam_memory[13][2] ;
 wire \cam_memory[13][3] ;
 wire \cam_memory[13][4] ;
 wire \cam_memory[13][5] ;
 wire \cam_memory[13][6] ;
 wire \cam_memory[13][7] ;
 wire \cam_memory[14][0] ;
 wire \cam_memory[14][1] ;
 wire \cam_memory[14][2] ;
 wire \cam_memory[14][3] ;
 wire \cam_memory[14][4] ;
 wire \cam_memory[14][5] ;
 wire \cam_memory[14][6] ;
 wire \cam_memory[14][7] ;
 wire \cam_memory[15][0] ;
 wire \cam_memory[15][1] ;
 wire \cam_memory[15][2] ;
 wire \cam_memory[15][3] ;
 wire \cam_memory[15][4] ;
 wire \cam_memory[15][5] ;
 wire \cam_memory[15][6] ;
 wire \cam_memory[15][7] ;
 wire \cam_memory[1][0] ;
 wire \cam_memory[1][1] ;
 wire \cam_memory[1][2] ;
 wire \cam_memory[1][3] ;
 wire \cam_memory[1][4] ;
 wire \cam_memory[1][5] ;
 wire \cam_memory[1][6] ;
 wire \cam_memory[1][7] ;
 wire \cam_memory[2][0] ;
 wire \cam_memory[2][1] ;
 wire \cam_memory[2][2] ;
 wire \cam_memory[2][3] ;
 wire \cam_memory[2][4] ;
 wire \cam_memory[2][5] ;
 wire \cam_memory[2][6] ;
 wire \cam_memory[2][7] ;
 wire \cam_memory[3][0] ;
 wire \cam_memory[3][1] ;
 wire \cam_memory[3][2] ;
 wire \cam_memory[3][3] ;
 wire \cam_memory[3][4] ;
 wire \cam_memory[3][5] ;
 wire \cam_memory[3][6] ;
 wire \cam_memory[3][7] ;
 wire \cam_memory[4][0] ;
 wire \cam_memory[4][1] ;
 wire \cam_memory[4][2] ;
 wire \cam_memory[4][3] ;
 wire \cam_memory[4][4] ;
 wire \cam_memory[4][5] ;
 wire \cam_memory[4][6] ;
 wire \cam_memory[4][7] ;
 wire \cam_memory[5][0] ;
 wire \cam_memory[5][1] ;
 wire \cam_memory[5][2] ;
 wire \cam_memory[5][3] ;
 wire \cam_memory[5][4] ;
 wire \cam_memory[5][5] ;
 wire \cam_memory[5][6] ;
 wire \cam_memory[5][7] ;
 wire \cam_memory[6][0] ;
 wire \cam_memory[6][1] ;
 wire \cam_memory[6][2] ;
 wire \cam_memory[6][3] ;
 wire \cam_memory[6][4] ;
 wire \cam_memory[6][5] ;
 wire \cam_memory[6][6] ;
 wire \cam_memory[6][7] ;
 wire \cam_memory[7][0] ;
 wire \cam_memory[7][1] ;
 wire \cam_memory[7][2] ;
 wire \cam_memory[7][3] ;
 wire \cam_memory[7][4] ;
 wire \cam_memory[7][5] ;
 wire \cam_memory[7][6] ;
 wire \cam_memory[7][7] ;
 wire \cam_memory[8][0] ;
 wire \cam_memory[8][1] ;
 wire \cam_memory[8][2] ;
 wire \cam_memory[8][3] ;
 wire \cam_memory[8][4] ;
 wire \cam_memory[8][5] ;
 wire \cam_memory[8][6] ;
 wire \cam_memory[8][7] ;
 wire \cam_memory[9][0] ;
 wire \cam_memory[9][1] ;
 wire \cam_memory[9][2] ;
 wire \cam_memory[9][3] ;
 wire \cam_memory[9][4] ;
 wire \cam_memory[9][5] ;
 wire \cam_memory[9][6] ;
 wire \cam_memory[9][7] ;
 wire \valid_bits[0] ;
 wire \valid_bits[10] ;
 wire \valid_bits[11] ;
 wire \valid_bits[12] ;
 wire \valid_bits[13] ;
 wire \valid_bits[14] ;
 wire \valid_bits[15] ;
 wire \valid_bits[1] ;
 wire \valid_bits[2] ;
 wire \valid_bits[3] ;
 wire \valid_bits[4] ;
 wire \valid_bits[5] ;
 wire \valid_bits[6] ;
 wire \valid_bits[7] ;
 wire \valid_bits[8] ;
 wire \valid_bits[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 INV_X1 _0932_ (.A(net1),
    .ZN(_0920_));
 INV_X1 _0933_ (.A(net2),
    .ZN(_0921_));
 BUF_X2 _0934_ (.A(write_data[0]),
    .Z(_0231_));
 BUF_X4 _0935_ (.A(_0231_),
    .Z(_0232_));
 BUF_X4 _0936_ (.A(write_addr[3]),
    .Z(_0233_));
 BUF_X8 _0937_ (.A(write_addr[2]),
    .Z(_0234_));
 BUF_X4 _0938_ (.A(write_enable),
    .Z(_0235_));
 BUF_X4 _0939_ (.A(rst_n),
    .Z(_0236_));
 NAND3_X4 _0940_ (.A1(_0235_),
    .A2(_0236_),
    .A3(_0922_),
    .ZN(_0237_));
 NOR3_X4 _0941_ (.A1(_0233_),
    .A2(_0234_),
    .A3(_0237_),
    .ZN(_0238_));
 BUF_X2 _0942_ (.A(_0238_),
    .Z(_0239_));
 NAND2_X1 _0943_ (.A1(_0232_),
    .A2(_0239_),
    .ZN(_0240_));
 CLKBUF_X3 _0944_ (.A(_0236_),
    .Z(_0241_));
 CLKBUF_X3 _0945_ (.A(_0241_),
    .Z(_0242_));
 CLKBUF_X3 _0946_ (.A(_0242_),
    .Z(_0243_));
 NAND2_X1 _0947_ (.A1(_0243_),
    .A2(\cam_memory[0][0] ),
    .ZN(_0244_));
 OAI21_X1 _0948_ (.A(_0240_),
    .B1(_0244_),
    .B2(_0239_),
    .ZN(_0000_));
 CLKBUF_X3 _0949_ (.A(write_data[1]),
    .Z(_0245_));
 BUF_X4 _0950_ (.A(_0245_),
    .Z(_0246_));
 NAND2_X1 _0951_ (.A1(_0246_),
    .A2(_0239_),
    .ZN(_0247_));
 NAND2_X1 _0952_ (.A1(_0243_),
    .A2(\cam_memory[0][1] ),
    .ZN(_0248_));
 OAI21_X1 _0953_ (.A(_0247_),
    .B1(_0248_),
    .B2(_0239_),
    .ZN(_0001_));
 BUF_X2 _0954_ (.A(write_data[2]),
    .Z(_0249_));
 BUF_X4 _0955_ (.A(_0249_),
    .Z(_0250_));
 NAND2_X1 _0956_ (.A1(_0250_),
    .A2(_0238_),
    .ZN(_0251_));
 NAND2_X1 _0957_ (.A1(_0243_),
    .A2(\cam_memory[0][2] ),
    .ZN(_0252_));
 OAI21_X1 _0958_ (.A(_0251_),
    .B1(_0252_),
    .B2(_0239_),
    .ZN(_0002_));
 BUF_X2 _0959_ (.A(write_data[3]),
    .Z(_0253_));
 BUF_X4 _0960_ (.A(_0253_),
    .Z(_0254_));
 NAND2_X1 _0961_ (.A1(_0254_),
    .A2(_0238_),
    .ZN(_0255_));
 NAND2_X1 _0962_ (.A1(_0243_),
    .A2(\cam_memory[0][3] ),
    .ZN(_0256_));
 OAI21_X1 _0963_ (.A(_0255_),
    .B1(_0256_),
    .B2(_0239_),
    .ZN(_0003_));
 CLKBUF_X3 _0964_ (.A(write_data[4]),
    .Z(_0257_));
 BUF_X4 _0965_ (.A(_0257_),
    .Z(_0258_));
 NAND2_X1 _0966_ (.A1(_0258_),
    .A2(_0238_),
    .ZN(_0259_));
 NAND2_X1 _0967_ (.A1(_0243_),
    .A2(\cam_memory[0][4] ),
    .ZN(_0260_));
 OAI21_X1 _0968_ (.A(_0259_),
    .B1(_0260_),
    .B2(_0239_),
    .ZN(_0004_));
 BUF_X2 _0969_ (.A(write_data[5]),
    .Z(_0261_));
 BUF_X4 _0970_ (.A(_0261_),
    .Z(_0262_));
 NAND2_X1 _0971_ (.A1(_0262_),
    .A2(_0238_),
    .ZN(_0263_));
 CLKBUF_X3 _0972_ (.A(_0242_),
    .Z(_0264_));
 NAND2_X1 _0973_ (.A1(_0264_),
    .A2(\cam_memory[0][5] ),
    .ZN(_0265_));
 OAI21_X1 _0974_ (.A(_0263_),
    .B1(_0265_),
    .B2(_0239_),
    .ZN(_0005_));
 CLKBUF_X3 _0975_ (.A(write_data[6]),
    .Z(_0266_));
 BUF_X4 _0976_ (.A(_0266_),
    .Z(_0267_));
 NAND2_X1 _0977_ (.A1(_0267_),
    .A2(_0238_),
    .ZN(_0268_));
 NAND2_X1 _0978_ (.A1(_0264_),
    .A2(\cam_memory[0][6] ),
    .ZN(_0269_));
 OAI21_X1 _0979_ (.A(_0268_),
    .B1(_0269_),
    .B2(_0239_),
    .ZN(_0006_));
 CLKBUF_X3 _0980_ (.A(write_data[7]),
    .Z(_0270_));
 BUF_X4 _0981_ (.A(_0270_),
    .Z(_0271_));
 NAND2_X1 _0982_ (.A1(_0271_),
    .A2(_0238_),
    .ZN(_0272_));
 NAND2_X1 _0983_ (.A1(_0264_),
    .A2(\cam_memory[0][7] ),
    .ZN(_0273_));
 OAI21_X1 _0984_ (.A(_0272_),
    .B1(_0273_),
    .B2(_0239_),
    .ZN(_0007_));
 INV_X1 _0985_ (.A(_0234_),
    .ZN(_0274_));
 NAND2_X2 _0986_ (.A1(_0233_),
    .A2(_0274_),
    .ZN(_0275_));
 NAND3_X4 _0987_ (.A1(_0926_),
    .A2(_0235_),
    .A3(_0236_),
    .ZN(_0276_));
 NOR2_X2 _0988_ (.A1(_0275_),
    .A2(_0276_),
    .ZN(_0277_));
 BUF_X2 _0989_ (.A(_0277_),
    .Z(_0278_));
 NAND2_X1 _0990_ (.A1(_0232_),
    .A2(_0278_),
    .ZN(_0279_));
 NAND2_X1 _0991_ (.A1(_0264_),
    .A2(\cam_memory[10][0] ),
    .ZN(_0280_));
 OAI21_X1 _0992_ (.A(_0279_),
    .B1(_0280_),
    .B2(_0278_),
    .ZN(_0008_));
 NAND2_X1 _0993_ (.A1(_0246_),
    .A2(_0278_),
    .ZN(_0281_));
 NAND2_X1 _0994_ (.A1(_0264_),
    .A2(\cam_memory[10][1] ),
    .ZN(_0282_));
 OAI21_X1 _0995_ (.A(_0281_),
    .B1(_0282_),
    .B2(_0278_),
    .ZN(_0009_));
 NAND2_X1 _0996_ (.A1(_0250_),
    .A2(_0277_),
    .ZN(_0283_));
 NAND2_X1 _0997_ (.A1(_0264_),
    .A2(\cam_memory[10][2] ),
    .ZN(_0284_));
 OAI21_X1 _0998_ (.A(_0283_),
    .B1(_0284_),
    .B2(_0278_),
    .ZN(_0010_));
 NAND2_X1 _0999_ (.A1(_0254_),
    .A2(_0277_),
    .ZN(_0285_));
 NAND2_X1 _1000_ (.A1(_0264_),
    .A2(\cam_memory[10][3] ),
    .ZN(_0286_));
 OAI21_X1 _1001_ (.A(_0285_),
    .B1(_0286_),
    .B2(_0278_),
    .ZN(_0011_));
 NAND2_X1 _1002_ (.A1(_0258_),
    .A2(_0277_),
    .ZN(_0287_));
 NAND2_X1 _1003_ (.A1(_0264_),
    .A2(\cam_memory[10][4] ),
    .ZN(_0288_));
 OAI21_X1 _1004_ (.A(_0287_),
    .B1(_0288_),
    .B2(_0278_),
    .ZN(_0012_));
 NAND2_X1 _1005_ (.A1(_0262_),
    .A2(_0277_),
    .ZN(_0289_));
 NAND2_X1 _1006_ (.A1(_0264_),
    .A2(\cam_memory[10][5] ),
    .ZN(_0290_));
 OAI21_X1 _1007_ (.A(_0289_),
    .B1(_0290_),
    .B2(_0278_),
    .ZN(_0013_));
 NAND2_X1 _1008_ (.A1(_0267_),
    .A2(_0277_),
    .ZN(_0291_));
 NAND2_X1 _1009_ (.A1(_0264_),
    .A2(\cam_memory[10][6] ),
    .ZN(_0292_));
 OAI21_X1 _1010_ (.A(_0291_),
    .B1(_0292_),
    .B2(_0278_),
    .ZN(_0014_));
 NAND2_X1 _1011_ (.A1(_0271_),
    .A2(_0277_),
    .ZN(_0293_));
 CLKBUF_X3 _1012_ (.A(_0242_),
    .Z(_0294_));
 NAND2_X1 _1013_ (.A1(_0294_),
    .A2(\cam_memory[10][7] ),
    .ZN(_0295_));
 OAI21_X1 _1014_ (.A(_0293_),
    .B1(_0295_),
    .B2(_0278_),
    .ZN(_0015_));
 BUF_X2 _1015_ (.A(_0930_),
    .Z(_0296_));
 NAND3_X4 _1016_ (.A1(_0235_),
    .A2(_0236_),
    .A3(_0296_),
    .ZN(_0297_));
 NOR2_X2 _1017_ (.A1(_0275_),
    .A2(_0297_),
    .ZN(_0298_));
 BUF_X2 _1018_ (.A(_0298_),
    .Z(_0299_));
 NAND2_X1 _1019_ (.A1(_0232_),
    .A2(_0299_),
    .ZN(_0300_));
 NAND2_X1 _1020_ (.A1(_0294_),
    .A2(\cam_memory[11][0] ),
    .ZN(_0301_));
 OAI21_X1 _1021_ (.A(_0300_),
    .B1(_0301_),
    .B2(_0299_),
    .ZN(_0016_));
 NAND2_X1 _1022_ (.A1(_0246_),
    .A2(_0299_),
    .ZN(_0302_));
 NAND2_X1 _1023_ (.A1(_0294_),
    .A2(\cam_memory[11][1] ),
    .ZN(_0303_));
 OAI21_X1 _1024_ (.A(_0302_),
    .B1(_0303_),
    .B2(_0299_),
    .ZN(_0017_));
 NAND2_X1 _1025_ (.A1(_0250_),
    .A2(_0298_),
    .ZN(_0304_));
 NAND2_X1 _1026_ (.A1(_0294_),
    .A2(\cam_memory[11][2] ),
    .ZN(_0305_));
 OAI21_X1 _1027_ (.A(_0304_),
    .B1(_0305_),
    .B2(_0299_),
    .ZN(_0018_));
 NAND2_X1 _1028_ (.A1(_0254_),
    .A2(_0298_),
    .ZN(_0306_));
 NAND2_X1 _1029_ (.A1(_0294_),
    .A2(\cam_memory[11][3] ),
    .ZN(_0307_));
 OAI21_X1 _1030_ (.A(_0306_),
    .B1(_0307_),
    .B2(_0299_),
    .ZN(_0019_));
 NAND2_X1 _1031_ (.A1(_0258_),
    .A2(_0298_),
    .ZN(_0308_));
 NAND2_X1 _1032_ (.A1(_0294_),
    .A2(\cam_memory[11][4] ),
    .ZN(_0309_));
 OAI21_X1 _1033_ (.A(_0308_),
    .B1(_0309_),
    .B2(_0299_),
    .ZN(_0020_));
 NAND2_X1 _1034_ (.A1(_0262_),
    .A2(_0298_),
    .ZN(_0310_));
 NAND2_X1 _1035_ (.A1(_0294_),
    .A2(\cam_memory[11][5] ),
    .ZN(_0311_));
 OAI21_X1 _1036_ (.A(_0310_),
    .B1(_0311_),
    .B2(_0299_),
    .ZN(_0021_));
 NAND2_X1 _1037_ (.A1(_0267_),
    .A2(_0298_),
    .ZN(_0312_));
 NAND2_X1 _1038_ (.A1(_0294_),
    .A2(\cam_memory[11][6] ),
    .ZN(_0313_));
 OAI21_X1 _1039_ (.A(_0312_),
    .B1(_0313_),
    .B2(_0299_),
    .ZN(_0022_));
 NAND2_X1 _1040_ (.A1(_0271_),
    .A2(_0298_),
    .ZN(_0314_));
 NAND2_X1 _1041_ (.A1(_0294_),
    .A2(\cam_memory[11][7] ),
    .ZN(_0315_));
 OAI21_X1 _1042_ (.A(_0314_),
    .B1(_0315_),
    .B2(_0299_),
    .ZN(_0023_));
 NAND2_X4 _1043_ (.A1(_0233_),
    .A2(_0234_),
    .ZN(_0316_));
 NOR2_X2 _1044_ (.A1(_0237_),
    .A2(_0316_),
    .ZN(_0317_));
 BUF_X2 _1045_ (.A(_0317_),
    .Z(_0318_));
 NAND2_X1 _1046_ (.A1(_0232_),
    .A2(_0318_),
    .ZN(_0319_));
 NAND2_X1 _1047_ (.A1(_0294_),
    .A2(\cam_memory[12][0] ),
    .ZN(_0320_));
 OAI21_X1 _1048_ (.A(_0319_),
    .B1(_0320_),
    .B2(_0318_),
    .ZN(_0024_));
 NAND2_X1 _1049_ (.A1(_0246_),
    .A2(_0318_),
    .ZN(_0321_));
 CLKBUF_X3 _1050_ (.A(_0242_),
    .Z(_0322_));
 NAND2_X1 _1051_ (.A1(_0322_),
    .A2(\cam_memory[12][1] ),
    .ZN(_0323_));
 OAI21_X1 _1052_ (.A(_0321_),
    .B1(_0323_),
    .B2(_0318_),
    .ZN(_0025_));
 NAND2_X1 _1053_ (.A1(_0250_),
    .A2(_0317_),
    .ZN(_0324_));
 NAND2_X1 _1054_ (.A1(_0322_),
    .A2(\cam_memory[12][2] ),
    .ZN(_0325_));
 OAI21_X1 _1055_ (.A(_0324_),
    .B1(_0325_),
    .B2(_0318_),
    .ZN(_0026_));
 NAND2_X1 _1056_ (.A1(_0254_),
    .A2(_0317_),
    .ZN(_0326_));
 NAND2_X1 _1057_ (.A1(_0322_),
    .A2(\cam_memory[12][3] ),
    .ZN(_0327_));
 OAI21_X1 _1058_ (.A(_0326_),
    .B1(_0327_),
    .B2(_0318_),
    .ZN(_0027_));
 NAND2_X1 _1059_ (.A1(_0258_),
    .A2(_0317_),
    .ZN(_0328_));
 NAND2_X1 _1060_ (.A1(_0322_),
    .A2(\cam_memory[12][4] ),
    .ZN(_0329_));
 OAI21_X1 _1061_ (.A(_0328_),
    .B1(_0329_),
    .B2(_0318_),
    .ZN(_0028_));
 NAND2_X1 _1062_ (.A1(_0262_),
    .A2(_0317_),
    .ZN(_0330_));
 NAND2_X1 _1063_ (.A1(_0322_),
    .A2(\cam_memory[12][5] ),
    .ZN(_0331_));
 OAI21_X1 _1064_ (.A(_0330_),
    .B1(_0331_),
    .B2(_0318_),
    .ZN(_0029_));
 NAND2_X1 _1065_ (.A1(_0267_),
    .A2(_0317_),
    .ZN(_0332_));
 NAND2_X1 _1066_ (.A1(_0322_),
    .A2(\cam_memory[12][6] ),
    .ZN(_0333_));
 OAI21_X1 _1067_ (.A(_0332_),
    .B1(_0333_),
    .B2(_0318_),
    .ZN(_0030_));
 NAND2_X1 _1068_ (.A1(_0271_),
    .A2(_0317_),
    .ZN(_0334_));
 NAND2_X1 _1069_ (.A1(_0322_),
    .A2(\cam_memory[12][7] ),
    .ZN(_0335_));
 OAI21_X1 _1070_ (.A(_0334_),
    .B1(_0335_),
    .B2(_0318_),
    .ZN(_0031_));
 BUF_X2 _1071_ (.A(_0928_),
    .Z(_0336_));
 NAND3_X4 _1072_ (.A1(_0235_),
    .A2(_0236_),
    .A3(_0336_),
    .ZN(_0337_));
 NOR2_X4 _1073_ (.A1(_0316_),
    .A2(_0337_),
    .ZN(_0338_));
 BUF_X2 _1074_ (.A(_0338_),
    .Z(_0339_));
 NAND2_X1 _1075_ (.A1(_0232_),
    .A2(_0339_),
    .ZN(_0340_));
 NAND2_X1 _1076_ (.A1(_0322_),
    .A2(\cam_memory[13][0] ),
    .ZN(_0341_));
 OAI21_X1 _1077_ (.A(_0340_),
    .B1(_0341_),
    .B2(_0339_),
    .ZN(_0032_));
 NAND2_X1 _1078_ (.A1(_0246_),
    .A2(_0339_),
    .ZN(_0342_));
 NAND2_X1 _1079_ (.A1(_0322_),
    .A2(\cam_memory[13][1] ),
    .ZN(_0343_));
 OAI21_X1 _1080_ (.A(_0342_),
    .B1(_0343_),
    .B2(_0339_),
    .ZN(_0033_));
 NAND2_X1 _1081_ (.A1(_0250_),
    .A2(_0338_),
    .ZN(_0344_));
 NAND2_X1 _1082_ (.A1(_0322_),
    .A2(\cam_memory[13][2] ),
    .ZN(_0345_));
 OAI21_X1 _1083_ (.A(_0344_),
    .B1(_0345_),
    .B2(_0339_),
    .ZN(_0034_));
 NAND2_X1 _1084_ (.A1(_0254_),
    .A2(_0338_),
    .ZN(_0346_));
 CLKBUF_X3 _1085_ (.A(_0242_),
    .Z(_0347_));
 NAND2_X1 _1086_ (.A1(_0347_),
    .A2(\cam_memory[13][3] ),
    .ZN(_0348_));
 OAI21_X1 _1087_ (.A(_0346_),
    .B1(_0348_),
    .B2(_0339_),
    .ZN(_0035_));
 NAND2_X1 _1088_ (.A1(_0258_),
    .A2(_0338_),
    .ZN(_0349_));
 NAND2_X1 _1089_ (.A1(_0347_),
    .A2(\cam_memory[13][4] ),
    .ZN(_0350_));
 OAI21_X1 _1090_ (.A(_0349_),
    .B1(_0350_),
    .B2(_0339_),
    .ZN(_0036_));
 NAND2_X1 _1091_ (.A1(_0262_),
    .A2(_0338_),
    .ZN(_0351_));
 NAND2_X1 _1092_ (.A1(_0347_),
    .A2(\cam_memory[13][5] ),
    .ZN(_0352_));
 OAI21_X1 _1093_ (.A(_0351_),
    .B1(_0352_),
    .B2(_0339_),
    .ZN(_0037_));
 NAND2_X1 _1094_ (.A1(_0267_),
    .A2(_0338_),
    .ZN(_0353_));
 NAND2_X1 _1095_ (.A1(_0347_),
    .A2(\cam_memory[13][6] ),
    .ZN(_0354_));
 OAI21_X1 _1096_ (.A(_0353_),
    .B1(_0354_),
    .B2(_0339_),
    .ZN(_0038_));
 NAND2_X1 _1097_ (.A1(_0271_),
    .A2(_0338_),
    .ZN(_0355_));
 NAND2_X1 _1098_ (.A1(_0347_),
    .A2(\cam_memory[13][7] ),
    .ZN(_0356_));
 OAI21_X1 _1099_ (.A(_0355_),
    .B1(_0356_),
    .B2(_0339_),
    .ZN(_0039_));
 NOR2_X2 _1100_ (.A1(_0276_),
    .A2(_0316_),
    .ZN(_0357_));
 BUF_X2 _1101_ (.A(_0357_),
    .Z(_0358_));
 NAND2_X1 _1102_ (.A1(_0232_),
    .A2(_0358_),
    .ZN(_0359_));
 NAND2_X1 _1103_ (.A1(_0347_),
    .A2(\cam_memory[14][0] ),
    .ZN(_0360_));
 OAI21_X1 _1104_ (.A(_0359_),
    .B1(_0360_),
    .B2(_0358_),
    .ZN(_0040_));
 NAND2_X1 _1105_ (.A1(_0246_),
    .A2(_0358_),
    .ZN(_0361_));
 NAND2_X1 _1106_ (.A1(_0347_),
    .A2(\cam_memory[14][1] ),
    .ZN(_0362_));
 OAI21_X1 _1107_ (.A(_0361_),
    .B1(_0362_),
    .B2(_0358_),
    .ZN(_0041_));
 NAND2_X1 _1108_ (.A1(_0250_),
    .A2(_0357_),
    .ZN(_0363_));
 NAND2_X1 _1109_ (.A1(_0347_),
    .A2(\cam_memory[14][2] ),
    .ZN(_0364_));
 OAI21_X1 _1110_ (.A(_0363_),
    .B1(_0364_),
    .B2(_0358_),
    .ZN(_0042_));
 NAND2_X1 _1111_ (.A1(_0254_),
    .A2(_0357_),
    .ZN(_0365_));
 NAND2_X1 _1112_ (.A1(_0347_),
    .A2(\cam_memory[14][3] ),
    .ZN(_0366_));
 OAI21_X1 _1113_ (.A(_0365_),
    .B1(_0366_),
    .B2(_0358_),
    .ZN(_0043_));
 NAND2_X1 _1114_ (.A1(_0258_),
    .A2(_0357_),
    .ZN(_0367_));
 NAND2_X1 _1115_ (.A1(_0347_),
    .A2(\cam_memory[14][4] ),
    .ZN(_0368_));
 OAI21_X1 _1116_ (.A(_0367_),
    .B1(_0368_),
    .B2(_0358_),
    .ZN(_0044_));
 NAND2_X1 _1117_ (.A1(_0262_),
    .A2(_0357_),
    .ZN(_0369_));
 CLKBUF_X3 _1118_ (.A(_0242_),
    .Z(_0370_));
 NAND2_X1 _1119_ (.A1(_0370_),
    .A2(\cam_memory[14][5] ),
    .ZN(_0371_));
 OAI21_X1 _1120_ (.A(_0369_),
    .B1(_0371_),
    .B2(_0358_),
    .ZN(_0045_));
 NAND2_X1 _1121_ (.A1(_0267_),
    .A2(_0357_),
    .ZN(_0372_));
 NAND2_X1 _1122_ (.A1(_0370_),
    .A2(\cam_memory[14][6] ),
    .ZN(_0373_));
 OAI21_X1 _1123_ (.A(_0372_),
    .B1(_0373_),
    .B2(_0358_),
    .ZN(_0046_));
 NAND2_X1 _1124_ (.A1(_0271_),
    .A2(_0357_),
    .ZN(_0374_));
 NAND2_X1 _1125_ (.A1(_0370_),
    .A2(\cam_memory[14][7] ),
    .ZN(_0375_));
 OAI21_X1 _1126_ (.A(_0374_),
    .B1(_0375_),
    .B2(_0358_),
    .ZN(_0047_));
 NOR2_X4 _1127_ (.A1(_0297_),
    .A2(_0316_),
    .ZN(_0376_));
 BUF_X2 _1128_ (.A(_0376_),
    .Z(_0377_));
 NAND2_X1 _1129_ (.A1(_0232_),
    .A2(_0377_),
    .ZN(_0378_));
 NAND2_X1 _1130_ (.A1(_0370_),
    .A2(\cam_memory[15][0] ),
    .ZN(_0379_));
 OAI21_X1 _1131_ (.A(_0378_),
    .B1(_0379_),
    .B2(_0377_),
    .ZN(_0048_));
 NAND2_X1 _1132_ (.A1(_0246_),
    .A2(_0377_),
    .ZN(_0380_));
 NAND2_X1 _1133_ (.A1(_0370_),
    .A2(\cam_memory[15][1] ),
    .ZN(_0381_));
 OAI21_X1 _1134_ (.A(_0380_),
    .B1(_0381_),
    .B2(_0377_),
    .ZN(_0049_));
 NAND2_X1 _1135_ (.A1(_0250_),
    .A2(_0376_),
    .ZN(_0382_));
 NAND2_X1 _1136_ (.A1(_0370_),
    .A2(\cam_memory[15][2] ),
    .ZN(_0383_));
 OAI21_X1 _1137_ (.A(_0382_),
    .B1(_0383_),
    .B2(_0377_),
    .ZN(_0050_));
 NAND2_X1 _1138_ (.A1(_0254_),
    .A2(_0376_),
    .ZN(_0384_));
 NAND2_X1 _1139_ (.A1(_0370_),
    .A2(\cam_memory[15][3] ),
    .ZN(_0385_));
 OAI21_X1 _1140_ (.A(_0384_),
    .B1(_0385_),
    .B2(_0377_),
    .ZN(_0051_));
 NAND2_X1 _1141_ (.A1(_0258_),
    .A2(_0376_),
    .ZN(_0386_));
 NAND2_X1 _1142_ (.A1(_0370_),
    .A2(\cam_memory[15][4] ),
    .ZN(_0387_));
 OAI21_X1 _1143_ (.A(_0386_),
    .B1(_0387_),
    .B2(_0377_),
    .ZN(_0052_));
 NAND2_X1 _1144_ (.A1(_0262_),
    .A2(_0376_),
    .ZN(_0388_));
 NAND2_X1 _1145_ (.A1(_0370_),
    .A2(\cam_memory[15][5] ),
    .ZN(_0389_));
 OAI21_X1 _1146_ (.A(_0388_),
    .B1(_0389_),
    .B2(_0377_),
    .ZN(_0053_));
 NAND2_X1 _1147_ (.A1(_0267_),
    .A2(_0376_),
    .ZN(_0390_));
 NAND2_X1 _1148_ (.A1(_0370_),
    .A2(\cam_memory[15][6] ),
    .ZN(_0391_));
 OAI21_X1 _1149_ (.A(_0390_),
    .B1(_0391_),
    .B2(_0377_),
    .ZN(_0054_));
 NAND2_X1 _1150_ (.A1(_0271_),
    .A2(_0376_),
    .ZN(_0392_));
 CLKBUF_X3 _1151_ (.A(_0241_),
    .Z(_0393_));
 NAND2_X1 _1152_ (.A1(_0393_),
    .A2(\cam_memory[15][7] ),
    .ZN(_0394_));
 OAI21_X1 _1153_ (.A(_0392_),
    .B1(_0394_),
    .B2(_0377_),
    .ZN(_0055_));
 NOR3_X4 _1154_ (.A1(_0233_),
    .A2(_0234_),
    .A3(_0337_),
    .ZN(_0395_));
 BUF_X2 _1155_ (.A(_0395_),
    .Z(_0396_));
 NAND2_X1 _1156_ (.A1(_0232_),
    .A2(_0396_),
    .ZN(_0397_));
 NAND2_X1 _1157_ (.A1(_0393_),
    .A2(\cam_memory[1][0] ),
    .ZN(_0398_));
 OAI21_X1 _1158_ (.A(_0397_),
    .B1(_0398_),
    .B2(_0396_),
    .ZN(_0056_));
 NAND2_X1 _1159_ (.A1(_0246_),
    .A2(_0396_),
    .ZN(_0399_));
 NAND2_X1 _1160_ (.A1(_0393_),
    .A2(\cam_memory[1][1] ),
    .ZN(_0400_));
 OAI21_X1 _1161_ (.A(_0399_),
    .B1(_0400_),
    .B2(_0396_),
    .ZN(_0057_));
 NAND2_X1 _1162_ (.A1(_0250_),
    .A2(_0395_),
    .ZN(_0401_));
 NAND2_X1 _1163_ (.A1(_0393_),
    .A2(\cam_memory[1][2] ),
    .ZN(_0402_));
 OAI21_X1 _1164_ (.A(_0401_),
    .B1(_0402_),
    .B2(_0396_),
    .ZN(_0058_));
 NAND2_X1 _1165_ (.A1(_0254_),
    .A2(_0395_),
    .ZN(_0403_));
 NAND2_X1 _1166_ (.A1(_0393_),
    .A2(\cam_memory[1][3] ),
    .ZN(_0404_));
 OAI21_X1 _1167_ (.A(_0403_),
    .B1(_0404_),
    .B2(_0396_),
    .ZN(_0059_));
 NAND2_X1 _1168_ (.A1(_0258_),
    .A2(_0395_),
    .ZN(_0405_));
 NAND2_X1 _1169_ (.A1(_0393_),
    .A2(\cam_memory[1][4] ),
    .ZN(_0406_));
 OAI21_X1 _1170_ (.A(_0405_),
    .B1(_0406_),
    .B2(_0396_),
    .ZN(_0060_));
 NAND2_X1 _1171_ (.A1(_0262_),
    .A2(_0395_),
    .ZN(_0407_));
 NAND2_X1 _1172_ (.A1(_0393_),
    .A2(\cam_memory[1][5] ),
    .ZN(_0408_));
 OAI21_X1 _1173_ (.A(_0407_),
    .B1(_0408_),
    .B2(_0396_),
    .ZN(_0061_));
 NAND2_X1 _1174_ (.A1(_0267_),
    .A2(_0395_),
    .ZN(_0409_));
 NAND2_X1 _1175_ (.A1(_0393_),
    .A2(\cam_memory[1][6] ),
    .ZN(_0410_));
 OAI21_X1 _1176_ (.A(_0409_),
    .B1(_0410_),
    .B2(_0396_),
    .ZN(_0062_));
 NAND2_X1 _1177_ (.A1(_0271_),
    .A2(_0395_),
    .ZN(_0411_));
 NAND2_X1 _1178_ (.A1(_0393_),
    .A2(\cam_memory[1][7] ),
    .ZN(_0412_));
 OAI21_X1 _1179_ (.A(_0411_),
    .B1(_0412_),
    .B2(_0396_),
    .ZN(_0063_));
 NOR3_X4 _1180_ (.A1(_0233_),
    .A2(_0234_),
    .A3(_0276_),
    .ZN(_0413_));
 BUF_X2 _1181_ (.A(_0413_),
    .Z(_0414_));
 NAND2_X1 _1182_ (.A1(_0232_),
    .A2(_0414_),
    .ZN(_0415_));
 NAND2_X1 _1183_ (.A1(_0393_),
    .A2(\cam_memory[2][0] ),
    .ZN(_0416_));
 OAI21_X1 _1184_ (.A(_0415_),
    .B1(_0416_),
    .B2(_0414_),
    .ZN(_0064_));
 NAND2_X1 _1185_ (.A1(_0246_),
    .A2(_0414_),
    .ZN(_0417_));
 CLKBUF_X3 _1186_ (.A(_0241_),
    .Z(_0418_));
 NAND2_X1 _1187_ (.A1(_0418_),
    .A2(\cam_memory[2][1] ),
    .ZN(_0419_));
 OAI21_X1 _1188_ (.A(_0417_),
    .B1(_0419_),
    .B2(_0414_),
    .ZN(_0065_));
 NAND2_X1 _1189_ (.A1(_0250_),
    .A2(_0413_),
    .ZN(_0420_));
 NAND2_X1 _1190_ (.A1(_0418_),
    .A2(\cam_memory[2][2] ),
    .ZN(_0421_));
 OAI21_X1 _1191_ (.A(_0420_),
    .B1(_0421_),
    .B2(_0414_),
    .ZN(_0066_));
 NAND2_X1 _1192_ (.A1(_0254_),
    .A2(_0413_),
    .ZN(_0422_));
 NAND2_X1 _1193_ (.A1(_0418_),
    .A2(\cam_memory[2][3] ),
    .ZN(_0423_));
 OAI21_X1 _1194_ (.A(_0422_),
    .B1(_0423_),
    .B2(_0414_),
    .ZN(_0067_));
 NAND2_X1 _1195_ (.A1(_0258_),
    .A2(_0413_),
    .ZN(_0424_));
 NAND2_X1 _1196_ (.A1(_0418_),
    .A2(\cam_memory[2][4] ),
    .ZN(_0425_));
 OAI21_X1 _1197_ (.A(_0424_),
    .B1(_0425_),
    .B2(_0414_),
    .ZN(_0068_));
 NAND2_X1 _1198_ (.A1(_0262_),
    .A2(_0413_),
    .ZN(_0426_));
 NAND2_X1 _1199_ (.A1(_0418_),
    .A2(\cam_memory[2][5] ),
    .ZN(_0427_));
 OAI21_X1 _1200_ (.A(_0426_),
    .B1(_0427_),
    .B2(_0414_),
    .ZN(_0069_));
 NAND2_X1 _1201_ (.A1(_0267_),
    .A2(_0413_),
    .ZN(_0428_));
 NAND2_X1 _1202_ (.A1(_0418_),
    .A2(\cam_memory[2][6] ),
    .ZN(_0429_));
 OAI21_X1 _1203_ (.A(_0428_),
    .B1(_0429_),
    .B2(_0414_),
    .ZN(_0070_));
 NAND2_X1 _1204_ (.A1(_0271_),
    .A2(_0413_),
    .ZN(_0430_));
 NAND2_X1 _1205_ (.A1(_0418_),
    .A2(\cam_memory[2][7] ),
    .ZN(_0431_));
 OAI21_X1 _1206_ (.A(_0430_),
    .B1(_0431_),
    .B2(_0414_),
    .ZN(_0071_));
 NOR3_X4 _1207_ (.A1(_0233_),
    .A2(_0234_),
    .A3(_0297_),
    .ZN(_0432_));
 BUF_X2 _1208_ (.A(_0432_),
    .Z(_0433_));
 NAND2_X1 _1209_ (.A1(_0232_),
    .A2(_0433_),
    .ZN(_0434_));
 NAND2_X1 _1210_ (.A1(_0418_),
    .A2(\cam_memory[3][0] ),
    .ZN(_0435_));
 OAI21_X1 _1211_ (.A(_0434_),
    .B1(_0435_),
    .B2(_0433_),
    .ZN(_0072_));
 NAND2_X1 _1212_ (.A1(_0246_),
    .A2(_0433_),
    .ZN(_0436_));
 NAND2_X1 _1213_ (.A1(_0418_),
    .A2(\cam_memory[3][1] ),
    .ZN(_0437_));
 OAI21_X1 _1214_ (.A(_0436_),
    .B1(_0437_),
    .B2(_0433_),
    .ZN(_0073_));
 NAND2_X1 _1215_ (.A1(_0250_),
    .A2(_0432_),
    .ZN(_0438_));
 NAND2_X1 _1216_ (.A1(_0418_),
    .A2(\cam_memory[3][2] ),
    .ZN(_0439_));
 OAI21_X1 _1217_ (.A(_0438_),
    .B1(_0439_),
    .B2(_0433_),
    .ZN(_0074_));
 NAND2_X1 _1218_ (.A1(_0254_),
    .A2(_0432_),
    .ZN(_0440_));
 CLKBUF_X3 _1219_ (.A(_0241_),
    .Z(_0441_));
 NAND2_X1 _1220_ (.A1(_0441_),
    .A2(\cam_memory[3][3] ),
    .ZN(_0442_));
 OAI21_X1 _1221_ (.A(_0440_),
    .B1(_0442_),
    .B2(_0433_),
    .ZN(_0075_));
 NAND2_X1 _1222_ (.A1(_0258_),
    .A2(_0432_),
    .ZN(_0443_));
 NAND2_X1 _1223_ (.A1(_0441_),
    .A2(\cam_memory[3][4] ),
    .ZN(_0444_));
 OAI21_X1 _1224_ (.A(_0443_),
    .B1(_0444_),
    .B2(_0433_),
    .ZN(_0076_));
 NAND2_X1 _1225_ (.A1(_0262_),
    .A2(_0432_),
    .ZN(_0445_));
 NAND2_X1 _1226_ (.A1(_0441_),
    .A2(\cam_memory[3][5] ),
    .ZN(_0446_));
 OAI21_X1 _1227_ (.A(_0445_),
    .B1(_0446_),
    .B2(_0433_),
    .ZN(_0077_));
 NAND2_X1 _1228_ (.A1(_0267_),
    .A2(_0432_),
    .ZN(_0447_));
 NAND2_X1 _1229_ (.A1(_0441_),
    .A2(\cam_memory[3][6] ),
    .ZN(_0448_));
 OAI21_X1 _1230_ (.A(_0447_),
    .B1(_0448_),
    .B2(_0433_),
    .ZN(_0078_));
 NAND2_X1 _1231_ (.A1(_0271_),
    .A2(_0432_),
    .ZN(_0449_));
 NAND2_X1 _1232_ (.A1(_0441_),
    .A2(\cam_memory[3][7] ),
    .ZN(_0450_));
 OAI21_X1 _1233_ (.A(_0449_),
    .B1(_0450_),
    .B2(_0433_),
    .ZN(_0079_));
 INV_X2 _1234_ (.A(_0233_),
    .ZN(_0451_));
 NAND2_X4 _1235_ (.A1(_0451_),
    .A2(_0234_),
    .ZN(_0452_));
 NOR2_X4 _1236_ (.A1(_0237_),
    .A2(_0452_),
    .ZN(_0453_));
 BUF_X2 _1237_ (.A(_0453_),
    .Z(_0454_));
 NAND2_X1 _1238_ (.A1(_0231_),
    .A2(_0454_),
    .ZN(_0455_));
 NAND2_X1 _1239_ (.A1(_0441_),
    .A2(\cam_memory[4][0] ),
    .ZN(_0456_));
 OAI21_X1 _1240_ (.A(_0455_),
    .B1(_0456_),
    .B2(_0454_),
    .ZN(_0080_));
 NAND2_X1 _1241_ (.A1(_0245_),
    .A2(_0454_),
    .ZN(_0457_));
 NAND2_X1 _1242_ (.A1(_0441_),
    .A2(\cam_memory[4][1] ),
    .ZN(_0458_));
 OAI21_X1 _1243_ (.A(_0457_),
    .B1(_0458_),
    .B2(_0454_),
    .ZN(_0081_));
 NAND2_X1 _1244_ (.A1(_0249_),
    .A2(_0453_),
    .ZN(_0459_));
 NAND2_X1 _1245_ (.A1(_0441_),
    .A2(\cam_memory[4][2] ),
    .ZN(_0460_));
 OAI21_X1 _1246_ (.A(_0459_),
    .B1(_0460_),
    .B2(_0454_),
    .ZN(_0082_));
 NAND2_X1 _1247_ (.A1(_0253_),
    .A2(_0453_),
    .ZN(_0461_));
 NAND2_X1 _1248_ (.A1(_0441_),
    .A2(\cam_memory[4][3] ),
    .ZN(_0462_));
 OAI21_X1 _1249_ (.A(_0461_),
    .B1(_0462_),
    .B2(_0454_),
    .ZN(_0083_));
 NAND2_X1 _1250_ (.A1(_0257_),
    .A2(_0453_),
    .ZN(_0463_));
 NAND2_X1 _1251_ (.A1(_0441_),
    .A2(\cam_memory[4][4] ),
    .ZN(_0464_));
 OAI21_X1 _1252_ (.A(_0463_),
    .B1(_0464_),
    .B2(_0454_),
    .ZN(_0084_));
 NAND2_X1 _1253_ (.A1(_0261_),
    .A2(_0453_),
    .ZN(_0465_));
 CLKBUF_X3 _1254_ (.A(_0241_),
    .Z(_0466_));
 NAND2_X1 _1255_ (.A1(_0466_),
    .A2(\cam_memory[4][5] ),
    .ZN(_0467_));
 OAI21_X1 _1256_ (.A(_0465_),
    .B1(_0467_),
    .B2(_0454_),
    .ZN(_0085_));
 NAND2_X1 _1257_ (.A1(_0266_),
    .A2(_0453_),
    .ZN(_0468_));
 NAND2_X1 _1258_ (.A1(_0466_),
    .A2(\cam_memory[4][6] ),
    .ZN(_0469_));
 OAI21_X1 _1259_ (.A(_0468_),
    .B1(_0469_),
    .B2(_0454_),
    .ZN(_0086_));
 NAND2_X1 _1260_ (.A1(_0270_),
    .A2(_0453_),
    .ZN(_0470_));
 NAND2_X1 _1261_ (.A1(_0466_),
    .A2(\cam_memory[4][7] ),
    .ZN(_0471_));
 OAI21_X1 _1262_ (.A(_0470_),
    .B1(_0471_),
    .B2(_0454_),
    .ZN(_0087_));
 NOR2_X4 _1263_ (.A1(_0337_),
    .A2(_0452_),
    .ZN(_0472_));
 BUF_X2 _1264_ (.A(_0472_),
    .Z(_0473_));
 NAND2_X1 _1265_ (.A1(_0231_),
    .A2(_0473_),
    .ZN(_0474_));
 NAND2_X1 _1266_ (.A1(_0466_),
    .A2(\cam_memory[5][0] ),
    .ZN(_0475_));
 OAI21_X1 _1267_ (.A(_0474_),
    .B1(_0475_),
    .B2(_0473_),
    .ZN(_0088_));
 NAND2_X1 _1268_ (.A1(_0245_),
    .A2(_0473_),
    .ZN(_0476_));
 NAND2_X1 _1269_ (.A1(_0466_),
    .A2(\cam_memory[5][1] ),
    .ZN(_0477_));
 OAI21_X1 _1270_ (.A(_0476_),
    .B1(_0477_),
    .B2(_0473_),
    .ZN(_0089_));
 NAND2_X1 _1271_ (.A1(_0249_),
    .A2(_0472_),
    .ZN(_0478_));
 NAND2_X1 _1272_ (.A1(_0466_),
    .A2(\cam_memory[5][2] ),
    .ZN(_0479_));
 OAI21_X1 _1273_ (.A(_0478_),
    .B1(_0479_),
    .B2(_0473_),
    .ZN(_0090_));
 NAND2_X1 _1274_ (.A1(_0253_),
    .A2(_0472_),
    .ZN(_0480_));
 NAND2_X1 _1275_ (.A1(_0466_),
    .A2(\cam_memory[5][3] ),
    .ZN(_0481_));
 OAI21_X1 _1276_ (.A(_0480_),
    .B1(_0481_),
    .B2(_0473_),
    .ZN(_0091_));
 NAND2_X1 _1277_ (.A1(_0257_),
    .A2(_0472_),
    .ZN(_0482_));
 NAND2_X1 _1278_ (.A1(_0466_),
    .A2(\cam_memory[5][4] ),
    .ZN(_0483_));
 OAI21_X1 _1279_ (.A(_0482_),
    .B1(_0483_),
    .B2(_0473_),
    .ZN(_0092_));
 NAND2_X1 _1280_ (.A1(_0261_),
    .A2(_0472_),
    .ZN(_0484_));
 NAND2_X1 _1281_ (.A1(_0466_),
    .A2(\cam_memory[5][5] ),
    .ZN(_0485_));
 OAI21_X1 _1282_ (.A(_0484_),
    .B1(_0485_),
    .B2(_0473_),
    .ZN(_0093_));
 NAND2_X1 _1283_ (.A1(_0266_),
    .A2(_0472_),
    .ZN(_0486_));
 NAND2_X1 _1284_ (.A1(_0466_),
    .A2(\cam_memory[5][6] ),
    .ZN(_0487_));
 OAI21_X1 _1285_ (.A(_0486_),
    .B1(_0487_),
    .B2(_0473_),
    .ZN(_0094_));
 NAND2_X1 _1286_ (.A1(_0270_),
    .A2(_0472_),
    .ZN(_0488_));
 BUF_X2 _1287_ (.A(_0241_),
    .Z(_0489_));
 NAND2_X1 _1288_ (.A1(_0489_),
    .A2(\cam_memory[5][7] ),
    .ZN(_0490_));
 OAI21_X1 _1289_ (.A(_0488_),
    .B1(_0490_),
    .B2(_0473_),
    .ZN(_0095_));
 NOR2_X4 _1290_ (.A1(_0276_),
    .A2(_0452_),
    .ZN(_0491_));
 BUF_X2 _1291_ (.A(_0491_),
    .Z(_0492_));
 NAND2_X1 _1292_ (.A1(_0231_),
    .A2(_0492_),
    .ZN(_0493_));
 NAND2_X1 _1293_ (.A1(_0489_),
    .A2(\cam_memory[6][0] ),
    .ZN(_0494_));
 OAI21_X1 _1294_ (.A(_0493_),
    .B1(_0494_),
    .B2(_0492_),
    .ZN(_0096_));
 NAND2_X1 _1295_ (.A1(_0245_),
    .A2(_0492_),
    .ZN(_0495_));
 NAND2_X1 _1296_ (.A1(_0489_),
    .A2(\cam_memory[6][1] ),
    .ZN(_0496_));
 OAI21_X1 _1297_ (.A(_0495_),
    .B1(_0496_),
    .B2(_0492_),
    .ZN(_0097_));
 NAND2_X1 _1298_ (.A1(_0249_),
    .A2(_0491_),
    .ZN(_0497_));
 NAND2_X1 _1299_ (.A1(_0489_),
    .A2(\cam_memory[6][2] ),
    .ZN(_0498_));
 OAI21_X1 _1300_ (.A(_0497_),
    .B1(_0498_),
    .B2(_0492_),
    .ZN(_0098_));
 NAND2_X1 _1301_ (.A1(_0253_),
    .A2(_0491_),
    .ZN(_0499_));
 NAND2_X1 _1302_ (.A1(_0489_),
    .A2(\cam_memory[6][3] ),
    .ZN(_0500_));
 OAI21_X1 _1303_ (.A(_0499_),
    .B1(_0500_),
    .B2(_0492_),
    .ZN(_0099_));
 NAND2_X1 _1304_ (.A1(_0257_),
    .A2(_0491_),
    .ZN(_0501_));
 NAND2_X1 _1305_ (.A1(_0489_),
    .A2(\cam_memory[6][4] ),
    .ZN(_0502_));
 OAI21_X1 _1306_ (.A(_0501_),
    .B1(_0502_),
    .B2(_0492_),
    .ZN(_0100_));
 NAND2_X1 _1307_ (.A1(_0261_),
    .A2(_0491_),
    .ZN(_0503_));
 NAND2_X1 _1308_ (.A1(_0489_),
    .A2(\cam_memory[6][5] ),
    .ZN(_0504_));
 OAI21_X1 _1309_ (.A(_0503_),
    .B1(_0504_),
    .B2(_0492_),
    .ZN(_0101_));
 NAND2_X1 _1310_ (.A1(_0266_),
    .A2(_0491_),
    .ZN(_0505_));
 NAND2_X1 _1311_ (.A1(_0489_),
    .A2(\cam_memory[6][6] ),
    .ZN(_0506_));
 OAI21_X1 _1312_ (.A(_0505_),
    .B1(_0506_),
    .B2(_0492_),
    .ZN(_0102_));
 NAND2_X1 _1313_ (.A1(_0270_),
    .A2(_0491_),
    .ZN(_0507_));
 NAND2_X1 _1314_ (.A1(_0489_),
    .A2(\cam_memory[6][7] ),
    .ZN(_0508_));
 OAI21_X1 _1315_ (.A(_0507_),
    .B1(_0508_),
    .B2(_0492_),
    .ZN(_0103_));
 NOR2_X4 _1316_ (.A1(_0297_),
    .A2(_0452_),
    .ZN(_0509_));
 BUF_X2 _1317_ (.A(_0509_),
    .Z(_0510_));
 NAND2_X1 _1318_ (.A1(_0231_),
    .A2(_0510_),
    .ZN(_0511_));
 NAND2_X1 _1319_ (.A1(_0489_),
    .A2(\cam_memory[7][0] ),
    .ZN(_0512_));
 OAI21_X1 _1320_ (.A(_0511_),
    .B1(_0512_),
    .B2(_0510_),
    .ZN(_0104_));
 NAND2_X1 _1321_ (.A1(_0245_),
    .A2(_0510_),
    .ZN(_0513_));
 CLKBUF_X3 _1322_ (.A(_0241_),
    .Z(_0514_));
 NAND2_X1 _1323_ (.A1(_0514_),
    .A2(\cam_memory[7][1] ),
    .ZN(_0515_));
 OAI21_X1 _1324_ (.A(_0513_),
    .B1(_0515_),
    .B2(_0510_),
    .ZN(_0105_));
 NAND2_X1 _1325_ (.A1(_0249_),
    .A2(_0509_),
    .ZN(_0516_));
 NAND2_X1 _1326_ (.A1(_0514_),
    .A2(\cam_memory[7][2] ),
    .ZN(_0517_));
 OAI21_X1 _1327_ (.A(_0516_),
    .B1(_0517_),
    .B2(_0510_),
    .ZN(_0106_));
 NAND2_X1 _1328_ (.A1(_0253_),
    .A2(_0509_),
    .ZN(_0518_));
 NAND2_X1 _1329_ (.A1(_0514_),
    .A2(\cam_memory[7][3] ),
    .ZN(_0519_));
 OAI21_X1 _1330_ (.A(_0518_),
    .B1(_0519_),
    .B2(_0510_),
    .ZN(_0107_));
 NAND2_X1 _1331_ (.A1(_0257_),
    .A2(_0509_),
    .ZN(_0520_));
 NAND2_X1 _1332_ (.A1(_0514_),
    .A2(\cam_memory[7][4] ),
    .ZN(_0521_));
 OAI21_X1 _1333_ (.A(_0520_),
    .B1(_0521_),
    .B2(_0510_),
    .ZN(_0108_));
 NAND2_X1 _1334_ (.A1(_0261_),
    .A2(_0509_),
    .ZN(_0522_));
 NAND2_X1 _1335_ (.A1(_0514_),
    .A2(\cam_memory[7][5] ),
    .ZN(_0523_));
 OAI21_X1 _1336_ (.A(_0522_),
    .B1(_0523_),
    .B2(_0510_),
    .ZN(_0109_));
 NAND2_X1 _1337_ (.A1(_0266_),
    .A2(_0509_),
    .ZN(_0524_));
 NAND2_X1 _1338_ (.A1(_0514_),
    .A2(\cam_memory[7][6] ),
    .ZN(_0525_));
 OAI21_X1 _1339_ (.A(_0524_),
    .B1(_0525_),
    .B2(_0510_),
    .ZN(_0110_));
 NAND2_X1 _1340_ (.A1(_0270_),
    .A2(_0509_),
    .ZN(_0526_));
 NAND2_X1 _1341_ (.A1(_0514_),
    .A2(\cam_memory[7][7] ),
    .ZN(_0527_));
 OAI21_X1 _1342_ (.A(_0526_),
    .B1(_0527_),
    .B2(_0510_),
    .ZN(_0111_));
 NOR2_X2 _1343_ (.A1(_0237_),
    .A2(_0275_),
    .ZN(_0528_));
 BUF_X2 _1344_ (.A(_0528_),
    .Z(_0529_));
 NAND2_X1 _1345_ (.A1(_0231_),
    .A2(_0529_),
    .ZN(_0530_));
 NAND2_X1 _1346_ (.A1(_0514_),
    .A2(\cam_memory[8][0] ),
    .ZN(_0531_));
 OAI21_X1 _1347_ (.A(_0530_),
    .B1(_0531_),
    .B2(_0529_),
    .ZN(_0112_));
 NAND2_X1 _1348_ (.A1(_0245_),
    .A2(_0529_),
    .ZN(_0532_));
 NAND2_X1 _1349_ (.A1(_0514_),
    .A2(\cam_memory[8][1] ),
    .ZN(_0533_));
 OAI21_X1 _1350_ (.A(_0532_),
    .B1(_0533_),
    .B2(_0529_),
    .ZN(_0113_));
 NAND2_X1 _1351_ (.A1(_0249_),
    .A2(_0528_),
    .ZN(_0534_));
 NAND2_X1 _1352_ (.A1(_0514_),
    .A2(\cam_memory[8][2] ),
    .ZN(_0535_));
 OAI21_X1 _1353_ (.A(_0534_),
    .B1(_0535_),
    .B2(_0529_),
    .ZN(_0114_));
 NAND2_X1 _1354_ (.A1(_0253_),
    .A2(_0528_),
    .ZN(_0536_));
 CLKBUF_X3 _1355_ (.A(_0241_),
    .Z(_0537_));
 NAND2_X1 _1356_ (.A1(_0537_),
    .A2(\cam_memory[8][3] ),
    .ZN(_0538_));
 OAI21_X1 _1357_ (.A(_0536_),
    .B1(_0538_),
    .B2(_0529_),
    .ZN(_0115_));
 NAND2_X1 _1358_ (.A1(_0257_),
    .A2(_0528_),
    .ZN(_0539_));
 NAND2_X1 _1359_ (.A1(_0537_),
    .A2(\cam_memory[8][4] ),
    .ZN(_0540_));
 OAI21_X1 _1360_ (.A(_0539_),
    .B1(_0540_),
    .B2(_0529_),
    .ZN(_0116_));
 NAND2_X1 _1361_ (.A1(_0261_),
    .A2(_0528_),
    .ZN(_0541_));
 NAND2_X1 _1362_ (.A1(_0537_),
    .A2(\cam_memory[8][5] ),
    .ZN(_0542_));
 OAI21_X1 _1363_ (.A(_0541_),
    .B1(_0542_),
    .B2(_0529_),
    .ZN(_0117_));
 NAND2_X1 _1364_ (.A1(_0266_),
    .A2(_0528_),
    .ZN(_0543_));
 NAND2_X1 _1365_ (.A1(_0537_),
    .A2(\cam_memory[8][6] ),
    .ZN(_0544_));
 OAI21_X1 _1366_ (.A(_0543_),
    .B1(_0544_),
    .B2(_0529_),
    .ZN(_0118_));
 NAND2_X1 _1367_ (.A1(_0270_),
    .A2(_0528_),
    .ZN(_0545_));
 NAND2_X1 _1368_ (.A1(_0537_),
    .A2(\cam_memory[8][7] ),
    .ZN(_0546_));
 OAI21_X1 _1369_ (.A(_0545_),
    .B1(_0546_),
    .B2(_0529_),
    .ZN(_0119_));
 NOR2_X2 _1370_ (.A1(_0275_),
    .A2(_0337_),
    .ZN(_0547_));
 BUF_X2 _1371_ (.A(_0547_),
    .Z(_0548_));
 NAND2_X1 _1372_ (.A1(_0231_),
    .A2(_0548_),
    .ZN(_0549_));
 NAND2_X1 _1373_ (.A1(_0537_),
    .A2(\cam_memory[9][0] ),
    .ZN(_0550_));
 OAI21_X1 _1374_ (.A(_0549_),
    .B1(_0550_),
    .B2(_0548_),
    .ZN(_0120_));
 NAND2_X1 _1375_ (.A1(_0245_),
    .A2(_0548_),
    .ZN(_0551_));
 NAND2_X1 _1376_ (.A1(_0537_),
    .A2(\cam_memory[9][1] ),
    .ZN(_0552_));
 OAI21_X1 _1377_ (.A(_0551_),
    .B1(_0552_),
    .B2(_0548_),
    .ZN(_0121_));
 NAND2_X1 _1378_ (.A1(_0249_),
    .A2(_0547_),
    .ZN(_0553_));
 NAND2_X1 _1379_ (.A1(_0537_),
    .A2(\cam_memory[9][2] ),
    .ZN(_0554_));
 OAI21_X1 _1380_ (.A(_0553_),
    .B1(_0554_),
    .B2(_0548_),
    .ZN(_0122_));
 NAND2_X1 _1381_ (.A1(_0253_),
    .A2(_0547_),
    .ZN(_0555_));
 NAND2_X1 _1382_ (.A1(_0537_),
    .A2(\cam_memory[9][3] ),
    .ZN(_0556_));
 OAI21_X1 _1383_ (.A(_0555_),
    .B1(_0556_),
    .B2(_0548_),
    .ZN(_0123_));
 NAND2_X1 _1384_ (.A1(_0257_),
    .A2(_0547_),
    .ZN(_0557_));
 NAND2_X1 _1385_ (.A1(_0537_),
    .A2(\cam_memory[9][4] ),
    .ZN(_0558_));
 OAI21_X1 _1386_ (.A(_0557_),
    .B1(_0558_),
    .B2(_0548_),
    .ZN(_0124_));
 NAND2_X1 _1387_ (.A1(_0261_),
    .A2(_0547_),
    .ZN(_0559_));
 NAND2_X1 _1388_ (.A1(_0242_),
    .A2(\cam_memory[9][5] ),
    .ZN(_0560_));
 OAI21_X1 _1389_ (.A(_0559_),
    .B1(_0560_),
    .B2(_0548_),
    .ZN(_0125_));
 NAND2_X1 _1390_ (.A1(_0266_),
    .A2(_0547_),
    .ZN(_0561_));
 NAND2_X1 _1391_ (.A1(_0242_),
    .A2(\cam_memory[9][6] ),
    .ZN(_0562_));
 OAI21_X1 _1392_ (.A(_0561_),
    .B1(_0562_),
    .B2(_0548_),
    .ZN(_0126_));
 NAND2_X1 _1393_ (.A1(_0270_),
    .A2(_0547_),
    .ZN(_0563_));
 NAND2_X1 _1394_ (.A1(_0242_),
    .A2(\cam_memory[9][7] ),
    .ZN(_0564_));
 OAI21_X1 _1395_ (.A(_0563_),
    .B1(_0564_),
    .B2(_0548_),
    .ZN(_0127_));
 CLKBUF_X2 _1396_ (.A(compare_enable),
    .Z(_0565_));
 AND2_X1 _1397_ (.A1(_0241_),
    .A2(_0565_),
    .ZN(_0133_));
 BUF_X4 _1398_ (.A(compare_data[0]),
    .Z(_0566_));
 BUF_X4 _1399_ (.A(_0566_),
    .Z(_0567_));
 XNOR2_X1 _1400_ (.A(_0567_),
    .B(\cam_memory[14][0] ),
    .ZN(_0568_));
 BUF_X4 _1401_ (.A(compare_data[6]),
    .Z(_0569_));
 XOR2_X1 _1402_ (.A(_0569_),
    .B(\cam_memory[14][6] ),
    .Z(_0570_));
 BUF_X4 _1403_ (.A(compare_data[3]),
    .Z(_0571_));
 XOR2_X1 _1404_ (.A(_0571_),
    .B(\cam_memory[14][3] ),
    .Z(_0572_));
 BUF_X4 _1405_ (.A(compare_data[7]),
    .Z(_0573_));
 XOR2_X1 _1406_ (.A(_0573_),
    .B(\cam_memory[14][7] ),
    .Z(_0574_));
 NOR3_X1 _1407_ (.A1(_0570_),
    .A2(_0572_),
    .A3(_0574_),
    .ZN(_0575_));
 BUF_X4 _1408_ (.A(compare_data[2]),
    .Z(_0576_));
 BUF_X8 _1409_ (.A(_0576_),
    .Z(_0577_));
 XOR2_X1 _1410_ (.A(_0577_),
    .B(\cam_memory[14][2] ),
    .Z(_0578_));
 BUF_X8 _1411_ (.A(compare_data[1]),
    .Z(_0579_));
 XOR2_X1 _1412_ (.A(_0579_),
    .B(\cam_memory[14][1] ),
    .Z(_0580_));
 BUF_X8 _1413_ (.A(compare_data[4]),
    .Z(_0581_));
 XOR2_X1 _1414_ (.A(_0581_),
    .B(\cam_memory[14][4] ),
    .Z(_0582_));
 BUF_X4 _1415_ (.A(compare_data[5]),
    .Z(_0583_));
 XOR2_X1 _1416_ (.A(_0583_),
    .B(\cam_memory[14][5] ),
    .Z(_0584_));
 NOR4_X1 _1417_ (.A1(_0578_),
    .A2(_0580_),
    .A3(_0582_),
    .A4(_0584_),
    .ZN(_0585_));
 AND4_X2 _1418_ (.A1(\valid_bits[14] ),
    .A2(_0568_),
    .A3(_0575_),
    .A4(_0585_),
    .ZN(_0586_));
 XNOR2_X1 _1419_ (.A(_0567_),
    .B(\cam_memory[15][0] ),
    .ZN(_0587_));
 XOR2_X1 _1420_ (.A(_0569_),
    .B(\cam_memory[15][6] ),
    .Z(_0588_));
 XOR2_X1 _1421_ (.A(_0571_),
    .B(\cam_memory[15][3] ),
    .Z(_0589_));
 XOR2_X1 _1422_ (.A(_0573_),
    .B(\cam_memory[15][7] ),
    .Z(_0590_));
 NOR3_X1 _1423_ (.A1(_0588_),
    .A2(_0589_),
    .A3(_0590_),
    .ZN(_0591_));
 XOR2_X1 _1424_ (.A(_0576_),
    .B(\cam_memory[15][2] ),
    .Z(_0592_));
 XOR2_X1 _1425_ (.A(_0579_),
    .B(\cam_memory[15][1] ),
    .Z(_0593_));
 XOR2_X1 _1426_ (.A(_0581_),
    .B(\cam_memory[15][4] ),
    .Z(_0594_));
 XOR2_X1 _1427_ (.A(_0583_),
    .B(\cam_memory[15][5] ),
    .Z(_0595_));
 NOR4_X1 _1428_ (.A1(_0592_),
    .A2(_0593_),
    .A3(_0594_),
    .A4(_0595_),
    .ZN(_0596_));
 AND4_X2 _1429_ (.A1(\valid_bits[15] ),
    .A2(_0587_),
    .A3(_0591_),
    .A4(_0596_),
    .ZN(_0597_));
 XNOR2_X1 _1430_ (.A(_0567_),
    .B(\cam_memory[12][0] ),
    .ZN(_0598_));
 XOR2_X2 _1431_ (.A(_0569_),
    .B(\cam_memory[12][6] ),
    .Z(_0599_));
 XOR2_X2 _1432_ (.A(_0583_),
    .B(\cam_memory[12][5] ),
    .Z(_0600_));
 XOR2_X2 _1433_ (.A(_0573_),
    .B(\cam_memory[12][7] ),
    .Z(_0601_));
 NOR3_X2 _1434_ (.A1(_0599_),
    .A2(_0600_),
    .A3(_0601_),
    .ZN(_0602_));
 XOR2_X2 _1435_ (.A(_0581_),
    .B(\cam_memory[12][4] ),
    .Z(_0603_));
 XOR2_X2 _1436_ (.A(_0576_),
    .B(\cam_memory[12][2] ),
    .Z(_0604_));
 XOR2_X2 _1437_ (.A(_0571_),
    .B(\cam_memory[12][3] ),
    .Z(_0605_));
 XOR2_X2 _1438_ (.A(_0579_),
    .B(\cam_memory[12][1] ),
    .Z(_0606_));
 NOR4_X2 _1439_ (.A1(_0603_),
    .A2(_0604_),
    .A3(_0605_),
    .A4(_0606_),
    .ZN(_0607_));
 AND4_X1 _1440_ (.A1(\valid_bits[12] ),
    .A2(_0598_),
    .A3(_0602_),
    .A4(_0607_),
    .ZN(_0608_));
 XNOR2_X1 _1441_ (.A(_0566_),
    .B(\cam_memory[13][0] ),
    .ZN(_0609_));
 XOR2_X1 _1442_ (.A(_0569_),
    .B(\cam_memory[13][6] ),
    .Z(_0610_));
 XOR2_X1 _1443_ (.A(_0583_),
    .B(\cam_memory[13][5] ),
    .Z(_0611_));
 XOR2_X1 _1444_ (.A(_0573_),
    .B(\cam_memory[13][7] ),
    .Z(_0612_));
 NOR3_X1 _1445_ (.A1(_0610_),
    .A2(_0611_),
    .A3(_0612_),
    .ZN(_0613_));
 XOR2_X1 _1446_ (.A(_0581_),
    .B(\cam_memory[13][4] ),
    .Z(_0614_));
 XOR2_X1 _1447_ (.A(_0576_),
    .B(\cam_memory[13][2] ),
    .Z(_0615_));
 XOR2_X1 _1448_ (.A(_0571_),
    .B(\cam_memory[13][3] ),
    .Z(_0616_));
 XOR2_X1 _1449_ (.A(_0579_),
    .B(\cam_memory[13][1] ),
    .Z(_0617_));
 NOR4_X1 _1450_ (.A1(_0614_),
    .A2(_0615_),
    .A3(_0616_),
    .A4(_0617_),
    .ZN(_0618_));
 AND4_X1 _1451_ (.A1(\valid_bits[13] ),
    .A2(_0609_),
    .A3(_0613_),
    .A4(_0618_),
    .ZN(_0619_));
 NOR4_X2 _1452_ (.A1(_0586_),
    .A2(_0597_),
    .A3(_0608_),
    .A4(_0619_),
    .ZN(_0620_));
 XNOR2_X1 _1453_ (.A(_0567_),
    .B(\cam_memory[10][0] ),
    .ZN(_0621_));
 BUF_X8 _1454_ (.A(_0583_),
    .Z(_0622_));
 XOR2_X2 _1455_ (.A(_0622_),
    .B(\cam_memory[10][5] ),
    .Z(_0623_));
 BUF_X16 _1456_ (.A(_0581_),
    .Z(_0624_));
 XOR2_X2 _1457_ (.A(_0624_),
    .B(\cam_memory[10][4] ),
    .Z(_0625_));
 BUF_X8 _1458_ (.A(_0573_),
    .Z(_0626_));
 XOR2_X2 _1459_ (.A(_0626_),
    .B(\cam_memory[10][7] ),
    .Z(_0627_));
 NOR3_X2 _1460_ (.A1(_0623_),
    .A2(_0625_),
    .A3(_0627_),
    .ZN(_0628_));
 BUF_X16 _1461_ (.A(_0571_),
    .Z(_0629_));
 XOR2_X2 _1462_ (.A(_0629_),
    .B(\cam_memory[10][3] ),
    .Z(_0630_));
 XOR2_X2 _1463_ (.A(_0579_),
    .B(\cam_memory[10][1] ),
    .Z(_0631_));
 XOR2_X2 _1464_ (.A(_0576_),
    .B(\cam_memory[10][2] ),
    .Z(_0632_));
 XOR2_X2 _1465_ (.A(_0569_),
    .B(\cam_memory[10][6] ),
    .Z(_0633_));
 NOR4_X2 _1466_ (.A1(_0630_),
    .A2(_0631_),
    .A3(_0632_),
    .A4(_0633_),
    .ZN(_0634_));
 AND4_X1 _1467_ (.A1(\valid_bits[10] ),
    .A2(_0621_),
    .A3(_0628_),
    .A4(_0634_),
    .ZN(_0635_));
 BUF_X16 _1468_ (.A(_0579_),
    .Z(_0636_));
 XNOR2_X1 _1469_ (.A(_0636_),
    .B(\cam_memory[11][1] ),
    .ZN(_0637_));
 BUF_X8 _1470_ (.A(_0569_),
    .Z(_0638_));
 XOR2_X1 _1471_ (.A(_0638_),
    .B(\cam_memory[11][6] ),
    .Z(_0639_));
 XOR2_X1 _1472_ (.A(_0583_),
    .B(\cam_memory[11][5] ),
    .Z(_0640_));
 XOR2_X1 _1473_ (.A(_0573_),
    .B(\cam_memory[11][7] ),
    .Z(_0641_));
 NOR3_X1 _1474_ (.A1(_0639_),
    .A2(_0640_),
    .A3(_0641_),
    .ZN(_0642_));
 XOR2_X1 _1475_ (.A(_0629_),
    .B(\cam_memory[11][3] ),
    .Z(_0643_));
 XOR2_X1 _1476_ (.A(_0566_),
    .B(\cam_memory[11][0] ),
    .Z(_0644_));
 XOR2_X1 _1477_ (.A(_0576_),
    .B(\cam_memory[11][2] ),
    .Z(_0645_));
 XOR2_X1 _1478_ (.A(_0581_),
    .B(\cam_memory[11][4] ),
    .Z(_0646_));
 NOR4_X1 _1479_ (.A1(_0643_),
    .A2(_0644_),
    .A3(_0645_),
    .A4(_0646_),
    .ZN(_0647_));
 AND4_X1 _1480_ (.A1(\valid_bits[11] ),
    .A2(_0637_),
    .A3(_0642_),
    .A4(_0647_),
    .ZN(_0648_));
 XNOR2_X1 _1481_ (.A(_0636_),
    .B(\cam_memory[9][1] ),
    .ZN(_0649_));
 XNOR2_X1 _1482_ (.A(_0626_),
    .B(\cam_memory[9][7] ),
    .ZN(_0650_));
 XNOR2_X1 _1483_ (.A(_0629_),
    .B(\cam_memory[9][3] ),
    .ZN(_0651_));
 NAND3_X1 _1484_ (.A1(_0649_),
    .A2(_0650_),
    .A3(_0651_),
    .ZN(_0652_));
 XNOR2_X1 _1485_ (.A(_0622_),
    .B(\cam_memory[9][5] ),
    .ZN(_0653_));
 XNOR2_X1 _1486_ (.A(_0577_),
    .B(\cam_memory[9][2] ),
    .ZN(_0654_));
 XNOR2_X1 _1487_ (.A(_0566_),
    .B(\cam_memory[9][0] ),
    .ZN(_0655_));
 XNOR2_X1 _1488_ (.A(_0624_),
    .B(\cam_memory[9][4] ),
    .ZN(_0656_));
 NAND4_X1 _1489_ (.A1(_0653_),
    .A2(_0654_),
    .A3(_0655_),
    .A4(_0656_),
    .ZN(_0657_));
 XNOR2_X1 _1490_ (.A(_0638_),
    .B(\cam_memory[9][6] ),
    .ZN(_0658_));
 NAND2_X1 _1491_ (.A1(\valid_bits[9] ),
    .A2(_0658_),
    .ZN(_0659_));
 XNOR2_X1 _1492_ (.A(_0577_),
    .B(\cam_memory[8][2] ),
    .ZN(_0660_));
 XNOR2_X1 _1493_ (.A(_0638_),
    .B(\cam_memory[8][6] ),
    .ZN(_0661_));
 XNOR2_X1 _1494_ (.A(_0583_),
    .B(\cam_memory[8][5] ),
    .ZN(_0662_));
 NAND3_X1 _1495_ (.A1(_0660_),
    .A2(_0661_),
    .A3(_0662_),
    .ZN(_0663_));
 XNOR2_X1 _1496_ (.A(_0573_),
    .B(\cam_memory[8][7] ),
    .ZN(_0664_));
 XNOR2_X1 _1497_ (.A(_0624_),
    .B(\cam_memory[8][4] ),
    .ZN(_0665_));
 XNOR2_X1 _1498_ (.A(_0571_),
    .B(\cam_memory[8][3] ),
    .ZN(_0666_));
 XNOR2_X1 _1499_ (.A(_0566_),
    .B(\cam_memory[8][0] ),
    .ZN(_0667_));
 NAND4_X2 _1500_ (.A1(_0664_),
    .A2(_0665_),
    .A3(_0666_),
    .A4(_0667_),
    .ZN(_0668_));
 XNOR2_X1 _1501_ (.A(_0636_),
    .B(\cam_memory[8][1] ),
    .ZN(_0669_));
 NAND2_X1 _1502_ (.A1(\valid_bits[8] ),
    .A2(_0669_),
    .ZN(_0670_));
 OAI33_X1 _1503_ (.A1(_0652_),
    .A2(_0657_),
    .A3(_0659_),
    .B1(_0663_),
    .B2(_0668_),
    .B3(_0670_),
    .ZN(_0671_));
 NOR3_X1 _1504_ (.A1(_0635_),
    .A2(_0648_),
    .A3(_0671_),
    .ZN(_0672_));
 NAND2_X1 _1505_ (.A1(_0620_),
    .A2(_0672_),
    .ZN(_0673_));
 XNOR2_X1 _1506_ (.A(_0567_),
    .B(\cam_memory[7][0] ),
    .ZN(_0674_));
 NAND2_X1 _1507_ (.A1(\valid_bits[7] ),
    .A2(_0674_),
    .ZN(_0675_));
 XNOR2_X1 _1508_ (.A(_0622_),
    .B(\cam_memory[7][5] ),
    .ZN(_0676_));
 XNOR2_X1 _1509_ (.A(_0638_),
    .B(\cam_memory[7][6] ),
    .ZN(_0677_));
 XNOR2_X1 _1510_ (.A(_0629_),
    .B(\cam_memory[7][3] ),
    .ZN(_0678_));
 NAND3_X1 _1511_ (.A1(_0676_),
    .A2(_0677_),
    .A3(_0678_),
    .ZN(_0679_));
 XNOR2_X1 _1512_ (.A(_0626_),
    .B(\cam_memory[7][7] ),
    .ZN(_0680_));
 XNOR2_X1 _1513_ (.A(_0636_),
    .B(\cam_memory[7][1] ),
    .ZN(_0681_));
 XNOR2_X1 _1514_ (.A(_0624_),
    .B(\cam_memory[7][4] ),
    .ZN(_0682_));
 XNOR2_X1 _1515_ (.A(_0577_),
    .B(\cam_memory[7][2] ),
    .ZN(_0683_));
 NAND4_X1 _1516_ (.A1(_0680_),
    .A2(_0681_),
    .A3(_0682_),
    .A4(_0683_),
    .ZN(_0684_));
 NOR3_X2 _1517_ (.A1(_0675_),
    .A2(_0679_),
    .A3(_0684_),
    .ZN(_0685_));
 XNOR2_X1 _1518_ (.A(_0567_),
    .B(\cam_memory[6][0] ),
    .ZN(_0686_));
 XOR2_X1 _1519_ (.A(_0577_),
    .B(\cam_memory[6][2] ),
    .Z(_0687_));
 XOR2_X1 _1520_ (.A(_0636_),
    .B(\cam_memory[6][1] ),
    .Z(_0688_));
 XOR2_X1 _1521_ (.A(_0571_),
    .B(\cam_memory[6][3] ),
    .Z(_0689_));
 XOR2_X1 _1522_ (.A(_0581_),
    .B(\cam_memory[6][4] ),
    .Z(_0690_));
 NOR4_X1 _1523_ (.A1(_0687_),
    .A2(_0688_),
    .A3(_0689_),
    .A4(_0690_),
    .ZN(_0691_));
 AND3_X1 _1524_ (.A1(\valid_bits[6] ),
    .A2(_0686_),
    .A3(_0691_),
    .ZN(_0692_));
 XOR2_X2 _1525_ (.A(_0638_),
    .B(\cam_memory[6][6] ),
    .Z(_0693_));
 XOR2_X2 _1526_ (.A(_0622_),
    .B(\cam_memory[6][5] ),
    .Z(_0694_));
 XOR2_X2 _1527_ (.A(_0626_),
    .B(\cam_memory[6][7] ),
    .Z(_0695_));
 NOR3_X2 _1528_ (.A1(_0693_),
    .A2(_0694_),
    .A3(_0695_),
    .ZN(_0696_));
 AOI21_X2 _1529_ (.A(_0685_),
    .B1(_0692_),
    .B2(_0696_),
    .ZN(_0697_));
 XNOR2_X1 _1530_ (.A(_0567_),
    .B(\cam_memory[4][0] ),
    .ZN(_0698_));
 XOR2_X2 _1531_ (.A(_0622_),
    .B(\cam_memory[4][5] ),
    .Z(_0699_));
 XOR2_X2 _1532_ (.A(_0624_),
    .B(\cam_memory[4][4] ),
    .Z(_0700_));
 XOR2_X2 _1533_ (.A(_0626_),
    .B(\cam_memory[4][7] ),
    .Z(_0701_));
 NOR3_X2 _1534_ (.A1(_0699_),
    .A2(_0700_),
    .A3(_0701_),
    .ZN(_0702_));
 XOR2_X2 _1535_ (.A(_0629_),
    .B(\cam_memory[4][3] ),
    .Z(_0703_));
 XOR2_X2 _1536_ (.A(_0579_),
    .B(\cam_memory[4][1] ),
    .Z(_0704_));
 XOR2_X2 _1537_ (.A(_0576_),
    .B(\cam_memory[4][2] ),
    .Z(_0705_));
 XOR2_X2 _1538_ (.A(_0569_),
    .B(\cam_memory[4][6] ),
    .Z(_0706_));
 NOR4_X2 _1539_ (.A1(_0703_),
    .A2(_0704_),
    .A3(_0705_),
    .A4(_0706_),
    .ZN(_0707_));
 AND4_X1 _1540_ (.A1(\valid_bits[4] ),
    .A2(_0698_),
    .A3(_0702_),
    .A4(_0707_),
    .ZN(_0708_));
 XNOR2_X1 _1541_ (.A(_0629_),
    .B(\cam_memory[5][3] ),
    .ZN(_0709_));
 NAND2_X1 _1542_ (.A1(\valid_bits[5] ),
    .A2(_0709_),
    .ZN(_0710_));
 XNOR2_X1 _1543_ (.A(_0626_),
    .B(\cam_memory[5][7] ),
    .ZN(_0711_));
 XNOR2_X1 _1544_ (.A(_0624_),
    .B(\cam_memory[5][4] ),
    .ZN(_0712_));
 XNOR2_X1 _1545_ (.A(_0638_),
    .B(\cam_memory[5][6] ),
    .ZN(_0713_));
 NAND3_X1 _1546_ (.A1(_0711_),
    .A2(_0712_),
    .A3(_0713_),
    .ZN(_0714_));
 XNOR2_X1 _1547_ (.A(_0622_),
    .B(\cam_memory[5][5] ),
    .ZN(_0715_));
 XNOR2_X1 _1548_ (.A(_0566_),
    .B(\cam_memory[5][0] ),
    .ZN(_0716_));
 XNOR2_X1 _1549_ (.A(_0577_),
    .B(\cam_memory[5][2] ),
    .ZN(_0717_));
 XNOR2_X1 _1550_ (.A(_0636_),
    .B(\cam_memory[5][1] ),
    .ZN(_0718_));
 NAND4_X1 _1551_ (.A1(_0715_),
    .A2(_0716_),
    .A3(_0717_),
    .A4(_0718_),
    .ZN(_0719_));
 NOR3_X1 _1552_ (.A1(_0710_),
    .A2(_0714_),
    .A3(_0719_),
    .ZN(_0720_));
 NOR2_X1 _1553_ (.A1(_0708_),
    .A2(_0720_),
    .ZN(_0721_));
 XNOR2_X1 _1554_ (.A(_0636_),
    .B(\cam_memory[3][1] ),
    .ZN(_0722_));
 XOR2_X1 _1555_ (.A(_0638_),
    .B(\cam_memory[3][6] ),
    .Z(_0723_));
 XOR2_X1 _1556_ (.A(_0622_),
    .B(\cam_memory[3][5] ),
    .Z(_0724_));
 XOR2_X1 _1557_ (.A(_0626_),
    .B(\cam_memory[3][7] ),
    .Z(_0725_));
 NOR3_X1 _1558_ (.A1(_0723_),
    .A2(_0724_),
    .A3(_0725_),
    .ZN(_0726_));
 XOR2_X1 _1559_ (.A(_0629_),
    .B(\cam_memory[3][3] ),
    .Z(_0727_));
 XOR2_X1 _1560_ (.A(_0566_),
    .B(\cam_memory[3][0] ),
    .Z(_0728_));
 XOR2_X1 _1561_ (.A(_0577_),
    .B(\cam_memory[3][2] ),
    .Z(_0729_));
 XOR2_X1 _1562_ (.A(_0624_),
    .B(\cam_memory[3][4] ),
    .Z(_0730_));
 NOR4_X1 _1563_ (.A1(_0727_),
    .A2(_0728_),
    .A3(_0729_),
    .A4(_0730_),
    .ZN(_0731_));
 AND4_X1 _1564_ (.A1(\valid_bits[3] ),
    .A2(_0722_),
    .A3(_0726_),
    .A4(_0731_),
    .ZN(_0732_));
 XNOR2_X1 _1565_ (.A(_0567_),
    .B(\cam_memory[2][0] ),
    .ZN(_0733_));
 XOR2_X1 _1566_ (.A(_0638_),
    .B(\cam_memory[2][6] ),
    .Z(_0734_));
 XOR2_X1 _1567_ (.A(_0622_),
    .B(\cam_memory[2][5] ),
    .Z(_0735_));
 NOR2_X1 _1568_ (.A1(_0734_),
    .A2(_0735_),
    .ZN(_0736_));
 XOR2_X1 _1569_ (.A(_0626_),
    .B(\cam_memory[2][7] ),
    .Z(_0737_));
 XOR2_X1 _1570_ (.A(_0624_),
    .B(\cam_memory[2][4] ),
    .Z(_0738_));
 XOR2_X1 _1571_ (.A(_0577_),
    .B(\cam_memory[2][2] ),
    .Z(_0739_));
 XOR2_X1 _1572_ (.A(_0629_),
    .B(\cam_memory[2][3] ),
    .Z(_0740_));
 NOR4_X1 _1573_ (.A1(_0737_),
    .A2(_0738_),
    .A3(_0739_),
    .A4(_0740_),
    .ZN(_0741_));
 AND3_X1 _1574_ (.A1(_0733_),
    .A2(_0736_),
    .A3(_0741_),
    .ZN(_0742_));
 XNOR2_X1 _1575_ (.A(_0636_),
    .B(\cam_memory[2][1] ),
    .ZN(_0743_));
 AND2_X1 _1576_ (.A1(\valid_bits[2] ),
    .A2(_0743_),
    .ZN(_0744_));
 AOI21_X1 _1577_ (.A(_0732_),
    .B1(_0742_),
    .B2(_0744_),
    .ZN(_0745_));
 XNOR2_X1 _1578_ (.A(_0577_),
    .B(\cam_memory[1][2] ),
    .ZN(_0746_));
 XNOR2_X1 _1579_ (.A(_0638_),
    .B(\cam_memory[1][6] ),
    .ZN(_0747_));
 XNOR2_X1 _1580_ (.A(_0622_),
    .B(\cam_memory[1][5] ),
    .ZN(_0748_));
 NAND3_X1 _1581_ (.A1(_0746_),
    .A2(_0747_),
    .A3(_0748_),
    .ZN(_0749_));
 XNOR2_X1 _1582_ (.A(_0626_),
    .B(\cam_memory[1][7] ),
    .ZN(_0750_));
 XNOR2_X1 _1583_ (.A(_0624_),
    .B(\cam_memory[1][4] ),
    .ZN(_0751_));
 XNOR2_X1 _1584_ (.A(_0629_),
    .B(\cam_memory[1][3] ),
    .ZN(_0752_));
 XNOR2_X1 _1585_ (.A(_0567_),
    .B(\cam_memory[1][0] ),
    .ZN(_0753_));
 NAND4_X1 _1586_ (.A1(_0750_),
    .A2(_0751_),
    .A3(_0752_),
    .A4(_0753_),
    .ZN(_0754_));
 XNOR2_X1 _1587_ (.A(_0636_),
    .B(\cam_memory[1][1] ),
    .ZN(_0755_));
 NAND2_X1 _1588_ (.A1(\valid_bits[1] ),
    .A2(_0755_),
    .ZN(_0756_));
 XNOR2_X1 _1589_ (.A(\cam_memory[0][0] ),
    .B(_0567_),
    .ZN(_0757_));
 XNOR2_X1 _1590_ (.A(\cam_memory[0][4] ),
    .B(_0624_),
    .ZN(_0758_));
 XNOR2_X1 _1591_ (.A(\cam_memory[0][6] ),
    .B(_0638_),
    .ZN(_0759_));
 NAND3_X1 _1592_ (.A1(_0757_),
    .A2(_0758_),
    .A3(_0759_),
    .ZN(_0760_));
 XNOR2_X1 _1593_ (.A(\cam_memory[0][7] ),
    .B(_0626_),
    .ZN(_0761_));
 XNOR2_X1 _1594_ (.A(\cam_memory[0][5] ),
    .B(_0622_),
    .ZN(_0762_));
 XNOR2_X1 _1595_ (.A(\cam_memory[0][3] ),
    .B(_0629_),
    .ZN(_0763_));
 XNOR2_X1 _1596_ (.A(\cam_memory[0][1] ),
    .B(_0636_),
    .ZN(_0764_));
 NAND4_X1 _1597_ (.A1(_0761_),
    .A2(_0762_),
    .A3(_0763_),
    .A4(_0764_),
    .ZN(_0765_));
 XNOR2_X1 _1598_ (.A(\cam_memory[0][2] ),
    .B(_0577_),
    .ZN(_0766_));
 NAND2_X1 _1599_ (.A1(\valid_bits[0] ),
    .A2(_0766_),
    .ZN(_0767_));
 OAI33_X1 _1600_ (.A1(_0749_),
    .A2(_0754_),
    .A3(_0756_),
    .B1(_0760_),
    .B2(_0765_),
    .B3(_0767_),
    .ZN(_0768_));
 INV_X1 _1601_ (.A(_0768_),
    .ZN(_0769_));
 NAND4_X1 _1602_ (.A1(_0697_),
    .A2(_0721_),
    .A3(_0745_),
    .A4(_0769_),
    .ZN(_0150_));
 OAI21_X1 _1603_ (.A(_0133_),
    .B1(_0673_),
    .B2(_0150_),
    .ZN(_0151_));
 INV_X1 _1604_ (.A(_0151_),
    .ZN(_0128_));
 INV_X1 _1605_ (.A(_0241_),
    .ZN(_0152_));
 NOR2_X1 _1606_ (.A1(_0152_),
    .A2(_0565_),
    .ZN(_0153_));
 NAND2_X1 _1607_ (.A1(net4),
    .A2(_0153_),
    .ZN(_0154_));
 NAND4_X2 _1608_ (.A1(\valid_bits[12] ),
    .A2(_0598_),
    .A3(_0602_),
    .A4(_0607_),
    .ZN(_0155_));
 NAND4_X2 _1609_ (.A1(\valid_bits[10] ),
    .A2(_0621_),
    .A3(_0628_),
    .A4(_0634_),
    .ZN(_0156_));
 NOR3_X1 _1610_ (.A1(_0652_),
    .A2(_0657_),
    .A3(_0659_),
    .ZN(_0157_));
 NAND3_X1 _1611_ (.A1(_0155_),
    .A2(_0156_),
    .A3(_0157_),
    .ZN(_0158_));
 AOI21_X1 _1612_ (.A(_0619_),
    .B1(_0648_),
    .B2(_0155_),
    .ZN(_0159_));
 AOI21_X1 _1613_ (.A(_0586_),
    .B1(_0158_),
    .B2(_0159_),
    .ZN(_0160_));
 NOR3_X1 _1614_ (.A1(_0663_),
    .A2(_0668_),
    .A3(_0670_),
    .ZN(_0161_));
 NAND4_X1 _1615_ (.A1(\valid_bits[6] ),
    .A2(_0686_),
    .A3(_0696_),
    .A4(_0691_),
    .ZN(_0162_));
 NOR2_X1 _1616_ (.A1(_0162_),
    .A2(_0685_),
    .ZN(_0163_));
 NAND2_X1 _1617_ (.A1(_0155_),
    .A2(_0156_),
    .ZN(_0164_));
 NOR4_X2 _1618_ (.A1(_0586_),
    .A2(_0161_),
    .A3(_0163_),
    .A4(_0164_),
    .ZN(_0165_));
 NAND4_X2 _1619_ (.A1(\valid_bits[4] ),
    .A2(_0698_),
    .A3(_0702_),
    .A4(_0707_),
    .ZN(_0166_));
 NAND4_X1 _1620_ (.A1(_0733_),
    .A2(_0736_),
    .A3(_0741_),
    .A4(_0744_),
    .ZN(_0167_));
 NOR3_X1 _1621_ (.A1(_0749_),
    .A2(_0754_),
    .A3(_0756_),
    .ZN(_0168_));
 OR3_X1 _1622_ (.A1(_0760_),
    .A2(_0765_),
    .A3(_0767_),
    .ZN(_0169_));
 OAI211_X2 _1623_ (.A(_0166_),
    .B(_0167_),
    .C1(_0168_),
    .C2(_0169_),
    .ZN(_0170_));
 NAND3_X1 _1624_ (.A1(_0674_),
    .A2(_0677_),
    .A3(_0678_),
    .ZN(_0171_));
 NAND4_X1 _1625_ (.A1(_0676_),
    .A2(_0681_),
    .A3(_0682_),
    .A4(_0683_),
    .ZN(_0172_));
 NAND2_X1 _1626_ (.A1(\valid_bits[7] ),
    .A2(_0680_),
    .ZN(_0173_));
 NAND3_X1 _1627_ (.A1(_0709_),
    .A2(_0712_),
    .A3(_0713_),
    .ZN(_0174_));
 NAND4_X1 _1628_ (.A1(_0711_),
    .A2(_0715_),
    .A3(_0716_),
    .A4(_0717_),
    .ZN(_0175_));
 NAND2_X1 _1629_ (.A1(\valid_bits[5] ),
    .A2(_0718_),
    .ZN(_0176_));
 OAI33_X1 _1630_ (.A1(_0171_),
    .A2(_0172_),
    .A3(_0173_),
    .B1(_0174_),
    .B2(_0175_),
    .B3(_0176_),
    .ZN(_0177_));
 AOI21_X1 _1631_ (.A(_0177_),
    .B1(_0732_),
    .B2(_0166_),
    .ZN(_0178_));
 NAND2_X1 _1632_ (.A1(_0170_),
    .A2(_0178_),
    .ZN(_0179_));
 AOI211_X2 _1633_ (.A(_0597_),
    .B(_0160_),
    .C1(_0165_),
    .C2(_0179_),
    .ZN(_0180_));
 OAI21_X1 _1634_ (.A(_0154_),
    .B1(_0180_),
    .B2(_0151_),
    .ZN(_0129_));
 NAND2_X1 _1635_ (.A1(net5),
    .A2(_0153_),
    .ZN(_0181_));
 NOR2_X1 _1636_ (.A1(_0608_),
    .A2(_0619_),
    .ZN(_0182_));
 OR3_X1 _1637_ (.A1(_0671_),
    .A2(_0708_),
    .A3(_0720_),
    .ZN(_0183_));
 AOI21_X1 _1638_ (.A(_0183_),
    .B1(_0768_),
    .B2(_0745_),
    .ZN(_0184_));
 NOR2_X1 _1639_ (.A1(_0635_),
    .A2(_0648_),
    .ZN(_0185_));
 OAI21_X1 _1640_ (.A(_0185_),
    .B1(_0671_),
    .B2(_0697_),
    .ZN(_0186_));
 OAI21_X1 _1641_ (.A(_0182_),
    .B1(_0184_),
    .B2(_0186_),
    .ZN(_0187_));
 NOR2_X1 _1642_ (.A1(_0586_),
    .A2(_0597_),
    .ZN(_0188_));
 AND2_X1 _1643_ (.A1(_0188_),
    .A2(_0181_),
    .ZN(_0189_));
 AOI22_X1 _1644_ (.A1(_0151_),
    .A2(_0181_),
    .B1(_0187_),
    .B2(_0189_),
    .ZN(_0130_));
 OAI21_X1 _1645_ (.A(_0242_),
    .B1(_0565_),
    .B2(net6),
    .ZN(_0190_));
 INV_X1 _1646_ (.A(_0620_),
    .ZN(_0191_));
 NAND2_X1 _1647_ (.A1(_0697_),
    .A2(_0721_),
    .ZN(_0192_));
 AOI21_X1 _1648_ (.A(_0191_),
    .B1(_0672_),
    .B2(_0192_),
    .ZN(_0193_));
 AOI21_X1 _1649_ (.A(_0190_),
    .B1(_0193_),
    .B2(_0565_),
    .ZN(_0131_));
 MUX2_X1 _1650_ (.A(net7),
    .B(_0673_),
    .S(_0565_),
    .Z(_0194_));
 AND2_X1 _1651_ (.A1(_0243_),
    .A2(_0194_),
    .ZN(_0132_));
 NOR3_X4 _1652_ (.A1(_0234_),
    .A2(net1),
    .A3(net2),
    .ZN(_0195_));
 XNOR2_X2 _1653_ (.A(_0233_),
    .B(_0195_),
    .ZN(_0196_));
 NAND3_X1 _1654_ (.A1(_0451_),
    .A2(_0274_),
    .A3(_0922_),
    .ZN(_0197_));
 NOR2_X2 _1655_ (.A1(net1),
    .A2(_0923_),
    .ZN(_0198_));
 NAND2_X1 _1656_ (.A1(_0235_),
    .A2(_0198_),
    .ZN(_0199_));
 NOR3_X1 _1657_ (.A1(_0196_),
    .A2(_0197_),
    .A3(_0199_),
    .ZN(_0200_));
 OAI21_X1 _1658_ (.A(_0243_),
    .B1(\valid_bits[0] ),
    .B2(_0200_),
    .ZN(_0201_));
 INV_X1 _1659_ (.A(_0201_),
    .ZN(_0134_));
 CLKBUF_X3 _1660_ (.A(_0152_),
    .Z(_0202_));
 XNOR2_X1 _1661_ (.A(_0234_),
    .B(_0922_),
    .ZN(_0203_));
 NAND2_X1 _1662_ (.A1(_0235_),
    .A2(_0203_),
    .ZN(_0204_));
 NOR2_X1 _1663_ (.A1(_0196_),
    .A2(_0204_),
    .ZN(_0205_));
 AOI21_X1 _1664_ (.A(\valid_bits[10] ),
    .B1(_0924_),
    .B2(_0205_),
    .ZN(_0206_));
 NOR2_X1 _1665_ (.A1(_0202_),
    .A2(_0206_),
    .ZN(_0135_));
 AOI21_X1 _1666_ (.A(\valid_bits[11] ),
    .B1(_0296_),
    .B2(_0205_),
    .ZN(_0207_));
 NOR2_X1 _1667_ (.A1(_0202_),
    .A2(_0207_),
    .ZN(_0136_));
 AOI21_X1 _1668_ (.A(\valid_bits[12] ),
    .B1(_0198_),
    .B2(_0205_),
    .ZN(_0208_));
 NOR2_X1 _1669_ (.A1(_0202_),
    .A2(_0208_),
    .ZN(_0137_));
 INV_X1 _1670_ (.A(_0203_),
    .ZN(_0209_));
 NAND2_X1 _1671_ (.A1(_0235_),
    .A2(_0209_),
    .ZN(_0210_));
 NOR2_X1 _1672_ (.A1(_0196_),
    .A2(_0210_),
    .ZN(_0211_));
 AOI21_X1 _1673_ (.A(\valid_bits[13] ),
    .B1(_0336_),
    .B2(_0211_),
    .ZN(_0212_));
 NOR2_X1 _1674_ (.A1(_0202_),
    .A2(_0212_),
    .ZN(_0138_));
 AOI21_X1 _1675_ (.A(\valid_bits[14] ),
    .B1(_0924_),
    .B2(_0211_),
    .ZN(_0213_));
 NOR2_X1 _1676_ (.A1(_0202_),
    .A2(_0213_),
    .ZN(_0139_));
 AOI21_X1 _1677_ (.A(\valid_bits[15] ),
    .B1(_0296_),
    .B2(_0211_),
    .ZN(_0214_));
 NOR2_X1 _1678_ (.A1(_0202_),
    .A2(_0214_),
    .ZN(_0140_));
 XNOR2_X2 _1679_ (.A(_0451_),
    .B(_0195_),
    .ZN(_0215_));
 NAND3_X1 _1680_ (.A1(_0235_),
    .A2(_0336_),
    .A3(_0203_),
    .ZN(_0216_));
 NOR2_X1 _1681_ (.A1(_0215_),
    .A2(_0216_),
    .ZN(_0217_));
 OAI21_X1 _1682_ (.A(_0243_),
    .B1(\valid_bits[1] ),
    .B2(_0217_),
    .ZN(_0218_));
 INV_X1 _1683_ (.A(_0218_),
    .ZN(_0141_));
 NOR2_X1 _1684_ (.A1(_0215_),
    .A2(_0204_),
    .ZN(_0219_));
 AOI21_X1 _1685_ (.A(\valid_bits[2] ),
    .B1(_0924_),
    .B2(_0219_),
    .ZN(_0220_));
 NOR2_X1 _1686_ (.A1(_0202_),
    .A2(_0220_),
    .ZN(_0142_));
 AOI21_X1 _1687_ (.A(\valid_bits[3] ),
    .B1(_0296_),
    .B2(_0219_),
    .ZN(_0221_));
 NOR2_X1 _1688_ (.A1(_0202_),
    .A2(_0221_),
    .ZN(_0143_));
 AOI21_X1 _1689_ (.A(\valid_bits[4] ),
    .B1(_0198_),
    .B2(_0219_),
    .ZN(_0222_));
 NOR2_X1 _1690_ (.A1(_0202_),
    .A2(_0222_),
    .ZN(_0144_));
 NOR2_X1 _1691_ (.A1(_0215_),
    .A2(_0210_),
    .ZN(_0223_));
 AOI21_X1 _1692_ (.A(\valid_bits[5] ),
    .B1(_0336_),
    .B2(_0223_),
    .ZN(_0224_));
 NOR2_X1 _1693_ (.A1(_0202_),
    .A2(_0224_),
    .ZN(_0145_));
 AOI21_X1 _1694_ (.A(\valid_bits[6] ),
    .B1(_0924_),
    .B2(_0223_),
    .ZN(_0225_));
 NOR2_X1 _1695_ (.A1(_0152_),
    .A2(_0225_),
    .ZN(_0146_));
 AOI21_X1 _1696_ (.A(\valid_bits[7] ),
    .B1(_0296_),
    .B2(_0223_),
    .ZN(_0226_));
 NOR2_X1 _1697_ (.A1(_0152_),
    .A2(_0226_),
    .ZN(_0147_));
 AND3_X1 _1698_ (.A1(_0197_),
    .A2(_0198_),
    .A3(_0223_),
    .ZN(_0227_));
 OAI21_X1 _1699_ (.A(_0243_),
    .B1(\valid_bits[8] ),
    .B2(_0227_),
    .ZN(_0228_));
 INV_X1 _1700_ (.A(_0228_),
    .ZN(_0148_));
 NOR2_X1 _1701_ (.A1(_0196_),
    .A2(_0216_),
    .ZN(_0229_));
 OAI21_X1 _1702_ (.A(_0243_),
    .B1(\valid_bits[9] ),
    .B2(_0229_),
    .ZN(_0230_));
 INV_X1 _1703_ (.A(_0230_),
    .ZN(_0149_));
 HA_X1 _1704_ (.A(_0920_),
    .B(_0921_),
    .CO(_0922_),
    .S(_0923_));
 HA_X1 _1705_ (.A(_0920_),
    .B(net2),
    .CO(_0924_),
    .S(_0925_));
 HA_X1 _1706_ (.A(_0920_),
    .B(net2),
    .CO(_0926_),
    .S(_0927_));
 HA_X1 _1707_ (.A(net1),
    .B(_0921_),
    .CO(_0928_),
    .S(_0929_));
 HA_X1 _1708_ (.A(net1),
    .B(net2),
    .CO(_0930_),
    .S(_0931_));
 DFF_X1 \cam_memory[0][0]$_SDFFCE_PN0P_  (.D(_0000_),
    .CK(clknet_4_8_0_clk),
    .Q(\cam_memory[0][0] ),
    .QN(_0919_));
 DFF_X1 \cam_memory[0][1]$_SDFFCE_PN0P_  (.D(_0001_),
    .CK(clknet_4_8_0_clk),
    .Q(\cam_memory[0][1] ),
    .QN(_0918_));
 DFF_X1 \cam_memory[0][2]$_SDFFCE_PN0P_  (.D(_0002_),
    .CK(clknet_4_8_0_clk),
    .Q(\cam_memory[0][2] ),
    .QN(_0917_));
 DFF_X1 \cam_memory[0][3]$_SDFFCE_PN0P_  (.D(_0003_),
    .CK(clknet_4_8_0_clk),
    .Q(\cam_memory[0][3] ),
    .QN(_0916_));
 DFF_X1 \cam_memory[0][4]$_SDFFCE_PN0P_  (.D(_0004_),
    .CK(clknet_4_8_0_clk),
    .Q(\cam_memory[0][4] ),
    .QN(_0915_));
 DFF_X1 \cam_memory[0][5]$_SDFFCE_PN0P_  (.D(_0005_),
    .CK(clknet_4_8_0_clk),
    .Q(\cam_memory[0][5] ),
    .QN(_0914_));
 DFF_X1 \cam_memory[0][6]$_SDFFCE_PN0P_  (.D(_0006_),
    .CK(clknet_4_8_0_clk),
    .Q(\cam_memory[0][6] ),
    .QN(_0913_));
 DFF_X1 \cam_memory[0][7]$_SDFFCE_PN0P_  (.D(_0007_),
    .CK(clknet_4_8_0_clk),
    .Q(\cam_memory[0][7] ),
    .QN(_0912_));
 DFF_X1 \cam_memory[10][0]$_SDFFCE_PN0P_  (.D(_0008_),
    .CK(clknet_4_2_0_clk),
    .Q(\cam_memory[10][0] ),
    .QN(_0911_));
 DFF_X1 \cam_memory[10][1]$_SDFFCE_PN0P_  (.D(_0009_),
    .CK(clknet_4_2_0_clk),
    .Q(\cam_memory[10][1] ),
    .QN(_0910_));
 DFF_X1 \cam_memory[10][2]$_SDFFCE_PN0P_  (.D(_0010_),
    .CK(clknet_4_2_0_clk),
    .Q(\cam_memory[10][2] ),
    .QN(_0909_));
 DFF_X1 \cam_memory[10][3]$_SDFFCE_PN0P_  (.D(_0011_),
    .CK(clknet_4_2_0_clk),
    .Q(\cam_memory[10][3] ),
    .QN(_0908_));
 DFF_X1 \cam_memory[10][4]$_SDFFCE_PN0P_  (.D(_0012_),
    .CK(clknet_4_2_0_clk),
    .Q(\cam_memory[10][4] ),
    .QN(_0907_));
 DFF_X1 \cam_memory[10][5]$_SDFFCE_PN0P_  (.D(_0013_),
    .CK(clknet_4_2_0_clk),
    .Q(\cam_memory[10][5] ),
    .QN(_0906_));
 DFF_X1 \cam_memory[10][6]$_SDFFCE_PN0P_  (.D(_0014_),
    .CK(clknet_4_2_0_clk),
    .Q(\cam_memory[10][6] ),
    .QN(_0905_));
 DFF_X1 \cam_memory[10][7]$_SDFFCE_PN0P_  (.D(_0015_),
    .CK(clknet_4_2_0_clk),
    .Q(\cam_memory[10][7] ),
    .QN(_0904_));
 DFF_X1 \cam_memory[11][0]$_SDFFCE_PN0P_  (.D(_0016_),
    .CK(clknet_4_4_0_clk),
    .Q(\cam_memory[11][0] ),
    .QN(_0903_));
 DFF_X1 \cam_memory[11][1]$_SDFFCE_PN0P_  (.D(_0017_),
    .CK(clknet_4_6_0_clk),
    .Q(\cam_memory[11][1] ),
    .QN(_0902_));
 DFF_X1 \cam_memory[11][2]$_SDFFCE_PN0P_  (.D(_0018_),
    .CK(clknet_4_4_0_clk),
    .Q(\cam_memory[11][2] ),
    .QN(_0901_));
 DFF_X1 \cam_memory[11][3]$_SDFFCE_PN0P_  (.D(_0019_),
    .CK(clknet_4_6_0_clk),
    .Q(\cam_memory[11][3] ),
    .QN(_0900_));
 DFF_X1 \cam_memory[11][4]$_SDFFCE_PN0P_  (.D(_0020_),
    .CK(clknet_4_4_0_clk),
    .Q(\cam_memory[11][4] ),
    .QN(_0899_));
 DFF_X1 \cam_memory[11][5]$_SDFFCE_PN0P_  (.D(_0021_),
    .CK(clknet_4_5_0_clk),
    .Q(\cam_memory[11][5] ),
    .QN(_0898_));
 DFF_X1 \cam_memory[11][6]$_SDFFCE_PN0P_  (.D(_0022_),
    .CK(clknet_4_6_0_clk),
    .Q(\cam_memory[11][6] ),
    .QN(_0897_));
 DFF_X1 \cam_memory[11][7]$_SDFFCE_PN0P_  (.D(_0023_),
    .CK(clknet_4_4_0_clk),
    .Q(\cam_memory[11][7] ),
    .QN(_0896_));
 DFF_X1 \cam_memory[12][0]$_SDFFCE_PN0P_  (.D(_0024_),
    .CK(clknet_4_3_0_clk),
    .Q(\cam_memory[12][0] ),
    .QN(_0895_));
 DFF_X1 \cam_memory[12][1]$_SDFFCE_PN0P_  (.D(_0025_),
    .CK(clknet_4_1_0_clk),
    .Q(\cam_memory[12][1] ),
    .QN(_0894_));
 DFF_X1 \cam_memory[12][2]$_SDFFCE_PN0P_  (.D(_0026_),
    .CK(clknet_4_1_0_clk),
    .Q(\cam_memory[12][2] ),
    .QN(_0893_));
 DFF_X1 \cam_memory[12][3]$_SDFFCE_PN0P_  (.D(_0027_),
    .CK(clknet_4_1_0_clk),
    .Q(\cam_memory[12][3] ),
    .QN(_0892_));
 DFF_X1 \cam_memory[12][4]$_SDFFCE_PN0P_  (.D(_0028_),
    .CK(clknet_4_1_0_clk),
    .Q(\cam_memory[12][4] ),
    .QN(_0891_));
 DFF_X1 \cam_memory[12][5]$_SDFFCE_PN0P_  (.D(_0029_),
    .CK(clknet_4_1_0_clk),
    .Q(\cam_memory[12][5] ),
    .QN(_0890_));
 DFF_X1 \cam_memory[12][6]$_SDFFCE_PN0P_  (.D(_0030_),
    .CK(clknet_4_1_0_clk),
    .Q(\cam_memory[12][6] ),
    .QN(_0889_));
 DFF_X1 \cam_memory[12][7]$_SDFFCE_PN0P_  (.D(_0031_),
    .CK(clknet_4_1_0_clk),
    .Q(\cam_memory[12][7] ),
    .QN(_0888_));
 DFF_X1 \cam_memory[13][0]$_SDFFCE_PN0P_  (.D(_0032_),
    .CK(clknet_4_4_0_clk),
    .Q(\cam_memory[13][0] ),
    .QN(_0887_));
 DFF_X1 \cam_memory[13][1]$_SDFFCE_PN0P_  (.D(_0033_),
    .CK(clknet_4_4_0_clk),
    .Q(\cam_memory[13][1] ),
    .QN(_0886_));
 DFF_X1 \cam_memory[13][2]$_SDFFCE_PN0P_  (.D(_0034_),
    .CK(clknet_4_4_0_clk),
    .Q(\cam_memory[13][2] ),
    .QN(_0885_));
 DFF_X1 \cam_memory[13][3]$_SDFFCE_PN0P_  (.D(_0035_),
    .CK(clknet_4_4_0_clk),
    .Q(\cam_memory[13][3] ),
    .QN(_0884_));
 DFF_X1 \cam_memory[13][4]$_SDFFCE_PN0P_  (.D(_0036_),
    .CK(clknet_4_4_0_clk),
    .Q(\cam_memory[13][4] ),
    .QN(_0883_));
 DFF_X1 \cam_memory[13][5]$_SDFFCE_PN0P_  (.D(_0037_),
    .CK(clknet_4_4_0_clk),
    .Q(\cam_memory[13][5] ),
    .QN(_0882_));
 DFF_X1 \cam_memory[13][6]$_SDFFCE_PN0P_  (.D(_0038_),
    .CK(clknet_4_5_0_clk),
    .Q(\cam_memory[13][6] ),
    .QN(_0881_));
 DFF_X1 \cam_memory[13][7]$_SDFFCE_PN0P_  (.D(_0039_),
    .CK(clknet_4_5_0_clk),
    .Q(\cam_memory[13][7] ),
    .QN(_0880_));
 DFF_X1 \cam_memory[14][0]$_SDFFCE_PN0P_  (.D(_0040_),
    .CK(clknet_4_3_0_clk),
    .Q(\cam_memory[14][0] ),
    .QN(_0879_));
 DFF_X1 \cam_memory[14][1]$_SDFFCE_PN0P_  (.D(_0041_),
    .CK(clknet_4_0_0_clk),
    .Q(\cam_memory[14][1] ),
    .QN(_0878_));
 DFF_X1 \cam_memory[14][2]$_SDFFCE_PN0P_  (.D(_0042_),
    .CK(clknet_4_3_0_clk),
    .Q(\cam_memory[14][2] ),
    .QN(_0877_));
 DFF_X1 \cam_memory[14][3]$_SDFFCE_PN0P_  (.D(_0043_),
    .CK(clknet_4_1_0_clk),
    .Q(\cam_memory[14][3] ),
    .QN(_0876_));
 DFF_X1 \cam_memory[14][4]$_SDFFCE_PN0P_  (.D(_0044_),
    .CK(clknet_4_1_0_clk),
    .Q(\cam_memory[14][4] ),
    .QN(_0875_));
 DFF_X1 \cam_memory[14][5]$_SDFFCE_PN0P_  (.D(_0045_),
    .CK(clknet_4_0_0_clk),
    .Q(\cam_memory[14][5] ),
    .QN(_0874_));
 DFF_X1 \cam_memory[14][6]$_SDFFCE_PN0P_  (.D(_0046_),
    .CK(clknet_4_0_0_clk),
    .Q(\cam_memory[14][6] ),
    .QN(_0873_));
 DFF_X1 \cam_memory[14][7]$_SDFFCE_PN0P_  (.D(_0047_),
    .CK(clknet_4_0_0_clk),
    .Q(\cam_memory[14][7] ),
    .QN(_0872_));
 DFF_X1 \cam_memory[15][0]$_SDFFCE_PN0P_  (.D(_0048_),
    .CK(clknet_4_2_0_clk),
    .Q(\cam_memory[15][0] ),
    .QN(_0871_));
 DFF_X1 \cam_memory[15][1]$_SDFFCE_PN0P_  (.D(_0049_),
    .CK(clknet_4_0_0_clk),
    .Q(\cam_memory[15][1] ),
    .QN(_0870_));
 DFF_X1 \cam_memory[15][2]$_SDFFCE_PN0P_  (.D(_0050_),
    .CK(clknet_4_0_0_clk),
    .Q(\cam_memory[15][2] ),
    .QN(_0869_));
 DFF_X1 \cam_memory[15][3]$_SDFFCE_PN0P_  (.D(_0051_),
    .CK(clknet_4_0_0_clk),
    .Q(\cam_memory[15][3] ),
    .QN(_0868_));
 DFF_X1 \cam_memory[15][4]$_SDFFCE_PN0P_  (.D(_0052_),
    .CK(clknet_4_0_0_clk),
    .Q(\cam_memory[15][4] ),
    .QN(_0867_));
 DFF_X1 \cam_memory[15][5]$_SDFFCE_PN0P_  (.D(_0053_),
    .CK(clknet_4_0_0_clk),
    .Q(\cam_memory[15][5] ),
    .QN(_0866_));
 DFF_X1 \cam_memory[15][6]$_SDFFCE_PN0P_  (.D(_0054_),
    .CK(clknet_4_0_0_clk),
    .Q(\cam_memory[15][6] ),
    .QN(_0865_));
 DFF_X1 \cam_memory[15][7]$_SDFFCE_PN0P_  (.D(_0055_),
    .CK(clknet_4_2_0_clk),
    .Q(\cam_memory[15][7] ),
    .QN(_0864_));
 DFF_X1 \cam_memory[1][0]$_SDFFCE_PN0P_  (.D(_0056_),
    .CK(clknet_4_8_0_clk),
    .Q(\cam_memory[1][0] ),
    .QN(_0863_));
 DFF_X1 \cam_memory[1][1]$_SDFFCE_PN0P_  (.D(_0057_),
    .CK(clknet_4_10_0_clk),
    .Q(\cam_memory[1][1] ),
    .QN(_0862_));
 DFF_X1 \cam_memory[1][2]$_SDFFCE_PN0P_  (.D(_0058_),
    .CK(clknet_4_10_0_clk),
    .Q(\cam_memory[1][2] ),
    .QN(_0861_));
 DFF_X1 \cam_memory[1][3]$_SDFFCE_PN0P_  (.D(_0059_),
    .CK(clknet_4_10_0_clk),
    .Q(\cam_memory[1][3] ),
    .QN(_0860_));
 DFF_X1 \cam_memory[1][4]$_SDFFCE_PN0P_  (.D(_0060_),
    .CK(clknet_4_10_0_clk),
    .Q(\cam_memory[1][4] ),
    .QN(_0859_));
 DFF_X1 \cam_memory[1][5]$_SDFFCE_PN0P_  (.D(_0061_),
    .CK(clknet_4_10_0_clk),
    .Q(\cam_memory[1][5] ),
    .QN(_0858_));
 DFF_X1 \cam_memory[1][6]$_SDFFCE_PN0P_  (.D(_0062_),
    .CK(clknet_4_10_0_clk),
    .Q(\cam_memory[1][6] ),
    .QN(_0857_));
 DFF_X1 \cam_memory[1][7]$_SDFFCE_PN0P_  (.D(_0063_),
    .CK(clknet_4_10_0_clk),
    .Q(\cam_memory[1][7] ),
    .QN(_0856_));
 DFF_X1 \cam_memory[2][0]$_SDFFCE_PN0P_  (.D(_0064_),
    .CK(clknet_4_9_0_clk),
    .Q(\cam_memory[2][0] ),
    .QN(_0855_));
 DFF_X1 \cam_memory[2][1]$_SDFFCE_PN0P_  (.D(_0065_),
    .CK(clknet_4_9_0_clk),
    .Q(\cam_memory[2][1] ),
    .QN(_0854_));
 DFF_X1 \cam_memory[2][2]$_SDFFCE_PN0P_  (.D(_0066_),
    .CK(clknet_4_11_0_clk),
    .Q(\cam_memory[2][2] ),
    .QN(_0853_));
 DFF_X1 \cam_memory[2][3]$_SDFFCE_PN0P_  (.D(_0067_),
    .CK(clknet_4_11_0_clk),
    .Q(\cam_memory[2][3] ),
    .QN(_0852_));
 DFF_X1 \cam_memory[2][4]$_SDFFCE_PN0P_  (.D(_0068_),
    .CK(clknet_4_11_0_clk),
    .Q(\cam_memory[2][4] ),
    .QN(_0851_));
 DFF_X1 \cam_memory[2][5]$_SDFFCE_PN0P_  (.D(_0069_),
    .CK(clknet_4_11_0_clk),
    .Q(\cam_memory[2][5] ),
    .QN(_0850_));
 DFF_X1 \cam_memory[2][6]$_SDFFCE_PN0P_  (.D(_0070_),
    .CK(clknet_4_11_0_clk),
    .Q(\cam_memory[2][6] ),
    .QN(_0849_));
 DFF_X1 \cam_memory[2][7]$_SDFFCE_PN0P_  (.D(_0071_),
    .CK(clknet_4_11_0_clk),
    .Q(\cam_memory[2][7] ),
    .QN(_0848_));
 DFF_X1 \cam_memory[3][0]$_SDFFCE_PN0P_  (.D(_0072_),
    .CK(clknet_4_14_0_clk),
    .Q(\cam_memory[3][0] ),
    .QN(_0847_));
 DFF_X1 \cam_memory[3][1]$_SDFFCE_PN0P_  (.D(_0073_),
    .CK(clknet_4_9_0_clk),
    .Q(\cam_memory[3][1] ),
    .QN(_0846_));
 DFF_X1 \cam_memory[3][2]$_SDFFCE_PN0P_  (.D(_0074_),
    .CK(clknet_4_11_0_clk),
    .Q(\cam_memory[3][2] ),
    .QN(_0845_));
 DFF_X1 \cam_memory[3][3]$_SDFFCE_PN0P_  (.D(_0075_),
    .CK(clknet_4_14_0_clk),
    .Q(\cam_memory[3][3] ),
    .QN(_0844_));
 DFF_X1 \cam_memory[3][4]$_SDFFCE_PN0P_  (.D(_0076_),
    .CK(clknet_4_14_0_clk),
    .Q(\cam_memory[3][4] ),
    .QN(_0843_));
 DFF_X1 \cam_memory[3][5]$_SDFFCE_PN0P_  (.D(_0077_),
    .CK(clknet_4_11_0_clk),
    .Q(\cam_memory[3][5] ),
    .QN(_0842_));
 DFF_X1 \cam_memory[3][6]$_SDFFCE_PN0P_  (.D(_0078_),
    .CK(clknet_4_14_0_clk),
    .Q(\cam_memory[3][6] ),
    .QN(_0841_));
 DFF_X1 \cam_memory[3][7]$_SDFFCE_PN0P_  (.D(_0079_),
    .CK(clknet_4_14_0_clk),
    .Q(\cam_memory[3][7] ),
    .QN(_0840_));
 DFF_X1 \cam_memory[4][0]$_SDFFCE_PN0P_  (.D(_0080_),
    .CK(clknet_4_12_0_clk),
    .Q(\cam_memory[4][0] ),
    .QN(_0839_));
 DFF_X1 \cam_memory[4][1]$_SDFFCE_PN0P_  (.D(_0081_),
    .CK(clknet_4_12_0_clk),
    .Q(\cam_memory[4][1] ),
    .QN(_0838_));
 DFF_X1 \cam_memory[4][2]$_SDFFCE_PN0P_  (.D(_0082_),
    .CK(clknet_4_12_0_clk),
    .Q(\cam_memory[4][2] ),
    .QN(_0837_));
 DFF_X1 \cam_memory[4][3]$_SDFFCE_PN0P_  (.D(_0083_),
    .CK(clknet_4_12_0_clk),
    .Q(\cam_memory[4][3] ),
    .QN(_0836_));
 DFF_X1 \cam_memory[4][4]$_SDFFCE_PN0P_  (.D(_0084_),
    .CK(clknet_4_14_0_clk),
    .Q(\cam_memory[4][4] ),
    .QN(_0835_));
 DFF_X1 \cam_memory[4][5]$_SDFFCE_PN0P_  (.D(_0085_),
    .CK(clknet_4_14_0_clk),
    .Q(\cam_memory[4][5] ),
    .QN(_0834_));
 DFF_X1 \cam_memory[4][6]$_SDFFCE_PN0P_  (.D(_0086_),
    .CK(clknet_4_12_0_clk),
    .Q(\cam_memory[4][6] ),
    .QN(_0833_));
 DFF_X1 \cam_memory[4][7]$_SDFFCE_PN0P_  (.D(_0087_),
    .CK(clknet_4_14_0_clk),
    .Q(\cam_memory[4][7] ),
    .QN(_0832_));
 DFF_X1 \cam_memory[5][0]$_SDFFCE_PN0P_  (.D(_0088_),
    .CK(clknet_4_12_0_clk),
    .Q(\cam_memory[5][0] ),
    .QN(_0831_));
 DFF_X1 \cam_memory[5][1]$_SDFFCE_PN0P_  (.D(_0089_),
    .CK(clknet_4_15_0_clk),
    .Q(\cam_memory[5][1] ),
    .QN(_0830_));
 DFF_X1 \cam_memory[5][2]$_SDFFCE_PN0P_  (.D(_0090_),
    .CK(clknet_4_14_0_clk),
    .Q(\cam_memory[5][2] ),
    .QN(_0829_));
 DFF_X1 \cam_memory[5][3]$_SDFFCE_PN0P_  (.D(_0091_),
    .CK(clknet_4_12_0_clk),
    .Q(\cam_memory[5][3] ),
    .QN(_0828_));
 DFF_X1 \cam_memory[5][4]$_SDFFCE_PN0P_  (.D(_0092_),
    .CK(clknet_4_15_0_clk),
    .Q(\cam_memory[5][4] ),
    .QN(_0827_));
 DFF_X1 \cam_memory[5][5]$_SDFFCE_PN0P_  (.D(_0093_),
    .CK(clknet_4_15_0_clk),
    .Q(\cam_memory[5][5] ),
    .QN(_0826_));
 DFF_X1 \cam_memory[5][6]$_SDFFCE_PN0P_  (.D(_0094_),
    .CK(clknet_4_15_0_clk),
    .Q(\cam_memory[5][6] ),
    .QN(_0825_));
 DFF_X1 \cam_memory[5][7]$_SDFFCE_PN0P_  (.D(_0095_),
    .CK(clknet_4_13_0_clk),
    .Q(\cam_memory[5][7] ),
    .QN(_0824_));
 DFF_X1 \cam_memory[6][0]$_SDFFCE_PN0P_  (.D(_0096_),
    .CK(clknet_4_13_0_clk),
    .Q(\cam_memory[6][0] ),
    .QN(_0823_));
 DFF_X1 \cam_memory[6][1]$_SDFFCE_PN0P_  (.D(_0097_),
    .CK(clknet_4_13_0_clk),
    .Q(\cam_memory[6][1] ),
    .QN(_0822_));
 DFF_X1 \cam_memory[6][2]$_SDFFCE_PN0P_  (.D(_0098_),
    .CK(clknet_4_7_0_clk),
    .Q(\cam_memory[6][2] ),
    .QN(_0821_));
 DFF_X1 \cam_memory[6][3]$_SDFFCE_PN0P_  (.D(_0099_),
    .CK(clknet_4_7_0_clk),
    .Q(\cam_memory[6][3] ),
    .QN(_0820_));
 DFF_X1 \cam_memory[6][4]$_SDFFCE_PN0P_  (.D(_0100_),
    .CK(clknet_4_7_0_clk),
    .Q(\cam_memory[6][4] ),
    .QN(_0819_));
 DFF_X1 \cam_memory[6][5]$_SDFFCE_PN0P_  (.D(_0101_),
    .CK(clknet_4_13_0_clk),
    .Q(\cam_memory[6][5] ),
    .QN(_0818_));
 DFF_X1 \cam_memory[6][6]$_SDFFCE_PN0P_  (.D(_0102_),
    .CK(clknet_4_13_0_clk),
    .Q(\cam_memory[6][6] ),
    .QN(_0817_));
 DFF_X1 \cam_memory[6][7]$_SDFFCE_PN0P_  (.D(_0103_),
    .CK(clknet_4_13_0_clk),
    .Q(\cam_memory[6][7] ),
    .QN(_0816_));
 DFF_X1 \cam_memory[7][0]$_SDFFCE_PN0P_  (.D(_0104_),
    .CK(clknet_4_13_0_clk),
    .Q(\cam_memory[7][0] ),
    .QN(_0815_));
 DFF_X1 \cam_memory[7][1]$_SDFFCE_PN0P_  (.D(_0105_),
    .CK(clknet_4_13_0_clk),
    .Q(\cam_memory[7][1] ),
    .QN(_0814_));
 DFF_X1 \cam_memory[7][2]$_SDFFCE_PN0P_  (.D(_0106_),
    .CK(clknet_4_13_0_clk),
    .Q(\cam_memory[7][2] ),
    .QN(_0813_));
 DFF_X1 \cam_memory[7][3]$_SDFFCE_PN0P_  (.D(_0107_),
    .CK(clknet_4_13_0_clk),
    .Q(\cam_memory[7][3] ),
    .QN(_0812_));
 DFF_X1 \cam_memory[7][4]$_SDFFCE_PN0P_  (.D(_0108_),
    .CK(clknet_4_15_0_clk),
    .Q(\cam_memory[7][4] ),
    .QN(_0811_));
 DFF_X1 \cam_memory[7][5]$_SDFFCE_PN0P_  (.D(_0109_),
    .CK(clknet_4_15_0_clk),
    .Q(\cam_memory[7][5] ),
    .QN(_0810_));
 DFF_X1 \cam_memory[7][6]$_SDFFCE_PN0P_  (.D(_0110_),
    .CK(clknet_4_15_0_clk),
    .Q(\cam_memory[7][6] ),
    .QN(_0809_));
 DFF_X1 \cam_memory[7][7]$_SDFFCE_PN0P_  (.D(_0111_),
    .CK(clknet_4_15_0_clk),
    .Q(\cam_memory[7][7] ),
    .QN(_0808_));
 DFF_X1 \cam_memory[8][0]$_SDFFCE_PN0P_  (.D(_0112_),
    .CK(clknet_4_5_0_clk),
    .Q(\cam_memory[8][0] ),
    .QN(_0807_));
 DFF_X1 \cam_memory[8][1]$_SDFFCE_PN0P_  (.D(_0113_),
    .CK(clknet_4_7_0_clk),
    .Q(\cam_memory[8][1] ),
    .QN(_0806_));
 DFF_X1 \cam_memory[8][2]$_SDFFCE_PN0P_  (.D(_0114_),
    .CK(clknet_4_7_0_clk),
    .Q(\cam_memory[8][2] ),
    .QN(_0805_));
 DFF_X1 \cam_memory[8][3]$_SDFFCE_PN0P_  (.D(_0115_),
    .CK(clknet_4_5_0_clk),
    .Q(\cam_memory[8][3] ),
    .QN(_0804_));
 DFF_X1 \cam_memory[8][4]$_SDFFCE_PN0P_  (.D(_0116_),
    .CK(clknet_4_5_0_clk),
    .Q(\cam_memory[8][4] ),
    .QN(_0803_));
 DFF_X1 \cam_memory[8][5]$_SDFFCE_PN0P_  (.D(_0117_),
    .CK(clknet_4_5_0_clk),
    .Q(\cam_memory[8][5] ),
    .QN(_0802_));
 DFF_X1 \cam_memory[8][6]$_SDFFCE_PN0P_  (.D(_0118_),
    .CK(clknet_4_7_0_clk),
    .Q(\cam_memory[8][6] ),
    .QN(_0801_));
 DFF_X1 \cam_memory[8][7]$_SDFFCE_PN0P_  (.D(_0119_),
    .CK(clknet_4_5_0_clk),
    .Q(\cam_memory[8][7] ),
    .QN(_0800_));
 DFF_X1 \cam_memory[9][0]$_SDFFCE_PN0P_  (.D(_0120_),
    .CK(clknet_4_7_0_clk),
    .Q(\cam_memory[9][0] ),
    .QN(_0799_));
 DFF_X1 \cam_memory[9][1]$_SDFFCE_PN0P_  (.D(_0121_),
    .CK(clknet_4_7_0_clk),
    .Q(\cam_memory[9][1] ),
    .QN(_0798_));
 DFF_X1 \cam_memory[9][2]$_SDFFCE_PN0P_  (.D(_0122_),
    .CK(clknet_4_7_0_clk),
    .Q(\cam_memory[9][2] ),
    .QN(_0797_));
 DFF_X1 \cam_memory[9][3]$_SDFFCE_PN0P_  (.D(_0123_),
    .CK(clknet_4_7_0_clk),
    .Q(\cam_memory[9][3] ),
    .QN(_0796_));
 DFF_X1 \cam_memory[9][4]$_SDFFCE_PN0P_  (.D(_0124_),
    .CK(clknet_4_7_0_clk),
    .Q(\cam_memory[9][4] ),
    .QN(_0795_));
 DFF_X1 \cam_memory[9][5]$_SDFFCE_PN0P_  (.D(_0125_),
    .CK(clknet_4_6_0_clk),
    .Q(\cam_memory[9][5] ),
    .QN(_0794_));
 DFF_X1 \cam_memory[9][6]$_SDFFCE_PN0P_  (.D(_0126_),
    .CK(clknet_4_6_0_clk),
    .Q(\cam_memory[9][6] ),
    .QN(_0793_));
 DFF_X1 \cam_memory[9][7]$_SDFFCE_PN0P_  (.D(_0127_),
    .CK(clknet_4_6_0_clk),
    .Q(\cam_memory[9][7] ),
    .QN(_0792_));
 DFF_X1 \match$_SDFF_PN0_  (.D(_0128_),
    .CK(clknet_4_14_0_clk),
    .Q(net3),
    .QN(_0791_));
 DFF_X1 \match_addr[0]$_SDFFE_PN0P_  (.D(_0129_),
    .CK(clknet_4_6_0_clk),
    .Q(net4),
    .QN(_0790_));
 DFF_X1 \match_addr[1]$_SDFFE_PN0P_  (.D(_0130_),
    .CK(clknet_4_6_0_clk),
    .Q(net5),
    .QN(_0789_));
 DFF_X1 \match_addr[2]$_SDFFE_PN0P_  (.D(_0131_),
    .CK(clknet_4_12_0_clk),
    .Q(net6),
    .QN(_0788_));
 DFF_X1 \match_addr[3]$_SDFFE_PN0P_  (.D(_0132_),
    .CK(clknet_4_9_0_clk),
    .Q(net7),
    .QN(_0787_));
 DFF_X1 \valid$_SDFF_PN0_  (.D(_0133_),
    .CK(clknet_4_14_0_clk),
    .Q(net8),
    .QN(_0786_));
 DFF_X1 \valid_bits[0]$_SDFFE_PN0P_  (.D(_0134_),
    .CK(clknet_4_8_0_clk),
    .Q(\valid_bits[0] ),
    .QN(_0785_));
 DFF_X1 \valid_bits[10]$_SDFFE_PN0P_  (.D(_0135_),
    .CK(clknet_4_3_0_clk),
    .Q(\valid_bits[10] ),
    .QN(_0784_));
 DFF_X1 \valid_bits[11]$_SDFFE_PN0P_  (.D(_0136_),
    .CK(clknet_4_3_0_clk),
    .Q(\valid_bits[11] ),
    .QN(_0783_));
 DFF_X1 \valid_bits[12]$_SDFFE_PN0P_  (.D(_0137_),
    .CK(clknet_4_3_0_clk),
    .Q(\valid_bits[12] ),
    .QN(_0782_));
 DFF_X1 \valid_bits[13]$_SDFFE_PN0P_  (.D(_0138_),
    .CK(clknet_4_3_0_clk),
    .Q(\valid_bits[13] ),
    .QN(_0781_));
 DFF_X1 \valid_bits[14]$_SDFFE_PN0P_  (.D(_0139_),
    .CK(clknet_4_3_0_clk),
    .Q(\valid_bits[14] ),
    .QN(_0780_));
 DFF_X1 \valid_bits[15]$_SDFFE_PN0P_  (.D(_0140_),
    .CK(clknet_4_3_0_clk),
    .Q(\valid_bits[15] ),
    .QN(_0779_));
 DFF_X1 \valid_bits[1]$_SDFFE_PN0P_  (.D(_0141_),
    .CK(clknet_4_8_0_clk),
    .Q(\valid_bits[1] ),
    .QN(_0778_));
 DFF_X1 \valid_bits[2]$_SDFFE_PN0P_  (.D(_0142_),
    .CK(clknet_4_9_0_clk),
    .Q(\valid_bits[2] ),
    .QN(_0777_));
 DFF_X1 \valid_bits[3]$_SDFFE_PN0P_  (.D(_0143_),
    .CK(clknet_4_9_0_clk),
    .Q(\valid_bits[3] ),
    .QN(_0776_));
 DFF_X1 \valid_bits[4]$_SDFFE_PN0P_  (.D(_0144_),
    .CK(clknet_4_9_0_clk),
    .Q(\valid_bits[4] ),
    .QN(_0775_));
 DFF_X1 \valid_bits[5]$_SDFFE_PN0P_  (.D(_0145_),
    .CK(clknet_4_9_0_clk),
    .Q(\valid_bits[5] ),
    .QN(_0774_));
 DFF_X1 \valid_bits[6]$_SDFFE_PN0P_  (.D(_0146_),
    .CK(clknet_4_9_0_clk),
    .Q(\valid_bits[6] ),
    .QN(_0773_));
 DFF_X1 \valid_bits[7]$_SDFFE_PN0P_  (.D(_0147_),
    .CK(clknet_4_9_0_clk),
    .Q(\valid_bits[7] ),
    .QN(_0772_));
 DFF_X1 \valid_bits[8]$_SDFFE_PN0P_  (.D(_0148_),
    .CK(clknet_4_3_0_clk),
    .Q(\valid_bits[8] ),
    .QN(_0771_));
 DFF_X1 \valid_bits[9]$_SDFFE_PN0P_  (.D(_0149_),
    .CK(clknet_4_3_0_clk),
    .Q(\valid_bits[9] ),
    .QN(_0770_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_77 ();
 CLKBUF_X3 input1 (.A(write_addr[0]),
    .Z(net1));
 CLKBUF_X3 input2 (.A(write_addr[1]),
    .Z(net2));
 BUF_X1 output3 (.A(net3),
    .Z(match));
 BUF_X1 output4 (.A(net4),
    .Z(match_addr[0]));
 BUF_X1 output5 (.A(net5),
    .Z(match_addr[1]));
 BUF_X1 output6 (.A(net6),
    .Z(match_addr[2]));
 BUF_X1 output7 (.A(net7),
    .Z(match_addr[3]));
 BUF_X1 output8 (.A(net8),
    .Z(valid));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 CLKBUF_X3 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 CLKBUF_X3 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 CLKBUF_X3 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 CLKBUF_X3 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 CLKBUF_X3 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 CLKBUF_X3 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 CLKBUF_X3 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 CLKBUF_X3 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 CLKBUF_X3 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 CLKBUF_X3 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 CLKBUF_X3 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 CLKBUF_X3 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 CLKBUF_X3 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 CLKBUF_X3 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 CLKBUF_X3 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 CLKBUF_X1 clkload0 (.A(clknet_4_0_0_clk));
 INV_X1 clkload1 (.A(clknet_4_1_0_clk));
 CLKBUF_X1 clkload2 (.A(clknet_4_2_0_clk));
 CLKBUF_X1 clkload3 (.A(clknet_4_4_0_clk));
 INV_X2 clkload4 (.A(clknet_4_5_0_clk));
 INV_X2 clkload5 (.A(clknet_4_6_0_clk));
 CLKBUF_X1 clkload6 (.A(clknet_4_9_0_clk));
 INV_X2 clkload7 (.A(clknet_4_10_0_clk));
 INV_X2 clkload8 (.A(clknet_4_11_0_clk));
 INV_X2 clkload9 (.A(clknet_4_12_0_clk));
 CLKBUF_X1 clkload10 (.A(clknet_4_13_0_clk));
 INV_X2 clkload11 (.A(clknet_4_15_0_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X16 FILLER_0_65 ();
 FILLCELL_X8 FILLER_0_81 ();
 FILLCELL_X4 FILLER_0_89 ();
 FILLCELL_X2 FILLER_0_93 ();
 FILLCELL_X1 FILLER_0_95 ();
 FILLCELL_X4 FILLER_0_99 ();
 FILLCELL_X2 FILLER_0_103 ();
 FILLCELL_X1 FILLER_0_105 ();
 FILLCELL_X16 FILLER_0_109 ();
 FILLCELL_X8 FILLER_0_125 ();
 FILLCELL_X2 FILLER_0_133 ();
 FILLCELL_X1 FILLER_0_135 ();
 FILLCELL_X16 FILLER_0_141 ();
 FILLCELL_X4 FILLER_0_157 ();
 FILLCELL_X4 FILLER_0_168 ();
 FILLCELL_X2 FILLER_0_172 ();
 FILLCELL_X1 FILLER_0_174 ();
 FILLCELL_X32 FILLER_0_188 ();
 FILLCELL_X32 FILLER_0_220 ();
 FILLCELL_X32 FILLER_0_252 ();
 FILLCELL_X8 FILLER_0_284 ();
 FILLCELL_X1 FILLER_0_292 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X8 FILLER_1_65 ();
 FILLCELL_X4 FILLER_1_73 ();
 FILLCELL_X2 FILLER_1_77 ();
 FILLCELL_X2 FILLER_1_107 ();
 FILLCELL_X2 FILLER_1_129 ();
 FILLCELL_X1 FILLER_1_131 ();
 FILLCELL_X4 FILLER_1_137 ();
 FILLCELL_X1 FILLER_1_141 ();
 FILLCELL_X8 FILLER_1_166 ();
 FILLCELL_X4 FILLER_1_174 ();
 FILLCELL_X4 FILLER_1_195 ();
 FILLCELL_X2 FILLER_1_199 ();
 FILLCELL_X32 FILLER_1_218 ();
 FILLCELL_X32 FILLER_1_250 ();
 FILLCELL_X8 FILLER_1_282 ();
 FILLCELL_X2 FILLER_1_290 ();
 FILLCELL_X1 FILLER_1_292 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X8 FILLER_2_65 ();
 FILLCELL_X4 FILLER_2_73 ();
 FILLCELL_X2 FILLER_2_77 ();
 FILLCELL_X1 FILLER_2_79 ();
 FILLCELL_X1 FILLER_2_114 ();
 FILLCELL_X2 FILLER_2_119 ();
 FILLCELL_X1 FILLER_2_146 ();
 FILLCELL_X8 FILLER_2_195 ();
 FILLCELL_X4 FILLER_2_203 ();
 FILLCELL_X1 FILLER_2_207 ();
 FILLCELL_X32 FILLER_2_218 ();
 FILLCELL_X32 FILLER_2_250 ();
 FILLCELL_X8 FILLER_2_282 ();
 FILLCELL_X2 FILLER_2_290 ();
 FILLCELL_X1 FILLER_2_292 ();
 FILLCELL_X4 FILLER_3_1 ();
 FILLCELL_X1 FILLER_3_5 ();
 FILLCELL_X32 FILLER_3_19 ();
 FILLCELL_X1 FILLER_3_51 ();
 FILLCELL_X16 FILLER_3_69 ();
 FILLCELL_X2 FILLER_3_85 ();
 FILLCELL_X1 FILLER_3_87 ();
 FILLCELL_X1 FILLER_3_95 ();
 FILLCELL_X2 FILLER_3_99 ();
 FILLCELL_X8 FILLER_3_131 ();
 FILLCELL_X2 FILLER_3_139 ();
 FILLCELL_X1 FILLER_3_141 ();
 FILLCELL_X2 FILLER_3_203 ();
 FILLCELL_X4 FILLER_3_211 ();
 FILLCELL_X2 FILLER_3_215 ();
 FILLCELL_X4 FILLER_3_234 ();
 FILLCELL_X1 FILLER_3_238 ();
 FILLCELL_X32 FILLER_3_246 ();
 FILLCELL_X8 FILLER_3_278 ();
 FILLCELL_X4 FILLER_3_286 ();
 FILLCELL_X2 FILLER_3_290 ();
 FILLCELL_X1 FILLER_3_292 ();
 FILLCELL_X4 FILLER_4_1 ();
 FILLCELL_X1 FILLER_4_5 ();
 FILLCELL_X8 FILLER_4_40 ();
 FILLCELL_X2 FILLER_4_54 ();
 FILLCELL_X2 FILLER_4_64 ();
 FILLCELL_X16 FILLER_4_72 ();
 FILLCELL_X4 FILLER_4_88 ();
 FILLCELL_X4 FILLER_4_108 ();
 FILLCELL_X2 FILLER_4_112 ();
 FILLCELL_X1 FILLER_4_114 ();
 FILLCELL_X16 FILLER_4_124 ();
 FILLCELL_X8 FILLER_4_140 ();
 FILLCELL_X2 FILLER_4_148 ();
 FILLCELL_X1 FILLER_4_150 ();
 FILLCELL_X1 FILLER_4_158 ();
 FILLCELL_X2 FILLER_4_162 ();
 FILLCELL_X1 FILLER_4_168 ();
 FILLCELL_X2 FILLER_4_172 ();
 FILLCELL_X4 FILLER_4_179 ();
 FILLCELL_X1 FILLER_4_183 ();
 FILLCELL_X1 FILLER_4_188 ();
 FILLCELL_X2 FILLER_4_192 ();
 FILLCELL_X1 FILLER_4_197 ();
 FILLCELL_X1 FILLER_4_229 ();
 FILLCELL_X1 FILLER_4_236 ();
 FILLCELL_X32 FILLER_4_254 ();
 FILLCELL_X4 FILLER_4_286 ();
 FILLCELL_X2 FILLER_4_290 ();
 FILLCELL_X1 FILLER_4_292 ();
 FILLCELL_X8 FILLER_5_1 ();
 FILLCELL_X2 FILLER_5_9 ();
 FILLCELL_X1 FILLER_5_11 ();
 FILLCELL_X2 FILLER_5_42 ();
 FILLCELL_X8 FILLER_5_78 ();
 FILLCELL_X2 FILLER_5_90 ();
 FILLCELL_X8 FILLER_5_95 ();
 FILLCELL_X1 FILLER_5_103 ();
 FILLCELL_X4 FILLER_5_107 ();
 FILLCELL_X1 FILLER_5_111 ();
 FILLCELL_X4 FILLER_5_119 ();
 FILLCELL_X2 FILLER_5_123 ();
 FILLCELL_X1 FILLER_5_125 ();
 FILLCELL_X16 FILLER_5_129 ();
 FILLCELL_X8 FILLER_5_145 ();
 FILLCELL_X2 FILLER_5_163 ();
 FILLCELL_X1 FILLER_5_165 ();
 FILLCELL_X1 FILLER_5_169 ();
 FILLCELL_X8 FILLER_5_174 ();
 FILLCELL_X2 FILLER_5_185 ();
 FILLCELL_X1 FILLER_5_187 ();
 FILLCELL_X16 FILLER_5_194 ();
 FILLCELL_X2 FILLER_5_210 ();
 FILLCELL_X1 FILLER_5_221 ();
 FILLCELL_X4 FILLER_5_225 ();
 FILLCELL_X4 FILLER_5_239 ();
 FILLCELL_X2 FILLER_5_249 ();
 FILLCELL_X32 FILLER_5_254 ();
 FILLCELL_X4 FILLER_5_286 ();
 FILLCELL_X2 FILLER_5_290 ();
 FILLCELL_X1 FILLER_5_292 ();
 FILLCELL_X16 FILLER_6_1 ();
 FILLCELL_X8 FILLER_6_17 ();
 FILLCELL_X4 FILLER_6_25 ();
 FILLCELL_X1 FILLER_6_29 ();
 FILLCELL_X8 FILLER_6_39 ();
 FILLCELL_X1 FILLER_6_54 ();
 FILLCELL_X4 FILLER_6_64 ();
 FILLCELL_X2 FILLER_6_68 ();
 FILLCELL_X1 FILLER_6_70 ();
 FILLCELL_X2 FILLER_6_98 ();
 FILLCELL_X1 FILLER_6_107 ();
 FILLCELL_X4 FILLER_6_137 ();
 FILLCELL_X2 FILLER_6_141 ();
 FILLCELL_X1 FILLER_6_143 ();
 FILLCELL_X1 FILLER_6_190 ();
 FILLCELL_X16 FILLER_6_195 ();
 FILLCELL_X4 FILLER_6_211 ();
 FILLCELL_X1 FILLER_6_215 ();
 FILLCELL_X4 FILLER_6_220 ();
 FILLCELL_X4 FILLER_6_235 ();
 FILLCELL_X2 FILLER_6_239 ();
 FILLCELL_X1 FILLER_6_241 ();
 FILLCELL_X16 FILLER_6_263 ();
 FILLCELL_X8 FILLER_6_279 ();
 FILLCELL_X4 FILLER_6_287 ();
 FILLCELL_X2 FILLER_6_291 ();
 FILLCELL_X4 FILLER_7_1 ();
 FILLCELL_X2 FILLER_7_5 ();
 FILLCELL_X1 FILLER_7_24 ();
 FILLCELL_X2 FILLER_7_35 ();
 FILLCELL_X1 FILLER_7_37 ();
 FILLCELL_X1 FILLER_7_41 ();
 FILLCELL_X4 FILLER_7_46 ();
 FILLCELL_X4 FILLER_7_54 ();
 FILLCELL_X2 FILLER_7_61 ();
 FILLCELL_X2 FILLER_7_69 ();
 FILLCELL_X1 FILLER_7_117 ();
 FILLCELL_X1 FILLER_7_124 ();
 FILLCELL_X8 FILLER_7_143 ();
 FILLCELL_X2 FILLER_7_169 ();
 FILLCELL_X16 FILLER_7_177 ();
 FILLCELL_X4 FILLER_7_193 ();
 FILLCELL_X2 FILLER_7_197 ();
 FILLCELL_X1 FILLER_7_199 ();
 FILLCELL_X4 FILLER_7_205 ();
 FILLCELL_X1 FILLER_7_209 ();
 FILLCELL_X8 FILLER_7_230 ();
 FILLCELL_X1 FILLER_7_238 ();
 FILLCELL_X2 FILLER_7_245 ();
 FILLCELL_X16 FILLER_7_263 ();
 FILLCELL_X8 FILLER_7_279 ();
 FILLCELL_X4 FILLER_7_287 ();
 FILLCELL_X2 FILLER_7_291 ();
 FILLCELL_X4 FILLER_8_1 ();
 FILLCELL_X2 FILLER_8_5 ();
 FILLCELL_X1 FILLER_8_24 ();
 FILLCELL_X2 FILLER_8_28 ();
 FILLCELL_X2 FILLER_8_34 ();
 FILLCELL_X2 FILLER_8_41 ();
 FILLCELL_X1 FILLER_8_43 ();
 FILLCELL_X2 FILLER_8_65 ();
 FILLCELL_X2 FILLER_8_72 ();
 FILLCELL_X2 FILLER_8_81 ();
 FILLCELL_X8 FILLER_8_105 ();
 FILLCELL_X2 FILLER_8_113 ();
 FILLCELL_X4 FILLER_8_130 ();
 FILLCELL_X1 FILLER_8_134 ();
 FILLCELL_X8 FILLER_8_148 ();
 FILLCELL_X2 FILLER_8_156 ();
 FILLCELL_X1 FILLER_8_158 ();
 FILLCELL_X1 FILLER_8_211 ();
 FILLCELL_X1 FILLER_8_216 ();
 FILLCELL_X4 FILLER_8_220 ();
 FILLCELL_X4 FILLER_8_244 ();
 FILLCELL_X1 FILLER_8_248 ();
 FILLCELL_X16 FILLER_8_266 ();
 FILLCELL_X8 FILLER_8_282 ();
 FILLCELL_X2 FILLER_8_290 ();
 FILLCELL_X1 FILLER_8_292 ();
 FILLCELL_X16 FILLER_9_1 ();
 FILLCELL_X4 FILLER_9_17 ();
 FILLCELL_X16 FILLER_9_33 ();
 FILLCELL_X1 FILLER_9_49 ();
 FILLCELL_X4 FILLER_9_53 ();
 FILLCELL_X1 FILLER_9_57 ();
 FILLCELL_X8 FILLER_9_64 ();
 FILLCELL_X4 FILLER_9_72 ();
 FILLCELL_X2 FILLER_9_76 ();
 FILLCELL_X1 FILLER_9_78 ();
 FILLCELL_X8 FILLER_9_84 ();
 FILLCELL_X1 FILLER_9_92 ();
 FILLCELL_X32 FILLER_9_98 ();
 FILLCELL_X8 FILLER_9_130 ();
 FILLCELL_X4 FILLER_9_138 ();
 FILLCELL_X4 FILLER_9_162 ();
 FILLCELL_X2 FILLER_9_166 ();
 FILLCELL_X1 FILLER_9_168 ();
 FILLCELL_X4 FILLER_9_175 ();
 FILLCELL_X2 FILLER_9_179 ();
 FILLCELL_X16 FILLER_9_207 ();
 FILLCELL_X8 FILLER_9_223 ();
 FILLCELL_X4 FILLER_9_231 ();
 FILLCELL_X1 FILLER_9_250 ();
 FILLCELL_X32 FILLER_9_261 ();
 FILLCELL_X2 FILLER_10_1 ();
 FILLCELL_X1 FILLER_10_3 ();
 FILLCELL_X1 FILLER_10_31 ();
 FILLCELL_X16 FILLER_10_38 ();
 FILLCELL_X4 FILLER_10_64 ();
 FILLCELL_X1 FILLER_10_68 ();
 FILLCELL_X16 FILLER_10_79 ();
 FILLCELL_X8 FILLER_10_117 ();
 FILLCELL_X4 FILLER_10_125 ();
 FILLCELL_X2 FILLER_10_129 ();
 FILLCELL_X1 FILLER_10_131 ();
 FILLCELL_X4 FILLER_10_146 ();
 FILLCELL_X1 FILLER_10_150 ();
 FILLCELL_X32 FILLER_10_212 ();
 FILLCELL_X8 FILLER_10_244 ();
 FILLCELL_X2 FILLER_10_252 ();
 FILLCELL_X1 FILLER_10_254 ();
 FILLCELL_X32 FILLER_10_258 ();
 FILLCELL_X2 FILLER_10_290 ();
 FILLCELL_X1 FILLER_10_292 ();
 FILLCELL_X8 FILLER_11_1 ();
 FILLCELL_X4 FILLER_11_9 ();
 FILLCELL_X2 FILLER_11_13 ();
 FILLCELL_X2 FILLER_11_44 ();
 FILLCELL_X1 FILLER_11_69 ();
 FILLCELL_X8 FILLER_11_87 ();
 FILLCELL_X2 FILLER_11_95 ();
 FILLCELL_X1 FILLER_11_97 ();
 FILLCELL_X1 FILLER_11_120 ();
 FILLCELL_X1 FILLER_11_155 ();
 FILLCELL_X8 FILLER_11_196 ();
 FILLCELL_X4 FILLER_11_204 ();
 FILLCELL_X1 FILLER_11_208 ();
 FILLCELL_X1 FILLER_11_213 ();
 FILLCELL_X4 FILLER_11_217 ();
 FILLCELL_X1 FILLER_11_221 ();
 FILLCELL_X8 FILLER_11_239 ();
 FILLCELL_X1 FILLER_11_247 ();
 FILLCELL_X1 FILLER_11_251 ();
 FILLCELL_X1 FILLER_11_264 ();
 FILLCELL_X16 FILLER_11_269 ();
 FILLCELL_X8 FILLER_11_285 ();
 FILLCELL_X16 FILLER_12_1 ();
 FILLCELL_X1 FILLER_12_29 ();
 FILLCELL_X1 FILLER_12_36 ();
 FILLCELL_X2 FILLER_12_41 ();
 FILLCELL_X2 FILLER_12_77 ();
 FILLCELL_X1 FILLER_12_79 ();
 FILLCELL_X8 FILLER_12_86 ();
 FILLCELL_X4 FILLER_12_94 ();
 FILLCELL_X2 FILLER_12_98 ();
 FILLCELL_X4 FILLER_12_121 ();
 FILLCELL_X2 FILLER_12_125 ();
 FILLCELL_X2 FILLER_12_170 ();
 FILLCELL_X1 FILLER_12_172 ();
 FILLCELL_X1 FILLER_12_186 ();
 FILLCELL_X4 FILLER_12_201 ();
 FILLCELL_X1 FILLER_12_219 ();
 FILLCELL_X1 FILLER_12_223 ();
 FILLCELL_X1 FILLER_12_228 ();
 FILLCELL_X2 FILLER_12_232 ();
 FILLCELL_X1 FILLER_12_266 ();
 FILLCELL_X8 FILLER_12_284 ();
 FILLCELL_X1 FILLER_12_292 ();
 FILLCELL_X4 FILLER_13_1 ();
 FILLCELL_X1 FILLER_13_5 ();
 FILLCELL_X4 FILLER_13_37 ();
 FILLCELL_X2 FILLER_13_41 ();
 FILLCELL_X1 FILLER_13_43 ();
 FILLCELL_X2 FILLER_13_51 ();
 FILLCELL_X1 FILLER_13_56 ();
 FILLCELL_X1 FILLER_13_61 ();
 FILLCELL_X1 FILLER_13_68 ();
 FILLCELL_X1 FILLER_13_73 ();
 FILLCELL_X4 FILLER_13_77 ();
 FILLCELL_X4 FILLER_13_87 ();
 FILLCELL_X2 FILLER_13_91 ();
 FILLCELL_X8 FILLER_13_117 ();
 FILLCELL_X2 FILLER_13_125 ();
 FILLCELL_X1 FILLER_13_127 ();
 FILLCELL_X2 FILLER_13_161 ();
 FILLCELL_X1 FILLER_13_163 ();
 FILLCELL_X2 FILLER_13_167 ();
 FILLCELL_X2 FILLER_13_195 ();
 FILLCELL_X1 FILLER_13_197 ();
 FILLCELL_X1 FILLER_13_229 ();
 FILLCELL_X2 FILLER_13_248 ();
 FILLCELL_X1 FILLER_13_254 ();
 FILLCELL_X2 FILLER_13_258 ();
 FILLCELL_X1 FILLER_13_266 ();
 FILLCELL_X16 FILLER_13_274 ();
 FILLCELL_X2 FILLER_13_290 ();
 FILLCELL_X1 FILLER_13_292 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X8 FILLER_14_33 ();
 FILLCELL_X2 FILLER_14_58 ();
 FILLCELL_X2 FILLER_14_63 ();
 FILLCELL_X1 FILLER_14_65 ();
 FILLCELL_X8 FILLER_14_90 ();
 FILLCELL_X2 FILLER_14_101 ();
 FILLCELL_X8 FILLER_14_107 ();
 FILLCELL_X2 FILLER_14_115 ();
 FILLCELL_X4 FILLER_14_120 ();
 FILLCELL_X8 FILLER_14_128 ();
 FILLCELL_X4 FILLER_14_136 ();
 FILLCELL_X2 FILLER_14_140 ();
 FILLCELL_X1 FILLER_14_163 ();
 FILLCELL_X1 FILLER_14_167 ();
 FILLCELL_X1 FILLER_14_171 ();
 FILLCELL_X2 FILLER_14_176 ();
 FILLCELL_X4 FILLER_14_202 ();
 FILLCELL_X1 FILLER_14_233 ();
 FILLCELL_X2 FILLER_14_237 ();
 FILLCELL_X4 FILLER_14_256 ();
 FILLCELL_X1 FILLER_14_260 ();
 FILLCELL_X2 FILLER_14_273 ();
 FILLCELL_X1 FILLER_14_275 ();
 FILLCELL_X16 FILLER_15_1 ();
 FILLCELL_X2 FILLER_15_23 ();
 FILLCELL_X2 FILLER_15_28 ();
 FILLCELL_X1 FILLER_15_30 ();
 FILLCELL_X8 FILLER_15_41 ();
 FILLCELL_X4 FILLER_15_49 ();
 FILLCELL_X2 FILLER_15_53 ();
 FILLCELL_X1 FILLER_15_55 ();
 FILLCELL_X8 FILLER_15_59 ();
 FILLCELL_X2 FILLER_15_67 ();
 FILLCELL_X16 FILLER_15_74 ();
 FILLCELL_X4 FILLER_15_90 ();
 FILLCELL_X1 FILLER_15_94 ();
 FILLCELL_X8 FILLER_15_129 ();
 FILLCELL_X1 FILLER_15_139 ();
 FILLCELL_X1 FILLER_15_142 ();
 FILLCELL_X4 FILLER_15_151 ();
 FILLCELL_X1 FILLER_15_155 ();
 FILLCELL_X2 FILLER_15_161 ();
 FILLCELL_X1 FILLER_15_163 ();
 FILLCELL_X16 FILLER_15_181 ();
 FILLCELL_X4 FILLER_15_197 ();
 FILLCELL_X1 FILLER_15_201 ();
 FILLCELL_X1 FILLER_15_211 ();
 FILLCELL_X8 FILLER_15_222 ();
 FILLCELL_X4 FILLER_15_230 ();
 FILLCELL_X1 FILLER_15_240 ();
 FILLCELL_X32 FILLER_15_244 ();
 FILLCELL_X16 FILLER_15_276 ();
 FILLCELL_X1 FILLER_15_292 ();
 FILLCELL_X8 FILLER_16_1 ();
 FILLCELL_X4 FILLER_16_9 ();
 FILLCELL_X1 FILLER_16_13 ();
 FILLCELL_X2 FILLER_16_18 ();
 FILLCELL_X2 FILLER_16_24 ();
 FILLCELL_X2 FILLER_16_29 ();
 FILLCELL_X4 FILLER_16_48 ();
 FILLCELL_X2 FILLER_16_52 ();
 FILLCELL_X1 FILLER_16_58 ();
 FILLCELL_X4 FILLER_16_62 ();
 FILLCELL_X16 FILLER_16_75 ();
 FILLCELL_X8 FILLER_16_91 ();
 FILLCELL_X2 FILLER_16_102 ();
 FILLCELL_X2 FILLER_16_108 ();
 FILLCELL_X4 FILLER_16_115 ();
 FILLCELL_X1 FILLER_16_119 ();
 FILLCELL_X2 FILLER_16_127 ();
 FILLCELL_X16 FILLER_16_146 ();
 FILLCELL_X8 FILLER_16_162 ();
 FILLCELL_X2 FILLER_16_170 ();
 FILLCELL_X1 FILLER_16_172 ();
 FILLCELL_X1 FILLER_16_181 ();
 FILLCELL_X8 FILLER_16_199 ();
 FILLCELL_X4 FILLER_16_207 ();
 FILLCELL_X1 FILLER_16_211 ();
 FILLCELL_X16 FILLER_16_216 ();
 FILLCELL_X4 FILLER_16_232 ();
 FILLCELL_X2 FILLER_16_236 ();
 FILLCELL_X1 FILLER_16_238 ();
 FILLCELL_X32 FILLER_16_242 ();
 FILLCELL_X16 FILLER_16_274 ();
 FILLCELL_X2 FILLER_16_290 ();
 FILLCELL_X1 FILLER_16_292 ();
 FILLCELL_X2 FILLER_17_1 ();
 FILLCELL_X1 FILLER_17_3 ();
 FILLCELL_X2 FILLER_17_46 ();
 FILLCELL_X1 FILLER_17_48 ();
 FILLCELL_X1 FILLER_17_70 ();
 FILLCELL_X2 FILLER_17_78 ();
 FILLCELL_X16 FILLER_17_83 ();
 FILLCELL_X8 FILLER_17_99 ();
 FILLCELL_X4 FILLER_17_107 ();
 FILLCELL_X2 FILLER_17_128 ();
 FILLCELL_X1 FILLER_17_130 ();
 FILLCELL_X4 FILLER_17_148 ();
 FILLCELL_X2 FILLER_17_152 ();
 FILLCELL_X1 FILLER_17_154 ();
 FILLCELL_X8 FILLER_17_187 ();
 FILLCELL_X4 FILLER_17_195 ();
 FILLCELL_X16 FILLER_17_223 ();
 FILLCELL_X32 FILLER_17_246 ();
 FILLCELL_X8 FILLER_17_278 ();
 FILLCELL_X4 FILLER_17_286 ();
 FILLCELL_X2 FILLER_17_290 ();
 FILLCELL_X1 FILLER_17_292 ();
 FILLCELL_X2 FILLER_18_1 ();
 FILLCELL_X1 FILLER_18_3 ();
 FILLCELL_X4 FILLER_18_21 ();
 FILLCELL_X2 FILLER_18_25 ();
 FILLCELL_X1 FILLER_18_36 ();
 FILLCELL_X2 FILLER_18_41 ();
 FILLCELL_X8 FILLER_18_53 ();
 FILLCELL_X4 FILLER_18_61 ();
 FILLCELL_X1 FILLER_18_65 ();
 FILLCELL_X4 FILLER_18_75 ();
 FILLCELL_X4 FILLER_18_83 ();
 FILLCELL_X2 FILLER_18_87 ();
 FILLCELL_X1 FILLER_18_89 ();
 FILLCELL_X1 FILLER_18_93 ();
 FILLCELL_X16 FILLER_18_109 ();
 FILLCELL_X8 FILLER_18_125 ();
 FILLCELL_X4 FILLER_18_133 ();
 FILLCELL_X2 FILLER_18_137 ();
 FILLCELL_X4 FILLER_18_144 ();
 FILLCELL_X1 FILLER_18_148 ();
 FILLCELL_X2 FILLER_18_166 ();
 FILLCELL_X1 FILLER_18_168 ();
 FILLCELL_X2 FILLER_18_176 ();
 FILLCELL_X8 FILLER_18_198 ();
 FILLCELL_X2 FILLER_18_206 ();
 FILLCELL_X1 FILLER_18_208 ();
 FILLCELL_X2 FILLER_18_215 ();
 FILLCELL_X1 FILLER_18_227 ();
 FILLCELL_X2 FILLER_18_231 ();
 FILLCELL_X1 FILLER_18_233 ();
 FILLCELL_X4 FILLER_18_258 ();
 FILLCELL_X8 FILLER_18_279 ();
 FILLCELL_X4 FILLER_18_287 ();
 FILLCELL_X2 FILLER_18_291 ();
 FILLCELL_X8 FILLER_19_1 ();
 FILLCELL_X4 FILLER_19_9 ();
 FILLCELL_X1 FILLER_19_13 ();
 FILLCELL_X4 FILLER_19_30 ();
 FILLCELL_X2 FILLER_19_34 ();
 FILLCELL_X8 FILLER_19_59 ();
 FILLCELL_X2 FILLER_19_67 ();
 FILLCELL_X1 FILLER_19_69 ();
 FILLCELL_X4 FILLER_19_96 ();
 FILLCELL_X1 FILLER_19_100 ();
 FILLCELL_X16 FILLER_19_107 ();
 FILLCELL_X2 FILLER_19_123 ();
 FILLCELL_X32 FILLER_19_128 ();
 FILLCELL_X1 FILLER_19_160 ();
 FILLCELL_X32 FILLER_19_167 ();
 FILLCELL_X4 FILLER_19_199 ();
 FILLCELL_X1 FILLER_19_206 ();
 FILLCELL_X2 FILLER_19_217 ();
 FILLCELL_X1 FILLER_19_219 ();
 FILLCELL_X2 FILLER_19_237 ();
 FILLCELL_X4 FILLER_19_245 ();
 FILLCELL_X2 FILLER_19_249 ();
 FILLCELL_X1 FILLER_19_251 ();
 FILLCELL_X1 FILLER_19_255 ();
 FILLCELL_X16 FILLER_19_269 ();
 FILLCELL_X8 FILLER_19_285 ();
 FILLCELL_X4 FILLER_20_1 ();
 FILLCELL_X2 FILLER_20_5 ();
 FILLCELL_X8 FILLER_20_36 ();
 FILLCELL_X1 FILLER_20_44 ();
 FILLCELL_X16 FILLER_20_62 ();
 FILLCELL_X2 FILLER_20_78 ();
 FILLCELL_X1 FILLER_20_80 ();
 FILLCELL_X4 FILLER_20_106 ();
 FILLCELL_X1 FILLER_20_110 ();
 FILLCELL_X1 FILLER_20_115 ();
 FILLCELL_X2 FILLER_20_136 ();
 FILLCELL_X2 FILLER_20_174 ();
 FILLCELL_X32 FILLER_20_182 ();
 FILLCELL_X4 FILLER_20_214 ();
 FILLCELL_X1 FILLER_20_218 ();
 FILLCELL_X2 FILLER_20_222 ();
 FILLCELL_X1 FILLER_20_224 ();
 FILLCELL_X8 FILLER_20_236 ();
 FILLCELL_X4 FILLER_20_244 ();
 FILLCELL_X1 FILLER_20_254 ();
 FILLCELL_X2 FILLER_20_259 ();
 FILLCELL_X2 FILLER_20_270 ();
 FILLCELL_X16 FILLER_21_1 ();
 FILLCELL_X4 FILLER_21_17 ();
 FILLCELL_X1 FILLER_21_21 ();
 FILLCELL_X8 FILLER_21_25 ();
 FILLCELL_X2 FILLER_21_33 ();
 FILLCELL_X8 FILLER_21_38 ();
 FILLCELL_X4 FILLER_21_46 ();
 FILLCELL_X2 FILLER_21_50 ();
 FILLCELL_X32 FILLER_21_58 ();
 FILLCELL_X8 FILLER_21_90 ();
 FILLCELL_X4 FILLER_21_98 ();
 FILLCELL_X1 FILLER_21_152 ();
 FILLCELL_X1 FILLER_21_157 ();
 FILLCELL_X1 FILLER_21_165 ();
 FILLCELL_X2 FILLER_21_174 ();
 FILLCELL_X16 FILLER_21_181 ();
 FILLCELL_X8 FILLER_21_204 ();
 FILLCELL_X4 FILLER_21_212 ();
 FILLCELL_X2 FILLER_21_216 ();
 FILLCELL_X1 FILLER_21_237 ();
 FILLCELL_X4 FILLER_21_241 ();
 FILLCELL_X2 FILLER_21_245 ();
 FILLCELL_X1 FILLER_21_247 ();
 FILLCELL_X2 FILLER_21_251 ();
 FILLCELL_X1 FILLER_21_253 ();
 FILLCELL_X16 FILLER_21_257 ();
 FILLCELL_X1 FILLER_22_1 ();
 FILLCELL_X8 FILLER_22_9 ();
 FILLCELL_X2 FILLER_22_17 ();
 FILLCELL_X1 FILLER_22_19 ();
 FILLCELL_X2 FILLER_22_30 ();
 FILLCELL_X2 FILLER_22_52 ();
 FILLCELL_X1 FILLER_22_54 ();
 FILLCELL_X2 FILLER_22_61 ();
 FILLCELL_X4 FILLER_22_75 ();
 FILLCELL_X1 FILLER_22_79 ();
 FILLCELL_X1 FILLER_22_83 ();
 FILLCELL_X2 FILLER_22_88 ();
 FILLCELL_X2 FILLER_22_100 ();
 FILLCELL_X1 FILLER_22_102 ();
 FILLCELL_X4 FILLER_22_109 ();
 FILLCELL_X1 FILLER_22_113 ();
 FILLCELL_X4 FILLER_22_146 ();
 FILLCELL_X8 FILLER_22_160 ();
 FILLCELL_X2 FILLER_22_168 ();
 FILLCELL_X2 FILLER_22_173 ();
 FILLCELL_X1 FILLER_22_175 ();
 FILLCELL_X2 FILLER_22_184 ();
 FILLCELL_X1 FILLER_22_186 ();
 FILLCELL_X4 FILLER_22_202 ();
 FILLCELL_X1 FILLER_22_212 ();
 FILLCELL_X2 FILLER_22_230 ();
 FILLCELL_X1 FILLER_22_232 ();
 FILLCELL_X8 FILLER_22_240 ();
 FILLCELL_X4 FILLER_22_248 ();
 FILLCELL_X4 FILLER_23_1 ();
 FILLCELL_X1 FILLER_23_37 ();
 FILLCELL_X8 FILLER_23_45 ();
 FILLCELL_X2 FILLER_23_53 ();
 FILLCELL_X4 FILLER_23_78 ();
 FILLCELL_X1 FILLER_23_82 ();
 FILLCELL_X4 FILLER_23_100 ();
 FILLCELL_X2 FILLER_23_104 ();
 FILLCELL_X32 FILLER_23_112 ();
 FILLCELL_X16 FILLER_23_144 ();
 FILLCELL_X8 FILLER_23_160 ();
 FILLCELL_X4 FILLER_23_177 ();
 FILLCELL_X2 FILLER_23_181 ();
 FILLCELL_X8 FILLER_23_210 ();
 FILLCELL_X2 FILLER_23_218 ();
 FILLCELL_X4 FILLER_23_237 ();
 FILLCELL_X1 FILLER_23_241 ();
 FILLCELL_X32 FILLER_23_258 ();
 FILLCELL_X2 FILLER_23_290 ();
 FILLCELL_X1 FILLER_23_292 ();
 FILLCELL_X8 FILLER_24_1 ();
 FILLCELL_X2 FILLER_24_29 ();
 FILLCELL_X8 FILLER_24_36 ();
 FILLCELL_X4 FILLER_24_44 ();
 FILLCELL_X1 FILLER_24_51 ();
 FILLCELL_X1 FILLER_24_69 ();
 FILLCELL_X1 FILLER_24_76 ();
 FILLCELL_X1 FILLER_24_82 ();
 FILLCELL_X1 FILLER_24_87 ();
 FILLCELL_X1 FILLER_24_91 ();
 FILLCELL_X16 FILLER_24_98 ();
 FILLCELL_X4 FILLER_24_114 ();
 FILLCELL_X1 FILLER_24_121 ();
 FILLCELL_X8 FILLER_24_126 ();
 FILLCELL_X2 FILLER_24_134 ();
 FILLCELL_X16 FILLER_24_139 ();
 FILLCELL_X4 FILLER_24_155 ();
 FILLCELL_X2 FILLER_24_159 ();
 FILLCELL_X1 FILLER_24_170 ();
 FILLCELL_X1 FILLER_24_180 ();
 FILLCELL_X1 FILLER_24_218 ();
 FILLCELL_X2 FILLER_24_226 ();
 FILLCELL_X1 FILLER_24_228 ();
 FILLCELL_X1 FILLER_24_246 ();
 FILLCELL_X2 FILLER_24_256 ();
 FILLCELL_X8 FILLER_24_284 ();
 FILLCELL_X1 FILLER_24_292 ();
 FILLCELL_X16 FILLER_25_1 ();
 FILLCELL_X2 FILLER_25_17 ();
 FILLCELL_X8 FILLER_25_38 ();
 FILLCELL_X2 FILLER_25_46 ();
 FILLCELL_X1 FILLER_25_71 ();
 FILLCELL_X2 FILLER_25_75 ();
 FILLCELL_X8 FILLER_25_97 ();
 FILLCELL_X1 FILLER_25_131 ();
 FILLCELL_X16 FILLER_25_141 ();
 FILLCELL_X1 FILLER_25_187 ();
 FILLCELL_X8 FILLER_25_209 ();
 FILLCELL_X1 FILLER_25_217 ();
 FILLCELL_X2 FILLER_25_235 ();
 FILLCELL_X8 FILLER_25_244 ();
 FILLCELL_X4 FILLER_25_252 ();
 FILLCELL_X1 FILLER_25_266 ();
 FILLCELL_X16 FILLER_25_270 ();
 FILLCELL_X4 FILLER_25_286 ();
 FILLCELL_X2 FILLER_25_290 ();
 FILLCELL_X1 FILLER_25_292 ();
 FILLCELL_X4 FILLER_26_1 ();
 FILLCELL_X2 FILLER_26_5 ();
 FILLCELL_X1 FILLER_26_7 ();
 FILLCELL_X2 FILLER_26_25 ();
 FILLCELL_X1 FILLER_26_27 ();
 FILLCELL_X2 FILLER_26_35 ();
 FILLCELL_X1 FILLER_26_37 ();
 FILLCELL_X1 FILLER_26_42 ();
 FILLCELL_X8 FILLER_26_60 ();
 FILLCELL_X16 FILLER_26_72 ();
 FILLCELL_X8 FILLER_26_88 ();
 FILLCELL_X4 FILLER_26_96 ();
 FILLCELL_X2 FILLER_26_100 ();
 FILLCELL_X2 FILLER_26_106 ();
 FILLCELL_X2 FILLER_26_111 ();
 FILLCELL_X2 FILLER_26_117 ();
 FILLCELL_X8 FILLER_26_140 ();
 FILLCELL_X4 FILLER_26_148 ();
 FILLCELL_X2 FILLER_26_152 ();
 FILLCELL_X1 FILLER_26_154 ();
 FILLCELL_X1 FILLER_26_188 ();
 FILLCELL_X8 FILLER_26_192 ();
 FILLCELL_X4 FILLER_26_200 ();
 FILLCELL_X2 FILLER_26_208 ();
 FILLCELL_X1 FILLER_26_210 ();
 FILLCELL_X2 FILLER_26_214 ();
 FILLCELL_X4 FILLER_26_240 ();
 FILLCELL_X2 FILLER_26_248 ();
 FILLCELL_X8 FILLER_26_283 ();
 FILLCELL_X2 FILLER_26_291 ();
 FILLCELL_X2 FILLER_27_1 ();
 FILLCELL_X1 FILLER_27_3 ();
 FILLCELL_X16 FILLER_27_27 ();
 FILLCELL_X4 FILLER_27_43 ();
 FILLCELL_X2 FILLER_27_47 ();
 FILLCELL_X2 FILLER_27_56 ();
 FILLCELL_X8 FILLER_27_61 ();
 FILLCELL_X1 FILLER_27_69 ();
 FILLCELL_X2 FILLER_27_90 ();
 FILLCELL_X2 FILLER_27_109 ();
 FILLCELL_X2 FILLER_27_118 ();
 FILLCELL_X4 FILLER_27_130 ();
 FILLCELL_X8 FILLER_27_137 ();
 FILLCELL_X4 FILLER_27_145 ();
 FILLCELL_X2 FILLER_27_149 ();
 FILLCELL_X1 FILLER_27_151 ();
 FILLCELL_X1 FILLER_27_156 ();
 FILLCELL_X4 FILLER_27_161 ();
 FILLCELL_X2 FILLER_27_165 ();
 FILLCELL_X1 FILLER_27_167 ();
 FILLCELL_X1 FILLER_27_184 ();
 FILLCELL_X1 FILLER_27_189 ();
 FILLCELL_X4 FILLER_27_193 ();
 FILLCELL_X2 FILLER_27_197 ();
 FILLCELL_X1 FILLER_27_216 ();
 FILLCELL_X1 FILLER_27_223 ();
 FILLCELL_X2 FILLER_27_233 ();
 FILLCELL_X2 FILLER_27_242 ();
 FILLCELL_X1 FILLER_27_244 ();
 FILLCELL_X4 FILLER_27_252 ();
 FILLCELL_X2 FILLER_27_256 ();
 FILLCELL_X2 FILLER_27_271 ();
 FILLCELL_X16 FILLER_27_277 ();
 FILLCELL_X16 FILLER_28_1 ();
 FILLCELL_X1 FILLER_28_21 ();
 FILLCELL_X1 FILLER_28_39 ();
 FILLCELL_X2 FILLER_28_61 ();
 FILLCELL_X2 FILLER_28_69 ();
 FILLCELL_X1 FILLER_28_75 ();
 FILLCELL_X2 FILLER_28_83 ();
 FILLCELL_X4 FILLER_28_91 ();
 FILLCELL_X2 FILLER_28_95 ();
 FILLCELL_X1 FILLER_28_97 ();
 FILLCELL_X1 FILLER_28_110 ();
 FILLCELL_X1 FILLER_28_116 ();
 FILLCELL_X8 FILLER_28_140 ();
 FILLCELL_X4 FILLER_28_165 ();
 FILLCELL_X8 FILLER_28_189 ();
 FILLCELL_X2 FILLER_28_202 ();
 FILLCELL_X1 FILLER_28_204 ();
 FILLCELL_X8 FILLER_28_208 ();
 FILLCELL_X4 FILLER_28_219 ();
 FILLCELL_X2 FILLER_28_223 ();
 FILLCELL_X1 FILLER_28_225 ();
 FILLCELL_X1 FILLER_28_229 ();
 FILLCELL_X1 FILLER_28_235 ();
 FILLCELL_X4 FILLER_28_242 ();
 FILLCELL_X1 FILLER_28_246 ();
 FILLCELL_X1 FILLER_28_273 ();
 FILLCELL_X16 FILLER_28_277 ();
 FILLCELL_X8 FILLER_29_1 ();
 FILLCELL_X4 FILLER_29_9 ();
 FILLCELL_X1 FILLER_29_13 ();
 FILLCELL_X1 FILLER_29_37 ();
 FILLCELL_X2 FILLER_29_42 ();
 FILLCELL_X1 FILLER_29_44 ();
 FILLCELL_X1 FILLER_29_68 ();
 FILLCELL_X16 FILLER_29_75 ();
 FILLCELL_X8 FILLER_29_91 ();
 FILLCELL_X1 FILLER_29_102 ();
 FILLCELL_X1 FILLER_29_109 ();
 FILLCELL_X2 FILLER_29_119 ();
 FILLCELL_X2 FILLER_29_124 ();
 FILLCELL_X1 FILLER_29_126 ();
 FILLCELL_X32 FILLER_29_144 ();
 FILLCELL_X16 FILLER_29_176 ();
 FILLCELL_X8 FILLER_29_192 ();
 FILLCELL_X4 FILLER_29_200 ();
 FILLCELL_X1 FILLER_29_214 ();
 FILLCELL_X1 FILLER_29_221 ();
 FILLCELL_X1 FILLER_29_229 ();
 FILLCELL_X8 FILLER_29_283 ();
 FILLCELL_X2 FILLER_29_291 ();
 FILLCELL_X8 FILLER_30_1 ();
 FILLCELL_X1 FILLER_30_9 ();
 FILLCELL_X2 FILLER_30_27 ();
 FILLCELL_X2 FILLER_30_36 ();
 FILLCELL_X16 FILLER_30_44 ();
 FILLCELL_X8 FILLER_30_60 ();
 FILLCELL_X4 FILLER_30_68 ();
 FILLCELL_X1 FILLER_30_106 ();
 FILLCELL_X1 FILLER_30_110 ();
 FILLCELL_X2 FILLER_30_142 ();
 FILLCELL_X16 FILLER_30_147 ();
 FILLCELL_X8 FILLER_30_173 ();
 FILLCELL_X4 FILLER_30_181 ();
 FILLCELL_X2 FILLER_30_185 ();
 FILLCELL_X2 FILLER_30_195 ();
 FILLCELL_X1 FILLER_30_197 ();
 FILLCELL_X2 FILLER_30_219 ();
 FILLCELL_X1 FILLER_30_227 ();
 FILLCELL_X1 FILLER_30_238 ();
 FILLCELL_X1 FILLER_30_273 ();
 FILLCELL_X8 FILLER_30_281 ();
 FILLCELL_X4 FILLER_30_289 ();
 FILLCELL_X2 FILLER_31_1 ();
 FILLCELL_X4 FILLER_31_23 ();
 FILLCELL_X2 FILLER_31_27 ();
 FILLCELL_X2 FILLER_31_46 ();
 FILLCELL_X16 FILLER_31_56 ();
 FILLCELL_X8 FILLER_31_72 ();
 FILLCELL_X4 FILLER_31_80 ();
 FILLCELL_X1 FILLER_31_84 ();
 FILLCELL_X4 FILLER_31_106 ();
 FILLCELL_X2 FILLER_31_110 ();
 FILLCELL_X16 FILLER_31_142 ();
 FILLCELL_X2 FILLER_31_158 ();
 FILLCELL_X1 FILLER_31_160 ();
 FILLCELL_X1 FILLER_31_171 ();
 FILLCELL_X2 FILLER_31_178 ();
 FILLCELL_X1 FILLER_31_183 ();
 FILLCELL_X2 FILLER_31_187 ();
 FILLCELL_X1 FILLER_31_215 ();
 FILLCELL_X1 FILLER_31_219 ();
 FILLCELL_X1 FILLER_31_226 ();
 FILLCELL_X4 FILLER_31_234 ();
 FILLCELL_X2 FILLER_31_238 ();
 FILLCELL_X16 FILLER_31_246 ();
 FILLCELL_X4 FILLER_31_262 ();
 FILLCELL_X2 FILLER_31_266 ();
 FILLCELL_X8 FILLER_31_285 ();
 FILLCELL_X2 FILLER_32_1 ();
 FILLCELL_X1 FILLER_32_3 ();
 FILLCELL_X32 FILLER_32_11 ();
 FILLCELL_X4 FILLER_32_43 ();
 FILLCELL_X2 FILLER_32_47 ();
 FILLCELL_X8 FILLER_32_74 ();
 FILLCELL_X4 FILLER_32_82 ();
 FILLCELL_X1 FILLER_32_86 ();
 FILLCELL_X4 FILLER_32_107 ();
 FILLCELL_X2 FILLER_32_111 ();
 FILLCELL_X1 FILLER_32_113 ();
 FILLCELL_X8 FILLER_32_125 ();
 FILLCELL_X4 FILLER_32_133 ();
 FILLCELL_X2 FILLER_32_137 ();
 FILLCELL_X16 FILLER_32_144 ();
 FILLCELL_X8 FILLER_32_205 ();
 FILLCELL_X2 FILLER_32_213 ();
 FILLCELL_X4 FILLER_32_221 ();
 FILLCELL_X2 FILLER_32_249 ();
 FILLCELL_X32 FILLER_32_257 ();
 FILLCELL_X4 FILLER_32_289 ();
 FILLCELL_X4 FILLER_33_1 ();
 FILLCELL_X1 FILLER_33_5 ();
 FILLCELL_X1 FILLER_33_19 ();
 FILLCELL_X16 FILLER_33_27 ();
 FILLCELL_X8 FILLER_33_43 ();
 FILLCELL_X4 FILLER_33_51 ();
 FILLCELL_X2 FILLER_33_55 ();
 FILLCELL_X1 FILLER_33_57 ();
 FILLCELL_X16 FILLER_33_61 ();
 FILLCELL_X1 FILLER_33_77 ();
 FILLCELL_X2 FILLER_33_97 ();
 FILLCELL_X16 FILLER_33_115 ();
 FILLCELL_X1 FILLER_33_154 ();
 FILLCELL_X4 FILLER_33_161 ();
 FILLCELL_X2 FILLER_33_165 ();
 FILLCELL_X2 FILLER_33_177 ();
 FILLCELL_X8 FILLER_33_214 ();
 FILLCELL_X4 FILLER_33_222 ();
 FILLCELL_X2 FILLER_33_226 ();
 FILLCELL_X4 FILLER_33_240 ();
 FILLCELL_X1 FILLER_33_244 ();
 FILLCELL_X8 FILLER_33_251 ();
 FILLCELL_X16 FILLER_33_276 ();
 FILLCELL_X1 FILLER_33_292 ();
 FILLCELL_X16 FILLER_34_1 ();
 FILLCELL_X8 FILLER_34_17 ();
 FILLCELL_X4 FILLER_34_25 ();
 FILLCELL_X2 FILLER_34_29 ();
 FILLCELL_X1 FILLER_34_31 ();
 FILLCELL_X4 FILLER_34_85 ();
 FILLCELL_X1 FILLER_34_109 ();
 FILLCELL_X16 FILLER_34_113 ();
 FILLCELL_X4 FILLER_34_129 ();
 FILLCELL_X2 FILLER_34_133 ();
 FILLCELL_X8 FILLER_34_148 ();
 FILLCELL_X4 FILLER_34_156 ();
 FILLCELL_X16 FILLER_34_163 ();
 FILLCELL_X4 FILLER_34_179 ();
 FILLCELL_X2 FILLER_34_210 ();
 FILLCELL_X1 FILLER_34_212 ();
 FILLCELL_X4 FILLER_34_216 ();
 FILLCELL_X8 FILLER_34_240 ();
 FILLCELL_X2 FILLER_34_248 ();
 FILLCELL_X16 FILLER_34_274 ();
 FILLCELL_X2 FILLER_34_290 ();
 FILLCELL_X1 FILLER_34_292 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X4 FILLER_35_33 ();
 FILLCELL_X2 FILLER_35_66 ();
 FILLCELL_X8 FILLER_35_74 ();
 FILLCELL_X2 FILLER_35_86 ();
 FILLCELL_X1 FILLER_35_105 ();
 FILLCELL_X1 FILLER_35_110 ();
 FILLCELL_X1 FILLER_35_121 ();
 FILLCELL_X4 FILLER_35_125 ();
 FILLCELL_X2 FILLER_35_129 ();
 FILLCELL_X1 FILLER_35_131 ();
 FILLCELL_X8 FILLER_35_152 ();
 FILLCELL_X1 FILLER_35_164 ();
 FILLCELL_X2 FILLER_35_192 ();
 FILLCELL_X1 FILLER_35_194 ();
 FILLCELL_X2 FILLER_35_198 ();
 FILLCELL_X4 FILLER_35_223 ();
 FILLCELL_X8 FILLER_35_230 ();
 FILLCELL_X2 FILLER_35_249 ();
 FILLCELL_X16 FILLER_35_267 ();
 FILLCELL_X8 FILLER_35_283 ();
 FILLCELL_X2 FILLER_35_291 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X16 FILLER_36_33 ();
 FILLCELL_X4 FILLER_36_58 ();
 FILLCELL_X1 FILLER_36_62 ();
 FILLCELL_X8 FILLER_36_67 ();
 FILLCELL_X2 FILLER_36_75 ();
 FILLCELL_X1 FILLER_36_77 ();
 FILLCELL_X4 FILLER_36_85 ();
 FILLCELL_X2 FILLER_36_89 ();
 FILLCELL_X1 FILLER_36_91 ();
 FILLCELL_X1 FILLER_36_95 ();
 FILLCELL_X2 FILLER_36_127 ();
 FILLCELL_X1 FILLER_36_129 ();
 FILLCELL_X8 FILLER_36_147 ();
 FILLCELL_X1 FILLER_36_155 ();
 FILLCELL_X8 FILLER_36_173 ();
 FILLCELL_X2 FILLER_36_181 ();
 FILLCELL_X1 FILLER_36_183 ();
 FILLCELL_X8 FILLER_36_195 ();
 FILLCELL_X1 FILLER_36_203 ();
 FILLCELL_X2 FILLER_36_248 ();
 FILLCELL_X1 FILLER_36_250 ();
 FILLCELL_X32 FILLER_36_258 ();
 FILLCELL_X2 FILLER_36_290 ();
 FILLCELL_X1 FILLER_36_292 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X4 FILLER_37_33 ();
 FILLCELL_X2 FILLER_37_37 ();
 FILLCELL_X4 FILLER_37_60 ();
 FILLCELL_X2 FILLER_37_64 ();
 FILLCELL_X1 FILLER_37_66 ();
 FILLCELL_X16 FILLER_37_84 ();
 FILLCELL_X2 FILLER_37_100 ();
 FILLCELL_X1 FILLER_37_105 ();
 FILLCELL_X8 FILLER_37_109 ();
 FILLCELL_X1 FILLER_37_117 ();
 FILLCELL_X2 FILLER_37_121 ();
 FILLCELL_X2 FILLER_37_140 ();
 FILLCELL_X2 FILLER_37_156 ();
 FILLCELL_X1 FILLER_37_158 ();
 FILLCELL_X16 FILLER_37_163 ();
 FILLCELL_X1 FILLER_37_184 ();
 FILLCELL_X16 FILLER_37_189 ();
 FILLCELL_X8 FILLER_37_212 ();
 FILLCELL_X2 FILLER_37_224 ();
 FILLCELL_X1 FILLER_37_226 ();
 FILLCELL_X16 FILLER_37_266 ();
 FILLCELL_X8 FILLER_37_282 ();
 FILLCELL_X2 FILLER_37_290 ();
 FILLCELL_X1 FILLER_37_292 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X16 FILLER_38_33 ();
 FILLCELL_X4 FILLER_38_49 ();
 FILLCELL_X2 FILLER_38_53 ();
 FILLCELL_X1 FILLER_38_55 ();
 FILLCELL_X16 FILLER_38_63 ();
 FILLCELL_X4 FILLER_38_79 ();
 FILLCELL_X2 FILLER_38_83 ();
 FILLCELL_X32 FILLER_38_92 ();
 FILLCELL_X32 FILLER_38_124 ();
 FILLCELL_X2 FILLER_38_156 ();
 FILLCELL_X1 FILLER_38_158 ();
 FILLCELL_X4 FILLER_38_162 ();
 FILLCELL_X2 FILLER_38_166 ();
 FILLCELL_X1 FILLER_38_168 ();
 FILLCELL_X2 FILLER_38_172 ();
 FILLCELL_X8 FILLER_38_192 ();
 FILLCELL_X2 FILLER_38_200 ();
 FILLCELL_X1 FILLER_38_202 ();
 FILLCELL_X32 FILLER_38_207 ();
 FILLCELL_X32 FILLER_38_239 ();
 FILLCELL_X16 FILLER_38_271 ();
 FILLCELL_X4 FILLER_38_287 ();
 FILLCELL_X2 FILLER_38_291 ();
endmodule
