module fir_filter (clk,
    data_out_valid,
    data_valid,
    rst_n,
    data_in,
    data_out);
 input clk;
 output data_out_valid;
 input data_valid;
 input rst_n;
 input [7:0] data_in;
 output [18:0] data_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire \delay_line[0][0] ;
 wire \delay_line[0][1] ;
 wire \delay_line[0][2] ;
 wire \delay_line[0][3] ;
 wire \delay_line[0][4] ;
 wire \delay_line[0][5] ;
 wire \delay_line[0][6] ;
 wire \delay_line[0][7] ;
 wire \delay_line[1][0] ;
 wire \delay_line[1][1] ;
 wire \delay_line[1][2] ;
 wire \delay_line[1][3] ;
 wire \delay_line[1][4] ;
 wire \delay_line[1][5] ;
 wire \delay_line[1][6] ;
 wire \delay_line[1][7] ;
 wire \delay_line[2][0] ;
 wire \delay_line[2][1] ;
 wire \delay_line[2][2] ;
 wire \delay_line[2][3] ;
 wire \delay_line[2][4] ;
 wire \delay_line[2][5] ;
 wire \delay_line[2][6] ;
 wire \delay_line[2][7] ;
 wire \delay_line[3][0] ;
 wire \delay_line[3][1] ;
 wire \delay_line[3][2] ;
 wire \delay_line[3][3] ;
 wire \delay_line[3][4] ;
 wire \delay_line[3][5] ;
 wire \delay_line[3][6] ;
 wire \delay_line[3][7] ;
 wire \mac_result[0] ;
 wire \mac_result[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net31;

 sky130_fd_sc_hd__inv_1 _169_ (.A(_114_),
    .Y(_142_));
 sky130_fd_sc_hd__inv_1 _170_ (.A(_147_),
    .Y(_143_));
 sky130_fd_sc_hd__inv_1 _171_ (.A(_168_),
    .Y(_144_));
 sky130_fd_sc_hd__clkbuf_2 _172_ (.A(net10),
    .X(_051_));
 sky130_fd_sc_hd__buf_4 _173_ (.A(_051_),
    .X(_052_));
 sky130_fd_sc_hd__mux2_1 _174_ (.A0(\delay_line[0][0] ),
    .A1(net2),
    .S(_052_),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _175_ (.A0(\delay_line[0][1] ),
    .A1(net3),
    .S(_052_),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _176_ (.A0(\delay_line[0][2] ),
    .A1(net4),
    .S(_052_),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _177_ (.A0(\delay_line[0][3] ),
    .A1(net5),
    .S(_052_),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _178_ (.A0(\delay_line[0][4] ),
    .A1(net6),
    .S(_052_),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _179_ (.A0(\delay_line[0][5] ),
    .A1(net7),
    .S(_052_),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _180_ (.A0(\delay_line[0][6] ),
    .A1(net8),
    .S(_052_),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _181_ (.A0(\delay_line[0][7] ),
    .A1(net9),
    .S(_052_),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _182_ (.A0(\delay_line[1][0] ),
    .A1(\delay_line[0][0] ),
    .S(_052_),
    .X(_008_));
 sky130_fd_sc_hd__buf_4 _183_ (.A(_051_),
    .X(_053_));
 sky130_fd_sc_hd__mux2_1 _184_ (.A0(\delay_line[1][1] ),
    .A1(\delay_line[0][1] ),
    .S(_053_),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _185_ (.A0(\delay_line[1][2] ),
    .A1(\delay_line[0][2] ),
    .S(_053_),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _186_ (.A0(\delay_line[1][3] ),
    .A1(\delay_line[0][3] ),
    .S(_053_),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _187_ (.A0(\delay_line[1][4] ),
    .A1(\delay_line[0][4] ),
    .S(_053_),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _188_ (.A0(\delay_line[1][5] ),
    .A1(\delay_line[0][5] ),
    .S(_053_),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _189_ (.A0(\delay_line[1][6] ),
    .A1(\delay_line[0][6] ),
    .S(_053_),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _190_ (.A0(\delay_line[1][7] ),
    .A1(\delay_line[0][7] ),
    .S(_053_),
    .X(_015_));
 sky130_fd_sc_hd__mux2_1 _191_ (.A0(\delay_line[2][0] ),
    .A1(\delay_line[1][0] ),
    .S(_053_),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _192_ (.A0(\delay_line[2][1] ),
    .A1(\delay_line[1][1] ),
    .S(_053_),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _193_ (.A0(\delay_line[2][2] ),
    .A1(\delay_line[1][2] ),
    .S(_053_),
    .X(_018_));
 sky130_fd_sc_hd__buf_4 _194_ (.A(_051_),
    .X(_054_));
 sky130_fd_sc_hd__mux2_1 _195_ (.A0(\delay_line[2][3] ),
    .A1(\delay_line[1][3] ),
    .S(_054_),
    .X(_019_));
 sky130_fd_sc_hd__mux2_1 _196_ (.A0(\delay_line[2][4] ),
    .A1(\delay_line[1][4] ),
    .S(_054_),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _197_ (.A0(\delay_line[2][5] ),
    .A1(\delay_line[1][5] ),
    .S(_054_),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _198_ (.A0(\delay_line[2][6] ),
    .A1(\delay_line[1][6] ),
    .S(_054_),
    .X(_022_));
 sky130_fd_sc_hd__mux2_1 _199_ (.A0(\delay_line[2][7] ),
    .A1(\delay_line[1][7] ),
    .S(_054_),
    .X(_023_));
 sky130_fd_sc_hd__mux2_1 _200_ (.A0(\delay_line[3][0] ),
    .A1(\delay_line[2][0] ),
    .S(_054_),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _201_ (.A0(\delay_line[3][1] ),
    .A1(\delay_line[2][1] ),
    .S(_054_),
    .X(_025_));
 sky130_fd_sc_hd__mux2_1 _202_ (.A0(\delay_line[3][2] ),
    .A1(\delay_line[2][2] ),
    .S(_054_),
    .X(_026_));
 sky130_fd_sc_hd__mux2_1 _203_ (.A0(\delay_line[3][3] ),
    .A1(\delay_line[2][3] ),
    .S(_054_),
    .X(_027_));
 sky130_fd_sc_hd__mux2_1 _204_ (.A0(\delay_line[3][4] ),
    .A1(\delay_line[2][4] ),
    .S(_054_),
    .X(_028_));
 sky130_fd_sc_hd__buf_4 _205_ (.A(_051_),
    .X(_055_));
 sky130_fd_sc_hd__mux2_1 _206_ (.A0(\delay_line[3][5] ),
    .A1(\delay_line[2][5] ),
    .S(_055_),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _207_ (.A0(\delay_line[3][6] ),
    .A1(\delay_line[2][6] ),
    .S(_055_),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _208_ (.A0(\delay_line[3][7] ),
    .A1(\delay_line[2][7] ),
    .S(_055_),
    .X(_031_));
 sky130_fd_sc_hd__mux2_1 _209_ (.A0(net11),
    .A1(\mac_result[0] ),
    .S(_055_),
    .X(_032_));
 sky130_fd_sc_hd__inv_1 _210_ (.A(_055_),
    .Y(_056_));
 sky130_fd_sc_hd__a21o_1 _211_ (.A1(_160_),
    .A2(_157_),
    .B1(_159_),
    .X(_057_));
 sky130_fd_sc_hd__a211oi_1 _212_ (.A1(_149_),
    .A2(_168_),
    .B1(_148_),
    .C1(_151_),
    .Y(_058_));
 sky130_fd_sc_hd__o211ai_1 _213_ (.A1(_152_),
    .A2(_151_),
    .B1(_156_),
    .C1(_154_),
    .Y(_059_));
 sky130_fd_sc_hd__a21oi_1 _214_ (.A1(_156_),
    .A2(_153_),
    .B1(_155_),
    .Y(_060_));
 sky130_fd_sc_hd__o21ai_2 _215_ (.A1(_058_),
    .A2(_059_),
    .B1(_060_),
    .Y(_061_));
 sky130_fd_sc_hd__o21ai_0 _216_ (.A1(_158_),
    .A2(_157_),
    .B1(_160_),
    .Y(_062_));
 sky130_fd_sc_hd__nand2b_1 _217_ (.A_N(_159_),
    .B(_062_),
    .Y(_063_));
 sky130_fd_sc_hd__o2111ai_2 _218_ (.A1(_057_),
    .A2(_061_),
    .B1(_063_),
    .C1(_164_),
    .D1(_162_),
    .Y(_064_));
 sky130_fd_sc_hd__a21oi_1 _219_ (.A1(_164_),
    .A2(_161_),
    .B1(_163_),
    .Y(_065_));
 sky130_fd_sc_hd__a21boi_0 _220_ (.A1(_064_),
    .A2(_065_),
    .B1_N(_166_),
    .Y(_066_));
 sky130_fd_sc_hd__and3b_1 _221_ (.A_N(_166_),
    .B(_064_),
    .C(_065_),
    .X(_067_));
 sky130_fd_sc_hd__nand2_1 _222_ (.A(_056_),
    .B(net12),
    .Y(_068_));
 sky130_fd_sc_hd__o31ai_1 _223_ (.A1(_056_),
    .A2(_066_),
    .A3(_067_),
    .B1(_068_),
    .Y(_033_));
 sky130_fd_sc_hd__nor3b_1 _224_ (.A(_163_),
    .B(_165_),
    .C_N(_166_),
    .Y(_069_));
 sky130_fd_sc_hd__a21oi_1 _225_ (.A1(_162_),
    .A2(_057_),
    .B1(_161_),
    .Y(_070_));
 sky130_fd_sc_hd__nor2b_1 _226_ (.A(_145_),
    .B_N(_152_),
    .Y(_071_));
 sky130_fd_sc_hd__o211ai_1 _227_ (.A1(_151_),
    .A2(_071_),
    .B1(_154_),
    .C1(_156_),
    .Y(_072_));
 sky130_fd_sc_hd__nand3_1 _228_ (.A(_158_),
    .B(_160_),
    .C(_162_),
    .Y(_073_));
 sky130_fd_sc_hd__a21o_1 _229_ (.A1(_060_),
    .A2(_072_),
    .B1(_073_),
    .X(_074_));
 sky130_fd_sc_hd__inv_1 _230_ (.A(_164_),
    .Y(_075_));
 sky130_fd_sc_hd__inv_1 _231_ (.A(_165_),
    .Y(_076_));
 sky130_fd_sc_hd__o21ai_1 _232_ (.A1(_166_),
    .A2(_076_),
    .B1(_051_),
    .Y(_077_));
 sky130_fd_sc_hd__a21o_1 _233_ (.A1(_075_),
    .A2(_069_),
    .B1(_077_),
    .X(_078_));
 sky130_fd_sc_hd__a31oi_2 _234_ (.A1(_069_),
    .A2(_070_),
    .A3(_074_),
    .B1(_078_),
    .Y(_079_));
 sky130_fd_sc_hd__buf_2 _235_ (.A(_051_),
    .X(_080_));
 sky130_fd_sc_hd__nor2_1 _236_ (.A(_080_),
    .B(net13),
    .Y(_081_));
 sky130_fd_sc_hd__nor2_1 _237_ (.A(_079_),
    .B(_081_),
    .Y(_034_));
 sky130_fd_sc_hd__nand2_1 _238_ (.A(_164_),
    .B(_161_),
    .Y(_082_));
 sky130_fd_sc_hd__a31oi_2 _239_ (.A1(_064_),
    .A2(_082_),
    .A3(_069_),
    .B1(_077_),
    .Y(_083_));
 sky130_fd_sc_hd__nor2_1 _240_ (.A(_080_),
    .B(net14),
    .Y(_084_));
 sky130_fd_sc_hd__nor2_1 _241_ (.A(_083_),
    .B(_084_),
    .Y(_035_));
 sky130_fd_sc_hd__nor2_1 _242_ (.A(_080_),
    .B(net15),
    .Y(_085_));
 sky130_fd_sc_hd__nor2_1 _243_ (.A(_079_),
    .B(_085_),
    .Y(_036_));
 sky130_fd_sc_hd__nor2_1 _244_ (.A(_080_),
    .B(net16),
    .Y(_086_));
 sky130_fd_sc_hd__nor2_1 _245_ (.A(_083_),
    .B(_086_),
    .Y(_037_));
 sky130_fd_sc_hd__nor2_1 _246_ (.A(_080_),
    .B(net17),
    .Y(_087_));
 sky130_fd_sc_hd__nor2_1 _247_ (.A(_079_),
    .B(_087_),
    .Y(_038_));
 sky130_fd_sc_hd__nor2_1 _248_ (.A(_080_),
    .B(net18),
    .Y(_088_));
 sky130_fd_sc_hd__nor2_1 _249_ (.A(_083_),
    .B(_088_),
    .Y(_039_));
 sky130_fd_sc_hd__nor2_1 _250_ (.A(_080_),
    .B(net19),
    .Y(_089_));
 sky130_fd_sc_hd__nor2_1 _251_ (.A(_079_),
    .B(_089_),
    .Y(_040_));
 sky130_fd_sc_hd__nor2_1 _252_ (.A(_080_),
    .B(net20),
    .Y(_090_));
 sky130_fd_sc_hd__nor2_1 _253_ (.A(_083_),
    .B(_090_),
    .Y(_041_));
 sky130_fd_sc_hd__mux2_1 _254_ (.A0(net21),
    .A1(\mac_result[1] ),
    .S(_055_),
    .X(_042_));
 sky130_fd_sc_hd__nand2_1 _255_ (.A(_056_),
    .B(net22),
    .Y(_091_));
 sky130_fd_sc_hd__o21ai_0 _256_ (.A1(_146_),
    .A2(_056_),
    .B1(_091_),
    .Y(_043_));
 sky130_fd_sc_hd__xnor2_1 _257_ (.A(_152_),
    .B(_145_),
    .Y(_092_));
 sky130_fd_sc_hd__mux2_1 _258_ (.A0(net23),
    .A1(_092_),
    .S(_055_),
    .X(_044_));
 sky130_fd_sc_hd__a21o_1 _259_ (.A1(_149_),
    .A2(_168_),
    .B1(_148_),
    .X(_093_));
 sky130_fd_sc_hd__a21oi_1 _260_ (.A1(_152_),
    .A2(_093_),
    .B1(_151_),
    .Y(_094_));
 sky130_fd_sc_hd__xnor2_1 _261_ (.A(_154_),
    .B(_094_),
    .Y(_095_));
 sky130_fd_sc_hd__mux2_1 _262_ (.A0(net24),
    .A1(_095_),
    .S(_055_),
    .X(_045_));
 sky130_fd_sc_hd__o21a_1 _263_ (.A1(_151_),
    .A2(_071_),
    .B1(_154_),
    .X(_096_));
 sky130_fd_sc_hd__nor2_1 _264_ (.A(_153_),
    .B(_096_),
    .Y(_097_));
 sky130_fd_sc_hd__xnor2_1 _265_ (.A(_156_),
    .B(_097_),
    .Y(_098_));
 sky130_fd_sc_hd__mux2_1 _266_ (.A0(net25),
    .A1(_098_),
    .S(_055_),
    .X(_046_));
 sky130_fd_sc_hd__xor2_1 _267_ (.A(_158_),
    .B(_061_),
    .X(_099_));
 sky130_fd_sc_hd__mux2_1 _268_ (.A0(net26),
    .A1(_099_),
    .S(_055_),
    .X(_047_));
 sky130_fd_sc_hd__a21boi_0 _269_ (.A1(_060_),
    .A2(_072_),
    .B1_N(_158_),
    .Y(_100_));
 sky130_fd_sc_hd__o21ai_0 _270_ (.A1(_157_),
    .A2(_100_),
    .B1(_160_),
    .Y(_101_));
 sky130_fd_sc_hd__or3_1 _271_ (.A(_160_),
    .B(_157_),
    .C(_100_),
    .X(_102_));
 sky130_fd_sc_hd__nor2b_1 _272_ (.A(_051_),
    .B_N(net27),
    .Y(_103_));
 sky130_fd_sc_hd__a31o_1 _273_ (.A1(_052_),
    .A2(_101_),
    .A3(_102_),
    .B1(_103_),
    .X(_048_));
 sky130_fd_sc_hd__o21ai_0 _274_ (.A1(_057_),
    .A2(_061_),
    .B1(_063_),
    .Y(_104_));
 sky130_fd_sc_hd__xor2_1 _275_ (.A(_162_),
    .B(_104_),
    .X(_105_));
 sky130_fd_sc_hd__nor2_1 _276_ (.A(_080_),
    .B(net28),
    .Y(_106_));
 sky130_fd_sc_hd__a21oi_1 _277_ (.A1(_080_),
    .A2(_105_),
    .B1(_106_),
    .Y(_049_));
 sky130_fd_sc_hd__and3_1 _278_ (.A(_075_),
    .B(_070_),
    .C(_074_),
    .X(_107_));
 sky130_fd_sc_hd__a21oi_1 _279_ (.A1(_070_),
    .A2(_074_),
    .B1(_075_),
    .Y(_108_));
 sky130_fd_sc_hd__nand2_1 _280_ (.A(_056_),
    .B(net29),
    .Y(_109_));
 sky130_fd_sc_hd__o31ai_1 _281_ (.A1(_056_),
    .A2(_107_),
    .A3(_108_),
    .B1(_109_),
    .Y(_050_));
 sky130_fd_sc_hd__fa_1 _282_ (.A(\delay_line[0][2] ),
    .B(\delay_line[1][1] ),
    .CIN(\delay_line[2][1] ),
    .COUT(_110_),
    .SUM(_111_));
 sky130_fd_sc_hd__fa_1 _283_ (.A(\delay_line[3][2] ),
    .B(_111_),
    .CIN(_112_),
    .COUT(_113_),
    .SUM(_114_));
 sky130_fd_sc_hd__fa_1 _284_ (.A(\delay_line[0][1] ),
    .B(\delay_line[1][0] ),
    .CIN(\delay_line[2][0] ),
    .COUT(_112_),
    .SUM(_115_));
 sky130_fd_sc_hd__fa_1 _285_ (.A(\delay_line[0][3] ),
    .B(\delay_line[1][2] ),
    .CIN(\delay_line[2][2] ),
    .COUT(_116_),
    .SUM(_117_));
 sky130_fd_sc_hd__fa_1 _286_ (.A(\delay_line[3][3] ),
    .B(_117_),
    .CIN(_110_),
    .COUT(_118_),
    .SUM(_119_));
 sky130_fd_sc_hd__fa_1 _287_ (.A(\delay_line[0][4] ),
    .B(\delay_line[1][3] ),
    .CIN(\delay_line[2][3] ),
    .COUT(_120_),
    .SUM(_121_));
 sky130_fd_sc_hd__fa_1 _288_ (.A(\delay_line[3][4] ),
    .B(_121_),
    .CIN(_116_),
    .COUT(_122_),
    .SUM(_123_));
 sky130_fd_sc_hd__fa_1 _289_ (.A(\delay_line[0][5] ),
    .B(\delay_line[1][4] ),
    .CIN(\delay_line[2][4] ),
    .COUT(_124_),
    .SUM(_125_));
 sky130_fd_sc_hd__fa_1 _290_ (.A(\delay_line[3][5] ),
    .B(_125_),
    .CIN(_120_),
    .COUT(_126_),
    .SUM(_127_));
 sky130_fd_sc_hd__fa_1 _291_ (.A(\delay_line[0][6] ),
    .B(\delay_line[1][5] ),
    .CIN(\delay_line[2][5] ),
    .COUT(_128_),
    .SUM(_129_));
 sky130_fd_sc_hd__fa_1 _292_ (.A(\delay_line[3][6] ),
    .B(_129_),
    .CIN(_124_),
    .COUT(_130_),
    .SUM(_131_));
 sky130_fd_sc_hd__fa_1 _293_ (.A(\delay_line[0][7] ),
    .B(\delay_line[1][6] ),
    .CIN(\delay_line[2][6] ),
    .COUT(_132_),
    .SUM(_133_));
 sky130_fd_sc_hd__fa_1 _294_ (.A(\delay_line[3][7] ),
    .B(_133_),
    .CIN(_128_),
    .COUT(_134_),
    .SUM(_135_));
 sky130_fd_sc_hd__fa_1 _295_ (.A(\delay_line[0][7] ),
    .B(\delay_line[1][7] ),
    .CIN(\delay_line[2][7] ),
    .COUT(_136_),
    .SUM(_137_));
 sky130_fd_sc_hd__fa_1 _296_ (.A(\delay_line[3][7] ),
    .B(_137_),
    .CIN(_132_),
    .COUT(_138_),
    .SUM(_139_));
 sky130_fd_sc_hd__fa_1 _297_ (.A(\delay_line[3][7] ),
    .B(_137_),
    .CIN(_136_),
    .COUT(_140_),
    .SUM(_141_));
 sky130_fd_sc_hd__fa_1 _298_ (.A(_142_),
    .B(_143_),
    .CIN(_144_),
    .COUT(_145_),
    .SUM(_146_));
 sky130_fd_sc_hd__ha_1 _299_ (.A(_114_),
    .B(_147_),
    .COUT(_148_),
    .SUM(_149_));
 sky130_fd_sc_hd__ha_1 _300_ (.A(\delay_line[3][1] ),
    .B(_115_),
    .COUT(_147_),
    .SUM(_150_));
 sky130_fd_sc_hd__ha_1 _301_ (.A(_119_),
    .B(_113_),
    .COUT(_151_),
    .SUM(_152_));
 sky130_fd_sc_hd__ha_1 _302_ (.A(_123_),
    .B(_118_),
    .COUT(_153_),
    .SUM(_154_));
 sky130_fd_sc_hd__ha_1 _303_ (.A(_127_),
    .B(_122_),
    .COUT(_155_),
    .SUM(_156_));
 sky130_fd_sc_hd__ha_1 _304_ (.A(_131_),
    .B(_126_),
    .COUT(_157_),
    .SUM(_158_));
 sky130_fd_sc_hd__ha_1 _305_ (.A(_135_),
    .B(_130_),
    .COUT(_159_),
    .SUM(_160_));
 sky130_fd_sc_hd__ha_1 _306_ (.A(_139_),
    .B(_134_),
    .COUT(_161_),
    .SUM(_162_));
 sky130_fd_sc_hd__ha_1 _307_ (.A(_141_),
    .B(_138_),
    .COUT(_163_),
    .SUM(_164_));
 sky130_fd_sc_hd__ha_1 _308_ (.A(_141_),
    .B(_140_),
    .COUT(_165_),
    .SUM(_166_));
 sky130_fd_sc_hd__ha_1 _309_ (.A(\delay_line[0][0] ),
    .B(\delay_line[3][0] ),
    .COUT(_167_),
    .SUM(\mac_result[0] ));
 sky130_fd_sc_hd__ha_1 _310_ (.A(_150_),
    .B(_167_),
    .COUT(_168_),
    .SUM(\mac_result[1] ));
 sky130_fd_sc_hd__dfrtp_1 \data_out_valid$_DFF_PN0_  (.D(net10),
    .Q(net30),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[0][0]$_DFFE_PN0P_  (.D(_000_),
    .Q(\delay_line[0][0] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[0][1]$_DFFE_PN0P_  (.D(_001_),
    .Q(\delay_line[0][1] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[0][2]$_DFFE_PN0P_  (.D(_002_),
    .Q(\delay_line[0][2] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[0][3]$_DFFE_PN0P_  (.D(_003_),
    .Q(\delay_line[0][3] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[0][4]$_DFFE_PN0P_  (.D(_004_),
    .Q(\delay_line[0][4] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[0][5]$_DFFE_PN0P_  (.D(_005_),
    .Q(\delay_line[0][5] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[0][6]$_DFFE_PN0P_  (.D(_006_),
    .Q(\delay_line[0][6] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[0][7]$_DFFE_PN0P_  (.D(_007_),
    .Q(\delay_line[0][7] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[1][0]$_DFFE_PN0P_  (.D(_008_),
    .Q(\delay_line[1][0] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[1][1]$_DFFE_PN0P_  (.D(_009_),
    .Q(\delay_line[1][1] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[1][2]$_DFFE_PN0P_  (.D(_010_),
    .Q(\delay_line[1][2] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[1][3]$_DFFE_PN0P_  (.D(_011_),
    .Q(\delay_line[1][3] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[1][4]$_DFFE_PN0P_  (.D(_012_),
    .Q(\delay_line[1][4] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[1][5]$_DFFE_PN0P_  (.D(_013_),
    .Q(\delay_line[1][5] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[1][6]$_DFFE_PN0P_  (.D(_014_),
    .Q(\delay_line[1][6] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[1][7]$_DFFE_PN0P_  (.D(_015_),
    .Q(\delay_line[1][7] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[2][0]$_DFFE_PN0P_  (.D(_016_),
    .Q(\delay_line[2][0] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[2][1]$_DFFE_PN0P_  (.D(_017_),
    .Q(\delay_line[2][1] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[2][2]$_DFFE_PN0P_  (.D(_018_),
    .Q(\delay_line[2][2] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[2][3]$_DFFE_PN0P_  (.D(_019_),
    .Q(\delay_line[2][3] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[2][4]$_DFFE_PN0P_  (.D(_020_),
    .Q(\delay_line[2][4] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[2][5]$_DFFE_PN0P_  (.D(_021_),
    .Q(\delay_line[2][5] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[2][6]$_DFFE_PN0P_  (.D(_022_),
    .Q(\delay_line[2][6] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[2][7]$_DFFE_PN0P_  (.D(_023_),
    .Q(\delay_line[2][7] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[3][0]$_DFFE_PN0P_  (.D(_024_),
    .Q(\delay_line[3][0] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[3][1]$_DFFE_PN0P_  (.D(_025_),
    .Q(\delay_line[3][1] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[3][2]$_DFFE_PN0P_  (.D(_026_),
    .Q(\delay_line[3][2] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[3][3]$_DFFE_PN0P_  (.D(_027_),
    .Q(\delay_line[3][3] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[3][4]$_DFFE_PN0P_  (.D(_028_),
    .Q(\delay_line[3][4] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[3][5]$_DFFE_PN0P_  (.D(_029_),
    .Q(\delay_line[3][5] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \delay_line[3][6]$_DFFE_PN0P_  (.D(_030_),
    .Q(\delay_line[3][6] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \delay_line[3][7]$_DFFE_PN0P_  (.D(_031_),
    .Q(\delay_line[3][7] ),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[0]$_DFFE_PN0P_  (.D(_032_),
    .Q(net11),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[10]$_DFFE_PN0P_  (.D(_033_),
    .Q(net12),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[11]$_DFFE_PN0P_  (.D(_034_),
    .Q(net13),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[12]$_DFFE_PN0P_  (.D(_035_),
    .Q(net14),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[13]$_DFFE_PN0P_  (.D(_036_),
    .Q(net15),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[14]$_DFFE_PN0P_  (.D(_037_),
    .Q(net16),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[15]$_DFFE_PN0P_  (.D(_038_),
    .Q(net17),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[16]$_DFFE_PN0P_  (.D(_039_),
    .Q(net18),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[17]$_DFFE_PN0P_  (.D(_040_),
    .Q(net19),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[18]$_DFFE_PN0P_  (.D(_041_),
    .Q(net20),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[1]$_DFFE_PN0P_  (.D(_042_),
    .Q(net21),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[2]$_DFFE_PN0P_  (.D(_043_),
    .Q(net22),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[3]$_DFFE_PN0P_  (.D(_044_),
    .Q(net23),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[4]$_DFFE_PN0P_  (.D(_045_),
    .Q(net24),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[5]$_DFFE_PN0P_  (.D(_046_),
    .Q(net25),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[6]$_DFFE_PN0P_  (.D(_047_),
    .Q(net26),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[7]$_DFFE_PN0P_  (.D(_048_),
    .Q(net27),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[8]$_DFFE_PN0P_  (.D(_049_),
    .Q(net28),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \result[9]$_DFFE_PN0P_  (.D(_050_),
    .Q(net29),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__buf_12 hold1 (.A(net31),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_51 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(data_in[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(data_in[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(data_in[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(data_in[3]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(data_in[4]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(data_in[5]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(data_in[6]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(data_in[7]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(data_valid),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 output10 (.A(net11),
    .X(data_out[0]));
 sky130_fd_sc_hd__clkbuf_1 output11 (.A(net12),
    .X(data_out[10]));
 sky130_fd_sc_hd__clkbuf_1 output12 (.A(net13),
    .X(data_out[11]));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net14),
    .X(data_out[12]));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net15),
    .X(data_out[13]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net16),
    .X(data_out[14]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net17),
    .X(data_out[15]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net18),
    .X(data_out[16]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net19),
    .X(data_out[17]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net20),
    .X(data_out[18]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net21),
    .X(data_out[1]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net22),
    .X(data_out[2]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net23),
    .X(data_out[3]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net24),
    .X(data_out[4]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net25),
    .X(data_out[5]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net26),
    .X(data_out[6]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net27),
    .X(data_out[7]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net28),
    .X(data_out[8]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net29),
    .X(data_out[9]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net30),
    .X(data_out_valid));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload0 (.A(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload1 (.A(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload2 (.A(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net31));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_30 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_30 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_38 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_42 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_34 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_43 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_4 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_26 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_149 ();
endmodule
