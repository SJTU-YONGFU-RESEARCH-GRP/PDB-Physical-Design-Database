module spi_master (clk,
    rst_n,
    rx_valid,
    spi_clk,
    spi_cs_n,
    spi_miso,
    spi_mosi,
    tx_ready,
    tx_valid,
    rx_data,
    tx_data);
 input clk;
 input rst_n;
 output rx_valid;
 output spi_clk;
 output spi_cs_n;
 input spi_miso;
 output spi_mosi;
 output tx_ready;
 input tx_valid;
 output [7:0] rx_data;
 input [7:0] tx_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire \bit_count[0] ;
 wire \bit_count[1] ;
 wire \bit_count[2] ;
 wire \bit_count[3] ;
 wire \debug_miso_samples[0] ;
 wire \debug_miso_samples[1] ;
 wire \debug_miso_samples[2] ;
 wire \debug_miso_samples[3] ;
 wire \debug_miso_samples[4] ;
 wire \debug_miso_samples[5] ;
 wire \debug_miso_samples[6] ;
 wire \debug_miso_samples[7] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \tx_shift[0] ;
 wire \tx_shift[1] ;
 wire \tx_shift[2] ;
 wire \tx_shift[3] ;
 wire \tx_shift[4] ;
 wire \tx_shift[5] ;
 wire \tx_shift[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net26;

 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _137_ (.I(\bit_count[3] ),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _138_ (.A1(\bit_count[2] ),
    .A2(_117_),
    .A3(_132_),
    .ZN(_118_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _139_ (.I(_118_),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _140_ (.A1(\bit_count[2] ),
    .A2(\bit_count[1] ),
    .A3(\bit_count[0] ),
    .ZN(_134_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _141_ (.A1(\bit_count[3] ),
    .A2(_134_),
    .Z(_126_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _142_ (.A1(\bit_count[2] ),
    .A2(_117_),
    .A3(_132_),
    .ZN(_129_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _143_ (.I(\state[1] ),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _144_ (.I(net22),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _145_ (.A1(_034_),
    .A2(_035_),
    .Z(_036_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _146_ (.I(\bit_count[0] ),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _147_ (.I0(net22),
    .I1(_036_),
    .S(_037_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_4 _148_ (.A1(\state[0] ),
    .A2(net12),
    .B(_034_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _149_ (.A1(\state[0] ),
    .A2(_038_),
    .B1(_039_),
    .B2(\bit_count[0] ),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _150_ (.I(_040_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 _151_ (.I(\state[0] ),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _152_ (.A1(net22),
    .A2(\bit_count[1] ),
    .B1(_133_),
    .B2(_036_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _153_ (.A1(\bit_count[1] ),
    .A2(_039_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _154_ (.A1(_041_),
    .A2(_042_),
    .B(_043_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _155_ (.A1(\state[1] ),
    .A2(\bit_count[2] ),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _156_ (.A1(_035_),
    .A2(_132_),
    .Z(_045_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _157_ (.I0(\bit_count[2] ),
    .I1(_044_),
    .S(_045_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _158_ (.A1(\bit_count[2] ),
    .A2(_039_),
    .B1(_046_),
    .B2(\state[0] ),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _159_ (.I(_047_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _160_ (.I(net12),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _161_ (.A1(_041_),
    .A2(_048_),
    .B(\state[1] ),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _162_ (.A1(net22),
    .A2(\bit_count[3] ),
    .B1(_136_),
    .B2(_036_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _163_ (.A1(_117_),
    .A2(_049_),
    .B1(_050_),
    .B2(_041_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _164_ (.I(\debug_miso_samples[0] ),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _165_ (.I(_131_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _166_ (.A1(_120_),
    .A2(_128_),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _167_ (.A1(_130_),
    .A2(_135_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _168_ (.A1(_052_),
    .A2(_127_),
    .A3(_053_),
    .A4(_054_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _169_ (.A1(_120_),
    .A2(_128_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _170_ (.A1(_130_),
    .A2(_135_),
    .Z(_057_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _171_ (.A1(_052_),
    .A2(_127_),
    .A3(_056_),
    .A4(_057_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _172_ (.A1(\bit_count[2] ),
    .A2(_132_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _173_ (.A1(_124_),
    .A2(_121_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _174_ (.A1(\bit_count[0] ),
    .A2(_059_),
    .A3(_060_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _175_ (.I(_133_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _176_ (.A1(_120_),
    .A2(_062_),
    .A3(_136_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _177_ (.A1(_055_),
    .A2(_058_),
    .B(_061_),
    .C(_063_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _178_ (.A1(_034_),
    .A2(\state[0] ),
    .A3(_035_),
    .Z(_065_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _179_ (.A1(\state[0] ),
    .A2(net22),
    .Z(_066_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _180_ (.A1(\state[1] ),
    .A2(_066_),
    .Z(_067_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _181_ (.A1(_064_),
    .A2(_065_),
    .B(_067_),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _182_ (.A1(net3),
    .A2(_065_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _183_ (.A1(_051_),
    .A2(_068_),
    .B1(_069_),
    .B2(_064_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _184_ (.A1(\debug_miso_samples[1] ),
    .A2(_067_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _185_ (.I(_136_),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_4 _186_ (.A1(_055_),
    .A2(_058_),
    .B(_133_),
    .C(_071_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _187_ (.A1(_124_),
    .A2(_121_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _188_ (.A1(\bit_count[0] ),
    .A2(_120_),
    .A3(_059_),
    .A4(_073_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _189_ (.A1(_072_),
    .A2(_074_),
    .B(\debug_miso_samples[1] ),
    .C(_065_),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _190_ (.A1(_069_),
    .A2(_072_),
    .A3(_074_),
    .Z(_076_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _191_ (.A1(_070_),
    .A2(_075_),
    .A3(_076_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _192_ (.A1(\debug_miso_samples[2] ),
    .A2(_067_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _193_ (.A1(_037_),
    .A2(_120_),
    .A3(_059_),
    .A4(_073_),
    .Z(_078_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _194_ (.A1(_072_),
    .A2(_078_),
    .B(\debug_miso_samples[2] ),
    .C(_065_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _195_ (.A1(_069_),
    .A2(_072_),
    .A3(_078_),
    .Z(_080_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _196_ (.A1(_077_),
    .A2(_079_),
    .A3(_080_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _197_ (.A1(_055_),
    .A2(_058_),
    .B(_071_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _198_ (.A1(_133_),
    .A2(_069_),
    .A3(_081_),
    .Z(_082_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _199_ (.A1(_035_),
    .A2(_062_),
    .B(_041_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _200_ (.A1(\state[1] ),
    .A2(_074_),
    .A3(_083_),
    .Z(_084_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _201_ (.A1(_034_),
    .A2(_041_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _202_ (.A1(_081_),
    .A2(_084_),
    .B(_085_),
    .C(\debug_miso_samples[3] ),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _203_ (.A1(_074_),
    .A2(_082_),
    .B(_086_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _204_ (.A1(_133_),
    .A2(_067_),
    .A3(_078_),
    .Z(_087_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _205_ (.A1(_081_),
    .A2(_087_),
    .B(_085_),
    .C(\debug_miso_samples[4] ),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _206_ (.A1(_078_),
    .A2(_082_),
    .B(_088_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _207_ (.A1(\debug_miso_samples[5] ),
    .A2(_067_),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _208_ (.I(_120_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu9t5v0__nand4_4 _209_ (.A1(_037_),
    .A2(_090_),
    .A3(_059_),
    .A4(_060_),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _210_ (.A1(_072_),
    .A2(_091_),
    .B(\debug_miso_samples[5] ),
    .C(_065_),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _211_ (.A1(_069_),
    .A2(_072_),
    .A3(_091_),
    .Z(_093_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _212_ (.A1(_089_),
    .A2(_092_),
    .A3(_093_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _213_ (.A1(\debug_miso_samples[6] ),
    .A2(_067_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _214_ (.A1(\bit_count[0] ),
    .A2(_059_),
    .A3(_060_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _215_ (.A1(\debug_miso_samples[6] ),
    .A2(_065_),
    .Z(_096_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _216_ (.A1(_120_),
    .A2(_095_),
    .A3(_072_),
    .B(_096_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _217_ (.A1(_120_),
    .A2(_095_),
    .A3(_069_),
    .A4(_072_),
    .Z(_098_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _218_ (.A1(_094_),
    .A2(_097_),
    .A3(_098_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _219_ (.A1(\state[1] ),
    .A2(_083_),
    .A3(_091_),
    .Z(_099_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _220_ (.A1(_081_),
    .A2(_099_),
    .B(_085_),
    .C(\debug_miso_samples[7] ),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _221_ (.A1(_082_),
    .A2(_091_),
    .B(_100_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _222_ (.A1(\state[1] ),
    .A2(_041_),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _223_ (.I0(\debug_miso_samples[0] ),
    .I1(net13),
    .S(_101_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _224_ (.I0(\debug_miso_samples[1] ),
    .I1(net14),
    .S(_101_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _225_ (.I0(\debug_miso_samples[2] ),
    .I1(net15),
    .S(_101_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _226_ (.I0(\debug_miso_samples[3] ),
    .I1(net16),
    .S(_101_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _227_ (.I0(\debug_miso_samples[4] ),
    .I1(net17),
    .S(_101_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _228_ (.I0(\debug_miso_samples[5] ),
    .I1(net18),
    .S(_101_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _229_ (.I0(\debug_miso_samples[6] ),
    .I1(net19),
    .S(_101_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _230_ (.I0(\debug_miso_samples[7] ),
    .I1(net20),
    .S(_101_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _231_ (.I0(\state[1] ),
    .I1(net21),
    .S(\state[0] ),
    .Z(_020_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _232_ (.A1(\state[1] ),
    .A2(net22),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _233_ (.A1(\state[0] ),
    .A2(_102_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _234_ (.A1(_034_),
    .A2(net12),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _235_ (.I0(net23),
    .I1(_103_),
    .S(_041_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _236_ (.A1(_034_),
    .A2(\state[0] ),
    .Z(_104_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _237_ (.I0(net11),
    .I1(\tx_shift[6] ),
    .S(_104_),
    .Z(_105_));
 gf180mcu_fd_sc_mcu9t5v0__aoi22_2 _238_ (.A1(_041_),
    .A2(net12),
    .B1(_119_),
    .B2(_066_),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_4 _239_ (.A1(\state[1] ),
    .A2(_106_),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _240_ (.I0(net24),
    .I1(_105_),
    .S(_107_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _241_ (.A1(\state[0] ),
    .A2(_035_),
    .A3(_123_),
    .Z(_108_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _242_ (.A1(_039_),
    .A2(_108_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _243_ (.A1(_123_),
    .A2(_065_),
    .Z(_025_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _244_ (.I0(_048_),
    .I1(net25),
    .S(_085_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _245_ (.I(\tx_shift[0] ),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _246_ (.A1(net12),
    .A2(net4),
    .ZN(_110_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _247_ (.A1(_109_),
    .A2(_107_),
    .B1(_110_),
    .B2(_085_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _248_ (.I0(net5),
    .I1(\tx_shift[0] ),
    .S(_104_),
    .Z(_111_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _249_ (.I0(\tx_shift[1] ),
    .I1(_111_),
    .S(_107_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _250_ (.I0(net6),
    .I1(\tx_shift[1] ),
    .S(_104_),
    .Z(_112_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _251_ (.I0(\tx_shift[2] ),
    .I1(_112_),
    .S(_107_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _252_ (.I0(net7),
    .I1(\tx_shift[2] ),
    .S(_104_),
    .Z(_113_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _253_ (.I0(\tx_shift[3] ),
    .I1(_113_),
    .S(_107_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _254_ (.I0(net8),
    .I1(\tx_shift[3] ),
    .S(_104_),
    .Z(_114_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _255_ (.I0(\tx_shift[4] ),
    .I1(_114_),
    .S(_107_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _256_ (.I0(net9),
    .I1(\tx_shift[4] ),
    .S(_104_),
    .Z(_115_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _257_ (.I0(\tx_shift[5] ),
    .I1(_115_),
    .S(_107_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _258_ (.I0(net10),
    .I1(\tx_shift[5] ),
    .S(_104_),
    .Z(_116_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _259_ (.I0(\tx_shift[6] ),
    .I1(_116_),
    .S(_107_),
    .Z(_033_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _260_ (.A(_117_),
    .B(_118_),
    .CO(_119_),
    .S(_120_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _261_ (.A(\bit_count[3] ),
    .B(_118_),
    .CO(_121_),
    .S(_122_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _262_ (.A(\bit_count[3] ),
    .B(_123_),
    .CO(_124_),
    .S(_125_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _263_ (.A(_117_),
    .B(_126_),
    .CO(_127_),
    .S(_128_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _264_ (.A(_117_),
    .B(_129_),
    .CO(_130_),
    .S(_131_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _265_ (.A(\bit_count[0] ),
    .B(\bit_count[1] ),
    .CO(_132_),
    .S(_133_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _266_ (.A(_117_),
    .B(_134_),
    .CO(_135_),
    .S(_136_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_count[0]$_DFFE_PN0P_  (.D(_000_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\bit_count[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_count[1]$_DFFE_PN0P_  (.D(_001_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\bit_count[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_count[2]$_DFFE_PN0P_  (.D(_002_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\bit_count[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_count[3]$_DFFE_PN0P_  (.D(_003_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\bit_count[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \debug_miso_samples[0]$_DFFE_PN0P_  (.D(_004_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\debug_miso_samples[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \debug_miso_samples[1]$_DFFE_PN0P_  (.D(_005_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\debug_miso_samples[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \debug_miso_samples[2]$_DFFE_PN0P_  (.D(_006_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\debug_miso_samples[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \debug_miso_samples[3]$_DFFE_PN0P_  (.D(_007_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\debug_miso_samples[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \debug_miso_samples[4]$_DFFE_PN0P_  (.D(_008_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\debug_miso_samples[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \debug_miso_samples[5]$_DFFE_PN0P_  (.D(_009_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\debug_miso_samples[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \debug_miso_samples[6]$_DFFE_PN0P_  (.D(_010_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\debug_miso_samples[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \debug_miso_samples[7]$_DFFE_PN0P_  (.D(_011_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\debug_miso_samples[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[0]$_DFFE_PN0P_  (.D(_012_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net13));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[1]$_DFFE_PN0P_  (.D(_013_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net14));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[2]$_DFFE_PN0P_  (.D(_014_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net15));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[3]$_DFFE_PN0P_  (.D(_015_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net16));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[4]$_DFFE_PN0P_  (.D(_016_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net17));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[5]$_DFFE_PN0P_  (.D(_017_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[6]$_DFFE_PN0P_  (.D(_018_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[7]$_DFFE_PN0P_  (.D(_019_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_valid$_DFFE_PN0P_  (.D(_020_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \spi_clk$_DFFE_PN0P_  (.D(_021_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \spi_cs_n$_DFFE_PN1P_  (.D(_022_),
    .SETN(net2),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \spi_mosi$_DFFE_PN0P_  (.D(_023_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \state[0]$_DFFE_PN0P_  (.D(_024_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\state[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \state[1]$_DFFE_PN0P_  (.D(_025_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\state[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \tx_ready$_DFFE_PN1P_  (.D(_026_),
    .SETN(net2),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[0]$_DFFE_PN0P_  (.D(_027_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\tx_shift[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[1]$_DFFE_PN0P_  (.D(_028_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\tx_shift[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[2]$_DFFE_PN0P_  (.D(_029_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[3]$_DFFE_PN0P_  (.D(_030_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[4]$_DFFE_PN0P_  (.D(_031_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[5]$_DFFE_PN0P_  (.D(_032_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift[6]$_DFFE_PN0P_  (.D(_033_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift[6] ));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 hold1 (.I(net2),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_52 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_26_Left_53 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_54 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_55 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_56 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_57 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_58 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_59 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_60 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_61 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_62 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_63 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_64 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_65 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_66 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_26_67 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input1 (.I(net26),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input2 (.I(spi_miso),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(tx_data[0]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(tx_data[1]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(tx_data[2]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(tx_data[3]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(tx_data[4]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(tx_data[5]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(tx_data[6]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(tx_data[7]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__buf_3 input11 (.I(tx_valid),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output12 (.I(net13),
    .Z(rx_data[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output13 (.I(net14),
    .Z(rx_data[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output14 (.I(net15),
    .Z(rx_data[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output15 (.I(net16),
    .Z(rx_data[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output16 (.I(net17),
    .Z(rx_data[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output17 (.I(net18),
    .Z(rx_data[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output18 (.I(net19),
    .Z(rx_data[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output19 (.I(net20),
    .Z(rx_data[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output20 (.I(net21),
    .Z(rx_valid));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output21 (.I(net22),
    .Z(spi_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output22 (.I(net23),
    .Z(spi_cs_n));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output23 (.I(net24),
    .Z(spi_mosi));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output24 (.I(net25),
    .Z(tx_ready));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__inv_4 clkload0 (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload1 (.I(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 clkload2 (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_138 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_133 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_183 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_2_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_3_242 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_3_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_234 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_156 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_190 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_5_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_119 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_167 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_162 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_159 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_9_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_9_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_245 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_49 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_11_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_205 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_52 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_38 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_72 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_76 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_115 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_158 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_137 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_194 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_202 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_61 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_65 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_210 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_230 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_16_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_214 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_32 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_48 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_17_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_191 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_231 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_6 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_24 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_91 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_160 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_53 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_77 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_217 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_10 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_14 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_16 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_248 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_40 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_56 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_79 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_81 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_185 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_201 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_247 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_251 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_153 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_215 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_246 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_23_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_23_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_249 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_252 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_112 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_145 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_181 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_54 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_26_207 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_26_209 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_26_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_26_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_26_249 ();
endmodule
