module axi_stream_interface (clk,
    m_tdest,
    m_tid,
    m_tlast,
    m_tready,
    m_tuser,
    m_tvalid,
    rst_n,
    s_tdest,
    s_tid,
    s_tlast,
    s_tready,
    s_tuser,
    s_tvalid,
    m_tdata,
    m_tkeep,
    m_tstrb,
    s_tdata,
    s_tkeep,
    s_tstrb);
 input clk;
 output m_tdest;
 output m_tid;
 output m_tlast;
 input m_tready;
 output m_tuser;
 output m_tvalid;
 input rst_n;
 input s_tdest;
 input s_tid;
 input s_tlast;
 output s_tready;
 input s_tuser;
 input s_tvalid;
 output [31:0] m_tdata;
 output [3:0] m_tkeep;
 output [3:0] m_tstrb;
 input [31:0] s_tdata;
 input [3:0] s_tkeep;
 input [3:0] s_tstrb;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;

 sky130_fd_sc_hd__clkbuf_1 _00_ (.A(s_tdata[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 _01_ (.A(s_tdata[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 _02_ (.A(s_tdata[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 _03_ (.A(s_tdata[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 _04_ (.A(s_tdata[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 _05_ (.A(s_tdata[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 _06_ (.A(s_tdata[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 _07_ (.A(s_tdata[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 _08_ (.A(s_tdata[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 _09_ (.A(s_tdata[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 _10_ (.A(s_tdata[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 _11_ (.A(s_tdata[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 _12_ (.A(s_tdata[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 _13_ (.A(s_tdata[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 _14_ (.A(s_tdata[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 _15_ (.A(s_tdata[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 _16_ (.A(s_tdata[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 _17_ (.A(s_tdata[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 _18_ (.A(s_tdata[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 _19_ (.A(s_tdata[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 _20_ (.A(s_tdata[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 _21_ (.A(s_tdata[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 _22_ (.A(s_tdata[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 _23_ (.A(s_tdata[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 _24_ (.A(s_tdata[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 _25_ (.A(s_tdata[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 _26_ (.A(s_tdata[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 _27_ (.A(s_tdata[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 _28_ (.A(s_tdata[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 _29_ (.A(s_tdata[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 _30_ (.A(s_tdata[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 _31_ (.A(s_tdata[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 _32_ (.A(s_tdest),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 _33_ (.A(s_tid),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 _34_ (.A(s_tkeep[0]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 _35_ (.A(s_tkeep[1]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 _36_ (.A(s_tkeep[2]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 _37_ (.A(s_tkeep[3]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 _38_ (.A(s_tlast),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 _39_ (.A(s_tstrb[0]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 _40_ (.A(s_tstrb[1]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 _41_ (.A(s_tstrb[2]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 _42_ (.A(s_tstrb[3]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 _43_ (.A(s_tuser),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 _44_ (.A(s_tvalid),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 _45_ (.A(m_tready),
    .X(net46));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_15 ();
 sky130_fd_sc_hd__clkbuf_1 output1 (.A(net1),
    .X(m_tdata[0]));
 sky130_fd_sc_hd__clkbuf_1 output2 (.A(net2),
    .X(m_tdata[10]));
 sky130_fd_sc_hd__clkbuf_1 output3 (.A(net3),
    .X(m_tdata[11]));
 sky130_fd_sc_hd__clkbuf_1 output4 (.A(net4),
    .X(m_tdata[12]));
 sky130_fd_sc_hd__clkbuf_1 output5 (.A(net5),
    .X(m_tdata[13]));
 sky130_fd_sc_hd__clkbuf_1 output6 (.A(net6),
    .X(m_tdata[14]));
 sky130_fd_sc_hd__clkbuf_1 output7 (.A(net7),
    .X(m_tdata[15]));
 sky130_fd_sc_hd__clkbuf_1 output8 (.A(net8),
    .X(m_tdata[16]));
 sky130_fd_sc_hd__clkbuf_1 output9 (.A(net9),
    .X(m_tdata[17]));
 sky130_fd_sc_hd__clkbuf_1 output10 (.A(net10),
    .X(m_tdata[18]));
 sky130_fd_sc_hd__clkbuf_1 output11 (.A(net11),
    .X(m_tdata[19]));
 sky130_fd_sc_hd__clkbuf_1 output12 (.A(net12),
    .X(m_tdata[1]));
 sky130_fd_sc_hd__clkbuf_1 output13 (.A(net13),
    .X(m_tdata[20]));
 sky130_fd_sc_hd__clkbuf_1 output14 (.A(net14),
    .X(m_tdata[21]));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net15),
    .X(m_tdata[22]));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net16),
    .X(m_tdata[23]));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net17),
    .X(m_tdata[24]));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net18),
    .X(m_tdata[25]));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net19),
    .X(m_tdata[26]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net20),
    .X(m_tdata[27]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net21),
    .X(m_tdata[28]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net22),
    .X(m_tdata[29]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net23),
    .X(m_tdata[2]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net24),
    .X(m_tdata[30]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net25),
    .X(m_tdata[31]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net26),
    .X(m_tdata[3]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net27),
    .X(m_tdata[4]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net28),
    .X(m_tdata[5]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net29),
    .X(m_tdata[6]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net30),
    .X(m_tdata[7]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net31),
    .X(m_tdata[8]));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(net32),
    .X(m_tdata[9]));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net33),
    .X(m_tdest));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net34),
    .X(m_tid));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(net35),
    .X(m_tkeep[0]));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net36),
    .X(m_tkeep[1]));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(net37),
    .X(m_tkeep[2]));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net38),
    .X(m_tkeep[3]));
 sky130_fd_sc_hd__clkbuf_1 output39 (.A(net39),
    .X(m_tlast));
 sky130_fd_sc_hd__clkbuf_1 output40 (.A(net40),
    .X(m_tstrb[0]));
 sky130_fd_sc_hd__clkbuf_1 output41 (.A(net41),
    .X(m_tstrb[1]));
 sky130_fd_sc_hd__clkbuf_1 output42 (.A(net42),
    .X(m_tstrb[2]));
 sky130_fd_sc_hd__clkbuf_1 output43 (.A(net43),
    .X(m_tstrb[3]));
 sky130_fd_sc_hd__clkbuf_1 output44 (.A(net44),
    .X(m_tuser));
 sky130_fd_sc_hd__clkbuf_1 output45 (.A(net45),
    .X(m_tvalid));
 sky130_fd_sc_hd__clkbuf_1 output46 (.A(net46),
    .X(s_tready));
 sky130_fd_sc_hd__fill_1 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_85 ();
endmodule
