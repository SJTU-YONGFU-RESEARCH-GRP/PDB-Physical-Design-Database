module onehot_decoder_register (clk,
    enable,
    rst_n,
    binary_in,
    onehot_out);
 input clk;
 input enable;
 input rst_n;
 input [3:0] binary_in;
 output [15:0] onehot_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 INV_X1 _063_ (.A(net6),
    .ZN(_016_));
 INV_X2 _064_ (.A(net5),
    .ZN(_017_));
 BUF_X4 _065_ (.A(rst_n),
    .Z(_018_));
 NAND2_X2 _066_ (.A1(_017_),
    .A2(_018_),
    .ZN(_019_));
 BUF_X4 _067_ (.A(_019_),
    .Z(_020_));
 INV_X1 _068_ (.A(net1),
    .ZN(_021_));
 INV_X1 _069_ (.A(net2),
    .ZN(_022_));
 NAND3_X2 _070_ (.A1(_021_),
    .A2(_022_),
    .A3(_018_),
    .ZN(_023_));
 OR3_X2 _071_ (.A1(net4),
    .A2(net3),
    .A3(_017_),
    .ZN(_024_));
 OAI22_X1 _072_ (.A1(_016_),
    .A2(_020_),
    .B1(_023_),
    .B2(_024_),
    .ZN(_000_));
 NAND3_X1 _073_ (.A1(_017_),
    .A2(net7),
    .A3(_018_),
    .ZN(_025_));
 NAND3_X2 _074_ (.A1(_021_),
    .A2(net2),
    .A3(_018_),
    .ZN(_026_));
 INV_X1 _075_ (.A(net3),
    .ZN(_027_));
 NAND3_X2 _076_ (.A1(net4),
    .A2(_027_),
    .A3(net5),
    .ZN(_028_));
 OAI21_X1 _077_ (.A(_025_),
    .B1(_026_),
    .B2(_028_),
    .ZN(_001_));
 INV_X1 _078_ (.A(net8),
    .ZN(_029_));
 NAND3_X2 _079_ (.A1(net1),
    .A2(net2),
    .A3(_018_),
    .ZN(_030_));
 OAI22_X1 _080_ (.A1(_029_),
    .A2(_020_),
    .B1(_028_),
    .B2(_030_),
    .ZN(_002_));
 INV_X1 _081_ (.A(net9),
    .ZN(_031_));
 NAND3_X2 _082_ (.A1(net4),
    .A2(net3),
    .A3(net5),
    .ZN(_032_));
 OAI22_X1 _083_ (.A1(_031_),
    .A2(_020_),
    .B1(_023_),
    .B2(_032_),
    .ZN(_003_));
 INV_X1 _084_ (.A(net10),
    .ZN(_033_));
 NAND3_X2 _085_ (.A1(net1),
    .A2(_022_),
    .A3(_018_),
    .ZN(_034_));
 OAI22_X1 _086_ (.A1(_033_),
    .A2(_020_),
    .B1(_032_),
    .B2(_034_),
    .ZN(_004_));
 INV_X1 _087_ (.A(net11),
    .ZN(_035_));
 OAI22_X1 _088_ (.A1(_035_),
    .A2(_020_),
    .B1(_026_),
    .B2(_032_),
    .ZN(_005_));
 INV_X1 _089_ (.A(net12),
    .ZN(_036_));
 OAI22_X1 _090_ (.A1(_036_),
    .A2(_020_),
    .B1(_030_),
    .B2(_032_),
    .ZN(_006_));
 INV_X1 _091_ (.A(net13),
    .ZN(_037_));
 OAI22_X1 _092_ (.A1(_037_),
    .A2(_020_),
    .B1(_024_),
    .B2(_034_),
    .ZN(_007_));
 NAND3_X1 _093_ (.A1(_017_),
    .A2(net14),
    .A3(_018_),
    .ZN(_038_));
 OAI21_X1 _094_ (.A(_038_),
    .B1(_026_),
    .B2(_024_),
    .ZN(_008_));
 INV_X1 _095_ (.A(net15),
    .ZN(_039_));
 OAI22_X1 _096_ (.A1(_039_),
    .A2(_020_),
    .B1(_024_),
    .B2(_030_),
    .ZN(_009_));
 INV_X1 _097_ (.A(net16),
    .ZN(_040_));
 OR3_X2 _098_ (.A1(net4),
    .A2(_027_),
    .A3(_017_),
    .ZN(_041_));
 OAI22_X1 _099_ (.A1(_040_),
    .A2(_020_),
    .B1(_023_),
    .B2(_041_),
    .ZN(_010_));
 INV_X1 _100_ (.A(net17),
    .ZN(_042_));
 OAI22_X1 _101_ (.A1(_042_),
    .A2(_020_),
    .B1(_034_),
    .B2(_041_),
    .ZN(_011_));
 INV_X1 _102_ (.A(net18),
    .ZN(_043_));
 OAI22_X1 _103_ (.A1(_043_),
    .A2(_019_),
    .B1(_026_),
    .B2(_041_),
    .ZN(_012_));
 INV_X1 _104_ (.A(net19),
    .ZN(_044_));
 OAI22_X1 _105_ (.A1(_044_),
    .A2(_019_),
    .B1(_030_),
    .B2(_041_),
    .ZN(_013_));
 NAND3_X1 _106_ (.A1(_017_),
    .A2(net20),
    .A3(_018_),
    .ZN(_045_));
 OAI21_X1 _107_ (.A(_045_),
    .B1(_028_),
    .B2(_023_),
    .ZN(_014_));
 INV_X1 _108_ (.A(net21),
    .ZN(_046_));
 OAI22_X1 _109_ (.A1(_046_),
    .A2(_019_),
    .B1(_028_),
    .B2(_034_),
    .ZN(_015_));
 DFF_X1 \onehot_out[0]$_SDFFE_PN0P_  (.D(_000_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net6),
    .QN(_062_));
 DFF_X1 \onehot_out[10]$_SDFFE_PN0P_  (.D(_001_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net7),
    .QN(_061_));
 DFF_X1 \onehot_out[11]$_SDFFE_PN0P_  (.D(_002_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net8),
    .QN(_060_));
 DFF_X1 \onehot_out[12]$_SDFFE_PN0P_  (.D(_003_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net9),
    .QN(_059_));
 DFF_X1 \onehot_out[13]$_SDFFE_PN0P_  (.D(_004_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net10),
    .QN(_058_));
 DFF_X1 \onehot_out[14]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net11),
    .QN(_057_));
 DFF_X1 \onehot_out[15]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net12),
    .QN(_056_));
 DFF_X1 \onehot_out[1]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net13),
    .QN(_055_));
 DFF_X1 \onehot_out[2]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net14),
    .QN(_054_));
 DFF_X1 \onehot_out[3]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net15),
    .QN(_053_));
 DFF_X1 \onehot_out[4]$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net16),
    .QN(_052_));
 DFF_X1 \onehot_out[5]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net17),
    .QN(_051_));
 DFF_X1 \onehot_out[6]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net18),
    .QN(_050_));
 DFF_X1 \onehot_out[7]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net19),
    .QN(_049_));
 DFF_X1 \onehot_out[8]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net20),
    .QN(_048_));
 DFF_X1 \onehot_out[9]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net21),
    .QN(_047_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_71 ();
 BUF_X1 input1 (.A(binary_in[0]),
    .Z(net1));
 CLKBUF_X2 input2 (.A(binary_in[1]),
    .Z(net2));
 BUF_X1 input3 (.A(binary_in[2]),
    .Z(net3));
 CLKBUF_X2 input4 (.A(binary_in[3]),
    .Z(net4));
 BUF_X2 input5 (.A(enable),
    .Z(net5));
 BUF_X1 output6 (.A(net6),
    .Z(onehot_out[0]));
 BUF_X1 output7 (.A(net7),
    .Z(onehot_out[10]));
 BUF_X1 output8 (.A(net8),
    .Z(onehot_out[11]));
 BUF_X1 output9 (.A(net9),
    .Z(onehot_out[12]));
 BUF_X1 output10 (.A(net10),
    .Z(onehot_out[13]));
 BUF_X1 output11 (.A(net11),
    .Z(onehot_out[14]));
 BUF_X1 output12 (.A(net12),
    .Z(onehot_out[15]));
 BUF_X1 output13 (.A(net13),
    .Z(onehot_out[1]));
 BUF_X1 output14 (.A(net14),
    .Z(onehot_out[2]));
 BUF_X1 output15 (.A(net15),
    .Z(onehot_out[3]));
 BUF_X1 output16 (.A(net16),
    .Z(onehot_out[4]));
 BUF_X1 output17 (.A(net17),
    .Z(onehot_out[5]));
 BUF_X1 output18 (.A(net18),
    .Z(onehot_out[6]));
 BUF_X1 output19 (.A(net19),
    .Z(onehot_out[7]));
 BUF_X1 output20 (.A(net20),
    .Z(onehot_out[8]));
 BUF_X1 output21 (.A(net21),
    .Z(onehot_out[9]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X16 FILLER_0_97 ();
 FILLCELL_X2 FILLER_0_113 ();
 FILLCELL_X8 FILLER_0_118 ();
 FILLCELL_X4 FILLER_0_126 ();
 FILLCELL_X2 FILLER_0_137 ();
 FILLCELL_X4 FILLER_0_146 ();
 FILLCELL_X1 FILLER_0_150 ();
 FILLCELL_X32 FILLER_0_154 ();
 FILLCELL_X32 FILLER_0_186 ();
 FILLCELL_X32 FILLER_0_218 ();
 FILLCELL_X16 FILLER_0_250 ();
 FILLCELL_X2 FILLER_0_266 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X16 FILLER_1_97 ();
 FILLCELL_X1 FILLER_1_113 ();
 FILLCELL_X32 FILLER_1_117 ();
 FILLCELL_X8 FILLER_1_149 ();
 FILLCELL_X4 FILLER_1_157 ();
 FILLCELL_X2 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_166 ();
 FILLCELL_X32 FILLER_1_198 ();
 FILLCELL_X32 FILLER_1_230 ();
 FILLCELL_X4 FILLER_1_262 ();
 FILLCELL_X2 FILLER_1_266 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X8 FILLER_2_257 ();
 FILLCELL_X2 FILLER_2_265 ();
 FILLCELL_X1 FILLER_2_267 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X8 FILLER_3_257 ();
 FILLCELL_X2 FILLER_3_265 ();
 FILLCELL_X1 FILLER_3_267 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X8 FILLER_4_257 ();
 FILLCELL_X2 FILLER_4_265 ();
 FILLCELL_X1 FILLER_4_267 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X8 FILLER_5_257 ();
 FILLCELL_X2 FILLER_5_265 ();
 FILLCELL_X1 FILLER_5_267 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X32 FILLER_6_225 ();
 FILLCELL_X8 FILLER_6_257 ();
 FILLCELL_X2 FILLER_6_265 ();
 FILLCELL_X1 FILLER_6_267 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X32 FILLER_7_193 ();
 FILLCELL_X32 FILLER_7_225 ();
 FILLCELL_X8 FILLER_7_257 ();
 FILLCELL_X2 FILLER_7_265 ();
 FILLCELL_X1 FILLER_7_267 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X32 FILLER_8_193 ();
 FILLCELL_X32 FILLER_8_225 ();
 FILLCELL_X8 FILLER_8_257 ();
 FILLCELL_X2 FILLER_8_265 ();
 FILLCELL_X1 FILLER_8_267 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X32 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_225 ();
 FILLCELL_X8 FILLER_9_257 ();
 FILLCELL_X2 FILLER_9_265 ();
 FILLCELL_X1 FILLER_9_267 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X4 FILLER_10_97 ();
 FILLCELL_X2 FILLER_10_101 ();
 FILLCELL_X1 FILLER_10_103 ();
 FILLCELL_X4 FILLER_10_123 ();
 FILLCELL_X2 FILLER_10_127 ();
 FILLCELL_X2 FILLER_10_146 ();
 FILLCELL_X32 FILLER_10_167 ();
 FILLCELL_X32 FILLER_10_199 ();
 FILLCELL_X32 FILLER_10_231 ();
 FILLCELL_X4 FILLER_10_263 ();
 FILLCELL_X1 FILLER_10_267 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X16 FILLER_11_97 ();
 FILLCELL_X2 FILLER_11_113 ();
 FILLCELL_X1 FILLER_11_115 ();
 FILLCELL_X8 FILLER_11_121 ();
 FILLCELL_X2 FILLER_11_129 ();
 FILLCELL_X8 FILLER_11_138 ();
 FILLCELL_X4 FILLER_11_146 ();
 FILLCELL_X2 FILLER_11_150 ();
 FILLCELL_X1 FILLER_11_152 ();
 FILLCELL_X32 FILLER_11_177 ();
 FILLCELL_X16 FILLER_11_209 ();
 FILLCELL_X4 FILLER_11_225 ();
 FILLCELL_X32 FILLER_11_232 ();
 FILLCELL_X4 FILLER_11_264 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X16 FILLER_12_116 ();
 FILLCELL_X4 FILLER_12_132 ();
 FILLCELL_X2 FILLER_12_136 ();
 FILLCELL_X16 FILLER_12_143 ();
 FILLCELL_X2 FILLER_12_159 ();
 FILLCELL_X32 FILLER_12_166 ();
 FILLCELL_X32 FILLER_12_198 ();
 FILLCELL_X32 FILLER_12_230 ();
 FILLCELL_X4 FILLER_12_262 ();
 FILLCELL_X2 FILLER_12_266 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X16 FILLER_13_97 ();
 FILLCELL_X8 FILLER_13_118 ();
 FILLCELL_X4 FILLER_13_126 ();
 FILLCELL_X2 FILLER_13_130 ();
 FILLCELL_X1 FILLER_13_132 ();
 FILLCELL_X32 FILLER_13_157 ();
 FILLCELL_X32 FILLER_13_189 ();
 FILLCELL_X32 FILLER_13_221 ();
 FILLCELL_X8 FILLER_13_253 ();
 FILLCELL_X4 FILLER_13_261 ();
 FILLCELL_X2 FILLER_13_265 ();
 FILLCELL_X1 FILLER_13_267 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X8 FILLER_14_129 ();
 FILLCELL_X4 FILLER_14_137 ();
 FILLCELL_X2 FILLER_14_141 ();
 FILLCELL_X4 FILLER_14_148 ();
 FILLCELL_X32 FILLER_14_154 ();
 FILLCELL_X32 FILLER_14_186 ();
 FILLCELL_X32 FILLER_14_218 ();
 FILLCELL_X16 FILLER_14_250 ();
 FILLCELL_X2 FILLER_14_266 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X16 FILLER_15_129 ();
 FILLCELL_X8 FILLER_15_145 ();
 FILLCELL_X4 FILLER_15_153 ();
 FILLCELL_X2 FILLER_15_157 ();
 FILLCELL_X1 FILLER_15_159 ();
 FILLCELL_X32 FILLER_15_184 ();
 FILLCELL_X16 FILLER_15_216 ();
 FILLCELL_X1 FILLER_15_232 ();
 FILLCELL_X32 FILLER_15_236 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X8 FILLER_16_97 ();
 FILLCELL_X4 FILLER_16_105 ();
 FILLCELL_X2 FILLER_16_109 ();
 FILLCELL_X1 FILLER_16_111 ();
 FILLCELL_X8 FILLER_16_116 ();
 FILLCELL_X4 FILLER_16_124 ();
 FILLCELL_X1 FILLER_16_128 ();
 FILLCELL_X32 FILLER_16_140 ();
 FILLCELL_X32 FILLER_16_172 ();
 FILLCELL_X32 FILLER_16_204 ();
 FILLCELL_X32 FILLER_16_236 ();
 FILLCELL_X16 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_20 ();
 FILLCELL_X32 FILLER_17_52 ();
 FILLCELL_X8 FILLER_17_84 ();
 FILLCELL_X2 FILLER_17_92 ();
 FILLCELL_X1 FILLER_17_94 ();
 FILLCELL_X8 FILLER_17_116 ();
 FILLCELL_X4 FILLER_17_124 ();
 FILLCELL_X2 FILLER_17_128 ();
 FILLCELL_X1 FILLER_17_130 ();
 FILLCELL_X32 FILLER_17_144 ();
 FILLCELL_X32 FILLER_17_176 ();
 FILLCELL_X32 FILLER_17_208 ();
 FILLCELL_X16 FILLER_17_240 ();
 FILLCELL_X8 FILLER_17_256 ();
 FILLCELL_X4 FILLER_17_264 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X8 FILLER_18_129 ();
 FILLCELL_X2 FILLER_18_137 ();
 FILLCELL_X8 FILLER_18_144 ();
 FILLCELL_X4 FILLER_18_152 ();
 FILLCELL_X2 FILLER_18_156 ();
 FILLCELL_X1 FILLER_18_158 ();
 FILLCELL_X32 FILLER_18_183 ();
 FILLCELL_X8 FILLER_18_215 ();
 FILLCELL_X4 FILLER_18_223 ();
 FILLCELL_X2 FILLER_18_227 ();
 FILLCELL_X1 FILLER_18_229 ();
 FILLCELL_X32 FILLER_18_233 ();
 FILLCELL_X2 FILLER_18_265 ();
 FILLCELL_X1 FILLER_18_267 ();
 FILLCELL_X4 FILLER_19_1 ();
 FILLCELL_X2 FILLER_19_5 ();
 FILLCELL_X32 FILLER_19_10 ();
 FILLCELL_X32 FILLER_19_42 ();
 FILLCELL_X16 FILLER_19_74 ();
 FILLCELL_X4 FILLER_19_90 ();
 FILLCELL_X8 FILLER_19_119 ();
 FILLCELL_X4 FILLER_19_127 ();
 FILLCELL_X32 FILLER_19_138 ();
 FILLCELL_X32 FILLER_19_170 ();
 FILLCELL_X32 FILLER_19_202 ();
 FILLCELL_X32 FILLER_19_234 ();
 FILLCELL_X2 FILLER_19_266 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X8 FILLER_20_65 ();
 FILLCELL_X4 FILLER_20_73 ();
 FILLCELL_X2 FILLER_20_77 ();
 FILLCELL_X1 FILLER_20_79 ();
 FILLCELL_X16 FILLER_20_87 ();
 FILLCELL_X4 FILLER_20_103 ();
 FILLCELL_X2 FILLER_20_107 ();
 FILLCELL_X1 FILLER_20_109 ();
 FILLCELL_X8 FILLER_20_114 ();
 FILLCELL_X4 FILLER_20_133 ();
 FILLCELL_X32 FILLER_20_142 ();
 FILLCELL_X32 FILLER_20_174 ();
 FILLCELL_X32 FILLER_20_206 ();
 FILLCELL_X16 FILLER_20_238 ();
 FILLCELL_X8 FILLER_20_254 ();
 FILLCELL_X4 FILLER_20_262 ();
 FILLCELL_X2 FILLER_20_266 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X16 FILLER_21_65 ();
 FILLCELL_X8 FILLER_21_81 ();
 FILLCELL_X4 FILLER_21_89 ();
 FILLCELL_X2 FILLER_21_93 ();
 FILLCELL_X8 FILLER_21_116 ();
 FILLCELL_X4 FILLER_21_124 ();
 FILLCELL_X16 FILLER_21_142 ();
 FILLCELL_X4 FILLER_21_158 ();
 FILLCELL_X32 FILLER_21_186 ();
 FILLCELL_X32 FILLER_21_218 ();
 FILLCELL_X4 FILLER_21_250 ();
 FILLCELL_X1 FILLER_21_254 ();
 FILLCELL_X8 FILLER_21_258 ();
 FILLCELL_X2 FILLER_21_266 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X4 FILLER_22_129 ();
 FILLCELL_X2 FILLER_22_133 ();
 FILLCELL_X1 FILLER_22_135 ();
 FILLCELL_X32 FILLER_22_143 ();
 FILLCELL_X32 FILLER_22_175 ();
 FILLCELL_X32 FILLER_22_207 ();
 FILLCELL_X16 FILLER_22_239 ();
 FILLCELL_X8 FILLER_22_255 ();
 FILLCELL_X4 FILLER_22_263 ();
 FILLCELL_X1 FILLER_22_267 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X16 FILLER_23_97 ();
 FILLCELL_X4 FILLER_23_113 ();
 FILLCELL_X2 FILLER_23_117 ();
 FILLCELL_X4 FILLER_23_124 ();
 FILLCELL_X2 FILLER_23_128 ();
 FILLCELL_X1 FILLER_23_130 ();
 FILLCELL_X4 FILLER_23_136 ();
 FILLCELL_X1 FILLER_23_150 ();
 FILLCELL_X4 FILLER_23_158 ();
 FILLCELL_X2 FILLER_23_162 ();
 FILLCELL_X1 FILLER_23_164 ();
 FILLCELL_X32 FILLER_23_167 ();
 FILLCELL_X32 FILLER_23_199 ();
 FILLCELL_X32 FILLER_23_231 ();
 FILLCELL_X4 FILLER_23_263 ();
 FILLCELL_X1 FILLER_23_267 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X4 FILLER_24_97 ();
 FILLCELL_X2 FILLER_24_101 ();
 FILLCELL_X8 FILLER_24_122 ();
 FILLCELL_X2 FILLER_24_130 ();
 FILLCELL_X1 FILLER_24_132 ();
 FILLCELL_X8 FILLER_24_135 ();
 FILLCELL_X1 FILLER_24_160 ();
 FILLCELL_X32 FILLER_24_178 ();
 FILLCELL_X32 FILLER_24_210 ();
 FILLCELL_X16 FILLER_24_242 ();
 FILLCELL_X8 FILLER_24_258 ();
 FILLCELL_X2 FILLER_24_266 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X16 FILLER_25_97 ();
 FILLCELL_X8 FILLER_25_113 ();
 FILLCELL_X2 FILLER_25_121 ();
 FILLCELL_X32 FILLER_25_140 ();
 FILLCELL_X32 FILLER_25_172 ();
 FILLCELL_X32 FILLER_25_204 ();
 FILLCELL_X32 FILLER_25_236 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X32 FILLER_26_97 ();
 FILLCELL_X32 FILLER_26_129 ();
 FILLCELL_X32 FILLER_26_161 ();
 FILLCELL_X32 FILLER_26_193 ();
 FILLCELL_X32 FILLER_26_225 ();
 FILLCELL_X8 FILLER_26_257 ();
 FILLCELL_X2 FILLER_26_265 ();
 FILLCELL_X1 FILLER_26_267 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X32 FILLER_27_129 ();
 FILLCELL_X32 FILLER_27_161 ();
 FILLCELL_X32 FILLER_27_193 ();
 FILLCELL_X32 FILLER_27_225 ();
 FILLCELL_X8 FILLER_27_257 ();
 FILLCELL_X2 FILLER_27_265 ();
 FILLCELL_X1 FILLER_27_267 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X32 FILLER_28_129 ();
 FILLCELL_X32 FILLER_28_161 ();
 FILLCELL_X32 FILLER_28_193 ();
 FILLCELL_X32 FILLER_28_225 ();
 FILLCELL_X8 FILLER_28_257 ();
 FILLCELL_X2 FILLER_28_265 ();
 FILLCELL_X1 FILLER_28_267 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X32 FILLER_29_129 ();
 FILLCELL_X32 FILLER_29_161 ();
 FILLCELL_X32 FILLER_29_193 ();
 FILLCELL_X32 FILLER_29_225 ();
 FILLCELL_X8 FILLER_29_257 ();
 FILLCELL_X2 FILLER_29_265 ();
 FILLCELL_X1 FILLER_29_267 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X32 FILLER_30_129 ();
 FILLCELL_X32 FILLER_30_161 ();
 FILLCELL_X32 FILLER_30_193 ();
 FILLCELL_X32 FILLER_30_225 ();
 FILLCELL_X8 FILLER_30_257 ();
 FILLCELL_X2 FILLER_30_265 ();
 FILLCELL_X1 FILLER_30_267 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X32 FILLER_31_129 ();
 FILLCELL_X32 FILLER_31_161 ();
 FILLCELL_X32 FILLER_31_193 ();
 FILLCELL_X32 FILLER_31_225 ();
 FILLCELL_X8 FILLER_31_257 ();
 FILLCELL_X2 FILLER_31_265 ();
 FILLCELL_X1 FILLER_31_267 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X32 FILLER_32_129 ();
 FILLCELL_X32 FILLER_32_161 ();
 FILLCELL_X32 FILLER_32_193 ();
 FILLCELL_X32 FILLER_32_225 ();
 FILLCELL_X8 FILLER_32_257 ();
 FILLCELL_X2 FILLER_32_265 ();
 FILLCELL_X1 FILLER_32_267 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X32 FILLER_33_129 ();
 FILLCELL_X32 FILLER_33_161 ();
 FILLCELL_X32 FILLER_33_193 ();
 FILLCELL_X32 FILLER_33_225 ();
 FILLCELL_X8 FILLER_33_257 ();
 FILLCELL_X2 FILLER_33_265 ();
 FILLCELL_X1 FILLER_33_267 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X16 FILLER_34_132 ();
 FILLCELL_X4 FILLER_34_148 ();
 FILLCELL_X2 FILLER_34_152 ();
 FILLCELL_X16 FILLER_34_157 ();
 FILLCELL_X4 FILLER_34_173 ();
 FILLCELL_X32 FILLER_34_180 ();
 FILLCELL_X32 FILLER_34_212 ();
 FILLCELL_X16 FILLER_34_244 ();
 FILLCELL_X8 FILLER_34_260 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X32 FILLER_35_33 ();
 FILLCELL_X32 FILLER_35_65 ();
 FILLCELL_X8 FILLER_35_97 ();
 FILLCELL_X4 FILLER_35_105 ();
 FILLCELL_X1 FILLER_35_109 ();
 FILLCELL_X2 FILLER_35_113 ();
 FILLCELL_X8 FILLER_35_118 ();
 FILLCELL_X1 FILLER_35_126 ();
 FILLCELL_X2 FILLER_35_131 ();
 FILLCELL_X1 FILLER_35_133 ();
 FILLCELL_X32 FILLER_35_137 ();
 FILLCELL_X32 FILLER_35_169 ();
 FILLCELL_X32 FILLER_35_201 ();
 FILLCELL_X32 FILLER_35_233 ();
 FILLCELL_X2 FILLER_35_265 ();
 FILLCELL_X1 FILLER_35_267 ();
endmodule
