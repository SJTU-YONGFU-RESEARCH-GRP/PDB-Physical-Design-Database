module configurable_kogge_stone_adder (cin,
    cout,
    a,
    b,
    sum);
 input cin;
 output cout;
 input [31:0] a;
 input [31:0] b;
 output [31:0] sum;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;

 sky130_fd_sc_hd__inv_1 _319_ (.A(net1),
    .Y(_251_));
 sky130_fd_sc_hd__inv_1 _320_ (.A(net33),
    .Y(_252_));
 sky130_fd_sc_hd__inv_1 _321_ (.A(net65),
    .Y(_253_));
 sky130_fd_sc_hd__inv_1 _322_ (.A(_256_),
    .Y(_000_));
 sky130_fd_sc_hd__and3_1 _323_ (.A(_258_),
    .B(_260_),
    .C(_262_),
    .X(_001_));
 sky130_fd_sc_hd__clkbuf_2 _324_ (.A(_264_),
    .X(_002_));
 sky130_fd_sc_hd__buf_2 _325_ (.A(_266_),
    .X(_003_));
 sky130_fd_sc_hd__buf_2 _326_ (.A(_272_),
    .X(_004_));
 sky130_fd_sc_hd__buf_2 _327_ (.A(_274_),
    .X(_005_));
 sky130_fd_sc_hd__a21o_1 _328_ (.A1(_276_),
    .A2(_277_),
    .B1(_275_),
    .X(_006_));
 sky130_fd_sc_hd__a21o_1 _329_ (.A1(_005_),
    .A2(_006_),
    .B1(_273_),
    .X(_007_));
 sky130_fd_sc_hd__a21oi_1 _330_ (.A1(_284_),
    .A2(_285_),
    .B1(_283_),
    .Y(_008_));
 sky130_fd_sc_hd__nand2_1 _331_ (.A(_280_),
    .B(_282_),
    .Y(_009_));
 sky130_fd_sc_hd__a21oi_1 _332_ (.A1(_280_),
    .A2(_281_),
    .B1(_279_),
    .Y(_010_));
 sky130_fd_sc_hd__o21ai_1 _333_ (.A1(_008_),
    .A2(_009_),
    .B1(_010_),
    .Y(_011_));
 sky130_fd_sc_hd__nand2_1 _334_ (.A(_276_),
    .B(_278_),
    .Y(_012_));
 sky130_fd_sc_hd__nand2_1 _335_ (.A(_004_),
    .B(_005_),
    .Y(_013_));
 sky130_fd_sc_hd__nor2_1 _336_ (.A(_012_),
    .B(_013_),
    .Y(_014_));
 sky130_fd_sc_hd__a221oi_2 _337_ (.A1(_004_),
    .A2(_007_),
    .B1(_011_),
    .B2(_014_),
    .C1(_271_),
    .Y(_015_));
 sky130_fd_sc_hd__a21o_1 _338_ (.A1(_298_),
    .A2(_299_),
    .B1(_297_),
    .X(_016_));
 sky130_fd_sc_hd__buf_2 _339_ (.A(_293_),
    .X(_017_));
 sky130_fd_sc_hd__a211oi_1 _340_ (.A1(_296_),
    .A2(_016_),
    .B1(_295_),
    .C1(_017_),
    .Y(_018_));
 sky130_fd_sc_hd__nor2_1 _341_ (.A(_301_),
    .B(_303_),
    .Y(_019_));
 sky130_fd_sc_hd__buf_6 _342_ (.A(_304_),
    .X(_020_));
 sky130_fd_sc_hd__o21ai_0 _343_ (.A1(_306_),
    .A2(_305_),
    .B1(_020_),
    .Y(_021_));
 sky130_fd_sc_hd__o21ai_0 _344_ (.A1(_302_),
    .A2(_301_),
    .B1(_300_),
    .Y(_022_));
 sky130_fd_sc_hd__nand2_1 _345_ (.A(_296_),
    .B(_298_),
    .Y(_023_));
 sky130_fd_sc_hd__a211o_1 _346_ (.A1(_019_),
    .A2(_021_),
    .B1(_022_),
    .C1(_023_),
    .X(_024_));
 sky130_fd_sc_hd__nor2_1 _347_ (.A(_294_),
    .B(_017_),
    .Y(_025_));
 sky130_fd_sc_hd__a21oi_2 _348_ (.A1(_018_),
    .A2(_024_),
    .B1(_025_),
    .Y(_026_));
 sky130_fd_sc_hd__a211o_1 _349_ (.A1(_020_),
    .A2(_305_),
    .B1(_303_),
    .C1(_301_),
    .X(_027_));
 sky130_fd_sc_hd__a2111oi_2 _350_ (.A1(_296_),
    .A2(_016_),
    .B1(_027_),
    .C1(_017_),
    .D1(_295_),
    .Y(_028_));
 sky130_fd_sc_hd__nand2_1 _351_ (.A(_308_),
    .B(_310_),
    .Y(_029_));
 sky130_fd_sc_hd__a21oi_1 _352_ (.A1(_312_),
    .A2(_313_),
    .B1(_311_),
    .Y(_030_));
 sky130_fd_sc_hd__a21oi_1 _353_ (.A1(_316_),
    .A2(_317_),
    .B1(_315_),
    .Y(_031_));
 sky130_fd_sc_hd__nand4_1 _354_ (.A(_312_),
    .B(_308_),
    .C(_310_),
    .D(_314_),
    .Y(_032_));
 sky130_fd_sc_hd__a21oi_1 _355_ (.A1(_308_),
    .A2(_309_),
    .B1(_307_),
    .Y(_033_));
 sky130_fd_sc_hd__o221a_1 _356_ (.A1(_029_),
    .A2(_030_),
    .B1(_031_),
    .B2(_032_),
    .C1(_033_),
    .X(_034_));
 sky130_fd_sc_hd__clkbuf_4 _357_ (.A(_292_),
    .X(_035_));
 sky130_fd_sc_hd__clkbuf_2 _358_ (.A(_286_),
    .X(_036_));
 sky130_fd_sc_hd__clkbuf_2 _359_ (.A(_288_),
    .X(_037_));
 sky130_fd_sc_hd__clkbuf_2 _360_ (.A(_290_),
    .X(_038_));
 sky130_fd_sc_hd__and4_1 _361_ (.A(_284_),
    .B(_036_),
    .C(_037_),
    .D(_038_),
    .X(_039_));
 sky130_fd_sc_hd__nand2_1 _362_ (.A(_035_),
    .B(_039_),
    .Y(_040_));
 sky130_fd_sc_hd__a21oi_1 _363_ (.A1(_028_),
    .A2(_034_),
    .B1(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__nand2_1 _364_ (.A(_284_),
    .B(_036_),
    .Y(_042_));
 sky130_fd_sc_hd__a21oi_1 _365_ (.A1(_037_),
    .A2(_289_),
    .B1(_287_),
    .Y(_043_));
 sky130_fd_sc_hd__nand2_1 _366_ (.A(_291_),
    .B(_039_),
    .Y(_044_));
 sky130_fd_sc_hd__o21ai_0 _367_ (.A1(_042_),
    .A2(_043_),
    .B1(_044_),
    .Y(_045_));
 sky130_fd_sc_hd__a21oi_2 _368_ (.A1(_026_),
    .A2(_041_),
    .B1(_045_),
    .Y(_046_));
 sky130_fd_sc_hd__nor2_1 _369_ (.A(_267_),
    .B(_269_),
    .Y(_047_));
 sky130_fd_sc_hd__nor2_1 _370_ (.A(_009_),
    .B(_012_),
    .Y(_048_));
 sky130_fd_sc_hd__nand3_1 _371_ (.A(_004_),
    .B(_005_),
    .C(_048_),
    .Y(_049_));
 sky130_fd_sc_hd__clkbuf_2 _372_ (.A(_270_),
    .X(_050_));
 sky130_fd_sc_hd__o21ai_0 _373_ (.A1(_050_),
    .A2(_269_),
    .B1(_268_),
    .Y(_051_));
 sky130_fd_sc_hd__inv_1 _374_ (.A(_267_),
    .Y(_052_));
 sky130_fd_sc_hd__a32o_1 _375_ (.A1(_015_),
    .A2(_049_),
    .A3(_047_),
    .B1(_051_),
    .B2(_052_),
    .X(_053_));
 sky130_fd_sc_hd__a31oi_2 _376_ (.A1(_015_),
    .A2(_046_),
    .A3(_047_),
    .B1(_053_),
    .Y(_054_));
 sky130_fd_sc_hd__a21o_1 _377_ (.A1(_003_),
    .A2(_054_),
    .B1(_265_),
    .X(_055_));
 sky130_fd_sc_hd__a21o_1 _378_ (.A1(_002_),
    .A2(_055_),
    .B1(_263_),
    .X(_056_));
 sky130_fd_sc_hd__nor2_1 _379_ (.A(_265_),
    .B(_054_),
    .Y(_057_));
 sky130_fd_sc_hd__nand4_1 _380_ (.A(_005_),
    .B(_276_),
    .C(_278_),
    .D(_280_),
    .Y(_058_));
 sky130_fd_sc_hd__a21oi_1 _381_ (.A1(_038_),
    .A2(_291_),
    .B1(_289_),
    .Y(_059_));
 sky130_fd_sc_hd__nand2_1 _382_ (.A(_036_),
    .B(_037_),
    .Y(_060_));
 sky130_fd_sc_hd__a21oi_1 _383_ (.A1(_036_),
    .A2(_287_),
    .B1(_285_),
    .Y(_061_));
 sky130_fd_sc_hd__o21a_1 _384_ (.A1(_059_),
    .A2(_060_),
    .B1(_061_),
    .X(_062_));
 sky130_fd_sc_hd__nand2_1 _385_ (.A(_282_),
    .B(_284_),
    .Y(_063_));
 sky130_fd_sc_hd__a21oi_1 _386_ (.A1(_282_),
    .A2(_283_),
    .B1(_281_),
    .Y(_064_));
 sky130_fd_sc_hd__o21a_1 _387_ (.A1(_062_),
    .A2(_063_),
    .B1(_064_),
    .X(_065_));
 sky130_fd_sc_hd__nand2_1 _388_ (.A(_005_),
    .B(_276_),
    .Y(_066_));
 sky130_fd_sc_hd__a21oi_1 _389_ (.A1(_278_),
    .A2(_279_),
    .B1(_277_),
    .Y(_067_));
 sky130_fd_sc_hd__a21oi_1 _390_ (.A1(_005_),
    .A2(_275_),
    .B1(_273_),
    .Y(_068_));
 sky130_fd_sc_hd__o21ai_0 _391_ (.A1(_066_),
    .A2(_067_),
    .B1(_068_),
    .Y(_069_));
 sky130_fd_sc_hd__nor2_1 _392_ (.A(_271_),
    .B(_069_),
    .Y(_070_));
 sky130_fd_sc_hd__o21ai_0 _393_ (.A1(_058_),
    .A2(_065_),
    .B1(_070_),
    .Y(_071_));
 sky130_fd_sc_hd__o21a_1 _394_ (.A1(_004_),
    .A2(_271_),
    .B1(_050_),
    .X(_072_));
 sky130_fd_sc_hd__a21o_1 _395_ (.A1(_071_),
    .A2(_072_),
    .B1(_269_),
    .X(_073_));
 sky130_fd_sc_hd__a211oi_1 _396_ (.A1(_306_),
    .A2(_307_),
    .B1(_305_),
    .C1(_303_),
    .Y(_074_));
 sky130_fd_sc_hd__o21ai_0 _397_ (.A1(_020_),
    .A2(_303_),
    .B1(_302_),
    .Y(_075_));
 sky130_fd_sc_hd__nor3_1 _398_ (.A(_297_),
    .B(_299_),
    .C(_301_),
    .Y(_076_));
 sky130_fd_sc_hd__o21a_1 _399_ (.A1(_074_),
    .A2(_075_),
    .B1(_076_),
    .X(_077_));
 sky130_fd_sc_hd__o21a_1 _400_ (.A1(_300_),
    .A2(_299_),
    .B1(_298_),
    .X(_078_));
 sky130_fd_sc_hd__o21ai_1 _401_ (.A1(_297_),
    .A2(_078_),
    .B1(_296_),
    .Y(_079_));
 sky130_fd_sc_hd__and4_1 _402_ (.A(_302_),
    .B(_020_),
    .C(_306_),
    .D(_308_),
    .X(_080_));
 sky130_fd_sc_hd__o211ai_2 _403_ (.A1(_297_),
    .A2(_078_),
    .B1(_080_),
    .C1(_296_),
    .Y(_081_));
 sky130_fd_sc_hd__inv_1 _404_ (.A(_310_),
    .Y(_082_));
 sky130_fd_sc_hd__nand3_1 _405_ (.A(_312_),
    .B(_310_),
    .C(_314_),
    .Y(_083_));
 sky130_fd_sc_hd__inv_1 _406_ (.A(_309_),
    .Y(_084_));
 sky130_fd_sc_hd__o221a_2 _407_ (.A1(_082_),
    .A2(_030_),
    .B1(_031_),
    .B2(_083_),
    .C1(_084_),
    .X(_085_));
 sky130_fd_sc_hd__inv_1 _408_ (.A(_295_),
    .Y(_086_));
 sky130_fd_sc_hd__o221ai_4 _409_ (.A1(_077_),
    .A2(_079_),
    .B1(_081_),
    .B2(_085_),
    .C1(_086_),
    .Y(_087_));
 sky130_fd_sc_hd__a21oi_2 _410_ (.A1(_294_),
    .A2(_087_),
    .B1(_017_),
    .Y(_088_));
 sky130_fd_sc_hd__nand4_2 _411_ (.A(_036_),
    .B(_037_),
    .C(_038_),
    .D(_035_),
    .Y(_089_));
 sky130_fd_sc_hd__nand4_1 _412_ (.A(_278_),
    .B(_280_),
    .C(_282_),
    .D(_284_),
    .Y(_090_));
 sky130_fd_sc_hd__nand4_1 _413_ (.A(_050_),
    .B(_004_),
    .C(_005_),
    .D(_276_),
    .Y(_091_));
 sky130_fd_sc_hd__or2_1 _414_ (.A(_090_),
    .B(_091_),
    .X(_092_));
 sky130_fd_sc_hd__nor3_1 _415_ (.A(_088_),
    .B(_089_),
    .C(_092_),
    .Y(_093_));
 sky130_fd_sc_hd__nand4_1 _416_ (.A(_262_),
    .B(_002_),
    .C(_003_),
    .D(_268_),
    .Y(_094_));
 sky130_fd_sc_hd__or3_1 _417_ (.A(_089_),
    .B(_092_),
    .C(_094_),
    .X(_095_));
 sky130_fd_sc_hd__nand2_1 _418_ (.A(_278_),
    .B(_280_),
    .Y(_096_));
 sky130_fd_sc_hd__o21a_1 _419_ (.A1(_096_),
    .A2(_064_),
    .B1(_067_),
    .X(_097_));
 sky130_fd_sc_hd__o22ai_1 _420_ (.A1(_062_),
    .A2(_092_),
    .B1(_097_),
    .B2(_091_),
    .Y(_098_));
 sky130_fd_sc_hd__a21o_1 _421_ (.A1(_003_),
    .A2(_267_),
    .B1(_265_),
    .X(_099_));
 sky130_fd_sc_hd__inv_1 _422_ (.A(_004_),
    .Y(_100_));
 sky130_fd_sc_hd__o21bai_1 _423_ (.A1(_100_),
    .A2(_068_),
    .B1_N(_271_),
    .Y(_101_));
 sky130_fd_sc_hd__or3_1 _424_ (.A(_261_),
    .B(_263_),
    .C(_269_),
    .X(_102_));
 sky130_fd_sc_hd__a221o_1 _425_ (.A1(_002_),
    .A2(_099_),
    .B1(_101_),
    .B2(_050_),
    .C1(_102_),
    .X(_103_));
 sky130_fd_sc_hd__inv_1 _426_ (.A(_263_),
    .Y(_104_));
 sky130_fd_sc_hd__o21a_1 _427_ (.A1(_268_),
    .A2(_267_),
    .B1(_003_),
    .X(_105_));
 sky130_fd_sc_hd__o21ai_0 _428_ (.A1(_265_),
    .A2(_105_),
    .B1(_002_),
    .Y(_106_));
 sky130_fd_sc_hd__a21boi_0 _429_ (.A1(_104_),
    .A2(_106_),
    .B1_N(_262_),
    .Y(_107_));
 sky130_fd_sc_hd__o22ai_1 _430_ (.A1(_098_),
    .A2(_103_),
    .B1(_107_),
    .B2(_261_),
    .Y(_108_));
 sky130_fd_sc_hd__o21ai_0 _431_ (.A1(_088_),
    .A2(_095_),
    .B1(_108_),
    .Y(_109_));
 sky130_fd_sc_hd__nand2_1 _432_ (.A(_028_),
    .B(_034_),
    .Y(_110_));
 sky130_fd_sc_hd__a31o_1 _433_ (.A1(_035_),
    .A2(_110_),
    .A3(_026_),
    .B1(_291_),
    .X(_111_));
 sky130_fd_sc_hd__o21ai_2 _434_ (.A1(_042_),
    .A2(_043_),
    .B1(_008_),
    .Y(_112_));
 sky130_fd_sc_hd__nor2_1 _435_ (.A(_010_),
    .B(_012_),
    .Y(_113_));
 sky130_fd_sc_hd__a211oi_2 _436_ (.A1(_048_),
    .A2(_112_),
    .B1(_113_),
    .C1(_006_),
    .Y(_114_));
 sky130_fd_sc_hd__o21ai_0 _437_ (.A1(_003_),
    .A2(_265_),
    .B1(_002_),
    .Y(_115_));
 sky130_fd_sc_hd__nand2_1 _438_ (.A(_260_),
    .B(_262_),
    .Y(_116_));
 sky130_fd_sc_hd__a21oi_1 _439_ (.A1(_104_),
    .A2(_115_),
    .B1(_116_),
    .Y(_117_));
 sky130_fd_sc_hd__nand2_1 _440_ (.A(_268_),
    .B(_050_),
    .Y(_118_));
 sky130_fd_sc_hd__nor2_1 _441_ (.A(_013_),
    .B(_118_),
    .Y(_119_));
 sky130_fd_sc_hd__nand2_1 _442_ (.A(_117_),
    .B(_119_),
    .Y(_120_));
 sky130_fd_sc_hd__a21oi_1 _443_ (.A1(_004_),
    .A2(_273_),
    .B1(_271_),
    .Y(_121_));
 sky130_fd_sc_hd__a2111oi_0 _444_ (.A1(_268_),
    .A2(_269_),
    .B1(_267_),
    .C1(_265_),
    .D1(_263_),
    .Y(_122_));
 sky130_fd_sc_hd__o21ai_0 _445_ (.A1(_121_),
    .A2(_118_),
    .B1(_122_),
    .Y(_123_));
 sky130_fd_sc_hd__a21o_1 _446_ (.A1(_260_),
    .A2(_261_),
    .B1(_259_),
    .X(_124_));
 sky130_fd_sc_hd__a21oi_1 _447_ (.A1(_117_),
    .A2(_123_),
    .B1(_124_),
    .Y(_125_));
 sky130_fd_sc_hd__o21ai_0 _448_ (.A1(_114_),
    .A2(_120_),
    .B1(_125_),
    .Y(_126_));
 sky130_fd_sc_hd__nor2_1 _449_ (.A(_111_),
    .B(_126_),
    .Y(_127_));
 sky130_fd_sc_hd__nor4b_1 _450_ (.A(_073_),
    .B(_093_),
    .C(_109_),
    .D_N(_127_),
    .Y(_128_));
 sky130_fd_sc_hd__a31oi_4 _451_ (.A1(_035_),
    .A2(_110_),
    .A3(_026_),
    .B1(_291_),
    .Y(_129_));
 sky130_fd_sc_hd__nand2_1 _452_ (.A(_039_),
    .B(_048_),
    .Y(_130_));
 sky130_fd_sc_hd__o21ai_2 _453_ (.A1(_129_),
    .A2(_130_),
    .B1(_114_),
    .Y(_131_));
 sky130_fd_sc_hd__o21bai_1 _454_ (.A1(_009_),
    .A2(_046_),
    .B1_N(_011_),
    .Y(_132_));
 sky130_fd_sc_hd__nor2b_1 _455_ (.A(_254_),
    .B_N(_318_),
    .Y(_133_));
 sky130_fd_sc_hd__o2111a_1 _456_ (.A1(_317_),
    .A2(_133_),
    .B1(_314_),
    .C1(_312_),
    .D1(_316_),
    .X(_134_));
 sky130_fd_sc_hd__nand2_1 _457_ (.A(_312_),
    .B(_313_),
    .Y(_135_));
 sky130_fd_sc_hd__nand3_1 _458_ (.A(_312_),
    .B(_314_),
    .C(_315_),
    .Y(_136_));
 sky130_fd_sc_hd__nand2_1 _459_ (.A(_135_),
    .B(_136_),
    .Y(_137_));
 sky130_fd_sc_hd__nor3_2 _460_ (.A(_311_),
    .B(_134_),
    .C(_137_),
    .Y(_138_));
 sky130_fd_sc_hd__o221ai_2 _461_ (.A1(_029_),
    .A2(_030_),
    .B1(_031_),
    .B2(_032_),
    .C1(_033_),
    .Y(_139_));
 sky130_fd_sc_hd__nor3_1 _462_ (.A(_305_),
    .B(_309_),
    .C(_139_),
    .Y(_140_));
 sky130_fd_sc_hd__inv_1 _463_ (.A(_308_),
    .Y(_141_));
 sky130_fd_sc_hd__nand2_1 _464_ (.A(_020_),
    .B(_306_),
    .Y(_142_));
 sky130_fd_sc_hd__nand2_1 _465_ (.A(_316_),
    .B(_318_),
    .Y(_143_));
 sky130_fd_sc_hd__or2_1 _466_ (.A(_083_),
    .B(_143_),
    .X(_144_));
 sky130_fd_sc_hd__nor3_1 _467_ (.A(_141_),
    .B(_142_),
    .C(_144_),
    .Y(_145_));
 sky130_fd_sc_hd__a21boi_2 _468_ (.A1(_138_),
    .A2(_140_),
    .B1_N(_145_),
    .Y(_146_));
 sky130_fd_sc_hd__nor2_1 _469_ (.A(_297_),
    .B(_078_),
    .Y(_147_));
 sky130_fd_sc_hd__o21ai_0 _470_ (.A1(_297_),
    .A2(_078_),
    .B1(_080_),
    .Y(_148_));
 sky130_fd_sc_hd__o22ai_2 _471_ (.A1(_147_),
    .A2(_077_),
    .B1(_085_),
    .B2(_148_),
    .Y(_149_));
 sky130_fd_sc_hd__o21bai_2 _472_ (.A1(_034_),
    .A2(_142_),
    .B1_N(_027_),
    .Y(_150_));
 sky130_fd_sc_hd__nor3_2 _473_ (.A(_299_),
    .B(_149_),
    .C(_150_),
    .Y(_151_));
 sky130_fd_sc_hd__nor2_1 _474_ (.A(_291_),
    .B(_087_),
    .Y(_152_));
 sky130_fd_sc_hd__nand4bb_2 _475_ (.A_N(_017_),
    .B_N(_146_),
    .C(_151_),
    .D(_152_),
    .Y(_153_));
 sky130_fd_sc_hd__a21o_1 _476_ (.A1(_294_),
    .A2(_087_),
    .B1(_017_),
    .X(_154_));
 sky130_fd_sc_hd__nor2_1 _477_ (.A(_089_),
    .B(_090_),
    .Y(_155_));
 sky130_fd_sc_hd__o21ai_0 _478_ (.A1(_062_),
    .A2(_090_),
    .B1(_097_),
    .Y(_156_));
 sky130_fd_sc_hd__a21o_1 _479_ (.A1(_154_),
    .A2(_155_),
    .B1(_156_),
    .X(_157_));
 sky130_fd_sc_hd__nand2_1 _480_ (.A(_037_),
    .B(_038_),
    .Y(_158_));
 sky130_fd_sc_hd__nand2_1 _481_ (.A(_036_),
    .B(_035_),
    .Y(_159_));
 sky130_fd_sc_hd__nor2_1 _482_ (.A(_158_),
    .B(_159_),
    .Y(_160_));
 sky130_fd_sc_hd__nand4_1 _483_ (.A(_302_),
    .B(_020_),
    .C(_306_),
    .D(_308_),
    .Y(_161_));
 sky130_fd_sc_hd__nand4_1 _484_ (.A(_294_),
    .B(_296_),
    .C(_298_),
    .D(_300_),
    .Y(_162_));
 sky130_fd_sc_hd__nor4_2 _485_ (.A(_083_),
    .B(_161_),
    .C(_143_),
    .D(_162_),
    .Y(_163_));
 sky130_fd_sc_hd__nand2_2 _486_ (.A(_160_),
    .B(_163_),
    .Y(_164_));
 sky130_fd_sc_hd__nor2_1 _487_ (.A(_092_),
    .B(_164_),
    .Y(_165_));
 sky130_fd_sc_hd__o41ai_2 _488_ (.A1(_131_),
    .A2(_132_),
    .A3(_153_),
    .A4(_157_),
    .B1(_165_),
    .Y(_166_));
 sky130_fd_sc_hd__nand3_1 _489_ (.A(_057_),
    .B(_128_),
    .C(_166_),
    .Y(_167_));
 sky130_fd_sc_hd__nand4_1 _490_ (.A(_003_),
    .B(_268_),
    .C(_050_),
    .D(_004_),
    .Y(_168_));
 sky130_fd_sc_hd__nor4_2 _491_ (.A(_058_),
    .B(_063_),
    .C(_164_),
    .D(_168_),
    .Y(_169_));
 sky130_fd_sc_hd__and3_1 _492_ (.A(_002_),
    .B(_001_),
    .C(_169_),
    .X(_170_));
 sky130_fd_sc_hd__a21o_1 _493_ (.A1(_258_),
    .A2(_124_),
    .B1(_257_),
    .X(_171_));
 sky130_fd_sc_hd__a221oi_2 _494_ (.A1(_001_),
    .A2(_056_),
    .B1(_167_),
    .B2(_170_),
    .C1(_171_),
    .Y(_172_));
 sky130_fd_sc_hd__o21bai_1 _495_ (.A1(_000_),
    .A2(_172_),
    .B1_N(_255_),
    .Y(net66));
 sky130_fd_sc_hd__nand3_2 _496_ (.A(_300_),
    .B(_302_),
    .C(_145_),
    .Y(_173_));
 sky130_fd_sc_hd__nand2b_1 _497_ (.A_N(_022_),
    .B(_150_),
    .Y(_174_));
 sky130_fd_sc_hd__a2bb2oi_1 _498_ (.A1_N(_146_),
    .A2_N(_150_),
    .B1(_173_),
    .B2(_174_),
    .Y(_175_));
 sky130_fd_sc_hd__nor2_1 _499_ (.A(_299_),
    .B(_175_),
    .Y(_176_));
 sky130_fd_sc_hd__xnor2_1 _500_ (.A(_298_),
    .B(_176_),
    .Y(net68));
 sky130_fd_sc_hd__nor3b_1 _501_ (.A(_176_),
    .B(_173_),
    .C_N(_298_),
    .Y(_177_));
 sky130_fd_sc_hd__nor2_1 _502_ (.A(_149_),
    .B(_177_),
    .Y(_178_));
 sky130_fd_sc_hd__xnor2_1 _503_ (.A(_296_),
    .B(_178_),
    .Y(net69));
 sky130_fd_sc_hd__nor2_1 _504_ (.A(_305_),
    .B(_139_),
    .Y(_179_));
 sky130_fd_sc_hd__a211o_1 _505_ (.A1(_084_),
    .A2(_138_),
    .B1(_144_),
    .C1(_141_),
    .X(_180_));
 sky130_fd_sc_hd__a311oi_4 _506_ (.A1(_179_),
    .A2(_151_),
    .A3(_180_),
    .B1(_173_),
    .C1(_023_),
    .Y(_181_));
 sky130_fd_sc_hd__nor2_1 _507_ (.A(_087_),
    .B(_181_),
    .Y(_182_));
 sky130_fd_sc_hd__xnor2_1 _508_ (.A(_294_),
    .B(_182_),
    .Y(net70));
 sky130_fd_sc_hd__or3_1 _509_ (.A(_161_),
    .B(_144_),
    .C(_162_),
    .X(_183_));
 sky130_fd_sc_hd__o21ai_0 _510_ (.A1(_183_),
    .A2(_182_),
    .B1(_088_),
    .Y(_184_));
 sky130_fd_sc_hd__xor2_1 _511_ (.A(_035_),
    .B(_184_),
    .X(net71));
 sky130_fd_sc_hd__nand2_1 _512_ (.A(_035_),
    .B(_163_),
    .Y(_185_));
 sky130_fd_sc_hd__nor3_1 _513_ (.A(_017_),
    .B(_087_),
    .C(_181_),
    .Y(_186_));
 sky130_fd_sc_hd__o21ai_1 _514_ (.A1(_185_),
    .A2(_186_),
    .B1(_129_),
    .Y(_187_));
 sky130_fd_sc_hd__xor2_1 _515_ (.A(_038_),
    .B(_187_),
    .X(net72));
 sky130_fd_sc_hd__a21oi_1 _516_ (.A1(_038_),
    .A2(_187_),
    .B1(_289_),
    .Y(_188_));
 sky130_fd_sc_hd__xnor2_1 _517_ (.A(_037_),
    .B(_188_),
    .Y(net73));
 sky130_fd_sc_hd__nor2_1 _518_ (.A(_185_),
    .B(_186_),
    .Y(_189_));
 sky130_fd_sc_hd__nor3_1 _519_ (.A(_038_),
    .B(_287_),
    .C(_289_),
    .Y(_190_));
 sky130_fd_sc_hd__nor2_1 _520_ (.A(_037_),
    .B(_287_),
    .Y(_191_));
 sky130_fd_sc_hd__nor2_1 _521_ (.A(_190_),
    .B(_191_),
    .Y(_192_));
 sky130_fd_sc_hd__o41ai_1 _522_ (.A1(_287_),
    .A2(_289_),
    .A3(_111_),
    .A4(_189_),
    .B1(_192_),
    .Y(_193_));
 sky130_fd_sc_hd__xnor2_1 _523_ (.A(_036_),
    .B(_193_),
    .Y(net74));
 sky130_fd_sc_hd__a2111oi_0 _524_ (.A1(_035_),
    .A2(_017_),
    .B1(_087_),
    .C1(_181_),
    .D1(_291_),
    .Y(_194_));
 sky130_fd_sc_hd__o21ai_0 _525_ (.A1(_183_),
    .A2(_194_),
    .B1(_088_),
    .Y(_195_));
 sky130_fd_sc_hd__o21ai_0 _526_ (.A1(_129_),
    .A2(_164_),
    .B1(_062_),
    .Y(_196_));
 sky130_fd_sc_hd__a21oi_1 _527_ (.A1(_160_),
    .A2(_195_),
    .B1(_196_),
    .Y(_197_));
 sky130_fd_sc_hd__xnor2_1 _528_ (.A(_284_),
    .B(_197_),
    .Y(net75));
 sky130_fd_sc_hd__o41ai_1 _529_ (.A1(_017_),
    .A2(_111_),
    .A3(_087_),
    .A4(_181_),
    .B1(_160_),
    .Y(_198_));
 sky130_fd_sc_hd__nor3_1 _530_ (.A(_111_),
    .B(_112_),
    .C(_196_),
    .Y(_199_));
 sky130_fd_sc_hd__a21oi_1 _531_ (.A1(_035_),
    .A2(_163_),
    .B1(_112_),
    .Y(_200_));
 sky130_fd_sc_hd__nand2_1 _532_ (.A(_129_),
    .B(_200_),
    .Y(_201_));
 sky130_fd_sc_hd__o21ai_0 _533_ (.A1(_039_),
    .A2(_112_),
    .B1(_201_),
    .Y(_202_));
 sky130_fd_sc_hd__a21oi_1 _534_ (.A1(_198_),
    .A2(_199_),
    .B1(_202_),
    .Y(_203_));
 sky130_fd_sc_hd__xor2_1 _535_ (.A(_282_),
    .B(_203_),
    .X(net76));
 sky130_fd_sc_hd__nor2_1 _536_ (.A(_063_),
    .B(_164_),
    .Y(_204_));
 sky130_fd_sc_hd__o31ai_1 _537_ (.A1(_063_),
    .A2(_088_),
    .A3(_089_),
    .B1(_065_),
    .Y(_205_));
 sky130_fd_sc_hd__a21oi_1 _538_ (.A1(_204_),
    .A2(_203_),
    .B1(_205_),
    .Y(_206_));
 sky130_fd_sc_hd__xnor2_1 _539_ (.A(_280_),
    .B(_206_),
    .Y(net77));
 sky130_fd_sc_hd__xnor2_1 _540_ (.A(_316_),
    .B(_254_),
    .Y(net78));
 sky130_fd_sc_hd__nor4_1 _541_ (.A(_009_),
    .B(_042_),
    .C(_158_),
    .D(_185_),
    .Y(_207_));
 sky130_fd_sc_hd__a21oi_1 _542_ (.A1(_153_),
    .A2(_207_),
    .B1(_132_),
    .Y(_208_));
 sky130_fd_sc_hd__xnor2_1 _543_ (.A(_278_),
    .B(_208_),
    .Y(net79));
 sky130_fd_sc_hd__nor2_1 _544_ (.A(_090_),
    .B(_164_),
    .Y(_209_));
 sky130_fd_sc_hd__and2_0 _545_ (.A(_207_),
    .B(_209_),
    .X(_210_));
 sky130_fd_sc_hd__a22oi_1 _546_ (.A1(_132_),
    .A2(_209_),
    .B1(_210_),
    .B2(_153_),
    .Y(_211_));
 sky130_fd_sc_hd__nor2b_1 _547_ (.A(_157_),
    .B_N(_211_),
    .Y(_212_));
 sky130_fd_sc_hd__xnor2_1 _548_ (.A(_276_),
    .B(_212_),
    .Y(net80));
 sky130_fd_sc_hd__nor2_1 _549_ (.A(_131_),
    .B(_157_),
    .Y(_213_));
 sky130_fd_sc_hd__nand2_1 _550_ (.A(_208_),
    .B(_213_),
    .Y(_214_));
 sky130_fd_sc_hd__nand4_2 _551_ (.A(_035_),
    .B(_039_),
    .C(_048_),
    .D(_163_),
    .Y(_215_));
 sky130_fd_sc_hd__o211ai_1 _552_ (.A1(_129_),
    .A2(_130_),
    .B1(_215_),
    .C1(_114_),
    .Y(_216_));
 sky130_fd_sc_hd__nand2_1 _553_ (.A(_214_),
    .B(_216_),
    .Y(_217_));
 sky130_fd_sc_hd__xnor2_1 _554_ (.A(_005_),
    .B(_217_),
    .Y(net81));
 sky130_fd_sc_hd__nor3_1 _555_ (.A(_131_),
    .B(_157_),
    .C(_205_),
    .Y(_218_));
 sky130_fd_sc_hd__nand2_1 _556_ (.A(_211_),
    .B(_218_),
    .Y(_219_));
 sky130_fd_sc_hd__a21oi_1 _557_ (.A1(_204_),
    .A2(_216_),
    .B1(_205_),
    .Y(_220_));
 sky130_fd_sc_hd__nor2_1 _558_ (.A(_058_),
    .B(_220_),
    .Y(_221_));
 sky130_fd_sc_hd__a21oi_1 _559_ (.A1(_219_),
    .A2(_221_),
    .B1(_069_),
    .Y(_222_));
 sky130_fd_sc_hd__xnor2_1 _560_ (.A(_004_),
    .B(_222_),
    .Y(net82));
 sky130_fd_sc_hd__nor3_1 _561_ (.A(_013_),
    .B(_215_),
    .C(_220_),
    .Y(_223_));
 sky130_fd_sc_hd__o21ai_0 _562_ (.A1(_046_),
    .A2(_049_),
    .B1(_015_),
    .Y(_224_));
 sky130_fd_sc_hd__a21oi_1 _563_ (.A1(_219_),
    .A2(_223_),
    .B1(_224_),
    .Y(_225_));
 sky130_fd_sc_hd__xnor2_1 _564_ (.A(_050_),
    .B(_225_),
    .Y(net83));
 sky130_fd_sc_hd__nor2_1 _565_ (.A(_073_),
    .B(_093_),
    .Y(_226_));
 sky130_fd_sc_hd__nand2_1 _566_ (.A(_226_),
    .B(_166_),
    .Y(_227_));
 sky130_fd_sc_hd__xor2_1 _567_ (.A(_268_),
    .B(_227_),
    .X(net84));
 sky130_fd_sc_hd__nor3_1 _568_ (.A(_013_),
    .B(_118_),
    .C(_215_),
    .Y(_228_));
 sky130_fd_sc_hd__a21oi_1 _569_ (.A1(_227_),
    .A2(_228_),
    .B1(_054_),
    .Y(_229_));
 sky130_fd_sc_hd__xnor2_1 _570_ (.A(_003_),
    .B(_229_),
    .Y(net85));
 sky130_fd_sc_hd__nand3_1 _571_ (.A(_057_),
    .B(_226_),
    .C(_166_),
    .Y(_230_));
 sky130_fd_sc_hd__o21ai_0 _572_ (.A1(_055_),
    .A2(_169_),
    .B1(_230_),
    .Y(_231_));
 sky130_fd_sc_hd__xnor2_1 _573_ (.A(_002_),
    .B(_231_),
    .Y(net86));
 sky130_fd_sc_hd__nand3_1 _574_ (.A(_002_),
    .B(_003_),
    .C(_119_),
    .Y(_232_));
 sky130_fd_sc_hd__nor2_1 _575_ (.A(_215_),
    .B(_232_),
    .Y(_233_));
 sky130_fd_sc_hd__o21a_1 _576_ (.A1(_055_),
    .A2(_169_),
    .B1(_233_),
    .X(_234_));
 sky130_fd_sc_hd__a21oi_1 _577_ (.A1(_230_),
    .A2(_234_),
    .B1(_056_),
    .Y(_235_));
 sky130_fd_sc_hd__xnor2_1 _578_ (.A(_262_),
    .B(_235_),
    .Y(net87));
 sky130_fd_sc_hd__nor2_1 _579_ (.A(_095_),
    .B(_183_),
    .Y(_236_));
 sky130_fd_sc_hd__a21oi_1 _580_ (.A1(_230_),
    .A2(_236_),
    .B1(_109_),
    .Y(_237_));
 sky130_fd_sc_hd__xnor2_1 _581_ (.A(_260_),
    .B(_237_),
    .Y(net88));
 sky130_fd_sc_hd__o21ai_0 _582_ (.A1(_317_),
    .A2(_133_),
    .B1(_316_),
    .Y(_238_));
 sky130_fd_sc_hd__nand2b_1 _583_ (.A_N(_315_),
    .B(_238_),
    .Y(_239_));
 sky130_fd_sc_hd__xor2_1 _584_ (.A(_314_),
    .B(_239_),
    .X(net89));
 sky130_fd_sc_hd__a2111oi_0 _585_ (.A1(_129_),
    .A2(_185_),
    .B1(_232_),
    .C1(_130_),
    .D1(_116_),
    .Y(_240_));
 sky130_fd_sc_hd__o21ai_1 _586_ (.A1(_126_),
    .A2(_240_),
    .B1(_167_),
    .Y(_241_));
 sky130_fd_sc_hd__xnor2_1 _587_ (.A(_258_),
    .B(_241_),
    .Y(net90));
 sky130_fd_sc_hd__xnor2_1 _588_ (.A(_256_),
    .B(_172_),
    .Y(net91));
 sky130_fd_sc_hd__a211oi_1 _589_ (.A1(_314_),
    .A2(_239_),
    .B1(_313_),
    .C1(_312_),
    .Y(_242_));
 sky130_fd_sc_hd__nor3_1 _590_ (.A(_134_),
    .B(_137_),
    .C(_242_),
    .Y(net92));
 sky130_fd_sc_hd__xnor2_1 _591_ (.A(_310_),
    .B(_138_),
    .Y(net93));
 sky130_fd_sc_hd__o21ai_0 _592_ (.A1(_144_),
    .A2(_138_),
    .B1(_085_),
    .Y(_243_));
 sky130_fd_sc_hd__xnor2_1 _593_ (.A(_141_),
    .B(_243_),
    .Y(net94));
 sky130_fd_sc_hd__nand2_1 _594_ (.A(_034_),
    .B(_180_),
    .Y(_244_));
 sky130_fd_sc_hd__xor2_1 _595_ (.A(_306_),
    .B(_244_),
    .X(net95));
 sky130_fd_sc_hd__a21oi_1 _596_ (.A1(_306_),
    .A2(_244_),
    .B1(_305_),
    .Y(_245_));
 sky130_fd_sc_hd__xnor2_1 _597_ (.A(_020_),
    .B(_245_),
    .Y(net96));
 sky130_fd_sc_hd__nor2_1 _598_ (.A(_034_),
    .B(_142_),
    .Y(_246_));
 sky130_fd_sc_hd__a2111oi_2 _599_ (.A1(_020_),
    .A2(_305_),
    .B1(_146_),
    .C1(_246_),
    .D1(_303_),
    .Y(_247_));
 sky130_fd_sc_hd__xnor2_1 _600_ (.A(_302_),
    .B(_247_),
    .Y(net97));
 sky130_fd_sc_hd__o21ai_0 _601_ (.A1(_144_),
    .A2(_247_),
    .B1(_085_),
    .Y(_248_));
 sky130_fd_sc_hd__nor2_1 _602_ (.A(_074_),
    .B(_075_),
    .Y(_249_));
 sky130_fd_sc_hd__a2111oi_0 _603_ (.A1(_080_),
    .A2(_248_),
    .B1(_300_),
    .C1(_301_),
    .D1(_249_),
    .Y(_250_));
 sky130_fd_sc_hd__nor2_1 _604_ (.A(_175_),
    .B(_250_),
    .Y(net98));
 sky130_fd_sc_hd__fa_1 _605_ (.A(_251_),
    .B(_252_),
    .CIN(_253_),
    .COUT(_254_),
    .SUM(net67));
 sky130_fd_sc_hd__ha_1 _606_ (.A(net25),
    .B(net57),
    .COUT(_255_),
    .SUM(_256_));
 sky130_fd_sc_hd__ha_1 _607_ (.A(net24),
    .B(net56),
    .COUT(_257_),
    .SUM(_258_));
 sky130_fd_sc_hd__ha_1 _608_ (.A(net22),
    .B(net54),
    .COUT(_259_),
    .SUM(_260_));
 sky130_fd_sc_hd__ha_1 _609_ (.A(net21),
    .B(net53),
    .COUT(_261_),
    .SUM(_262_));
 sky130_fd_sc_hd__ha_1 _610_ (.A(net20),
    .B(net52),
    .COUT(_263_),
    .SUM(_264_));
 sky130_fd_sc_hd__ha_1 _611_ (.A(net19),
    .B(net51),
    .COUT(_265_),
    .SUM(_266_));
 sky130_fd_sc_hd__ha_2 _612_ (.A(net18),
    .B(net50),
    .COUT(_267_),
    .SUM(_268_));
 sky130_fd_sc_hd__ha_1 _613_ (.A(net17),
    .B(net49),
    .COUT(_269_),
    .SUM(_270_));
 sky130_fd_sc_hd__ha_1 _614_ (.A(net16),
    .B(net48),
    .COUT(_271_),
    .SUM(_272_));
 sky130_fd_sc_hd__ha_1 _615_ (.A(net15),
    .B(net47),
    .COUT(_273_),
    .SUM(_274_));
 sky130_fd_sc_hd__ha_1 _616_ (.A(net14),
    .B(net46),
    .COUT(_275_),
    .SUM(_276_));
 sky130_fd_sc_hd__ha_2 _617_ (.A(net13),
    .B(net45),
    .COUT(_277_),
    .SUM(_278_));
 sky130_fd_sc_hd__ha_1 _618_ (.A(net11),
    .B(net43),
    .COUT(_279_),
    .SUM(_280_));
 sky130_fd_sc_hd__ha_1 _619_ (.A(net10),
    .B(net42),
    .COUT(_281_),
    .SUM(_282_));
 sky130_fd_sc_hd__ha_2 _620_ (.A(net9),
    .B(net41),
    .COUT(_283_),
    .SUM(_284_));
 sky130_fd_sc_hd__ha_1 _621_ (.A(net8),
    .B(net40),
    .COUT(_285_),
    .SUM(_286_));
 sky130_fd_sc_hd__ha_1 _622_ (.A(net7),
    .B(net39),
    .COUT(_287_),
    .SUM(_288_));
 sky130_fd_sc_hd__ha_1 _623_ (.A(net6),
    .B(net38),
    .COUT(_289_),
    .SUM(_290_));
 sky130_fd_sc_hd__ha_2 _624_ (.A(net5),
    .B(net37),
    .COUT(_291_),
    .SUM(_292_));
 sky130_fd_sc_hd__ha_1 _625_ (.A(net4),
    .B(net36),
    .COUT(_293_),
    .SUM(_294_));
 sky130_fd_sc_hd__ha_2 _626_ (.A(net3),
    .B(net35),
    .COUT(_295_),
    .SUM(_296_));
 sky130_fd_sc_hd__ha_1 _627_ (.A(net2),
    .B(net34),
    .COUT(_297_),
    .SUM(_298_));
 sky130_fd_sc_hd__ha_1 _628_ (.A(net32),
    .B(net64),
    .COUT(_299_),
    .SUM(_300_));
 sky130_fd_sc_hd__ha_2 _629_ (.A(net31),
    .B(net63),
    .COUT(_301_),
    .SUM(_302_));
 sky130_fd_sc_hd__ha_1 _630_ (.A(net30),
    .B(net62),
    .COUT(_303_),
    .SUM(_304_));
 sky130_fd_sc_hd__ha_2 _631_ (.A(net29),
    .B(net61),
    .COUT(_305_),
    .SUM(_306_));
 sky130_fd_sc_hd__ha_1 _632_ (.A(net28),
    .B(net60),
    .COUT(_307_),
    .SUM(_308_));
 sky130_fd_sc_hd__ha_1 _633_ (.A(net27),
    .B(net59),
    .COUT(_309_),
    .SUM(_310_));
 sky130_fd_sc_hd__ha_1 _634_ (.A(net26),
    .B(net58),
    .COUT(_311_),
    .SUM(_312_));
 sky130_fd_sc_hd__ha_1 _635_ (.A(net23),
    .B(net55),
    .COUT(_313_),
    .SUM(_314_));
 sky130_fd_sc_hd__ha_1 _636_ (.A(net12),
    .B(net44),
    .COUT(_315_),
    .SUM(_316_));
 sky130_fd_sc_hd__ha_1 _637_ (.A(net1),
    .B(net33),
    .COUT(_317_),
    .SUM(_318_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_47 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(a[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(a[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(a[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(a[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(a[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(a[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(a[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(a[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(a[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(a[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(a[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(a[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(a[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(a[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(a[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(a[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(a[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(a[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(a[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(a[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(a[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(a[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(a[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(a[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(a[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(a[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(a[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(a[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(a[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(a[8]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(a[9]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(b[0]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(b[10]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(b[11]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(b[12]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(b[13]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(b[14]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(b[15]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(b[16]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(b[17]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(b[18]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(b[19]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(b[1]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(b[20]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(b[21]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(b[22]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(b[23]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(b[24]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(b[25]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(b[26]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(b[27]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(b[28]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(b[29]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(b[2]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(b[30]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(b[31]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(b[3]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(b[4]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(b[5]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(b[6]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(b[7]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(b[8]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(b[9]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(cin),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 output66 (.A(net66),
    .X(cout));
 sky130_fd_sc_hd__clkbuf_1 output67 (.A(net67),
    .X(sum[0]));
 sky130_fd_sc_hd__clkbuf_1 output68 (.A(net68),
    .X(sum[10]));
 sky130_fd_sc_hd__clkbuf_1 output69 (.A(net69),
    .X(sum[11]));
 sky130_fd_sc_hd__clkbuf_1 output70 (.A(net70),
    .X(sum[12]));
 sky130_fd_sc_hd__clkbuf_1 output71 (.A(net71),
    .X(sum[13]));
 sky130_fd_sc_hd__clkbuf_1 output72 (.A(net72),
    .X(sum[14]));
 sky130_fd_sc_hd__clkbuf_1 output73 (.A(net73),
    .X(sum[15]));
 sky130_fd_sc_hd__clkbuf_1 output74 (.A(net74),
    .X(sum[16]));
 sky130_fd_sc_hd__clkbuf_1 output75 (.A(net75),
    .X(sum[17]));
 sky130_fd_sc_hd__clkbuf_1 output76 (.A(net76),
    .X(sum[18]));
 sky130_fd_sc_hd__clkbuf_1 output77 (.A(net77),
    .X(sum[19]));
 sky130_fd_sc_hd__clkbuf_1 output78 (.A(net78),
    .X(sum[1]));
 sky130_fd_sc_hd__clkbuf_1 output79 (.A(net79),
    .X(sum[20]));
 sky130_fd_sc_hd__clkbuf_1 output80 (.A(net80),
    .X(sum[21]));
 sky130_fd_sc_hd__clkbuf_1 output81 (.A(net81),
    .X(sum[22]));
 sky130_fd_sc_hd__clkbuf_1 output82 (.A(net82),
    .X(sum[23]));
 sky130_fd_sc_hd__clkbuf_1 output83 (.A(net83),
    .X(sum[24]));
 sky130_fd_sc_hd__clkbuf_1 output84 (.A(net84),
    .X(sum[25]));
 sky130_fd_sc_hd__clkbuf_1 output85 (.A(net85),
    .X(sum[26]));
 sky130_fd_sc_hd__clkbuf_1 output86 (.A(net86),
    .X(sum[27]));
 sky130_fd_sc_hd__clkbuf_1 output87 (.A(net87),
    .X(sum[28]));
 sky130_fd_sc_hd__clkbuf_1 output88 (.A(net88),
    .X(sum[29]));
 sky130_fd_sc_hd__clkbuf_1 output89 (.A(net89),
    .X(sum[2]));
 sky130_fd_sc_hd__clkbuf_1 output90 (.A(net90),
    .X(sum[30]));
 sky130_fd_sc_hd__clkbuf_1 output91 (.A(net91),
    .X(sum[31]));
 sky130_fd_sc_hd__clkbuf_1 output92 (.A(net92),
    .X(sum[3]));
 sky130_fd_sc_hd__clkbuf_1 output93 (.A(net93),
    .X(sum[4]));
 sky130_fd_sc_hd__clkbuf_1 output94 (.A(net94),
    .X(sum[5]));
 sky130_fd_sc_hd__clkbuf_1 output95 (.A(net95),
    .X(sum[6]));
 sky130_fd_sc_hd__clkbuf_1 output96 (.A(net96),
    .X(sum[7]));
 sky130_fd_sc_hd__clkbuf_1 output97 (.A(net97),
    .X(sum[8]));
 sky130_fd_sc_hd__clkbuf_1 output98 (.A(net98),
    .X(sum[9]));
 sky130_fd_sc_hd__fill_1 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_30 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_36 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_11 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_25 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_84 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_35 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_23 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_53 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_9 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_11 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_131 ();
endmodule
