module riscv (clk,
    memread,
    memwrite,
    reset,
    suspend,
    aluout,
    instr,
    pc,
    readdata,
    writedata);
 input clk;
 output memread;
 output memwrite;
 input reset;
 output suspend;
 output [31:0] aluout;
 input [31:0] instr;
 output [31:0] pc;
 input [31:0] readdata;
 output [31:0] writedata;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire clknet_leaf_40_clk;
 wire _0035_;
 wire _0036_;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_37_clk;
 wire _0040_;
 wire clknet_leaf_36_clk;
 wire _0042_;
 wire clknet_leaf_35_clk;
 wire _0044_;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_24_clk;
 wire _0056_;
 wire _0057_;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_22_clk;
 wire _0060_;
 wire _0061_;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_20_clk;
 wire _0064_;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_16_clk;
 wire _0069_;
 wire _0070_;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_14_clk;
 wire _0073_;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_10_clk;
 wire _0077_;
 wire clknet_leaf_9_clk;
 wire _0079_;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_5_clk;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire clknet_leaf_4_clk;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire clknet_leaf_3_clk;
 wire _0094_;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_1_clk;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire net192;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire net191;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire net190;
 wire net189;
 wire net188;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire net187;
 wire _0134_;
 wire _0135_;
 wire net186;
 wire _0137_;
 wire net185;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire net184;
 wire net183;
 wire _0146_;
 wire net182;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire net181;
 wire net180;
 wire _0154_;
 wire net179;
 wire net178;
 wire _0157_;
 wire _0158_;
 wire net702;
 wire net813;
 wire net739;
 wire net172;
 wire net173;
 wire net822;
 wire _0165_;
 wire _0166_;
 wire net815;
 wire net166;
 wire net809;
 wire net821;
 wire net803;
 wire _0172_;
 wire _0173_;
 wire net801;
 wire net799;
 wire net798;
 wire net806;
 wire net794;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire net791;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire net786;
 wire net785;
 wire net783;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire net789;
 wire net773;
 wire net774;
 wire net816;
 wire net825;
 wire net814;
 wire _0200_;
 wire _0201_;
 wire net772;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire net768;
 wire _0207_;
 wire _0208_;
 wire net765;
 wire net764;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire net777;
 wire net742;
 wire _0216_;
 wire _0217_;
 wire net697;
 wire net741;
 wire net749;
 wire _0221_;
 wire _0222_;
 wire net770;
 wire _0224_;
 wire net817;
 wire net716;
 wire net717;
 wire net823;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire net754;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire net758;
 wire net808;
 wire net810;
 wire net760;
 wire net782;
 wire _0244_;
 wire net780;
 wire net793;
 wire net775;
 wire _0248_;
 wire _0249_;
 wire net761;
 wire net763;
 wire net767;
 wire net820;
 wire _0254_;
 wire _0255_;
 wire net756;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire net252;
 wire net752;
 wire net753;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire net750;
 wire net743;
 wire net751;
 wire net224;
 wire net788;
 wire _0271_;
 wire net781;
 wire net748;
 wire net740;
 wire _0275_;
 wire net737;
 wire net736;
 wire net735;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire net734;
 wire net733;
 wire _0284_;
 wire net732;
 wire net731;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire net730;
 wire net729;
 wire _0296_;
 wire net728;
 wire _0298_;
 wire net727;
 wire net726;
 wire _0301_;
 wire net725;
 wire _0303_;
 wire _0304_;
 wire net724;
 wire net723;
 wire _0307_;
 wire net722;
 wire net721;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire net719;
 wire net718;
 wire net744;
 wire net745;
 wire net715;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire net714;
 wire net713;
 wire net712;
 wire _0327_;
 wire net711;
 wire net710;
 wire net746;
 wire net709;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire net701;
 wire net703;
 wire net700;
 wire net698;
 wire net771;
 wire net708;
 wire _0347_;
 wire net705;
 wire _0349_;
 wire net797;
 wire _0351_;
 wire net175;
 wire net325;
 wire _0354_;
 wire net769;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire net755;
 wire net177;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire net695;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire net694;
 wire _0373_;
 wire net174;
 wire net169;
 wire _0376_;
 wire net819;
 wire net699;
 wire _0379_;
 wire _0380_;
 wire net165;
 wire net738;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire net696;
 wire net706;
 wire net818;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire net707;
 wire net812;
 wire net807;
 wire _0399_;
 wire _0400_;
 wire net747;
 wire _0402_;
 wire _0403_;
 wire net170;
 wire net824;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire net167;
 wire net168;
 wire _0415_;
 wire _0416_;
 wire net176;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire net757;
 wire net171;
 wire _0425_;
 wire net811;
 wire net826;
 wire _0428_;
 wire net802;
 wire net800;
 wire _0431_;
 wire net805;
 wire _0433_;
 wire net796;
 wire net759;
 wire _0436_;
 wire _0437_;
 wire net795;
 wire _0439_;
 wire net790;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire net784;
 wire _0451_;
 wire _0452_;
 wire net787;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire net792;
 wire net778;
 wire _0459_;
 wire _0460_;
 wire net776;
 wire net766;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0485_;
 wire _0486_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0553_;
 wire _0554_;
 wire _0556_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0581_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0590_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0765_;
 wire _0768_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1718_;
 wire _1719_;
 wire _1721_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1803_;
 wire _1805_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1813_;
 wire _1816_;
 wire _1817_;
 wire _1820_;
 wire _1821_;
 wire _1824_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1834_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1840_;
 wire _1841_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire net65;
 wire _1859_;
 wire net64;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire net63;
 wire net62;
 wire net61;
 wire _1867_;
 wire net60;
 wire _1869_;
 wire _1870_;
 wire net59;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire net58;
 wire net57;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire net56;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire net55;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire net54;
 wire _1902_;
 wire _1903_;
 wire net53;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire net52;
 wire _1914_;
 wire net51;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire net50;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire net49;
 wire net48;
 wire net47;
 wire _1928_;
 wire _1929_;
 wire net46;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire net45;
 wire _1949_;
 wire net44;
 wire _1951_;
 wire _1952_;
 wire net43;
 wire _1954_;
 wire _1955_;
 wire net42;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire net41;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire net40;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire net39;
 wire net38;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire net37;
 wire net36;
 wire net35;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire net34;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire net33;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire net32;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire net31;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire net30;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire net29;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire net28;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire net27;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire net26;
 wire _2627_;
 wire net25;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire net24;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire net23;
 wire _2648_;
 wire net22;
 wire net21;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire net20;
 wire _2661_;
 wire net19;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire net18;
 wire _2673_;
 wire net17;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire net16;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire net15;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire net14;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire net13;
 wire net12;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire net11;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire net10;
 wire net9;
 wire _3074_;
 wire net8;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire net7;
 wire _3090_;
 wire net6;
 wire net5;
 wire _3093_;
 wire net4;
 wire _3095_;
 wire net3;
 wire _3097_;
 wire net2;
 wire net1;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3179_;
 wire _3180_;
 wire _3182_;
 wire _3183_;
 wire net804;
 wire net720;
 wire clknet_leaf_0_clk;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire \dp.ISRmux.d0[10] ;
 wire \dp.ISRmux.d0[11] ;
 wire \dp.ISRmux.d0[12] ;
 wire \dp.ISRmux.d0[13] ;
 wire \dp.ISRmux.d0[14] ;
 wire \dp.ISRmux.d0[15] ;
 wire \dp.ISRmux.d0[16] ;
 wire \dp.ISRmux.d0[17] ;
 wire \dp.ISRmux.d0[18] ;
 wire \dp.ISRmux.d0[19] ;
 wire \dp.ISRmux.d0[20] ;
 wire \dp.ISRmux.d0[21] ;
 wire \dp.ISRmux.d0[22] ;
 wire \dp.ISRmux.d0[23] ;
 wire \dp.ISRmux.d0[24] ;
 wire \dp.ISRmux.d0[25] ;
 wire \dp.ISRmux.d0[26] ;
 wire \dp.ISRmux.d0[27] ;
 wire \dp.ISRmux.d0[28] ;
 wire \dp.ISRmux.d0[29] ;
 wire \dp.ISRmux.d0[2] ;
 wire \dp.ISRmux.d0[30] ;
 wire \dp.ISRmux.d0[31] ;
 wire \dp.ISRmux.d0[3] ;
 wire \dp.ISRmux.d0[4] ;
 wire \dp.ISRmux.d0[5] ;
 wire \dp.ISRmux.d0[6] ;
 wire \dp.ISRmux.d0[7] ;
 wire \dp.ISRmux.d0[8] ;
 wire \dp.ISRmux.d0[9] ;
 wire \dp.result2[0] ;
 wire \dp.result2[10] ;
 wire \dp.result2[11] ;
 wire \dp.result2[12] ;
 wire \dp.result2[13] ;
 wire \dp.result2[14] ;
 wire \dp.result2[15] ;
 wire \dp.result2[16] ;
 wire \dp.result2[17] ;
 wire \dp.result2[18] ;
 wire \dp.result2[19] ;
 wire \dp.result2[1] ;
 wire \dp.result2[20] ;
 wire \dp.result2[21] ;
 wire \dp.result2[22] ;
 wire \dp.result2[23] ;
 wire \dp.result2[24] ;
 wire \dp.result2[25] ;
 wire \dp.result2[26] ;
 wire \dp.result2[27] ;
 wire \dp.result2[28] ;
 wire \dp.result2[29] ;
 wire \dp.result2[2] ;
 wire \dp.result2[30] ;
 wire \dp.result2[31] ;
 wire \dp.result2[3] ;
 wire \dp.result2[4] ;
 wire \dp.result2[5] ;
 wire \dp.result2[6] ;
 wire \dp.result2[7] ;
 wire \dp.result2[8] ;
 wire \dp.result2[9] ;
 wire \dp.rf.rf[0][0] ;
 wire \dp.rf.rf[0][10] ;
 wire \dp.rf.rf[0][11] ;
 wire \dp.rf.rf[0][12] ;
 wire \dp.rf.rf[0][13] ;
 wire \dp.rf.rf[0][14] ;
 wire \dp.rf.rf[0][15] ;
 wire \dp.rf.rf[0][17] ;
 wire \dp.rf.rf[0][18] ;
 wire \dp.rf.rf[0][19] ;
 wire \dp.rf.rf[0][1] ;
 wire \dp.rf.rf[0][21] ;
 wire \dp.rf.rf[0][22] ;
 wire \dp.rf.rf[0][23] ;
 wire \dp.rf.rf[0][24] ;
 wire \dp.rf.rf[0][25] ;
 wire \dp.rf.rf[0][27] ;
 wire \dp.rf.rf[0][28] ;
 wire \dp.rf.rf[0][29] ;
 wire \dp.rf.rf[0][30] ;
 wire \dp.rf.rf[0][31] ;
 wire \dp.rf.rf[0][3] ;
 wire \dp.rf.rf[0][4] ;
 wire \dp.rf.rf[0][5] ;
 wire \dp.rf.rf[0][6] ;
 wire \dp.rf.rf[0][7] ;
 wire \dp.rf.rf[0][8] ;
 wire \dp.rf.rf[0][9] ;
 wire \dp.rf.rf[10][0] ;
 wire \dp.rf.rf[10][10] ;
 wire \dp.rf.rf[10][11] ;
 wire \dp.rf.rf[10][12] ;
 wire \dp.rf.rf[10][13] ;
 wire \dp.rf.rf[10][14] ;
 wire \dp.rf.rf[10][15] ;
 wire \dp.rf.rf[10][16] ;
 wire \dp.rf.rf[10][17] ;
 wire \dp.rf.rf[10][18] ;
 wire \dp.rf.rf[10][19] ;
 wire \dp.rf.rf[10][1] ;
 wire \dp.rf.rf[10][20] ;
 wire \dp.rf.rf[10][21] ;
 wire \dp.rf.rf[10][22] ;
 wire \dp.rf.rf[10][23] ;
 wire \dp.rf.rf[10][24] ;
 wire \dp.rf.rf[10][25] ;
 wire \dp.rf.rf[10][26] ;
 wire \dp.rf.rf[10][27] ;
 wire \dp.rf.rf[10][28] ;
 wire \dp.rf.rf[10][29] ;
 wire \dp.rf.rf[10][2] ;
 wire \dp.rf.rf[10][30] ;
 wire \dp.rf.rf[10][31] ;
 wire \dp.rf.rf[10][3] ;
 wire \dp.rf.rf[10][4] ;
 wire \dp.rf.rf[10][5] ;
 wire \dp.rf.rf[10][6] ;
 wire \dp.rf.rf[10][7] ;
 wire \dp.rf.rf[10][8] ;
 wire \dp.rf.rf[10][9] ;
 wire \dp.rf.rf[11][0] ;
 wire \dp.rf.rf[11][10] ;
 wire \dp.rf.rf[11][11] ;
 wire \dp.rf.rf[11][12] ;
 wire \dp.rf.rf[11][13] ;
 wire \dp.rf.rf[11][14] ;
 wire \dp.rf.rf[11][15] ;
 wire \dp.rf.rf[11][16] ;
 wire \dp.rf.rf[11][17] ;
 wire \dp.rf.rf[11][18] ;
 wire \dp.rf.rf[11][19] ;
 wire \dp.rf.rf[11][1] ;
 wire \dp.rf.rf[11][20] ;
 wire \dp.rf.rf[11][21] ;
 wire \dp.rf.rf[11][22] ;
 wire \dp.rf.rf[11][23] ;
 wire \dp.rf.rf[11][24] ;
 wire \dp.rf.rf[11][25] ;
 wire \dp.rf.rf[11][26] ;
 wire \dp.rf.rf[11][27] ;
 wire \dp.rf.rf[11][28] ;
 wire \dp.rf.rf[11][29] ;
 wire \dp.rf.rf[11][2] ;
 wire \dp.rf.rf[11][30] ;
 wire \dp.rf.rf[11][31] ;
 wire \dp.rf.rf[11][3] ;
 wire \dp.rf.rf[11][4] ;
 wire \dp.rf.rf[11][5] ;
 wire \dp.rf.rf[11][6] ;
 wire \dp.rf.rf[11][7] ;
 wire \dp.rf.rf[11][8] ;
 wire \dp.rf.rf[11][9] ;
 wire \dp.rf.rf[12][0] ;
 wire \dp.rf.rf[12][10] ;
 wire \dp.rf.rf[12][11] ;
 wire \dp.rf.rf[12][12] ;
 wire \dp.rf.rf[12][13] ;
 wire \dp.rf.rf[12][14] ;
 wire \dp.rf.rf[12][15] ;
 wire \dp.rf.rf[12][16] ;
 wire \dp.rf.rf[12][17] ;
 wire \dp.rf.rf[12][18] ;
 wire \dp.rf.rf[12][19] ;
 wire \dp.rf.rf[12][1] ;
 wire \dp.rf.rf[12][20] ;
 wire \dp.rf.rf[12][21] ;
 wire \dp.rf.rf[12][22] ;
 wire \dp.rf.rf[12][23] ;
 wire \dp.rf.rf[12][24] ;
 wire \dp.rf.rf[12][25] ;
 wire \dp.rf.rf[12][26] ;
 wire \dp.rf.rf[12][27] ;
 wire \dp.rf.rf[12][28] ;
 wire \dp.rf.rf[12][29] ;
 wire \dp.rf.rf[12][2] ;
 wire \dp.rf.rf[12][30] ;
 wire \dp.rf.rf[12][31] ;
 wire \dp.rf.rf[12][3] ;
 wire \dp.rf.rf[12][4] ;
 wire \dp.rf.rf[12][5] ;
 wire \dp.rf.rf[12][6] ;
 wire \dp.rf.rf[12][7] ;
 wire \dp.rf.rf[12][8] ;
 wire \dp.rf.rf[12][9] ;
 wire \dp.rf.rf[13][0] ;
 wire \dp.rf.rf[13][10] ;
 wire \dp.rf.rf[13][11] ;
 wire \dp.rf.rf[13][12] ;
 wire \dp.rf.rf[13][13] ;
 wire \dp.rf.rf[13][14] ;
 wire \dp.rf.rf[13][15] ;
 wire \dp.rf.rf[13][16] ;
 wire \dp.rf.rf[13][17] ;
 wire \dp.rf.rf[13][18] ;
 wire \dp.rf.rf[13][19] ;
 wire \dp.rf.rf[13][1] ;
 wire \dp.rf.rf[13][20] ;
 wire \dp.rf.rf[13][21] ;
 wire \dp.rf.rf[13][22] ;
 wire \dp.rf.rf[13][23] ;
 wire \dp.rf.rf[13][24] ;
 wire \dp.rf.rf[13][25] ;
 wire \dp.rf.rf[13][26] ;
 wire \dp.rf.rf[13][27] ;
 wire \dp.rf.rf[13][28] ;
 wire \dp.rf.rf[13][29] ;
 wire \dp.rf.rf[13][2] ;
 wire \dp.rf.rf[13][30] ;
 wire \dp.rf.rf[13][31] ;
 wire \dp.rf.rf[13][3] ;
 wire \dp.rf.rf[13][4] ;
 wire \dp.rf.rf[13][5] ;
 wire \dp.rf.rf[13][6] ;
 wire \dp.rf.rf[13][7] ;
 wire \dp.rf.rf[13][8] ;
 wire \dp.rf.rf[13][9] ;
 wire \dp.rf.rf[14][0] ;
 wire \dp.rf.rf[14][10] ;
 wire \dp.rf.rf[14][11] ;
 wire \dp.rf.rf[14][12] ;
 wire \dp.rf.rf[14][13] ;
 wire \dp.rf.rf[14][14] ;
 wire \dp.rf.rf[14][15] ;
 wire \dp.rf.rf[14][16] ;
 wire \dp.rf.rf[14][17] ;
 wire \dp.rf.rf[14][18] ;
 wire \dp.rf.rf[14][19] ;
 wire \dp.rf.rf[14][1] ;
 wire \dp.rf.rf[14][20] ;
 wire \dp.rf.rf[14][21] ;
 wire \dp.rf.rf[14][22] ;
 wire \dp.rf.rf[14][23] ;
 wire \dp.rf.rf[14][24] ;
 wire \dp.rf.rf[14][25] ;
 wire \dp.rf.rf[14][26] ;
 wire \dp.rf.rf[14][27] ;
 wire \dp.rf.rf[14][28] ;
 wire \dp.rf.rf[14][29] ;
 wire \dp.rf.rf[14][2] ;
 wire \dp.rf.rf[14][30] ;
 wire \dp.rf.rf[14][31] ;
 wire \dp.rf.rf[14][3] ;
 wire \dp.rf.rf[14][4] ;
 wire \dp.rf.rf[14][5] ;
 wire \dp.rf.rf[14][6] ;
 wire \dp.rf.rf[14][7] ;
 wire \dp.rf.rf[14][8] ;
 wire \dp.rf.rf[14][9] ;
 wire \dp.rf.rf[15][0] ;
 wire \dp.rf.rf[15][10] ;
 wire \dp.rf.rf[15][11] ;
 wire \dp.rf.rf[15][12] ;
 wire \dp.rf.rf[15][13] ;
 wire \dp.rf.rf[15][14] ;
 wire \dp.rf.rf[15][15] ;
 wire \dp.rf.rf[15][16] ;
 wire \dp.rf.rf[15][17] ;
 wire \dp.rf.rf[15][18] ;
 wire \dp.rf.rf[15][19] ;
 wire \dp.rf.rf[15][1] ;
 wire \dp.rf.rf[15][20] ;
 wire \dp.rf.rf[15][21] ;
 wire \dp.rf.rf[15][22] ;
 wire \dp.rf.rf[15][23] ;
 wire \dp.rf.rf[15][24] ;
 wire \dp.rf.rf[15][25] ;
 wire \dp.rf.rf[15][26] ;
 wire \dp.rf.rf[15][27] ;
 wire \dp.rf.rf[15][28] ;
 wire \dp.rf.rf[15][29] ;
 wire \dp.rf.rf[15][2] ;
 wire \dp.rf.rf[15][30] ;
 wire \dp.rf.rf[15][31] ;
 wire \dp.rf.rf[15][3] ;
 wire \dp.rf.rf[15][4] ;
 wire \dp.rf.rf[15][5] ;
 wire \dp.rf.rf[15][6] ;
 wire \dp.rf.rf[15][7] ;
 wire \dp.rf.rf[15][8] ;
 wire \dp.rf.rf[15][9] ;
 wire \dp.rf.rf[16][0] ;
 wire \dp.rf.rf[16][10] ;
 wire \dp.rf.rf[16][11] ;
 wire \dp.rf.rf[16][12] ;
 wire \dp.rf.rf[16][13] ;
 wire \dp.rf.rf[16][14] ;
 wire \dp.rf.rf[16][15] ;
 wire \dp.rf.rf[16][16] ;
 wire \dp.rf.rf[16][17] ;
 wire \dp.rf.rf[16][18] ;
 wire \dp.rf.rf[16][19] ;
 wire \dp.rf.rf[16][1] ;
 wire \dp.rf.rf[16][20] ;
 wire \dp.rf.rf[16][21] ;
 wire \dp.rf.rf[16][22] ;
 wire \dp.rf.rf[16][23] ;
 wire \dp.rf.rf[16][24] ;
 wire \dp.rf.rf[16][25] ;
 wire \dp.rf.rf[16][26] ;
 wire \dp.rf.rf[16][27] ;
 wire \dp.rf.rf[16][28] ;
 wire \dp.rf.rf[16][29] ;
 wire \dp.rf.rf[16][2] ;
 wire \dp.rf.rf[16][30] ;
 wire \dp.rf.rf[16][31] ;
 wire \dp.rf.rf[16][3] ;
 wire \dp.rf.rf[16][4] ;
 wire \dp.rf.rf[16][5] ;
 wire \dp.rf.rf[16][6] ;
 wire \dp.rf.rf[16][7] ;
 wire \dp.rf.rf[16][8] ;
 wire \dp.rf.rf[16][9] ;
 wire \dp.rf.rf[17][0] ;
 wire \dp.rf.rf[17][10] ;
 wire \dp.rf.rf[17][11] ;
 wire \dp.rf.rf[17][12] ;
 wire \dp.rf.rf[17][13] ;
 wire \dp.rf.rf[17][14] ;
 wire \dp.rf.rf[17][15] ;
 wire \dp.rf.rf[17][16] ;
 wire \dp.rf.rf[17][17] ;
 wire \dp.rf.rf[17][18] ;
 wire \dp.rf.rf[17][19] ;
 wire \dp.rf.rf[17][1] ;
 wire \dp.rf.rf[17][20] ;
 wire \dp.rf.rf[17][21] ;
 wire \dp.rf.rf[17][22] ;
 wire \dp.rf.rf[17][23] ;
 wire \dp.rf.rf[17][24] ;
 wire \dp.rf.rf[17][25] ;
 wire \dp.rf.rf[17][26] ;
 wire \dp.rf.rf[17][27] ;
 wire \dp.rf.rf[17][28] ;
 wire \dp.rf.rf[17][29] ;
 wire \dp.rf.rf[17][2] ;
 wire \dp.rf.rf[17][30] ;
 wire \dp.rf.rf[17][31] ;
 wire \dp.rf.rf[17][3] ;
 wire \dp.rf.rf[17][4] ;
 wire \dp.rf.rf[17][5] ;
 wire \dp.rf.rf[17][6] ;
 wire \dp.rf.rf[17][7] ;
 wire \dp.rf.rf[17][8] ;
 wire \dp.rf.rf[17][9] ;
 wire \dp.rf.rf[18][0] ;
 wire \dp.rf.rf[18][10] ;
 wire \dp.rf.rf[18][11] ;
 wire \dp.rf.rf[18][12] ;
 wire \dp.rf.rf[18][13] ;
 wire \dp.rf.rf[18][14] ;
 wire \dp.rf.rf[18][15] ;
 wire \dp.rf.rf[18][16] ;
 wire \dp.rf.rf[18][17] ;
 wire \dp.rf.rf[18][18] ;
 wire \dp.rf.rf[18][19] ;
 wire \dp.rf.rf[18][1] ;
 wire \dp.rf.rf[18][20] ;
 wire \dp.rf.rf[18][21] ;
 wire \dp.rf.rf[18][22] ;
 wire \dp.rf.rf[18][23] ;
 wire \dp.rf.rf[18][24] ;
 wire \dp.rf.rf[18][25] ;
 wire \dp.rf.rf[18][26] ;
 wire \dp.rf.rf[18][27] ;
 wire \dp.rf.rf[18][28] ;
 wire \dp.rf.rf[18][29] ;
 wire \dp.rf.rf[18][2] ;
 wire \dp.rf.rf[18][30] ;
 wire \dp.rf.rf[18][31] ;
 wire \dp.rf.rf[18][3] ;
 wire \dp.rf.rf[18][4] ;
 wire \dp.rf.rf[18][5] ;
 wire \dp.rf.rf[18][6] ;
 wire \dp.rf.rf[18][7] ;
 wire \dp.rf.rf[18][8] ;
 wire \dp.rf.rf[18][9] ;
 wire \dp.rf.rf[19][0] ;
 wire \dp.rf.rf[19][10] ;
 wire \dp.rf.rf[19][11] ;
 wire \dp.rf.rf[19][12] ;
 wire \dp.rf.rf[19][13] ;
 wire \dp.rf.rf[19][14] ;
 wire \dp.rf.rf[19][15] ;
 wire \dp.rf.rf[19][16] ;
 wire \dp.rf.rf[19][17] ;
 wire \dp.rf.rf[19][18] ;
 wire \dp.rf.rf[19][19] ;
 wire \dp.rf.rf[19][1] ;
 wire \dp.rf.rf[19][20] ;
 wire \dp.rf.rf[19][21] ;
 wire \dp.rf.rf[19][22] ;
 wire \dp.rf.rf[19][23] ;
 wire \dp.rf.rf[19][24] ;
 wire \dp.rf.rf[19][25] ;
 wire \dp.rf.rf[19][26] ;
 wire \dp.rf.rf[19][27] ;
 wire \dp.rf.rf[19][28] ;
 wire \dp.rf.rf[19][29] ;
 wire \dp.rf.rf[19][2] ;
 wire \dp.rf.rf[19][30] ;
 wire \dp.rf.rf[19][31] ;
 wire \dp.rf.rf[19][3] ;
 wire \dp.rf.rf[19][4] ;
 wire \dp.rf.rf[19][5] ;
 wire \dp.rf.rf[19][6] ;
 wire \dp.rf.rf[19][7] ;
 wire \dp.rf.rf[19][8] ;
 wire \dp.rf.rf[19][9] ;
 wire \dp.rf.rf[1][0] ;
 wire \dp.rf.rf[1][10] ;
 wire \dp.rf.rf[1][11] ;
 wire \dp.rf.rf[1][12] ;
 wire \dp.rf.rf[1][13] ;
 wire \dp.rf.rf[1][14] ;
 wire \dp.rf.rf[1][15] ;
 wire \dp.rf.rf[1][16] ;
 wire \dp.rf.rf[1][17] ;
 wire \dp.rf.rf[1][18] ;
 wire \dp.rf.rf[1][19] ;
 wire \dp.rf.rf[1][1] ;
 wire \dp.rf.rf[1][20] ;
 wire \dp.rf.rf[1][21] ;
 wire \dp.rf.rf[1][22] ;
 wire \dp.rf.rf[1][23] ;
 wire \dp.rf.rf[1][24] ;
 wire \dp.rf.rf[1][25] ;
 wire \dp.rf.rf[1][26] ;
 wire \dp.rf.rf[1][27] ;
 wire \dp.rf.rf[1][28] ;
 wire \dp.rf.rf[1][29] ;
 wire \dp.rf.rf[1][2] ;
 wire \dp.rf.rf[1][30] ;
 wire \dp.rf.rf[1][31] ;
 wire \dp.rf.rf[1][3] ;
 wire \dp.rf.rf[1][4] ;
 wire \dp.rf.rf[1][5] ;
 wire \dp.rf.rf[1][6] ;
 wire \dp.rf.rf[1][7] ;
 wire \dp.rf.rf[1][8] ;
 wire \dp.rf.rf[1][9] ;
 wire \dp.rf.rf[20][0] ;
 wire \dp.rf.rf[20][10] ;
 wire \dp.rf.rf[20][11] ;
 wire \dp.rf.rf[20][12] ;
 wire \dp.rf.rf[20][13] ;
 wire \dp.rf.rf[20][14] ;
 wire \dp.rf.rf[20][15] ;
 wire \dp.rf.rf[20][16] ;
 wire \dp.rf.rf[20][17] ;
 wire \dp.rf.rf[20][18] ;
 wire \dp.rf.rf[20][19] ;
 wire \dp.rf.rf[20][1] ;
 wire \dp.rf.rf[20][20] ;
 wire \dp.rf.rf[20][21] ;
 wire \dp.rf.rf[20][22] ;
 wire \dp.rf.rf[20][23] ;
 wire \dp.rf.rf[20][24] ;
 wire \dp.rf.rf[20][25] ;
 wire \dp.rf.rf[20][26] ;
 wire \dp.rf.rf[20][27] ;
 wire \dp.rf.rf[20][28] ;
 wire \dp.rf.rf[20][29] ;
 wire \dp.rf.rf[20][2] ;
 wire \dp.rf.rf[20][30] ;
 wire \dp.rf.rf[20][31] ;
 wire \dp.rf.rf[20][3] ;
 wire \dp.rf.rf[20][4] ;
 wire \dp.rf.rf[20][5] ;
 wire \dp.rf.rf[20][6] ;
 wire \dp.rf.rf[20][7] ;
 wire \dp.rf.rf[20][8] ;
 wire \dp.rf.rf[20][9] ;
 wire \dp.rf.rf[21][0] ;
 wire \dp.rf.rf[21][10] ;
 wire \dp.rf.rf[21][11] ;
 wire \dp.rf.rf[21][12] ;
 wire \dp.rf.rf[21][13] ;
 wire \dp.rf.rf[21][14] ;
 wire \dp.rf.rf[21][15] ;
 wire \dp.rf.rf[21][16] ;
 wire \dp.rf.rf[21][17] ;
 wire \dp.rf.rf[21][18] ;
 wire \dp.rf.rf[21][19] ;
 wire \dp.rf.rf[21][1] ;
 wire \dp.rf.rf[21][20] ;
 wire \dp.rf.rf[21][21] ;
 wire \dp.rf.rf[21][22] ;
 wire \dp.rf.rf[21][23] ;
 wire \dp.rf.rf[21][24] ;
 wire \dp.rf.rf[21][25] ;
 wire \dp.rf.rf[21][26] ;
 wire \dp.rf.rf[21][27] ;
 wire \dp.rf.rf[21][28] ;
 wire \dp.rf.rf[21][29] ;
 wire \dp.rf.rf[21][2] ;
 wire \dp.rf.rf[21][30] ;
 wire \dp.rf.rf[21][31] ;
 wire \dp.rf.rf[21][3] ;
 wire \dp.rf.rf[21][4] ;
 wire \dp.rf.rf[21][5] ;
 wire \dp.rf.rf[21][6] ;
 wire \dp.rf.rf[21][7] ;
 wire \dp.rf.rf[21][8] ;
 wire \dp.rf.rf[21][9] ;
 wire \dp.rf.rf[22][0] ;
 wire \dp.rf.rf[22][10] ;
 wire \dp.rf.rf[22][11] ;
 wire \dp.rf.rf[22][12] ;
 wire \dp.rf.rf[22][13] ;
 wire \dp.rf.rf[22][14] ;
 wire \dp.rf.rf[22][15] ;
 wire \dp.rf.rf[22][16] ;
 wire \dp.rf.rf[22][17] ;
 wire \dp.rf.rf[22][18] ;
 wire \dp.rf.rf[22][19] ;
 wire \dp.rf.rf[22][1] ;
 wire \dp.rf.rf[22][20] ;
 wire \dp.rf.rf[22][21] ;
 wire \dp.rf.rf[22][22] ;
 wire \dp.rf.rf[22][23] ;
 wire \dp.rf.rf[22][24] ;
 wire \dp.rf.rf[22][25] ;
 wire \dp.rf.rf[22][26] ;
 wire \dp.rf.rf[22][27] ;
 wire \dp.rf.rf[22][28] ;
 wire \dp.rf.rf[22][29] ;
 wire \dp.rf.rf[22][2] ;
 wire \dp.rf.rf[22][30] ;
 wire \dp.rf.rf[22][31] ;
 wire \dp.rf.rf[22][3] ;
 wire \dp.rf.rf[22][4] ;
 wire \dp.rf.rf[22][5] ;
 wire \dp.rf.rf[22][6] ;
 wire \dp.rf.rf[22][7] ;
 wire \dp.rf.rf[22][8] ;
 wire \dp.rf.rf[22][9] ;
 wire \dp.rf.rf[23][0] ;
 wire \dp.rf.rf[23][10] ;
 wire \dp.rf.rf[23][11] ;
 wire \dp.rf.rf[23][12] ;
 wire \dp.rf.rf[23][13] ;
 wire \dp.rf.rf[23][14] ;
 wire \dp.rf.rf[23][15] ;
 wire \dp.rf.rf[23][16] ;
 wire \dp.rf.rf[23][17] ;
 wire \dp.rf.rf[23][18] ;
 wire \dp.rf.rf[23][19] ;
 wire \dp.rf.rf[23][1] ;
 wire \dp.rf.rf[23][20] ;
 wire \dp.rf.rf[23][21] ;
 wire \dp.rf.rf[23][22] ;
 wire \dp.rf.rf[23][23] ;
 wire \dp.rf.rf[23][24] ;
 wire \dp.rf.rf[23][25] ;
 wire \dp.rf.rf[23][26] ;
 wire \dp.rf.rf[23][27] ;
 wire \dp.rf.rf[23][28] ;
 wire \dp.rf.rf[23][29] ;
 wire \dp.rf.rf[23][2] ;
 wire \dp.rf.rf[23][30] ;
 wire \dp.rf.rf[23][31] ;
 wire \dp.rf.rf[23][3] ;
 wire \dp.rf.rf[23][4] ;
 wire \dp.rf.rf[23][5] ;
 wire \dp.rf.rf[23][6] ;
 wire \dp.rf.rf[23][7] ;
 wire \dp.rf.rf[23][8] ;
 wire \dp.rf.rf[23][9] ;
 wire \dp.rf.rf[24][0] ;
 wire \dp.rf.rf[24][10] ;
 wire \dp.rf.rf[24][11] ;
 wire \dp.rf.rf[24][12] ;
 wire \dp.rf.rf[24][13] ;
 wire \dp.rf.rf[24][14] ;
 wire \dp.rf.rf[24][15] ;
 wire \dp.rf.rf[24][16] ;
 wire \dp.rf.rf[24][17] ;
 wire \dp.rf.rf[24][18] ;
 wire \dp.rf.rf[24][19] ;
 wire \dp.rf.rf[24][1] ;
 wire \dp.rf.rf[24][20] ;
 wire \dp.rf.rf[24][21] ;
 wire \dp.rf.rf[24][22] ;
 wire \dp.rf.rf[24][23] ;
 wire \dp.rf.rf[24][24] ;
 wire \dp.rf.rf[24][25] ;
 wire \dp.rf.rf[24][26] ;
 wire \dp.rf.rf[24][27] ;
 wire \dp.rf.rf[24][28] ;
 wire \dp.rf.rf[24][29] ;
 wire \dp.rf.rf[24][2] ;
 wire \dp.rf.rf[24][30] ;
 wire \dp.rf.rf[24][31] ;
 wire \dp.rf.rf[24][3] ;
 wire \dp.rf.rf[24][4] ;
 wire \dp.rf.rf[24][5] ;
 wire \dp.rf.rf[24][6] ;
 wire \dp.rf.rf[24][7] ;
 wire \dp.rf.rf[24][8] ;
 wire \dp.rf.rf[24][9] ;
 wire \dp.rf.rf[25][0] ;
 wire \dp.rf.rf[25][10] ;
 wire \dp.rf.rf[25][11] ;
 wire \dp.rf.rf[25][12] ;
 wire \dp.rf.rf[25][13] ;
 wire \dp.rf.rf[25][14] ;
 wire \dp.rf.rf[25][15] ;
 wire \dp.rf.rf[25][16] ;
 wire \dp.rf.rf[25][17] ;
 wire \dp.rf.rf[25][18] ;
 wire \dp.rf.rf[25][19] ;
 wire \dp.rf.rf[25][1] ;
 wire \dp.rf.rf[25][20] ;
 wire \dp.rf.rf[25][21] ;
 wire \dp.rf.rf[25][22] ;
 wire \dp.rf.rf[25][23] ;
 wire \dp.rf.rf[25][24] ;
 wire \dp.rf.rf[25][25] ;
 wire \dp.rf.rf[25][26] ;
 wire \dp.rf.rf[25][27] ;
 wire \dp.rf.rf[25][28] ;
 wire \dp.rf.rf[25][29] ;
 wire \dp.rf.rf[25][2] ;
 wire \dp.rf.rf[25][30] ;
 wire \dp.rf.rf[25][31] ;
 wire \dp.rf.rf[25][3] ;
 wire \dp.rf.rf[25][4] ;
 wire \dp.rf.rf[25][5] ;
 wire \dp.rf.rf[25][6] ;
 wire \dp.rf.rf[25][7] ;
 wire \dp.rf.rf[25][8] ;
 wire \dp.rf.rf[25][9] ;
 wire \dp.rf.rf[26][0] ;
 wire \dp.rf.rf[26][10] ;
 wire \dp.rf.rf[26][11] ;
 wire \dp.rf.rf[26][12] ;
 wire \dp.rf.rf[26][13] ;
 wire \dp.rf.rf[26][14] ;
 wire \dp.rf.rf[26][15] ;
 wire \dp.rf.rf[26][16] ;
 wire \dp.rf.rf[26][17] ;
 wire \dp.rf.rf[26][18] ;
 wire \dp.rf.rf[26][19] ;
 wire \dp.rf.rf[26][1] ;
 wire \dp.rf.rf[26][20] ;
 wire \dp.rf.rf[26][21] ;
 wire \dp.rf.rf[26][22] ;
 wire \dp.rf.rf[26][23] ;
 wire \dp.rf.rf[26][24] ;
 wire \dp.rf.rf[26][25] ;
 wire \dp.rf.rf[26][26] ;
 wire \dp.rf.rf[26][27] ;
 wire \dp.rf.rf[26][28] ;
 wire \dp.rf.rf[26][29] ;
 wire \dp.rf.rf[26][2] ;
 wire \dp.rf.rf[26][30] ;
 wire \dp.rf.rf[26][31] ;
 wire \dp.rf.rf[26][3] ;
 wire \dp.rf.rf[26][4] ;
 wire \dp.rf.rf[26][5] ;
 wire \dp.rf.rf[26][6] ;
 wire \dp.rf.rf[26][7] ;
 wire \dp.rf.rf[26][8] ;
 wire \dp.rf.rf[26][9] ;
 wire \dp.rf.rf[27][0] ;
 wire \dp.rf.rf[27][10] ;
 wire \dp.rf.rf[27][11] ;
 wire \dp.rf.rf[27][12] ;
 wire \dp.rf.rf[27][13] ;
 wire \dp.rf.rf[27][14] ;
 wire \dp.rf.rf[27][15] ;
 wire \dp.rf.rf[27][16] ;
 wire \dp.rf.rf[27][17] ;
 wire \dp.rf.rf[27][18] ;
 wire \dp.rf.rf[27][19] ;
 wire \dp.rf.rf[27][1] ;
 wire \dp.rf.rf[27][20] ;
 wire \dp.rf.rf[27][21] ;
 wire \dp.rf.rf[27][22] ;
 wire \dp.rf.rf[27][23] ;
 wire \dp.rf.rf[27][24] ;
 wire \dp.rf.rf[27][25] ;
 wire \dp.rf.rf[27][26] ;
 wire \dp.rf.rf[27][27] ;
 wire \dp.rf.rf[27][28] ;
 wire \dp.rf.rf[27][29] ;
 wire \dp.rf.rf[27][2] ;
 wire \dp.rf.rf[27][30] ;
 wire \dp.rf.rf[27][31] ;
 wire \dp.rf.rf[27][3] ;
 wire \dp.rf.rf[27][4] ;
 wire \dp.rf.rf[27][5] ;
 wire \dp.rf.rf[27][6] ;
 wire \dp.rf.rf[27][7] ;
 wire \dp.rf.rf[27][8] ;
 wire \dp.rf.rf[27][9] ;
 wire \dp.rf.rf[28][0] ;
 wire \dp.rf.rf[28][10] ;
 wire \dp.rf.rf[28][11] ;
 wire \dp.rf.rf[28][12] ;
 wire \dp.rf.rf[28][13] ;
 wire \dp.rf.rf[28][14] ;
 wire \dp.rf.rf[28][15] ;
 wire \dp.rf.rf[28][16] ;
 wire \dp.rf.rf[28][17] ;
 wire \dp.rf.rf[28][18] ;
 wire \dp.rf.rf[28][19] ;
 wire \dp.rf.rf[28][1] ;
 wire \dp.rf.rf[28][20] ;
 wire \dp.rf.rf[28][21] ;
 wire \dp.rf.rf[28][22] ;
 wire \dp.rf.rf[28][23] ;
 wire \dp.rf.rf[28][24] ;
 wire \dp.rf.rf[28][25] ;
 wire \dp.rf.rf[28][26] ;
 wire \dp.rf.rf[28][27] ;
 wire \dp.rf.rf[28][28] ;
 wire \dp.rf.rf[28][29] ;
 wire \dp.rf.rf[28][2] ;
 wire \dp.rf.rf[28][30] ;
 wire \dp.rf.rf[28][31] ;
 wire \dp.rf.rf[28][3] ;
 wire \dp.rf.rf[28][4] ;
 wire \dp.rf.rf[28][5] ;
 wire \dp.rf.rf[28][6] ;
 wire \dp.rf.rf[28][7] ;
 wire \dp.rf.rf[28][8] ;
 wire \dp.rf.rf[28][9] ;
 wire \dp.rf.rf[29][0] ;
 wire \dp.rf.rf[29][10] ;
 wire \dp.rf.rf[29][11] ;
 wire \dp.rf.rf[29][12] ;
 wire \dp.rf.rf[29][13] ;
 wire \dp.rf.rf[29][14] ;
 wire \dp.rf.rf[29][15] ;
 wire \dp.rf.rf[29][16] ;
 wire \dp.rf.rf[29][17] ;
 wire \dp.rf.rf[29][18] ;
 wire \dp.rf.rf[29][19] ;
 wire \dp.rf.rf[29][1] ;
 wire \dp.rf.rf[29][20] ;
 wire \dp.rf.rf[29][21] ;
 wire \dp.rf.rf[29][22] ;
 wire \dp.rf.rf[29][23] ;
 wire \dp.rf.rf[29][24] ;
 wire \dp.rf.rf[29][25] ;
 wire \dp.rf.rf[29][26] ;
 wire \dp.rf.rf[29][27] ;
 wire \dp.rf.rf[29][28] ;
 wire \dp.rf.rf[29][29] ;
 wire \dp.rf.rf[29][2] ;
 wire \dp.rf.rf[29][30] ;
 wire \dp.rf.rf[29][31] ;
 wire \dp.rf.rf[29][3] ;
 wire \dp.rf.rf[29][4] ;
 wire \dp.rf.rf[29][5] ;
 wire \dp.rf.rf[29][6] ;
 wire \dp.rf.rf[29][7] ;
 wire \dp.rf.rf[29][8] ;
 wire \dp.rf.rf[29][9] ;
 wire \dp.rf.rf[2][0] ;
 wire \dp.rf.rf[2][10] ;
 wire \dp.rf.rf[2][11] ;
 wire \dp.rf.rf[2][12] ;
 wire \dp.rf.rf[2][13] ;
 wire \dp.rf.rf[2][14] ;
 wire \dp.rf.rf[2][15] ;
 wire \dp.rf.rf[2][16] ;
 wire \dp.rf.rf[2][17] ;
 wire \dp.rf.rf[2][18] ;
 wire \dp.rf.rf[2][19] ;
 wire \dp.rf.rf[2][1] ;
 wire \dp.rf.rf[2][20] ;
 wire \dp.rf.rf[2][21] ;
 wire \dp.rf.rf[2][22] ;
 wire \dp.rf.rf[2][23] ;
 wire \dp.rf.rf[2][24] ;
 wire \dp.rf.rf[2][25] ;
 wire \dp.rf.rf[2][26] ;
 wire \dp.rf.rf[2][27] ;
 wire \dp.rf.rf[2][28] ;
 wire \dp.rf.rf[2][29] ;
 wire \dp.rf.rf[2][2] ;
 wire \dp.rf.rf[2][30] ;
 wire \dp.rf.rf[2][31] ;
 wire \dp.rf.rf[2][3] ;
 wire \dp.rf.rf[2][4] ;
 wire \dp.rf.rf[2][5] ;
 wire \dp.rf.rf[2][6] ;
 wire \dp.rf.rf[2][7] ;
 wire \dp.rf.rf[2][8] ;
 wire \dp.rf.rf[2][9] ;
 wire \dp.rf.rf[30][0] ;
 wire \dp.rf.rf[30][10] ;
 wire \dp.rf.rf[30][11] ;
 wire \dp.rf.rf[30][12] ;
 wire \dp.rf.rf[30][13] ;
 wire \dp.rf.rf[30][14] ;
 wire \dp.rf.rf[30][15] ;
 wire \dp.rf.rf[30][16] ;
 wire \dp.rf.rf[30][17] ;
 wire \dp.rf.rf[30][18] ;
 wire \dp.rf.rf[30][19] ;
 wire \dp.rf.rf[30][1] ;
 wire \dp.rf.rf[30][20] ;
 wire \dp.rf.rf[30][21] ;
 wire \dp.rf.rf[30][22] ;
 wire \dp.rf.rf[30][23] ;
 wire \dp.rf.rf[30][24] ;
 wire \dp.rf.rf[30][25] ;
 wire \dp.rf.rf[30][26] ;
 wire \dp.rf.rf[30][27] ;
 wire \dp.rf.rf[30][28] ;
 wire \dp.rf.rf[30][29] ;
 wire \dp.rf.rf[30][2] ;
 wire \dp.rf.rf[30][30] ;
 wire \dp.rf.rf[30][31] ;
 wire \dp.rf.rf[30][3] ;
 wire \dp.rf.rf[30][4] ;
 wire \dp.rf.rf[30][5] ;
 wire \dp.rf.rf[30][6] ;
 wire \dp.rf.rf[30][7] ;
 wire \dp.rf.rf[30][8] ;
 wire \dp.rf.rf[30][9] ;
 wire \dp.rf.rf[31][0] ;
 wire \dp.rf.rf[31][10] ;
 wire \dp.rf.rf[31][11] ;
 wire \dp.rf.rf[31][12] ;
 wire \dp.rf.rf[31][13] ;
 wire \dp.rf.rf[31][14] ;
 wire \dp.rf.rf[31][15] ;
 wire \dp.rf.rf[31][16] ;
 wire \dp.rf.rf[31][17] ;
 wire \dp.rf.rf[31][18] ;
 wire \dp.rf.rf[31][19] ;
 wire \dp.rf.rf[31][1] ;
 wire \dp.rf.rf[31][20] ;
 wire \dp.rf.rf[31][21] ;
 wire \dp.rf.rf[31][22] ;
 wire \dp.rf.rf[31][23] ;
 wire \dp.rf.rf[31][24] ;
 wire \dp.rf.rf[31][25] ;
 wire \dp.rf.rf[31][26] ;
 wire \dp.rf.rf[31][27] ;
 wire \dp.rf.rf[31][28] ;
 wire \dp.rf.rf[31][29] ;
 wire \dp.rf.rf[31][2] ;
 wire \dp.rf.rf[31][30] ;
 wire \dp.rf.rf[31][31] ;
 wire \dp.rf.rf[31][3] ;
 wire \dp.rf.rf[31][4] ;
 wire \dp.rf.rf[31][5] ;
 wire \dp.rf.rf[31][6] ;
 wire \dp.rf.rf[31][7] ;
 wire \dp.rf.rf[31][8] ;
 wire \dp.rf.rf[31][9] ;
 wire \dp.rf.rf[3][0] ;
 wire \dp.rf.rf[3][10] ;
 wire \dp.rf.rf[3][11] ;
 wire \dp.rf.rf[3][12] ;
 wire \dp.rf.rf[3][13] ;
 wire \dp.rf.rf[3][14] ;
 wire \dp.rf.rf[3][15] ;
 wire \dp.rf.rf[3][16] ;
 wire \dp.rf.rf[3][17] ;
 wire \dp.rf.rf[3][18] ;
 wire \dp.rf.rf[3][19] ;
 wire \dp.rf.rf[3][1] ;
 wire \dp.rf.rf[3][20] ;
 wire \dp.rf.rf[3][21] ;
 wire \dp.rf.rf[3][22] ;
 wire \dp.rf.rf[3][23] ;
 wire \dp.rf.rf[3][24] ;
 wire \dp.rf.rf[3][25] ;
 wire \dp.rf.rf[3][26] ;
 wire \dp.rf.rf[3][27] ;
 wire \dp.rf.rf[3][28] ;
 wire \dp.rf.rf[3][29] ;
 wire \dp.rf.rf[3][2] ;
 wire \dp.rf.rf[3][30] ;
 wire \dp.rf.rf[3][31] ;
 wire \dp.rf.rf[3][3] ;
 wire \dp.rf.rf[3][4] ;
 wire \dp.rf.rf[3][5] ;
 wire \dp.rf.rf[3][6] ;
 wire \dp.rf.rf[3][7] ;
 wire \dp.rf.rf[3][8] ;
 wire \dp.rf.rf[3][9] ;
 wire \dp.rf.rf[4][0] ;
 wire \dp.rf.rf[4][10] ;
 wire \dp.rf.rf[4][11] ;
 wire \dp.rf.rf[4][12] ;
 wire \dp.rf.rf[4][13] ;
 wire \dp.rf.rf[4][14] ;
 wire \dp.rf.rf[4][15] ;
 wire \dp.rf.rf[4][16] ;
 wire \dp.rf.rf[4][17] ;
 wire \dp.rf.rf[4][18] ;
 wire \dp.rf.rf[4][19] ;
 wire \dp.rf.rf[4][1] ;
 wire \dp.rf.rf[4][20] ;
 wire \dp.rf.rf[4][21] ;
 wire \dp.rf.rf[4][22] ;
 wire \dp.rf.rf[4][23] ;
 wire \dp.rf.rf[4][24] ;
 wire \dp.rf.rf[4][25] ;
 wire \dp.rf.rf[4][26] ;
 wire \dp.rf.rf[4][27] ;
 wire \dp.rf.rf[4][28] ;
 wire \dp.rf.rf[4][29] ;
 wire \dp.rf.rf[4][2] ;
 wire \dp.rf.rf[4][30] ;
 wire \dp.rf.rf[4][31] ;
 wire \dp.rf.rf[4][3] ;
 wire \dp.rf.rf[4][4] ;
 wire \dp.rf.rf[4][5] ;
 wire \dp.rf.rf[4][6] ;
 wire \dp.rf.rf[4][7] ;
 wire \dp.rf.rf[4][8] ;
 wire \dp.rf.rf[4][9] ;
 wire \dp.rf.rf[5][0] ;
 wire \dp.rf.rf[5][10] ;
 wire \dp.rf.rf[5][11] ;
 wire \dp.rf.rf[5][12] ;
 wire \dp.rf.rf[5][13] ;
 wire \dp.rf.rf[5][14] ;
 wire \dp.rf.rf[5][15] ;
 wire \dp.rf.rf[5][16] ;
 wire \dp.rf.rf[5][17] ;
 wire \dp.rf.rf[5][18] ;
 wire \dp.rf.rf[5][19] ;
 wire \dp.rf.rf[5][1] ;
 wire \dp.rf.rf[5][20] ;
 wire \dp.rf.rf[5][21] ;
 wire \dp.rf.rf[5][22] ;
 wire \dp.rf.rf[5][23] ;
 wire \dp.rf.rf[5][24] ;
 wire \dp.rf.rf[5][25] ;
 wire \dp.rf.rf[5][26] ;
 wire \dp.rf.rf[5][27] ;
 wire \dp.rf.rf[5][28] ;
 wire \dp.rf.rf[5][29] ;
 wire \dp.rf.rf[5][2] ;
 wire \dp.rf.rf[5][30] ;
 wire \dp.rf.rf[5][31] ;
 wire \dp.rf.rf[5][3] ;
 wire \dp.rf.rf[5][4] ;
 wire \dp.rf.rf[5][5] ;
 wire \dp.rf.rf[5][6] ;
 wire \dp.rf.rf[5][7] ;
 wire \dp.rf.rf[5][8] ;
 wire \dp.rf.rf[5][9] ;
 wire \dp.rf.rf[6][0] ;
 wire \dp.rf.rf[6][10] ;
 wire \dp.rf.rf[6][11] ;
 wire \dp.rf.rf[6][12] ;
 wire \dp.rf.rf[6][13] ;
 wire \dp.rf.rf[6][14] ;
 wire \dp.rf.rf[6][15] ;
 wire \dp.rf.rf[6][16] ;
 wire \dp.rf.rf[6][17] ;
 wire \dp.rf.rf[6][18] ;
 wire \dp.rf.rf[6][19] ;
 wire \dp.rf.rf[6][1] ;
 wire \dp.rf.rf[6][20] ;
 wire \dp.rf.rf[6][21] ;
 wire \dp.rf.rf[6][22] ;
 wire \dp.rf.rf[6][23] ;
 wire \dp.rf.rf[6][24] ;
 wire \dp.rf.rf[6][25] ;
 wire \dp.rf.rf[6][26] ;
 wire \dp.rf.rf[6][27] ;
 wire \dp.rf.rf[6][28] ;
 wire \dp.rf.rf[6][29] ;
 wire \dp.rf.rf[6][2] ;
 wire \dp.rf.rf[6][30] ;
 wire \dp.rf.rf[6][31] ;
 wire \dp.rf.rf[6][3] ;
 wire \dp.rf.rf[6][4] ;
 wire \dp.rf.rf[6][5] ;
 wire \dp.rf.rf[6][6] ;
 wire \dp.rf.rf[6][7] ;
 wire \dp.rf.rf[6][8] ;
 wire \dp.rf.rf[6][9] ;
 wire \dp.rf.rf[7][0] ;
 wire \dp.rf.rf[7][10] ;
 wire \dp.rf.rf[7][11] ;
 wire \dp.rf.rf[7][12] ;
 wire \dp.rf.rf[7][13] ;
 wire \dp.rf.rf[7][14] ;
 wire \dp.rf.rf[7][15] ;
 wire \dp.rf.rf[7][16] ;
 wire \dp.rf.rf[7][17] ;
 wire \dp.rf.rf[7][18] ;
 wire \dp.rf.rf[7][19] ;
 wire \dp.rf.rf[7][1] ;
 wire \dp.rf.rf[7][20] ;
 wire \dp.rf.rf[7][21] ;
 wire \dp.rf.rf[7][22] ;
 wire \dp.rf.rf[7][23] ;
 wire \dp.rf.rf[7][24] ;
 wire \dp.rf.rf[7][25] ;
 wire \dp.rf.rf[7][26] ;
 wire \dp.rf.rf[7][27] ;
 wire \dp.rf.rf[7][28] ;
 wire \dp.rf.rf[7][29] ;
 wire \dp.rf.rf[7][2] ;
 wire \dp.rf.rf[7][30] ;
 wire \dp.rf.rf[7][31] ;
 wire \dp.rf.rf[7][3] ;
 wire \dp.rf.rf[7][4] ;
 wire \dp.rf.rf[7][5] ;
 wire \dp.rf.rf[7][6] ;
 wire \dp.rf.rf[7][7] ;
 wire \dp.rf.rf[7][8] ;
 wire \dp.rf.rf[7][9] ;
 wire \dp.rf.rf[8][0] ;
 wire \dp.rf.rf[8][10] ;
 wire \dp.rf.rf[8][11] ;
 wire \dp.rf.rf[8][12] ;
 wire \dp.rf.rf[8][13] ;
 wire \dp.rf.rf[8][14] ;
 wire \dp.rf.rf[8][15] ;
 wire \dp.rf.rf[8][16] ;
 wire \dp.rf.rf[8][17] ;
 wire \dp.rf.rf[8][18] ;
 wire \dp.rf.rf[8][19] ;
 wire \dp.rf.rf[8][1] ;
 wire \dp.rf.rf[8][20] ;
 wire \dp.rf.rf[8][21] ;
 wire \dp.rf.rf[8][22] ;
 wire \dp.rf.rf[8][23] ;
 wire \dp.rf.rf[8][24] ;
 wire \dp.rf.rf[8][25] ;
 wire \dp.rf.rf[8][26] ;
 wire \dp.rf.rf[8][27] ;
 wire \dp.rf.rf[8][28] ;
 wire \dp.rf.rf[8][29] ;
 wire \dp.rf.rf[8][2] ;
 wire \dp.rf.rf[8][30] ;
 wire \dp.rf.rf[8][31] ;
 wire \dp.rf.rf[8][3] ;
 wire \dp.rf.rf[8][4] ;
 wire \dp.rf.rf[8][5] ;
 wire \dp.rf.rf[8][6] ;
 wire \dp.rf.rf[8][7] ;
 wire \dp.rf.rf[8][8] ;
 wire \dp.rf.rf[8][9] ;
 wire \dp.rf.rf[9][0] ;
 wire \dp.rf.rf[9][10] ;
 wire \dp.rf.rf[9][11] ;
 wire \dp.rf.rf[9][12] ;
 wire \dp.rf.rf[9][13] ;
 wire \dp.rf.rf[9][14] ;
 wire \dp.rf.rf[9][15] ;
 wire \dp.rf.rf[9][16] ;
 wire \dp.rf.rf[9][17] ;
 wire \dp.rf.rf[9][18] ;
 wire \dp.rf.rf[9][19] ;
 wire \dp.rf.rf[9][1] ;
 wire \dp.rf.rf[9][20] ;
 wire \dp.rf.rf[9][21] ;
 wire \dp.rf.rf[9][22] ;
 wire \dp.rf.rf[9][23] ;
 wire \dp.rf.rf[9][24] ;
 wire \dp.rf.rf[9][25] ;
 wire \dp.rf.rf[9][26] ;
 wire \dp.rf.rf[9][27] ;
 wire \dp.rf.rf[9][28] ;
 wire \dp.rf.rf[9][29] ;
 wire \dp.rf.rf[9][2] ;
 wire \dp.rf.rf[9][30] ;
 wire \dp.rf.rf[9][31] ;
 wire \dp.rf.rf[9][3] ;
 wire \dp.rf.rf[9][4] ;
 wire \dp.rf.rf[9][5] ;
 wire \dp.rf.rf[9][6] ;
 wire \dp.rf.rf[9][7] ;
 wire \dp.rf.rf[9][8] ;
 wire \dp.rf.rf[9][9] ;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_leaf_224_clk;
 wire clknet_leaf_225_clk;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_227_clk;
 wire clknet_leaf_228_clk;
 wire clknet_leaf_229_clk;
 wire clknet_leaf_230_clk;
 wire clknet_leaf_231_clk;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_233_clk;
 wire clknet_leaf_234_clk;
 wire clknet_leaf_235_clk;
 wire clknet_leaf_236_clk;
 wire clknet_leaf_237_clk;
 wire clknet_leaf_238_clk;
 wire clknet_leaf_239_clk;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_241_clk;
 wire clknet_leaf_242_clk;
 wire clknet_leaf_243_clk;
 wire clknet_leaf_244_clk;
 wire clknet_leaf_245_clk;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_247_clk;
 wire clknet_leaf_248_clk;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_250_clk;
 wire clknet_leaf_251_clk;
 wire clknet_leaf_254_clk;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_256_clk;
 wire clknet_leaf_257_clk;
 wire clknet_leaf_258_clk;
 wire clknet_leaf_259_clk;
 wire clknet_leaf_260_clk;
 wire clknet_leaf_262_clk;
 wire clknet_leaf_263_clk;
 wire clknet_leaf_264_clk;
 wire clknet_leaf_265_clk;
 wire clknet_leaf_266_clk;
 wire clknet_leaf_267_clk;
 wire clknet_leaf_268_clk;
 wire clknet_leaf_269_clk;
 wire clknet_leaf_270_clk;
 wire clknet_leaf_271_clk;
 wire clknet_leaf_272_clk;
 wire clknet_leaf_273_clk;
 wire clknet_leaf_274_clk;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_276_clk;
 wire clknet_leaf_277_clk;
 wire clknet_leaf_278_clk;
 wire clknet_leaf_279_clk;
 wire clknet_leaf_280_clk;
 wire clknet_leaf_281_clk;
 wire clknet_leaf_282_clk;
 wire clknet_leaf_283_clk;
 wire clknet_leaf_284_clk;
 wire clknet_leaf_285_clk;
 wire clknet_leaf_286_clk;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_288_clk;
 wire clknet_leaf_289_clk;
 wire clknet_leaf_290_clk;
 wire clknet_leaf_291_clk;
 wire clknet_leaf_292_clk;
 wire clknet_leaf_293_clk;
 wire clknet_leaf_294_clk;
 wire clknet_leaf_295_clk;
 wire clknet_leaf_296_clk;
 wire clknet_leaf_297_clk;
 wire clknet_leaf_298_clk;
 wire clknet_leaf_299_clk;
 wire clknet_leaf_300_clk;
 wire clknet_leaf_301_clk;
 wire clknet_leaf_302_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;
 wire net193;
 wire net308;
 wire net307;
 wire net298;
 wire net297;
 wire net292;
 wire net289;
 wire net286;
 wire net285;
 wire net284;
 wire net283;
 wire net281;
 wire net271;
 wire net270;
 wire net262;
 wire net256;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net321;
 wire net309;
 wire net258;
 wire net226;
 wire net225;
 wire net223;
 wire net222;
 wire net382;
 wire net314;
 wire net313;
 wire net312;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net253;
 wire net254;
 wire net255;
 wire net331;
 wire net257;
 wire net259;
 wire net260;
 wire net261;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net326;
 wire net327;
 wire net332;
 wire net334;
 wire net335;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net358;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net367;
 wire net368;
 wire net371;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net329;
 wire net330;
 wire [0:0] _3184_;
 wire [0:0] _3185_;
 wire [0:0] _3186_;
 wire [0:0] _3187_;
 wire [0:0] _3188_;
 wire [0:0] _3189_;
 wire [0:0] _3190_;
 wire [0:0] _3191_;
 wire [0:0] _3192_;
 wire [0:0] _3193_;
 wire [0:0] _3194_;
 wire [0:0] _3195_;
 wire [0:0] _3196_;
 wire [0:0] _3197_;
 wire [0:0] _3199_;
 wire [0:0] _3200_;
 wire [0:0] _3201_;
 wire [0:0] _3202_;
 wire [0:0] _3204_;
 wire [0:0] _3205_;
 wire [0:0] _3206_;
 wire [0:0] _3208_;
 wire [0:0] _3209_;
 wire [0:0] _3210_;
 wire [0:0] _3211_;
 wire [0:0] _3212_;
 wire [0:0] _3213_;
 wire [0:0] _3214_;
 wire [0:0] _3215_;
 wire [0:0] _3216_;
 wire [0:0] _3217_;
 wire [0:0] _3219_;
 wire [0:0] _3220_;
 wire [0:0] _3221_;
 wire [0:0] _3222_;
 wire [0:0] _3223_;
 wire [0:0] _3224_;
 wire [0:0] _3225_;
 wire [0:0] _3226_;
 wire [0:0] _3227_;
 wire [0:0] _3228_;
 wire [0:0] _3229_;
 wire [0:0] _3230_;
 wire [0:0] _3231_;
 wire [0:0] _3232_;
 wire [0:0] _3233_;
 wire [0:0] _3234_;
 wire [0:0] _3235_;
 wire [0:0] _3236_;
 wire [0:0] _3237_;
 wire [0:0] _3238_;
 wire [0:0] _3239_;
 wire [0:0] _3240_;
 wire [0:0] _3241_;
 wire [0:0] _3242_;
 wire [0:0] _3243_;
 wire [0:0] _3244_;
 wire [0:0] _3245_;
 wire [0:0] _3246_;
 wire [0:0] _3247_;
 wire [0:0] _3248_;
 wire [0:0] _3249_;
 wire [0:0] _3250_;
 wire [0:0] _3251_;
 wire [0:0] _3252_;
 wire [0:0] _3253_;
 wire [0:0] _3254_;
 wire [0:0] _3255_;
 wire [0:0] _3256_;
 wire [0:0] _3257_;
 wire [0:0] _3258_;
 wire [0:0] _3259_;
 wire [0:0] _3260_;
 wire [0:0] _3261_;
 wire [0:0] _3262_;
 wire [0:0] _3263_;
 wire [0:0] _3264_;
 wire [0:0] _3265_;
 wire [0:0] _3266_;
 wire [0:0] _3267_;
 wire [0:0] _3268_;
 wire [0:0] _3269_;
 wire [0:0] _3270_;
 wire [0:0] _3271_;
 wire [0:0] _3272_;
 wire [0:0] _3273_;
 wire [0:0] _3274_;
 wire [0:0] _3275_;
 wire [0:0] _3276_;
 wire [0:0] _3277_;
 wire [0:0] _3278_;
 wire [0:0] _3279_;
 wire [0:0] _3280_;
 wire [0:0] _3281_;
 wire [0:0] _3282_;
 wire [0:0] _3283_;
 wire [0:0] _3284_;
 wire [0:0] _3285_;
 wire [0:0] _3286_;
 wire [0:0] _3287_;
 wire [0:0] _3288_;
 wire [0:0] _3289_;
 wire [0:0] _3290_;
 wire [0:0] _3291_;
 wire [0:0] _3292_;
 wire [0:0] _3293_;
 wire [0:0] _3294_;
 wire [0:0] _3295_;
 wire [0:0] _3296_;
 wire [0:0] _3297_;
 wire [0:0] _3298_;
 wire [0:0] _3299_;
 wire [0:0] _3300_;
 wire [0:0] _3301_;
 wire [0:0] _3302_;
 wire [0:0] _3303_;
 wire [0:0] _3304_;
 wire [0:0] _3305_;
 wire [0:0] _3306_;
 wire [0:0] _3307_;
 wire [0:0] _3308_;
 wire [0:0] _3309_;
 wire [0:0] _3310_;
 wire [0:0] _3311_;
 wire [0:0] _3312_;
 wire [0:0] _3313_;
 wire [0:0] _3314_;
 wire [0:0] _3315_;
 wire [0:0] _3316_;
 wire [0:0] _3317_;
 wire [0:0] _3318_;
 wire [0:0] _3319_;
 wire [0:0] _3320_;
 wire [0:0] _3321_;
 wire [0:0] _3322_;
 wire [0:0] _3323_;
 wire [0:0] _3324_;
 wire [0:0] _3325_;
 wire [0:0] _3326_;
 wire [0:0] _3327_;
 wire [0:0] _3328_;
 wire [0:0] _3329_;
 wire [0:0] _3330_;
 wire [0:0] _3331_;
 wire [0:0] _3332_;
 wire [0:0] _3333_;
 wire [0:0] _3334_;
 wire [0:0] _3335_;
 wire [0:0] _3336_;
 wire [0:0] _3337_;
 wire [0:0] _3338_;
 wire [0:0] _3339_;
 wire [0:0] _3340_;
 wire [0:0] _3341_;
 wire [0:0] _3342_;
 wire [0:0] _3343_;
 wire [0:0] _3344_;
 wire [0:0] _3345_;
 wire [0:0] _3346_;
 wire [0:0] _3347_;
 wire [0:0] _3348_;
 wire [0:0] _3349_;
 wire [0:0] _3351_;
 wire [0:0] _3352_;
 wire [0:0] _3353_;
 wire [0:0] _3354_;
 wire [0:0] _3355_;
 wire [0:0] _3356_;
 wire [0:0] _3357_;
 wire [0:0] _3358_;
 wire [0:0] _3359_;
 wire [0:0] _3360_;
 wire [0:0] _3361_;
 wire [0:0] _3362_;
 wire [0:0] _3363_;
 wire [0:0] _3364_;
 wire [0:0] _3365_;
 wire [0:0] _3366_;
 wire [0:0] _3367_;
 wire [0:0] _3368_;
 wire [0:0] _3369_;
 wire [0:0] _3370_;
 wire [0:0] _3371_;
 wire [0:0] _3372_;
 wire [0:0] _3373_;
 wire [0:0] _3374_;
 wire [0:0] _3375_;
 wire [0:0] _3376_;
 wire [0:0] _3377_;
 wire [0:0] _3378_;
 wire [0:0] _3379_;
 wire [0:0] _3380_;
 wire [0:0] _3381_;
 wire [0:0] _3383_;
 wire [0:0] _3384_;
 wire [0:0] _3385_;
 wire [0:0] _3386_;
 wire [0:0] _3387_;
 wire [0:0] _3388_;
 wire [0:0] _3389_;
 wire [0:0] _3391_;
 wire [0:0] _3392_;
 wire [0:0] _3393_;
 wire [0:0] _3394_;
 wire [0:0] _3395_;
 wire [0:0] _3396_;
 wire [0:0] _3397_;
 wire [0:0] _3398_;
 wire [0:0] _3399_;
 wire [0:0] _3400_;
 wire [0:0] _3401_;
 wire [0:0] _3402_;
 wire [0:0] _3403_;
 wire [0:0] _3404_;
 wire [0:0] _3405_;
 wire [0:0] _3406_;
 wire [0:0] _3407_;
 wire [0:0] _3408_;
 wire [0:0] _3409_;
 wire [0:0] _3410_;
 wire [0:0] _3411_;
 wire [0:0] _3412_;
 wire [0:0] _3413_;
 wire [0:0] _3414_;
 wire [0:0] _3415_;
 wire [0:0] _3416_;
 wire [0:0] _3417_;
 wire [0:0] _3418_;
 wire [0:0] _3419_;
 wire [0:0] _3420_;
 wire [0:0] _3421_;
 wire [0:0] _3422_;
 wire [0:0] _3423_;
 wire [0:0] _3424_;
 wire [0:0] _3425_;
 wire [0:0] _3426_;
 wire [0:0] _3427_;
 wire [0:0] _3428_;
 wire [0:0] _3429_;
 wire [0:0] _3430_;
 wire [0:0] _3431_;
 wire [0:0] _3432_;
 wire [0:0] _3433_;
 wire [0:0] _3434_;
 wire [0:0] _3435_;
 wire [0:0] _3436_;
 wire [0:0] _3437_;
 wire [0:0] _3438_;
 wire [0:0] _3439_;
 wire [0:0] _3440_;
 wire [0:0] _3441_;
 wire [0:0] _3442_;
 wire [0:0] _3443_;
 wire [0:0] _3445_;
 wire [0:0] _3446_;
 wire [0:0] _3447_;
 wire [0:0] _3448_;
 wire [0:0] _3449_;
 wire [0:0] _3450_;
 wire [0:0] _3451_;
 wire [0:0] _3452_;
 wire [0:0] _3453_;
 wire [0:0] _3454_;
 wire [0:0] _3455_;
 wire [0:0] _3456_;
 wire [0:0] _3457_;
 wire [0:0] _3458_;
 wire [0:0] _3459_;
 wire [0:0] _3460_;
 wire [0:0] _3461_;
 wire [0:0] _3462_;
 wire [0:0] _3463_;
 wire [0:0] _3464_;
 wire [0:0] _3465_;
 wire [0:0] _3466_;
 wire [0:0] _3467_;
 wire [0:0] _3468_;
 wire [0:0] _3469_;
 wire [0:0] _3470_;
 wire [0:0] _3471_;
 wire [0:0] _3472_;
 wire [0:0] _3473_;
 wire [0:0] _3474_;
 wire [0:0] _3475_;
 wire [0:0] _3476_;
 wire [0:0] _3477_;
 wire [0:0] _3478_;
 wire [0:0] _3479_;
 wire [0:0] _3480_;
 wire [0:0] _3481_;
 wire [0:0] _3482_;
 wire [0:0] _3483_;
 wire [0:0] _3484_;
 wire [0:0] _3485_;
 wire [0:0] _3486_;
 wire [0:0] _3487_;
 wire [0:0] _3488_;
 wire [0:0] _3489_;
 wire [0:0] _3490_;
 wire [0:0] _3491_;
 wire [0:0] _3492_;
 wire [0:0] _3493_;
 wire [0:0] _3494_;
 wire [0:0] _3495_;
 wire [0:0] _3496_;
 wire [0:0] _3497_;
 wire [0:0] _3498_;
 wire [0:0] _3499_;
 wire [0:0] _3500_;
 wire [0:0] _3501_;
 wire [0:0] _3502_;
 wire [0:0] _3503_;
 wire [0:0] _3504_;
 wire [0:0] _3505_;
 wire [0:0] _3506_;
 wire [0:0] _3507_;
 wire [0:0] _3508_;
 wire [0:0] _3509_;
 wire [0:0] _3510_;
 wire [0:0] _3511_;
 wire [0:0] _3512_;
 wire [0:0] _3513_;
 wire [0:0] _3514_;
 wire [0:0] _3515_;
 wire [0:0] _3516_;
 wire [0:0] _3517_;
 wire [0:0] _3518_;
 wire [0:0] _3519_;
 wire [0:0] _3520_;
 wire [0:0] _3521_;
 wire [0:0] _3522_;
 wire [0:0] _3523_;
 wire [0:0] _3524_;
 wire [0:0] _3525_;
 wire [0:0] _3526_;
 wire [0:0] _3527_;
 wire [0:0] _3528_;
 wire [0:0] _3529_;
 wire [0:0] _3530_;
 wire [0:0] _3531_;
 wire [0:0] _3532_;
 wire [0:0] _3533_;
 wire [0:0] _3534_;
 wire [0:0] _3535_;
 wire [0:0] _3536_;
 wire [0:0] _3537_;
 wire [0:0] _3538_;
 wire [0:0] _3539_;
 wire [0:0] _3540_;
 wire [0:0] _3541_;
 wire [0:0] _3542_;
 wire [0:0] _3543_;
 wire [0:0] _3544_;
 wire [0:0] _3545_;
 wire [0:0] _3546_;
 wire [0:0] _3547_;
 wire [0:0] _3548_;
 wire [0:0] _3549_;
 wire [0:0] _3550_;
 wire [0:0] _3551_;
 wire [0:0] _3552_;
 wire [0:0] _3553_;
 wire [0:0] _3554_;
 wire [0:0] _3555_;
 wire [0:0] _3556_;
 wire [0:0] _3557_;
 wire [0:0] _3558_;
 wire [0:0] _3559_;
 wire [0:0] _3560_;
 wire [0:0] _3561_;
 wire [0:0] _3562_;
 wire [0:0] _3563_;
 wire [0:0] _3564_;
 wire [0:0] _3565_;
 wire [0:0] _3566_;
 wire [0:0] _3567_;
 wire [0:0] _3568_;
 wire [0:0] _3569_;
 wire [0:0] _3570_;

 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_365 ();
 sky130_fd_sc_hd__inv_6 _3573_ (.A(net29),
    .Y(_0035_));
 sky130_fd_sc_hd__nor2b_4 _3574_ (.A(net27),
    .B_N(net28),
    .Y(_0036_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_362 ();
 sky130_fd_sc_hd__nor4bb_1 _3578_ (.A(net26),
    .B(net23),
    .C_N(net1),
    .D_N(net12),
    .Y(_0040_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_361 ();
 sky130_fd_sc_hd__and2_4 _3580_ (.A(_0036_),
    .B(net803),
    .X(_0042_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_360 ();
 sky130_fd_sc_hd__nand2_8 _3582_ (.A(_0035_),
    .B(_0042_),
    .Y(_0044_));
 sky130_fd_sc_hd__clkinv_1 _3583_ (.A(_0044_),
    .Y(net99));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_349 ();
 sky130_fd_sc_hd__mux4_2 _3595_ (.A0(\dp.rf.rf[20][0] ),
    .A1(\dp.rf.rf[21][0] ),
    .A2(\dp.rf.rf[22][0] ),
    .A3(\dp.rf.rf[23][0] ),
    .S0(net823),
    .S1(net821),
    .X(_0056_));
 sky130_fd_sc_hd__mux4_2 _3596_ (.A0(\dp.rf.rf[28][0] ),
    .A1(\dp.rf.rf[29][0] ),
    .A2(\dp.rf.rf[30][0] ),
    .A3(\dp.rf.rf[31][0] ),
    .S0(net823),
    .S1(net821),
    .X(_0057_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_347 ();
 sky130_fd_sc_hd__mux2_4 _3599_ (.A0(_0056_),
    .A1(_0057_),
    .S(net16),
    .X(_0060_));
 sky130_fd_sc_hd__nand3_1 _3600_ (.A(net17),
    .B(net15),
    .C(_0060_),
    .Y(_0061_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_345 ();
 sky130_fd_sc_hd__nor2b_4 _3603_ (.A(net821),
    .B_N(net16),
    .Y(_0064_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_341 ();
 sky130_fd_sc_hd__mux2i_1 _3608_ (.A0(\dp.rf.rf[8][0] ),
    .A1(\dp.rf.rf[9][0] ),
    .S(net823),
    .Y(_0069_));
 sky130_fd_sc_hd__nand2_1 _3609_ (.A(_0064_),
    .B(_0069_),
    .Y(_0070_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_339 ();
 sky130_fd_sc_hd__nand2_2 _3612_ (.A(net821),
    .B(net16),
    .Y(_0073_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_336 ();
 sky130_fd_sc_hd__mux2_1 _3616_ (.A0(\dp.rf.rf[10][0] ),
    .A1(\dp.rf.rf[11][0] ),
    .S(net823),
    .X(_0077_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_335 ();
 sky130_fd_sc_hd__nor2b_4 _3618_ (.A(net16),
    .B_N(net821),
    .Y(_0079_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_331 ();
 sky130_fd_sc_hd__mux2i_1 _3623_ (.A0(\dp.rf.rf[2][0] ),
    .A1(\dp.rf.rf[3][0] ),
    .S(net823),
    .Y(_0084_));
 sky130_fd_sc_hd__a2bb2oi_1 _3624_ (.A1_N(_0073_),
    .A2_N(_0077_),
    .B1(_0079_),
    .B2(_0084_),
    .Y(_0085_));
 sky130_fd_sc_hd__nor2_2 _3625_ (.A(net821),
    .B(net16),
    .Y(_0086_));
 sky130_fd_sc_hd__mux2i_1 _3626_ (.A0(\dp.rf.rf[0][0] ),
    .A1(\dp.rf.rf[1][0] ),
    .S(net823),
    .Y(_0087_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_330 ();
 sky130_fd_sc_hd__or2_4 _3628_ (.A(net17),
    .B(net15),
    .X(_0089_));
 sky130_fd_sc_hd__a21oi_1 _3629_ (.A1(_0086_),
    .A2(_0087_),
    .B1(_0089_),
    .Y(_0090_));
 sky130_fd_sc_hd__nand3_2 _3630_ (.A(_0070_),
    .B(_0085_),
    .C(_0090_),
    .Y(_0091_));
 sky130_fd_sc_hd__clkinv_16 _3631_ (.A(net17),
    .Y(_0092_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_329 ();
 sky130_fd_sc_hd__nor2_4 _3633_ (.A(_0092_),
    .B(net15),
    .Y(_0094_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_327 ();
 sky130_fd_sc_hd__mux2_1 _3636_ (.A0(\dp.rf.rf[26][0] ),
    .A1(\dp.rf.rf[27][0] ),
    .S(net823),
    .X(_0097_));
 sky130_fd_sc_hd__mux2i_1 _3637_ (.A0(\dp.rf.rf[16][0] ),
    .A1(\dp.rf.rf[17][0] ),
    .S(net823),
    .Y(_0098_));
 sky130_fd_sc_hd__a2bb2oi_1 _3638_ (.A1_N(_0073_),
    .A2_N(_0097_),
    .B1(_0086_),
    .B2(_0098_),
    .Y(_0099_));
 sky130_fd_sc_hd__mux2i_1 _3639_ (.A0(\dp.rf.rf[18][0] ),
    .A1(\dp.rf.rf[19][0] ),
    .S(net823),
    .Y(_0100_));
 sky130_fd_sc_hd__mux2i_1 _3640_ (.A0(\dp.rf.rf[24][0] ),
    .A1(\dp.rf.rf[25][0] ),
    .S(net823),
    .Y(_0101_));
 sky130_fd_sc_hd__a22oi_1 _3641_ (.A1(_0079_),
    .A2(_0100_),
    .B1(_0101_),
    .B2(_0064_),
    .Y(_0102_));
 sky130_fd_sc_hd__mux4_2 _3642_ (.A0(\dp.rf.rf[4][0] ),
    .A1(\dp.rf.rf[5][0] ),
    .A2(\dp.rf.rf[6][0] ),
    .A3(\dp.rf.rf[7][0] ),
    .S0(net823),
    .S1(net821),
    .X(_0103_));
 sky130_fd_sc_hd__nor3b_1 _3643_ (.A(net17),
    .B(net16),
    .C_N(net15),
    .Y(_0104_));
 sky130_fd_sc_hd__and3b_1 _3644_ (.A_N(net17),
    .B(net15),
    .C(net16),
    .X(_0105_));
 sky130_fd_sc_hd__mux4_2 _3645_ (.A0(\dp.rf.rf[12][0] ),
    .A1(\dp.rf.rf[13][0] ),
    .A2(\dp.rf.rf[14][0] ),
    .A3(\dp.rf.rf[15][0] ),
    .S0(net823),
    .S1(net821),
    .X(_0106_));
 sky130_fd_sc_hd__a22o_1 _3646_ (.A1(_0103_),
    .A2(_0104_),
    .B1(_0105_),
    .B2(_0106_),
    .X(_0107_));
 sky130_fd_sc_hd__a31oi_2 _3647_ (.A1(_0094_),
    .A2(_0099_),
    .A3(_0102_),
    .B1(_0107_),
    .Y(_0108_));
 sky130_fd_sc_hd__nor2_4 _3648_ (.A(net17),
    .B(net817),
    .Y(_0109_));
 sky130_fd_sc_hd__nor3_4 _3649_ (.A(net14),
    .B(net13),
    .C(net818),
    .Y(_0110_));
 sky130_fd_sc_hd__and2_4 _3650_ (.A(_0109_),
    .B(_0110_),
    .X(_0111_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_326 ();
 sky130_fd_sc_hd__a31oi_4 _3652_ (.A1(_0061_),
    .A2(_0091_),
    .A3(_0108_),
    .B1(_0111_),
    .Y(net133));
 sky130_fd_sc_hd__nor2_1 _3653_ (.A(net28),
    .B(net29),
    .Y(_0113_));
 sky130_fd_sc_hd__nor2_1 _3654_ (.A(net26),
    .B(net23),
    .Y(_0114_));
 sky130_fd_sc_hd__o21ai_2 _3655_ (.A1(_0036_),
    .A2(_0113_),
    .B1(_0114_),
    .Y(_0115_));
 sky130_fd_sc_hd__nor3b_2 _3656_ (.A(net26),
    .B(net29),
    .C_N(net27),
    .Y(_0116_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_325 ();
 sky130_fd_sc_hd__and3b_4 _3658_ (.A_N(net27),
    .B(net28),
    .C(net29),
    .X(_0118_));
 sky130_fd_sc_hd__o21ai_2 _3659_ (.A1(net802),
    .A2(_0118_),
    .B1(net23),
    .Y(_0119_));
 sky130_fd_sc_hd__nand2_4 _3660_ (.A(net1),
    .B(net12),
    .Y(_0120_));
 sky130_fd_sc_hd__a21o_4 _3661_ (.A1(_0115_),
    .A2(_0119_),
    .B1(_0120_),
    .X(_0121_));
 sky130_fd_sc_hd__nand2_2 _3662_ (.A(net133),
    .B(_0121_),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_4 _3663_ (.A(net27),
    .Y(_0123_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_322 ();
 sky130_fd_sc_hd__nand2_2 _3667_ (.A(net28),
    .B(net816),
    .Y(_0127_));
 sky130_fd_sc_hd__nor3_1 _3668_ (.A(net815),
    .B(net5),
    .C(_0127_),
    .Y(_0128_));
 sky130_fd_sc_hd__a32oi_2 _3669_ (.A1(_0035_),
    .A2(net803),
    .A3(_0128_),
    .B1(_0127_),
    .B2(net5),
    .Y(_0129_));
 sky130_fd_sc_hd__nand2_4 _3670_ (.A(_0035_),
    .B(net803),
    .Y(_0130_));
 sky130_fd_sc_hd__nand2_1 _3671_ (.A(net5),
    .B(_0130_),
    .Y(_0131_));
 sky130_fd_sc_hd__o21ai_4 _3672_ (.A1(_0123_),
    .A2(_0129_),
    .B1(_0131_),
    .Y(_0132_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_321 ();
 sky130_fd_sc_hd__nand3_4 _3674_ (.A(net1),
    .B(net12),
    .C(net23),
    .Y(_0134_));
 sky130_fd_sc_hd__or3b_4 _3675_ (.A(net26),
    .B(net29),
    .C_N(net27),
    .X(_0135_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_320 ();
 sky130_fd_sc_hd__nor2_4 _3677_ (.A(_0134_),
    .B(_0135_),
    .Y(_0137_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_319 ();
 sky130_fd_sc_hd__and3_4 _3679_ (.A(net29),
    .B(_0036_),
    .C(net803),
    .X(_0139_));
 sky130_fd_sc_hd__nor3_4 _3680_ (.A(net814),
    .B(_0137_),
    .C(_0139_),
    .Y(_0140_));
 sky130_fd_sc_hd__a21bo_1 _3681_ (.A1(_0036_),
    .A2(net803),
    .B1_N(net13),
    .X(_0141_));
 sky130_fd_sc_hd__nand4_1 _3682_ (.A(_0035_),
    .B(net30),
    .C(_0036_),
    .D(net803),
    .Y(_0142_));
 sky130_fd_sc_hd__and3_4 _3683_ (.A(net1),
    .B(net12),
    .C(net23),
    .X(_0143_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_317 ();
 sky130_fd_sc_hd__and3_4 _3686_ (.A(net26),
    .B(_0143_),
    .C(_0118_),
    .X(_0146_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_316 ();
 sky130_fd_sc_hd__a211oi_4 _3688_ (.A1(_0141_),
    .A2(_0142_),
    .B1(_0137_),
    .C1(_0146_),
    .Y(_3449_[0]));
 sky130_fd_sc_hd__a21oi_4 _3689_ (.A1(_0115_),
    .A2(_0119_),
    .B1(_0120_),
    .Y(_0148_));
 sky130_fd_sc_hd__and2_4 _3690_ (.A(_3449_[0]),
    .B(_0148_),
    .X(_0149_));
 sky130_fd_sc_hd__a21oi_4 _3691_ (.A1(_0132_),
    .A2(_0140_),
    .B1(_0149_),
    .Y(_0150_));
 sky130_fd_sc_hd__nand2_8 _3692_ (.A(_0132_),
    .B(_0140_),
    .Y(_0151_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_314 ();
 sky130_fd_sc_hd__a21oi_4 _3695_ (.A1(_0121_),
    .A2(net133),
    .B1(_0149_),
    .Y(_0154_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_312 ();
 sky130_fd_sc_hd__nor2_1 _3698_ (.A(_0151_),
    .B(net768),
    .Y(_0157_));
 sky130_fd_sc_hd__a21oi_2 _3699_ (.A1(_0122_),
    .A2(_0150_),
    .B1(_0157_),
    .Y(_3195_[0]));
 sky130_fd_sc_hd__inv_1 _3700_ (.A(_3195_[0]),
    .Y(_3199_[0]));
 sky130_fd_sc_hd__inv_1 _3701_ (.A(\dp.rf.rf[0][0] ),
    .Y(_0158_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_306 ();
 sky130_fd_sc_hd__nor2_2 _3708_ (.A(net810),
    .B(net804),
    .Y(_0165_));
 sky130_fd_sc_hd__a21oi_4 _3709_ (.A1(_0143_),
    .A2(net802),
    .B1(_0165_),
    .Y(_0166_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_301 ();
 sky130_fd_sc_hd__mux2_1 _3715_ (.A0(\dp.rf.rf[1][0] ),
    .A1(\dp.rf.rf[5][0] ),
    .S(net9),
    .X(_0172_));
 sky130_fd_sc_hd__nor2b_4 _3716_ (.A(net812),
    .B_N(net804),
    .Y(_0173_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_296 ();
 sky130_fd_sc_hd__or2_4 _3722_ (.A(net808),
    .B(net10),
    .X(_0179_));
 sky130_fd_sc_hd__a221oi_1 _3723_ (.A1(net7),
    .A2(_0172_),
    .B1(net801),
    .B2(\dp.rf.rf[4][0] ),
    .C1(_0179_),
    .Y(_0180_));
 sky130_fd_sc_hd__o22ai_1 _3724_ (.A1(_0158_),
    .A2(_0166_),
    .B1(_0180_),
    .B2(_0137_),
    .Y(_0181_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_295 ();
 sky130_fd_sc_hd__or2_4 _3726_ (.A(net810),
    .B(net8),
    .X(_0183_));
 sky130_fd_sc_hd__nor3_2 _3727_ (.A(net805),
    .B(net10),
    .C(_0183_),
    .Y(_0184_));
 sky130_fd_sc_hd__nor3_4 _3728_ (.A(net11),
    .B(net799),
    .C(_0184_),
    .Y(_0185_));
 sky130_fd_sc_hd__clkinv_16 _3729_ (.A(net8),
    .Y(_0186_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_292 ();
 sky130_fd_sc_hd__mux4_2 _3733_ (.A0(\dp.rf.rf[2][0] ),
    .A1(\dp.rf.rf[3][0] ),
    .A2(\dp.rf.rf[6][0] ),
    .A3(\dp.rf.rf[7][0] ),
    .S0(net7),
    .S1(net9),
    .X(_0190_));
 sky130_fd_sc_hd__or3_1 _3734_ (.A(_0186_),
    .B(net10),
    .C(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__clkinv_16 _3735_ (.A(net10),
    .Y(_0192_));
 sky130_fd_sc_hd__a21oi_4 _3736_ (.A1(_0143_),
    .A2(net802),
    .B1(_0192_),
    .Y(_0193_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_286 ();
 sky130_fd_sc_hd__mux4_2 _3743_ (.A0(\dp.rf.rf[10][0] ),
    .A1(\dp.rf.rf[11][0] ),
    .A2(\dp.rf.rf[14][0] ),
    .A3(\dp.rf.rf[15][0] ),
    .S0(net7),
    .S1(net9),
    .X(_0200_));
 sky130_fd_sc_hd__nand2_1 _3744_ (.A(net8),
    .B(_0200_),
    .Y(_0201_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_285 ();
 sky130_fd_sc_hd__mux4_2 _3746_ (.A0(\dp.rf.rf[8][0] ),
    .A1(\dp.rf.rf[9][0] ),
    .A2(\dp.rf.rf[12][0] ),
    .A3(\dp.rf.rf[13][0] ),
    .S0(net7),
    .S1(net9),
    .X(_0203_));
 sky130_fd_sc_hd__nand2_1 _3747_ (.A(_0186_),
    .B(_0203_),
    .Y(_0204_));
 sky130_fd_sc_hd__nand3_1 _3748_ (.A(net797),
    .B(_0201_),
    .C(_0204_),
    .Y(_0205_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_284 ();
 sky130_fd_sc_hd__nor2_4 _3750_ (.A(net810),
    .B(net8),
    .Y(_0207_));
 sky130_fd_sc_hd__a21oi_4 _3751_ (.A1(_0143_),
    .A2(net802),
    .B1(_0207_),
    .Y(_0208_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_282 ();
 sky130_fd_sc_hd__nand2b_4 _3754_ (.A_N(net8),
    .B(net810),
    .Y(_0211_));
 sky130_fd_sc_hd__a211o_1 _3755_ (.A1(_0143_),
    .A2(net802),
    .B1(_0211_),
    .C1(\dp.rf.rf[25][0] ),
    .X(_0212_));
 sky130_fd_sc_hd__mux2i_1 _3756_ (.A0(\dp.rf.rf[26][0] ),
    .A1(\dp.rf.rf[27][0] ),
    .S(net7),
    .Y(_0213_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_280 ();
 sky130_fd_sc_hd__a21oi_1 _3759_ (.A1(net8),
    .A2(_0213_),
    .B1(net9),
    .Y(_0216_));
 sky130_fd_sc_hd__o211ai_1 _3760_ (.A1(\dp.rf.rf[24][0] ),
    .A2(_0208_),
    .B1(_0212_),
    .C1(_0216_),
    .Y(_0217_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_277 ();
 sky130_fd_sc_hd__mux4_2 _3764_ (.A0(\dp.rf.rf[28][0] ),
    .A1(\dp.rf.rf[29][0] ),
    .A2(\dp.rf.rf[30][0] ),
    .A3(\dp.rf.rf[31][0] ),
    .S0(net7),
    .S1(net8),
    .X(_0221_));
 sky130_fd_sc_hd__nand2_1 _3765_ (.A(net9),
    .B(_0221_),
    .Y(_0222_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_276 ();
 sky130_fd_sc_hd__o21ai_4 _3767_ (.A1(_0134_),
    .A2(_0135_),
    .B1(net11),
    .Y(_0224_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_272 ();
 sky130_fd_sc_hd__mux4_2 _3772_ (.A0(\dp.rf.rf[20][0] ),
    .A1(\dp.rf.rf[21][0] ),
    .A2(\dp.rf.rf[22][0] ),
    .A3(\dp.rf.rf[23][0] ),
    .S0(net7),
    .S1(net8),
    .X(_0229_));
 sky130_fd_sc_hd__nand2_1 _3773_ (.A(net9),
    .B(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__clkinvlp_4 _3774_ (.A(net9),
    .Y(_0231_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_271 ();
 sky130_fd_sc_hd__mux4_2 _3776_ (.A0(\dp.rf.rf[16][0] ),
    .A1(\dp.rf.rf[17][0] ),
    .A2(\dp.rf.rf[18][0] ),
    .A3(\dp.rf.rf[19][0] ),
    .S0(net7),
    .S1(net8),
    .X(_0233_));
 sky130_fd_sc_hd__nand2_1 _3777_ (.A(_0231_),
    .B(_0233_),
    .Y(_0234_));
 sky130_fd_sc_hd__and3_1 _3778_ (.A(_0192_),
    .B(_0230_),
    .C(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__a311oi_1 _3779_ (.A1(net797),
    .A2(_0217_),
    .A3(_0222_),
    .B1(net794),
    .C1(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__a41o_4 _3780_ (.A1(_0181_),
    .A2(net780),
    .A3(_0191_),
    .A4(_0205_),
    .B1(_0236_),
    .X(_3194_[0]));
 sky130_fd_sc_hd__inv_8 _3781_ (.A(_3194_[0]),
    .Y(_0237_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_270 ();
 sky130_fd_sc_hd__nor2_1 _3783_ (.A(\dp.rf.rf[24][31] ),
    .B(_0208_),
    .Y(_0238_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_265 ();
 sky130_fd_sc_hd__mux2i_1 _3789_ (.A0(\dp.rf.rf[26][31] ),
    .A1(\dp.rf.rf[27][31] ),
    .S(net810),
    .Y(_0244_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_262 ();
 sky130_fd_sc_hd__a21oi_1 _3793_ (.A1(net8),
    .A2(_0244_),
    .B1(net805),
    .Y(_0248_));
 sky130_fd_sc_hd__o31ai_1 _3794_ (.A1(\dp.rf.rf[25][31] ),
    .A2(net799),
    .A3(_0211_),
    .B1(_0248_),
    .Y(_0249_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_258 ();
 sky130_fd_sc_hd__mux4_2 _3799_ (.A0(\dp.rf.rf[28][31] ),
    .A1(\dp.rf.rf[29][31] ),
    .A2(\dp.rf.rf[30][31] ),
    .A3(\dp.rf.rf[31][31] ),
    .S0(net810),
    .S1(net8),
    .X(_0254_));
 sky130_fd_sc_hd__o21ai_4 _3800_ (.A1(_0134_),
    .A2(_0135_),
    .B1(net10),
    .Y(_0255_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_257 ();
 sky130_fd_sc_hd__a21oi_1 _3802_ (.A1(net805),
    .A2(_0254_),
    .B1(net793),
    .Y(_0257_));
 sky130_fd_sc_hd__o21ai_0 _3803_ (.A1(_0238_),
    .A2(_0249_),
    .B1(_0257_),
    .Y(_0258_));
 sky130_fd_sc_hd__a21oi_4 _3804_ (.A1(_0143_),
    .A2(net802),
    .B1(_0231_),
    .Y(_0259_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_254 ();
 sky130_fd_sc_hd__mux4_2 _3808_ (.A0(\dp.rf.rf[20][31] ),
    .A1(\dp.rf.rf[21][31] ),
    .A2(\dp.rf.rf[22][31] ),
    .A3(\dp.rf.rf[23][31] ),
    .S0(net810),
    .S1(net8),
    .X(_0263_));
 sky130_fd_sc_hd__nand2_1 _3809_ (.A(_0259_),
    .B(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__o21ai_4 _3810_ (.A1(_0134_),
    .A2(_0135_),
    .B1(_0192_),
    .Y(_0265_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_249 ();
 sky130_fd_sc_hd__mux2i_1 _3816_ (.A0(\dp.rf.rf[17][31] ),
    .A1(\dp.rf.rf[19][31] ),
    .S(net8),
    .Y(_0271_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_246 ();
 sky130_fd_sc_hd__nor3b_1 _3820_ (.A(\dp.rf.rf[18][31] ),
    .B(net810),
    .C_N(net8),
    .Y(_0275_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_243 ();
 sky130_fd_sc_hd__a211oi_1 _3824_ (.A1(net810),
    .A2(_0271_),
    .B1(_0275_),
    .C1(net805),
    .Y(_0279_));
 sky130_fd_sc_hd__a22oi_1 _3825_ (.A1(_0143_),
    .A2(net802),
    .B1(_0207_),
    .B2(_0192_),
    .Y(_0280_));
 sky130_fd_sc_hd__o22ai_1 _3826_ (.A1(net789),
    .A2(_0279_),
    .B1(_0280_),
    .B2(\dp.rf.rf[16][31] ),
    .Y(_0281_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_241 ();
 sky130_fd_sc_hd__a21oi_1 _3829_ (.A1(_0264_),
    .A2(_0281_),
    .B1(_0224_),
    .Y(_0284_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_239 ();
 sky130_fd_sc_hd__mux4_2 _3832_ (.A0(\dp.rf.rf[2][31] ),
    .A1(\dp.rf.rf[3][31] ),
    .A2(\dp.rf.rf[6][31] ),
    .A3(\dp.rf.rf[7][31] ),
    .S0(net810),
    .S1(net805),
    .X(_0287_));
 sky130_fd_sc_hd__nor2_1 _3833_ (.A(net789),
    .B(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__inv_1 _3834_ (.A(\dp.rf.rf[0][31] ),
    .Y(_0289_));
 sky130_fd_sc_hd__mux2_1 _3835_ (.A0(\dp.rf.rf[1][31] ),
    .A1(\dp.rf.rf[5][31] ),
    .S(net805),
    .X(_0290_));
 sky130_fd_sc_hd__a221oi_1 _3836_ (.A1(\dp.rf.rf[4][31] ),
    .A2(net801),
    .B1(_0290_),
    .B2(net810),
    .C1(_0179_),
    .Y(_0291_));
 sky130_fd_sc_hd__o22a_1 _3837_ (.A1(_0289_),
    .A2(_0166_),
    .B1(_0291_),
    .B2(net799),
    .X(_0292_));
 sky130_fd_sc_hd__or3_4 _3838_ (.A(net11),
    .B(net799),
    .C(_0184_),
    .X(_0293_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_237 ();
 sky130_fd_sc_hd__a211oi_1 _3841_ (.A1(net8),
    .A2(_0288_),
    .B1(_0292_),
    .C1(_0293_),
    .Y(_0296_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_236 ();
 sky130_fd_sc_hd__o21ai_4 _3843_ (.A1(_0134_),
    .A2(_0135_),
    .B1(net810),
    .Y(_0298_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_234 ();
 sky130_fd_sc_hd__a221oi_1 _3846_ (.A1(\dp.rf.rf[11][31] ),
    .A2(net810),
    .B1(_0298_),
    .B2(\dp.rf.rf[10][31] ),
    .C1(net792),
    .Y(_0301_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_233 ();
 sky130_fd_sc_hd__mux2_1 _3848_ (.A0(\dp.rf.rf[14][31] ),
    .A1(\dp.rf.rf[15][31] ),
    .S(net810),
    .X(_0303_));
 sky130_fd_sc_hd__a21oi_4 _3849_ (.A1(_0143_),
    .A2(net802),
    .B1(_0186_),
    .Y(_0304_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_231 ();
 sky130_fd_sc_hd__o21ai_0 _3852_ (.A1(net800),
    .A2(_0303_),
    .B1(net786),
    .Y(_0307_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_229 ();
 sky130_fd_sc_hd__mux4_2 _3855_ (.A0(\dp.rf.rf[8][31] ),
    .A1(\dp.rf.rf[9][31] ),
    .A2(\dp.rf.rf[12][31] ),
    .A3(\dp.rf.rf[13][31] ),
    .S0(net810),
    .S1(net805),
    .X(_0310_));
 sky130_fd_sc_hd__a21oi_1 _3856_ (.A1(_0186_),
    .A2(_0310_),
    .B1(net793),
    .Y(_0311_));
 sky130_fd_sc_hd__o21ai_2 _3857_ (.A1(_0301_),
    .A2(_0307_),
    .B1(_0311_),
    .Y(_0312_));
 sky130_fd_sc_hd__a22o_4 _3858_ (.A1(_0258_),
    .A2(_0284_),
    .B1(_0296_),
    .B2(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__inv_16 _3859_ (.A(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_223 ();
 sky130_fd_sc_hd__mux4_2 _3866_ (.A0(\dp.rf.rf[16][31] ),
    .A1(\dp.rf.rf[17][31] ),
    .A2(\dp.rf.rf[18][31] ),
    .A3(\dp.rf.rf[19][31] ),
    .S0(net826),
    .S1(net820),
    .X(_0320_));
 sky130_fd_sc_hd__mux4_2 _3867_ (.A0(\dp.rf.rf[20][31] ),
    .A1(\dp.rf.rf[21][31] ),
    .A2(\dp.rf.rf[22][31] ),
    .A3(\dp.rf.rf[23][31] ),
    .S0(net826),
    .S1(net820),
    .X(_0321_));
 sky130_fd_sc_hd__mux4_2 _3868_ (.A0(\dp.rf.rf[24][31] ),
    .A1(\dp.rf.rf[25][31] ),
    .A2(\dp.rf.rf[26][31] ),
    .A3(\dp.rf.rf[27][31] ),
    .S0(net826),
    .S1(net820),
    .X(_0322_));
 sky130_fd_sc_hd__mux4_2 _3869_ (.A0(\dp.rf.rf[28][31] ),
    .A1(\dp.rf.rf[29][31] ),
    .A2(\dp.rf.rf[30][31] ),
    .A3(\dp.rf.rf[31][31] ),
    .S0(net826),
    .S1(net820),
    .X(_0323_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_220 ();
 sky130_fd_sc_hd__mux4_2 _3873_ (.A0(_0320_),
    .A1(_0321_),
    .A2(_0322_),
    .A3(_0323_),
    .S0(net818),
    .S1(net817),
    .X(_0327_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_216 ();
 sky130_fd_sc_hd__mux4_2 _3878_ (.A0(\dp.rf.rf[0][31] ),
    .A1(\dp.rf.rf[1][31] ),
    .A2(\dp.rf.rf[2][31] ),
    .A3(\dp.rf.rf[3][31] ),
    .S0(net826),
    .S1(net820),
    .X(_0332_));
 sky130_fd_sc_hd__mux4_2 _3879_ (.A0(\dp.rf.rf[4][31] ),
    .A1(\dp.rf.rf[5][31] ),
    .A2(\dp.rf.rf[6][31] ),
    .A3(\dp.rf.rf[7][31] ),
    .S0(net826),
    .S1(net820),
    .X(_0333_));
 sky130_fd_sc_hd__mux4_2 _3880_ (.A0(\dp.rf.rf[8][31] ),
    .A1(\dp.rf.rf[9][31] ),
    .A2(\dp.rf.rf[10][31] ),
    .A3(\dp.rf.rf[11][31] ),
    .S0(net826),
    .S1(net820),
    .X(_0334_));
 sky130_fd_sc_hd__mux4_2 _3881_ (.A0(\dp.rf.rf[12][31] ),
    .A1(\dp.rf.rf[13][31] ),
    .A2(\dp.rf.rf[14][31] ),
    .A3(\dp.rf.rf[15][31] ),
    .S0(net826),
    .S1(net820),
    .X(_0335_));
 sky130_fd_sc_hd__mux4_2 _3882_ (.A0(_0332_),
    .A1(_0333_),
    .A2(_0334_),
    .A3(_0335_),
    .S0(net818),
    .S1(net817),
    .X(_0336_));
 sky130_fd_sc_hd__nor2_4 _3883_ (.A(net17),
    .B(_0111_),
    .Y(_0337_));
 sky130_fd_sc_hd__a22oi_2 _3884_ (.A1(net17),
    .A2(_0327_),
    .B1(_0336_),
    .B2(_0337_),
    .Y(_0338_));
 sky130_fd_sc_hd__nand2_1 _3885_ (.A(_0121_),
    .B(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__o21ai_2 _3886_ (.A1(net25),
    .A2(_0121_),
    .B1(_0339_),
    .Y(_0340_));
 sky130_fd_sc_hd__xor2_1 _3887_ (.A(_0151_),
    .B(_0340_),
    .X(_3202_[0]));
 sky130_fd_sc_hd__inv_1 _3888_ (.A(_3202_[0]),
    .Y(_3206_[0]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_210 ();
 sky130_fd_sc_hd__nand2_8 _3895_ (.A(_0143_),
    .B(net802),
    .Y(_0347_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_209 ();
 sky130_fd_sc_hd__and2_4 _3897_ (.A(net25),
    .B(_0347_),
    .X(_0349_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_208 ();
 sky130_fd_sc_hd__a21o_4 _3899_ (.A1(net816),
    .A2(net799),
    .B1(_0349_),
    .X(_3568_[0]));
 sky130_fd_sc_hd__nand2_8 _3900_ (.A(_0109_),
    .B(_0110_),
    .Y(_0351_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_206 ();
 sky130_fd_sc_hd__mux4_2 _3903_ (.A0(\dp.rf.rf[16][30] ),
    .A1(\dp.rf.rf[17][30] ),
    .A2(\dp.rf.rf[24][30] ),
    .A3(\dp.rf.rf[25][30] ),
    .S0(net826),
    .S1(net16),
    .X(_0354_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_205 ();
 sky130_fd_sc_hd__mux4_2 _3905_ (.A0(\dp.rf.rf[0][30] ),
    .A1(\dp.rf.rf[1][30] ),
    .A2(\dp.rf.rf[8][30] ),
    .A3(\dp.rf.rf[9][30] ),
    .S0(net13),
    .S1(net16),
    .X(_0356_));
 sky130_fd_sc_hd__mux4_2 _3906_ (.A0(\dp.rf.rf[18][30] ),
    .A1(\dp.rf.rf[19][30] ),
    .A2(\dp.rf.rf[26][30] ),
    .A3(\dp.rf.rf[27][30] ),
    .S0(net826),
    .S1(net16),
    .X(_0357_));
 sky130_fd_sc_hd__mux4_2 _3907_ (.A0(\dp.rf.rf[2][30] ),
    .A1(\dp.rf.rf[3][30] ),
    .A2(\dp.rf.rf[10][30] ),
    .A3(\dp.rf.rf[11][30] ),
    .S0(net826),
    .S1(net16),
    .X(_0358_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_203 ();
 sky130_fd_sc_hd__mux4_2 _3910_ (.A0(_0354_),
    .A1(_0356_),
    .A2(_0357_),
    .A3(_0358_),
    .S0(_0092_),
    .S1(net820),
    .X(_0361_));
 sky130_fd_sc_hd__mux4_2 _3911_ (.A0(\dp.rf.rf[4][30] ),
    .A1(\dp.rf.rf[5][30] ),
    .A2(\dp.rf.rf[6][30] ),
    .A3(\dp.rf.rf[7][30] ),
    .S0(net13),
    .S1(net820),
    .X(_0362_));
 sky130_fd_sc_hd__mux4_2 _3912_ (.A0(\dp.rf.rf[20][30] ),
    .A1(\dp.rf.rf[21][30] ),
    .A2(\dp.rf.rf[22][30] ),
    .A3(\dp.rf.rf[23][30] ),
    .S0(net826),
    .S1(net820),
    .X(_0363_));
 sky130_fd_sc_hd__mux4_2 _3913_ (.A0(\dp.rf.rf[12][30] ),
    .A1(\dp.rf.rf[13][30] ),
    .A2(\dp.rf.rf[14][30] ),
    .A3(\dp.rf.rf[15][30] ),
    .S0(net13),
    .S1(net820),
    .X(_0364_));
 sky130_fd_sc_hd__mux4_2 _3914_ (.A0(\dp.rf.rf[28][30] ),
    .A1(\dp.rf.rf[29][30] ),
    .A2(\dp.rf.rf[30][30] ),
    .A3(\dp.rf.rf[31][30] ),
    .S0(net826),
    .S1(net820),
    .X(_0365_));
 sky130_fd_sc_hd__mux4_2 _3915_ (.A0(_0362_),
    .A1(_0363_),
    .A2(_0364_),
    .A3(_0365_),
    .S0(net17),
    .S1(net16),
    .X(_0366_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_202 ();
 sky130_fd_sc_hd__mux2_4 _3917_ (.A0(_0361_),
    .A1(_0366_),
    .S(net818),
    .X(_0368_));
 sky130_fd_sc_hd__nand2_4 _3918_ (.A(_0351_),
    .B(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__nor2_1 _3919_ (.A(net782),
    .B(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__a21oi_1 _3920_ (.A1(net782),
    .A2(_3568_[0]),
    .B1(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__xor2_1 _3921_ (.A(_0151_),
    .B(_0371_),
    .X(_3211_[0]));
 sky130_fd_sc_hd__inv_1 _3922_ (.A(_3211_[0]),
    .Y(_3215_[0]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_201 ();
 sky130_fd_sc_hd__inv_1 _3924_ (.A(\dp.rf.rf[28][30] ),
    .Y(_0373_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_199 ();
 sky130_fd_sc_hd__mux2i_1 _3927_ (.A0(\dp.rf.rf[25][30] ),
    .A1(\dp.rf.rf[29][30] ),
    .S(net805),
    .Y(_0376_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_197 ();
 sky130_fd_sc_hd__a221oi_1 _3930_ (.A1(_0373_),
    .A2(net801),
    .B1(_0376_),
    .B2(net810),
    .C1(net8),
    .Y(_0379_));
 sky130_fd_sc_hd__o21ai_0 _3931_ (.A1(\dp.rf.rf[24][30] ),
    .A2(_0166_),
    .B1(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_195 ();
 sky130_fd_sc_hd__mux4_2 _3934_ (.A0(\dp.rf.rf[26][30] ),
    .A1(\dp.rf.rf[27][30] ),
    .A2(\dp.rf.rf[30][30] ),
    .A3(\dp.rf.rf[31][30] ),
    .S0(net810),
    .S1(net805),
    .X(_0383_));
 sky130_fd_sc_hd__nand2_1 _3935_ (.A(net786),
    .B(_0383_),
    .Y(_0384_));
 sky130_fd_sc_hd__nand3_2 _3936_ (.A(net10),
    .B(_0380_),
    .C(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__nor3_4 _3937_ (.A(net810),
    .B(net805),
    .C(net10),
    .Y(_0386_));
 sky130_fd_sc_hd__a21oi_1 _3938_ (.A1(\dp.rf.rf[18][30] ),
    .A2(net8),
    .B1(\dp.rf.rf[16][30] ),
    .Y(_0387_));
 sky130_fd_sc_hd__a21oi_1 _3939_ (.A1(_0386_),
    .A2(_0387_),
    .B1(_0224_),
    .Y(_0388_));
 sky130_fd_sc_hd__a21oi_4 _3940_ (.A1(_0143_),
    .A2(net802),
    .B1(net10),
    .Y(_0389_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_192 ();
 sky130_fd_sc_hd__mux4_2 _3944_ (.A0(\dp.rf.rf[18][30] ),
    .A1(\dp.rf.rf[19][30] ),
    .A2(\dp.rf.rf[22][30] ),
    .A3(\dp.rf.rf[23][30] ),
    .S0(net810),
    .S1(net805),
    .X(_0393_));
 sky130_fd_sc_hd__nand2_1 _3945_ (.A(net8),
    .B(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__nand2b_4 _3946_ (.A_N(net809),
    .B(net9),
    .Y(_0395_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_189 ();
 sky130_fd_sc_hd__mux2_1 _3950_ (.A0(\dp.rf.rf[17][30] ),
    .A1(\dp.rf.rf[21][30] ),
    .S(net805),
    .X(_0399_));
 sky130_fd_sc_hd__clkinv_16 _3951_ (.A(net809),
    .Y(_0400_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_188 ();
 sky130_fd_sc_hd__o221ai_1 _3953_ (.A1(\dp.rf.rf[20][30] ),
    .A2(_0395_),
    .B1(_0399_),
    .B2(_0400_),
    .C1(_0186_),
    .Y(_0402_));
 sky130_fd_sc_hd__nand3_2 _3954_ (.A(net785),
    .B(_0394_),
    .C(_0402_),
    .Y(_0403_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_186 ();
 sky130_fd_sc_hd__mux2_1 _3957_ (.A0(\dp.rf.rf[6][30] ),
    .A1(\dp.rf.rf[7][30] ),
    .S(net810),
    .X(_0406_));
 sky130_fd_sc_hd__o21ai_0 _3958_ (.A1(_0231_),
    .A2(_0406_),
    .B1(net786),
    .Y(_0407_));
 sky130_fd_sc_hd__a221oi_1 _3959_ (.A1(\dp.rf.rf[3][30] ),
    .A2(net810),
    .B1(_0298_),
    .B2(\dp.rf.rf[2][30] ),
    .C1(_0259_),
    .Y(_0408_));
 sky130_fd_sc_hd__inv_1 _3960_ (.A(\dp.rf.rf[4][30] ),
    .Y(_0409_));
 sky130_fd_sc_hd__mux2i_1 _3961_ (.A0(\dp.rf.rf[1][30] ),
    .A1(\dp.rf.rf[5][30] ),
    .S(net805),
    .Y(_0410_));
 sky130_fd_sc_hd__a221oi_1 _3962_ (.A1(_0409_),
    .A2(net801),
    .B1(_0410_),
    .B2(net810),
    .C1(net8),
    .Y(_0411_));
 sky130_fd_sc_hd__a21oi_4 _3963_ (.A1(_0143_),
    .A2(net802),
    .B1(_0386_),
    .Y(_0412_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_184 ();
 sky130_fd_sc_hd__o22ai_1 _3966_ (.A1(_0265_),
    .A2(_0411_),
    .B1(_0412_),
    .B2(\dp.rf.rf[0][30] ),
    .Y(_0415_));
 sky130_fd_sc_hd__o21ai_2 _3967_ (.A1(_0407_),
    .A2(_0408_),
    .B1(_0415_),
    .Y(_0416_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_183 ();
 sky130_fd_sc_hd__mux4_2 _3969_ (.A0(\dp.rf.rf[10][30] ),
    .A1(\dp.rf.rf[11][30] ),
    .A2(\dp.rf.rf[14][30] ),
    .A3(\dp.rf.rf[15][30] ),
    .S0(net810),
    .S1(net805),
    .X(_0418_));
 sky130_fd_sc_hd__nand2_1 _3970_ (.A(net8),
    .B(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__mux4_2 _3971_ (.A0(\dp.rf.rf[8][30] ),
    .A1(\dp.rf.rf[9][30] ),
    .A2(\dp.rf.rf[12][30] ),
    .A3(\dp.rf.rf[13][30] ),
    .S0(net810),
    .S1(net805),
    .X(_0420_));
 sky130_fd_sc_hd__nand2_1 _3972_ (.A(_0186_),
    .B(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__a31oi_2 _3973_ (.A1(_0193_),
    .A2(_0419_),
    .A3(_0421_),
    .B1(_0293_),
    .Y(_0422_));
 sky130_fd_sc_hd__a32oi_4 _3974_ (.A1(_0385_),
    .A2(_0388_),
    .A3(_0403_),
    .B1(_0416_),
    .B2(_0422_),
    .Y(_3214_[0]));
 sky130_fd_sc_hd__a21o_4 _3975_ (.A1(net22),
    .A2(net799),
    .B1(_0349_),
    .X(_3564_[0]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_181 ();
 sky130_fd_sc_hd__mux4_2 _3978_ (.A0(\dp.rf.rf[16][29] ),
    .A1(\dp.rf.rf[17][29] ),
    .A2(\dp.rf.rf[18][29] ),
    .A3(\dp.rf.rf[19][29] ),
    .S0(net825),
    .S1(net819),
    .X(_0425_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_179 ();
 sky130_fd_sc_hd__mux4_2 _3981_ (.A0(\dp.rf.rf[20][29] ),
    .A1(\dp.rf.rf[21][29] ),
    .A2(\dp.rf.rf[22][29] ),
    .A3(\dp.rf.rf[23][29] ),
    .S0(net825),
    .S1(net819),
    .X(_0428_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_177 ();
 sky130_fd_sc_hd__mux4_2 _3984_ (.A0(\dp.rf.rf[24][29] ),
    .A1(\dp.rf.rf[25][29] ),
    .A2(\dp.rf.rf[26][29] ),
    .A3(\dp.rf.rf[27][29] ),
    .S0(net825),
    .S1(net819),
    .X(_0431_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_176 ();
 sky130_fd_sc_hd__mux4_2 _3986_ (.A0(\dp.rf.rf[28][29] ),
    .A1(\dp.rf.rf[29][29] ),
    .A2(\dp.rf.rf[30][29] ),
    .A3(\dp.rf.rf[31][29] ),
    .S0(net825),
    .S1(net819),
    .X(_0433_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_174 ();
 sky130_fd_sc_hd__mux4_2 _3989_ (.A0(_0425_),
    .A1(_0428_),
    .A2(_0431_),
    .A3(_0433_),
    .S0(net15),
    .S1(net817),
    .X(_0436_));
 sky130_fd_sc_hd__nand2_1 _3990_ (.A(net17),
    .B(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_173 ();
 sky130_fd_sc_hd__mux4_2 _3992_ (.A0(\dp.rf.rf[0][29] ),
    .A1(\dp.rf.rf[1][29] ),
    .A2(\dp.rf.rf[2][29] ),
    .A3(\dp.rf.rf[3][29] ),
    .S0(net13),
    .S1(net14),
    .X(_0439_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_172 ();
 sky130_fd_sc_hd__mux4_2 _3994_ (.A0(\dp.rf.rf[4][29] ),
    .A1(\dp.rf.rf[5][29] ),
    .A2(\dp.rf.rf[6][29] ),
    .A3(\dp.rf.rf[7][29] ),
    .S0(net13),
    .S1(net14),
    .X(_0441_));
 sky130_fd_sc_hd__mux4_2 _3995_ (.A0(\dp.rf.rf[8][29] ),
    .A1(\dp.rf.rf[9][29] ),
    .A2(\dp.rf.rf[10][29] ),
    .A3(\dp.rf.rf[11][29] ),
    .S0(net13),
    .S1(net14),
    .X(_0442_));
 sky130_fd_sc_hd__mux4_2 _3996_ (.A0(\dp.rf.rf[12][29] ),
    .A1(\dp.rf.rf[13][29] ),
    .A2(\dp.rf.rf[14][29] ),
    .A3(\dp.rf.rf[15][29] ),
    .S0(net13),
    .S1(net14),
    .X(_0443_));
 sky130_fd_sc_hd__mux4_2 _3997_ (.A0(_0439_),
    .A1(_0441_),
    .A2(_0442_),
    .A3(_0443_),
    .S0(net15),
    .S1(net16),
    .X(_0444_));
 sky130_fd_sc_hd__nand2_2 _3998_ (.A(_0092_),
    .B(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__nand2_4 _3999_ (.A(_0437_),
    .B(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__nand2_8 _4000_ (.A(_0351_),
    .B(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__nor2_1 _4001_ (.A(net782),
    .B(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__a21oi_2 _4002_ (.A1(net782),
    .A2(_3564_[0]),
    .B1(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__xor2_1 _4003_ (.A(_0151_),
    .B(_0449_),
    .X(_3219_[0]));
 sky130_fd_sc_hd__inv_1 _4004_ (.A(_3219_[0]),
    .Y(_3223_[0]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_171 ();
 sky130_fd_sc_hd__mux2_1 _4006_ (.A0(\dp.rf.rf[1][29] ),
    .A1(\dp.rf.rf[5][29] ),
    .S(net804),
    .X(_0451_));
 sky130_fd_sc_hd__o22ai_1 _4007_ (.A1(\dp.rf.rf[4][29] ),
    .A2(_0395_),
    .B1(_0451_),
    .B2(_0400_),
    .Y(_0452_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_170 ();
 sky130_fd_sc_hd__mux4_2 _4009_ (.A0(\dp.rf.rf[2][29] ),
    .A1(\dp.rf.rf[3][29] ),
    .A2(\dp.rf.rf[6][29] ),
    .A3(\dp.rf.rf[7][29] ),
    .S0(net812),
    .S1(net804),
    .X(_0454_));
 sky130_fd_sc_hd__nand2_1 _4010_ (.A(net808),
    .B(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__o211ai_1 _4011_ (.A1(net808),
    .A2(_0452_),
    .B1(_0455_),
    .C1(_0389_),
    .Y(_0456_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_168 ();
 sky130_fd_sc_hd__mux4_2 _4014_ (.A0(\dp.rf.rf[10][29] ),
    .A1(\dp.rf.rf[11][29] ),
    .A2(\dp.rf.rf[14][29] ),
    .A3(\dp.rf.rf[15][29] ),
    .S0(net812),
    .S1(net804),
    .X(_0459_));
 sky130_fd_sc_hd__nand2_1 _4015_ (.A(net808),
    .B(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_166 ();
 sky130_fd_sc_hd__mux4_2 _4018_ (.A0(\dp.rf.rf[8][29] ),
    .A1(\dp.rf.rf[9][29] ),
    .A2(\dp.rf.rf[12][29] ),
    .A3(\dp.rf.rf[13][29] ),
    .S0(net812),
    .S1(net804),
    .X(_0463_));
 sky130_fd_sc_hd__nand2_1 _4019_ (.A(_0186_),
    .B(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__nand3_2 _4020_ (.A(net796),
    .B(_0460_),
    .C(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_165 ();
 sky130_fd_sc_hd__mux2_1 _4022_ (.A0(\dp.rf.rf[30][29] ),
    .A1(\dp.rf.rf[31][29] ),
    .S(net813),
    .X(_0467_));
 sky130_fd_sc_hd__inv_4 _4023_ (.A(net11),
    .Y(_0468_));
 sky130_fd_sc_hd__a211oi_4 _4024_ (.A1(_0143_),
    .A2(net802),
    .B1(_0186_),
    .C1(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__o21ai_0 _4025_ (.A1(net800),
    .A2(_0467_),
    .B1(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_163 ();
 sky130_fd_sc_hd__a221oi_1 _4028_ (.A1(\dp.rf.rf[27][29] ),
    .A2(net813),
    .B1(_0298_),
    .B2(\dp.rf.rf[26][29] ),
    .C1(_0259_),
    .Y(_0473_));
 sky130_fd_sc_hd__mux4_2 _4029_ (.A0(\dp.rf.rf[24][29] ),
    .A1(\dp.rf.rf[25][29] ),
    .A2(\dp.rf.rf[28][29] ),
    .A3(\dp.rf.rf[29][29] ),
    .S0(net813),
    .S1(net806),
    .X(_0474_));
 sky130_fd_sc_hd__a21oi_1 _4030_ (.A1(_0186_),
    .A2(_0474_),
    .B1(_0192_),
    .Y(_0475_));
 sky130_fd_sc_hd__o22ai_1 _4031_ (.A1(_0470_),
    .A2(_0473_),
    .B1(_0475_),
    .B2(net795),
    .Y(_0476_));
 sky130_fd_sc_hd__o21ai_4 _4032_ (.A1(_0134_),
    .A2(_0135_),
    .B1(net8),
    .Y(_0477_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_162 ();
 sky130_fd_sc_hd__nor2b_1 _4034_ (.A(net812),
    .B_N(\dp.rf.rf[22][29] ),
    .Y(_0479_));
 sky130_fd_sc_hd__a211oi_1 _4035_ (.A1(\dp.rf.rf[23][29] ),
    .A2(net812),
    .B1(net800),
    .C1(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__a221oi_1 _4036_ (.A1(\dp.rf.rf[19][29] ),
    .A2(net812),
    .B1(_0298_),
    .B2(\dp.rf.rf[18][29] ),
    .C1(_0259_),
    .Y(_0481_));
 sky130_fd_sc_hd__inv_1 _4037_ (.A(\dp.rf.rf[20][29] ),
    .Y(_0482_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_160 ();
 sky130_fd_sc_hd__mux2i_1 _4040_ (.A0(\dp.rf.rf[17][29] ),
    .A1(\dp.rf.rf[21][29] ),
    .S(net806),
    .Y(_0485_));
 sky130_fd_sc_hd__a221oi_1 _4041_ (.A1(_0482_),
    .A2(net801),
    .B1(_0485_),
    .B2(net812),
    .C1(net808),
    .Y(_0486_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_159 ();
 sky130_fd_sc_hd__o22ai_1 _4043_ (.A1(\dp.rf.rf[16][29] ),
    .A2(_0412_),
    .B1(_0486_),
    .B2(_0265_),
    .Y(_0488_));
 sky130_fd_sc_hd__o31ai_1 _4044_ (.A1(_0477_),
    .A2(_0480_),
    .A3(_0481_),
    .B1(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__a32o_4 _4045_ (.A1(net781),
    .A2(_0456_),
    .A3(_0465_),
    .B1(_0476_),
    .B2(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_158 ();
 sky130_fd_sc_hd__clkinvlp_4 _4047_ (.A(_0490_),
    .Y(_3222_[0]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_157 ();
 sky130_fd_sc_hd__a21o_4 _4049_ (.A1(net21),
    .A2(net799),
    .B1(_0349_),
    .X(_3560_[0]));
 sky130_fd_sc_hd__nand2_8 _4050_ (.A(_0092_),
    .B(_0351_),
    .Y(_0492_));
 sky130_fd_sc_hd__mux4_2 _4051_ (.A0(\dp.rf.rf[4][28] ),
    .A1(\dp.rf.rf[5][28] ),
    .A2(\dp.rf.rf[6][28] ),
    .A3(\dp.rf.rf[7][28] ),
    .S0(net13),
    .S1(net14),
    .X(_0493_));
 sky130_fd_sc_hd__mux4_2 _4052_ (.A0(\dp.rf.rf[12][28] ),
    .A1(\dp.rf.rf[13][28] ),
    .A2(\dp.rf.rf[14][28] ),
    .A3(\dp.rf.rf[15][28] ),
    .S0(net13),
    .S1(net14),
    .X(_0494_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_156 ();
 sky130_fd_sc_hd__mux2_4 _4054_ (.A0(_0493_),
    .A1(_0494_),
    .S(net16),
    .X(_0496_));
 sky130_fd_sc_hd__mux4_2 _4055_ (.A0(\dp.rf.rf[0][28] ),
    .A1(\dp.rf.rf[1][28] ),
    .A2(\dp.rf.rf[2][28] ),
    .A3(\dp.rf.rf[3][28] ),
    .S0(net13),
    .S1(net14),
    .X(_0497_));
 sky130_fd_sc_hd__mux4_2 _4056_ (.A0(\dp.rf.rf[8][28] ),
    .A1(\dp.rf.rf[9][28] ),
    .A2(\dp.rf.rf[10][28] ),
    .A3(\dp.rf.rf[11][28] ),
    .S0(net13),
    .S1(net14),
    .X(_0498_));
 sky130_fd_sc_hd__mux2i_1 _4057_ (.A0(_0497_),
    .A1(_0498_),
    .S(net16),
    .Y(_0499_));
 sky130_fd_sc_hd__nor2_1 _4058_ (.A(net15),
    .B(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__a21oi_4 _4059_ (.A1(net15),
    .A2(_0496_),
    .B1(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__mux4_2 _4060_ (.A0(\dp.rf.rf[16][28] ),
    .A1(\dp.rf.rf[17][28] ),
    .A2(\dp.rf.rf[18][28] ),
    .A3(\dp.rf.rf[19][28] ),
    .S0(net825),
    .S1(net819),
    .X(_0502_));
 sky130_fd_sc_hd__mux4_2 _4061_ (.A0(\dp.rf.rf[20][28] ),
    .A1(\dp.rf.rf[21][28] ),
    .A2(\dp.rf.rf[22][28] ),
    .A3(\dp.rf.rf[23][28] ),
    .S0(net825),
    .S1(net819),
    .X(_0503_));
 sky130_fd_sc_hd__mux4_2 _4062_ (.A0(\dp.rf.rf[24][28] ),
    .A1(\dp.rf.rf[25][28] ),
    .A2(\dp.rf.rf[26][28] ),
    .A3(\dp.rf.rf[27][28] ),
    .S0(net825),
    .S1(net819),
    .X(_0504_));
 sky130_fd_sc_hd__mux4_2 _4063_ (.A0(\dp.rf.rf[28][28] ),
    .A1(\dp.rf.rf[29][28] ),
    .A2(\dp.rf.rf[30][28] ),
    .A3(\dp.rf.rf[31][28] ),
    .S0(net825),
    .S1(net819),
    .X(_0505_));
 sky130_fd_sc_hd__mux4_2 _4064_ (.A0(_0502_),
    .A1(_0503_),
    .A2(_0504_),
    .A3(_0505_),
    .S0(net15),
    .S1(net817),
    .X(_0506_));
 sky130_fd_sc_hd__nand2_4 _4065_ (.A(net17),
    .B(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__o21ai_4 _4066_ (.A1(_0492_),
    .A2(_0501_),
    .B1(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__mux2_1 _4067_ (.A0(_3560_[0]),
    .A1(_0508_),
    .S(_0121_),
    .X(_0509_));
 sky130_fd_sc_hd__xnor2_1 _4068_ (.A(_0151_),
    .B(_0509_),
    .Y(_3227_[0]));
 sky130_fd_sc_hd__inv_1 _4069_ (.A(_3227_[0]),
    .Y(_3231_[0]));
 sky130_fd_sc_hd__mux4_2 _4070_ (.A0(\dp.rf.rf[24][28] ),
    .A1(\dp.rf.rf[25][28] ),
    .A2(\dp.rf.rf[28][28] ),
    .A3(\dp.rf.rf[29][28] ),
    .S0(net811),
    .S1(net807),
    .X(_0510_));
 sky130_fd_sc_hd__mux2i_1 _4071_ (.A0(\dp.rf.rf[30][28] ),
    .A1(\dp.rf.rf[31][28] ),
    .S(net811),
    .Y(_0511_));
 sky130_fd_sc_hd__mux2i_1 _4072_ (.A0(\dp.rf.rf[26][28] ),
    .A1(\dp.rf.rf[27][28] ),
    .S(net811),
    .Y(_0512_));
 sky130_fd_sc_hd__o21ai_4 _4073_ (.A1(_0134_),
    .A2(_0135_),
    .B1(net804),
    .Y(_0513_));
 sky130_fd_sc_hd__a221oi_1 _4074_ (.A1(net807),
    .A2(_0511_),
    .B1(_0512_),
    .B2(_0513_),
    .C1(_0186_),
    .Y(_0514_));
 sky130_fd_sc_hd__a211o_1 _4075_ (.A1(_0186_),
    .A2(_0510_),
    .B1(_0514_),
    .C1(_0192_),
    .X(_0515_));
 sky130_fd_sc_hd__mux4_2 _4076_ (.A0(\dp.rf.rf[16][28] ),
    .A1(\dp.rf.rf[17][28] ),
    .A2(\dp.rf.rf[20][28] ),
    .A3(\dp.rf.rf[21][28] ),
    .S0(net811),
    .S1(net806),
    .X(_0516_));
 sky130_fd_sc_hd__a21oi_1 _4077_ (.A1(_0186_),
    .A2(_0516_),
    .B1(net10),
    .Y(_0517_));
 sky130_fd_sc_hd__mux4_2 _4078_ (.A0(\dp.rf.rf[18][28] ),
    .A1(\dp.rf.rf[19][28] ),
    .A2(\dp.rf.rf[22][28] ),
    .A3(\dp.rf.rf[23][28] ),
    .S0(net811),
    .S1(net806),
    .X(_0518_));
 sky130_fd_sc_hd__nand2_1 _4079_ (.A(_0469_),
    .B(_0518_),
    .Y(_0519_));
 sky130_fd_sc_hd__o21ai_2 _4080_ (.A1(net795),
    .A2(_0517_),
    .B1(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__mux4_2 _4081_ (.A0(\dp.rf.rf[2][28] ),
    .A1(\dp.rf.rf[3][28] ),
    .A2(\dp.rf.rf[6][28] ),
    .A3(\dp.rf.rf[7][28] ),
    .S0(net813),
    .S1(net807),
    .X(_0521_));
 sky130_fd_sc_hd__nand2_1 _4082_ (.A(net808),
    .B(_0521_),
    .Y(_0522_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_155 ();
 sky130_fd_sc_hd__mux2_1 _4084_ (.A0(\dp.rf.rf[1][28] ),
    .A1(\dp.rf.rf[5][28] ),
    .S(net807),
    .X(_0524_));
 sky130_fd_sc_hd__o221ai_1 _4085_ (.A1(\dp.rf.rf[4][28] ),
    .A2(_0395_),
    .B1(_0524_),
    .B2(_0400_),
    .C1(_0186_),
    .Y(_0525_));
 sky130_fd_sc_hd__a31o_4 _4086_ (.A1(net785),
    .A2(_0522_),
    .A3(_0525_),
    .B1(_0293_),
    .X(_0526_));
 sky130_fd_sc_hd__mux2i_1 _4087_ (.A0(\dp.rf.rf[14][28] ),
    .A1(\dp.rf.rf[15][28] ),
    .S(net813),
    .Y(_0527_));
 sky130_fd_sc_hd__a21oi_1 _4088_ (.A1(net807),
    .A2(_0527_),
    .B1(_0477_),
    .Y(_0528_));
 sky130_fd_sc_hd__a221o_1 _4089_ (.A1(\dp.rf.rf[11][28] ),
    .A2(net813),
    .B1(net787),
    .B2(\dp.rf.rf[10][28] ),
    .C1(net792),
    .X(_0529_));
 sky130_fd_sc_hd__mux4_2 _4090_ (.A0(\dp.rf.rf[8][28] ),
    .A1(\dp.rf.rf[9][28] ),
    .A2(\dp.rf.rf[12][28] ),
    .A3(\dp.rf.rf[13][28] ),
    .S0(net813),
    .S1(net807),
    .X(_0530_));
 sky130_fd_sc_hd__a221oi_2 _4091_ (.A1(_0528_),
    .A2(_0529_),
    .B1(_0530_),
    .B2(_0186_),
    .C1(net793),
    .Y(_0531_));
 sky130_fd_sc_hd__o2bb2ai_4 _4092_ (.A1_N(_0515_),
    .A2_N(_0520_),
    .B1(_0526_),
    .B2(_0531_),
    .Y(_3226_[0]));
 sky130_fd_sc_hd__inv_6 _4093_ (.A(_3226_[0]),
    .Y(_3230_[0]));
 sky130_fd_sc_hd__a21o_4 _4094_ (.A1(net20),
    .A2(net799),
    .B1(_0349_),
    .X(_3556_[0]));
 sky130_fd_sc_hd__mux4_2 _4095_ (.A0(\dp.rf.rf[16][27] ),
    .A1(\dp.rf.rf[17][27] ),
    .A2(\dp.rf.rf[18][27] ),
    .A3(\dp.rf.rf[19][27] ),
    .S0(net826),
    .S1(net820),
    .X(_0532_));
 sky130_fd_sc_hd__mux4_2 _4096_ (.A0(\dp.rf.rf[20][27] ),
    .A1(\dp.rf.rf[21][27] ),
    .A2(\dp.rf.rf[22][27] ),
    .A3(\dp.rf.rf[23][27] ),
    .S0(net826),
    .S1(net820),
    .X(_0533_));
 sky130_fd_sc_hd__mux4_2 _4097_ (.A0(\dp.rf.rf[24][27] ),
    .A1(\dp.rf.rf[25][27] ),
    .A2(\dp.rf.rf[26][27] ),
    .A3(\dp.rf.rf[27][27] ),
    .S0(net825),
    .S1(net819),
    .X(_0534_));
 sky130_fd_sc_hd__mux4_2 _4098_ (.A0(\dp.rf.rf[28][27] ),
    .A1(\dp.rf.rf[29][27] ),
    .A2(\dp.rf.rf[30][27] ),
    .A3(\dp.rf.rf[31][27] ),
    .S0(net825),
    .S1(net819),
    .X(_0535_));
 sky130_fd_sc_hd__mux4_2 _4099_ (.A0(_0532_),
    .A1(_0533_),
    .A2(_0534_),
    .A3(_0535_),
    .S0(net15),
    .S1(net817),
    .X(_0536_));
 sky130_fd_sc_hd__mux4_2 _4100_ (.A0(\dp.rf.rf[0][27] ),
    .A1(\dp.rf.rf[1][27] ),
    .A2(\dp.rf.rf[2][27] ),
    .A3(\dp.rf.rf[3][27] ),
    .S0(net825),
    .S1(net819),
    .X(_0537_));
 sky130_fd_sc_hd__mux4_2 _4101_ (.A0(\dp.rf.rf[4][27] ),
    .A1(\dp.rf.rf[5][27] ),
    .A2(\dp.rf.rf[6][27] ),
    .A3(\dp.rf.rf[7][27] ),
    .S0(net13),
    .S1(net14),
    .X(_0538_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_154 ();
 sky130_fd_sc_hd__mux4_2 _4103_ (.A0(\dp.rf.rf[8][27] ),
    .A1(\dp.rf.rf[9][27] ),
    .A2(\dp.rf.rf[10][27] ),
    .A3(\dp.rf.rf[11][27] ),
    .S0(net13),
    .S1(net14),
    .X(_0540_));
 sky130_fd_sc_hd__mux4_2 _4104_ (.A0(\dp.rf.rf[12][27] ),
    .A1(\dp.rf.rf[13][27] ),
    .A2(\dp.rf.rf[14][27] ),
    .A3(\dp.rf.rf[15][27] ),
    .S0(net13),
    .S1(net14),
    .X(_0541_));
 sky130_fd_sc_hd__mux4_2 _4105_ (.A0(_0537_),
    .A1(_0538_),
    .A2(_0540_),
    .A3(_0541_),
    .S0(net15),
    .S1(net16),
    .X(_0542_));
 sky130_fd_sc_hd__a22o_4 _4106_ (.A1(net17),
    .A2(_0536_),
    .B1(_0542_),
    .B2(_0337_),
    .X(_0543_));
 sky130_fd_sc_hd__mux2_1 _4107_ (.A0(_3556_[0]),
    .A1(_0543_),
    .S(_0121_),
    .X(_0544_));
 sky130_fd_sc_hd__xnor2_1 _4108_ (.A(_0151_),
    .B(_0544_),
    .Y(_3235_[0]));
 sky130_fd_sc_hd__inv_1 _4109_ (.A(_3235_[0]),
    .Y(_3239_[0]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_152 ();
 sky130_fd_sc_hd__mux4_2 _4112_ (.A0(\dp.rf.rf[10][27] ),
    .A1(\dp.rf.rf[11][27] ),
    .A2(\dp.rf.rf[14][27] ),
    .A3(\dp.rf.rf[15][27] ),
    .S0(net811),
    .S1(net807),
    .X(_0547_));
 sky130_fd_sc_hd__nand2_1 _4113_ (.A(net808),
    .B(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__mux4_2 _4114_ (.A0(\dp.rf.rf[8][27] ),
    .A1(\dp.rf.rf[9][27] ),
    .A2(\dp.rf.rf[12][27] ),
    .A3(\dp.rf.rf[13][27] ),
    .S0(net811),
    .S1(net807),
    .X(_0549_));
 sky130_fd_sc_hd__nand2_1 _4115_ (.A(_0186_),
    .B(_0549_),
    .Y(_0550_));
 sky130_fd_sc_hd__a31oi_2 _4116_ (.A1(net796),
    .A2(_0548_),
    .A3(_0550_),
    .B1(_0293_),
    .Y(_0551_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_151 ();
 sky130_fd_sc_hd__mux2_1 _4118_ (.A0(\dp.rf.rf[6][27] ),
    .A1(\dp.rf.rf[7][27] ),
    .S(net811),
    .X(_0553_));
 sky130_fd_sc_hd__o21ai_0 _4119_ (.A1(net800),
    .A2(_0553_),
    .B1(net786),
    .Y(_0554_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_150 ();
 sky130_fd_sc_hd__a221oi_1 _4121_ (.A1(\dp.rf.rf[3][27] ),
    .A2(net811),
    .B1(net787),
    .B2(\dp.rf.rf[2][27] ),
    .C1(net792),
    .Y(_0556_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_149 ();
 sky130_fd_sc_hd__inv_1 _4123_ (.A(\dp.rf.rf[4][27] ),
    .Y(_0558_));
 sky130_fd_sc_hd__mux2i_1 _4124_ (.A0(\dp.rf.rf[1][27] ),
    .A1(\dp.rf.rf[5][27] ),
    .S(net807),
    .Y(_0559_));
 sky130_fd_sc_hd__a221oi_1 _4125_ (.A1(_0558_),
    .A2(net801),
    .B1(_0559_),
    .B2(net811),
    .C1(net808),
    .Y(_0560_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_148 ();
 sky130_fd_sc_hd__o22ai_1 _4127_ (.A1(\dp.rf.rf[0][27] ),
    .A2(_0412_),
    .B1(_0560_),
    .B2(net789),
    .Y(_0562_));
 sky130_fd_sc_hd__o21ai_2 _4128_ (.A1(_0554_),
    .A2(_0556_),
    .B1(_0562_),
    .Y(_0563_));
 sky130_fd_sc_hd__inv_1 _4129_ (.A(\dp.rf.rf[28][27] ),
    .Y(_0564_));
 sky130_fd_sc_hd__mux2i_1 _4130_ (.A0(\dp.rf.rf[25][27] ),
    .A1(\dp.rf.rf[29][27] ),
    .S(net806),
    .Y(_0565_));
 sky130_fd_sc_hd__a221oi_1 _4131_ (.A1(_0564_),
    .A2(net801),
    .B1(_0565_),
    .B2(net811),
    .C1(net808),
    .Y(_0566_));
 sky130_fd_sc_hd__o21ai_0 _4132_ (.A1(\dp.rf.rf[24][27] ),
    .A2(net798),
    .B1(_0566_),
    .Y(_0567_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_147 ();
 sky130_fd_sc_hd__mux4_2 _4134_ (.A0(\dp.rf.rf[26][27] ),
    .A1(\dp.rf.rf[27][27] ),
    .A2(\dp.rf.rf[30][27] ),
    .A3(\dp.rf.rf[31][27] ),
    .S0(net811),
    .S1(net806),
    .X(_0569_));
 sky130_fd_sc_hd__nand2_1 _4135_ (.A(net786),
    .B(_0569_),
    .Y(_0570_));
 sky130_fd_sc_hd__nand3_1 _4136_ (.A(net10),
    .B(_0567_),
    .C(_0570_),
    .Y(_0571_));
 sky130_fd_sc_hd__inv_1 _4137_ (.A(\dp.rf.rf[20][27] ),
    .Y(_0572_));
 sky130_fd_sc_hd__mux2i_1 _4138_ (.A0(\dp.rf.rf[17][27] ),
    .A1(\dp.rf.rf[21][27] ),
    .S(net806),
    .Y(_0573_));
 sky130_fd_sc_hd__a221oi_1 _4139_ (.A1(_0572_),
    .A2(net801),
    .B1(_0573_),
    .B2(net811),
    .C1(net808),
    .Y(_0574_));
 sky130_fd_sc_hd__o22ai_1 _4140_ (.A1(\dp.rf.rf[16][27] ),
    .A2(net798),
    .B1(_0574_),
    .B2(net799),
    .Y(_0575_));
 sky130_fd_sc_hd__mux4_2 _4141_ (.A0(\dp.rf.rf[18][27] ),
    .A1(\dp.rf.rf[19][27] ),
    .A2(\dp.rf.rf[22][27] ),
    .A3(\dp.rf.rf[23][27] ),
    .S0(net811),
    .S1(net806),
    .X(_0576_));
 sky130_fd_sc_hd__a21oi_1 _4142_ (.A1(net808),
    .A2(_0576_),
    .B1(net10),
    .Y(_0577_));
 sky130_fd_sc_hd__a21oi_1 _4143_ (.A1(_0575_),
    .A2(_0577_),
    .B1(net795),
    .Y(_0578_));
 sky130_fd_sc_hd__a22oi_2 _4144_ (.A1(_0551_),
    .A2(_0563_),
    .B1(_0571_),
    .B2(_0578_),
    .Y(_3238_[0]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_146 ();
 sky130_fd_sc_hd__a21o_4 _4146_ (.A1(net19),
    .A2(net799),
    .B1(_0349_),
    .X(_3552_[0]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_145 ();
 sky130_fd_sc_hd__mux4_2 _4148_ (.A0(\dp.rf.rf[16][26] ),
    .A1(\dp.rf.rf[17][26] ),
    .A2(\dp.rf.rf[18][26] ),
    .A3(\dp.rf.rf[19][26] ),
    .S0(net826),
    .S1(net820),
    .X(_0581_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_144 ();
 sky130_fd_sc_hd__mux4_2 _4150_ (.A0(\dp.rf.rf[24][26] ),
    .A1(\dp.rf.rf[25][26] ),
    .A2(\dp.rf.rf[26][26] ),
    .A3(\dp.rf.rf[27][26] ),
    .S0(net826),
    .S1(net820),
    .X(_0583_));
 sky130_fd_sc_hd__mux4_2 _4151_ (.A0(\dp.rf.rf[20][26] ),
    .A1(\dp.rf.rf[21][26] ),
    .A2(\dp.rf.rf[22][26] ),
    .A3(\dp.rf.rf[23][26] ),
    .S0(net826),
    .S1(net820),
    .X(_0584_));
 sky130_fd_sc_hd__mux4_2 _4152_ (.A0(\dp.rf.rf[28][26] ),
    .A1(\dp.rf.rf[29][26] ),
    .A2(\dp.rf.rf[30][26] ),
    .A3(\dp.rf.rf[31][26] ),
    .S0(net826),
    .S1(net820),
    .X(_0585_));
 sky130_fd_sc_hd__mux4_2 _4153_ (.A0(_0581_),
    .A1(_0583_),
    .A2(_0584_),
    .A3(_0585_),
    .S0(net16),
    .S1(net15),
    .X(_0586_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_141 ();
 sky130_fd_sc_hd__nand2_1 _4157_ (.A(net826),
    .B(\dp.rf.rf[1][26] ),
    .Y(_0590_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_140 ();
 sky130_fd_sc_hd__mux2i_1 _4159_ (.A0(\dp.rf.rf[2][26] ),
    .A1(\dp.rf.rf[3][26] ),
    .S(net826),
    .Y(_0592_));
 sky130_fd_sc_hd__mux2i_1 _4160_ (.A0(_0590_),
    .A1(_0592_),
    .S(net820),
    .Y(_0593_));
 sky130_fd_sc_hd__mux4_2 _4161_ (.A0(\dp.rf.rf[4][26] ),
    .A1(\dp.rf.rf[5][26] ),
    .A2(\dp.rf.rf[6][26] ),
    .A3(\dp.rf.rf[7][26] ),
    .S0(net826),
    .S1(net820),
    .X(_0594_));
 sky130_fd_sc_hd__mux4_2 _4162_ (.A0(\dp.rf.rf[8][26] ),
    .A1(\dp.rf.rf[9][26] ),
    .A2(\dp.rf.rf[10][26] ),
    .A3(\dp.rf.rf[11][26] ),
    .S0(net826),
    .S1(net820),
    .X(_0595_));
 sky130_fd_sc_hd__mux4_2 _4163_ (.A0(\dp.rf.rf[12][26] ),
    .A1(\dp.rf.rf[13][26] ),
    .A2(\dp.rf.rf[14][26] ),
    .A3(\dp.rf.rf[15][26] ),
    .S0(net826),
    .S1(net820),
    .X(_0596_));
 sky130_fd_sc_hd__mux4_2 _4164_ (.A0(_0593_),
    .A1(_0594_),
    .A2(_0595_),
    .A3(_0596_),
    .S0(net15),
    .S1(net16),
    .X(_0597_));
 sky130_fd_sc_hd__mux2i_4 _4165_ (.A0(_0586_),
    .A1(_0597_),
    .S(_0092_),
    .Y(_0598_));
 sky130_fd_sc_hd__nand2_1 _4166_ (.A(_0121_),
    .B(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__o21ai_2 _4167_ (.A1(_0121_),
    .A2(_3552_[0]),
    .B1(_0599_),
    .Y(_0600_));
 sky130_fd_sc_hd__xor2_1 _4168_ (.A(_0151_),
    .B(_0600_),
    .X(_3243_[0]));
 sky130_fd_sc_hd__inv_1 _4169_ (.A(_3243_[0]),
    .Y(_3247_[0]));
 sky130_fd_sc_hd__mux4_2 _4170_ (.A0(\dp.rf.rf[10][26] ),
    .A1(\dp.rf.rf[11][26] ),
    .A2(\dp.rf.rf[14][26] ),
    .A3(\dp.rf.rf[15][26] ),
    .S0(net810),
    .S1(net806),
    .X(_0601_));
 sky130_fd_sc_hd__mux4_2 _4171_ (.A0(\dp.rf.rf[8][26] ),
    .A1(\dp.rf.rf[9][26] ),
    .A2(\dp.rf.rf[12][26] ),
    .A3(\dp.rf.rf[13][26] ),
    .S0(net810),
    .S1(net806),
    .X(_0602_));
 sky130_fd_sc_hd__mux2i_2 _4172_ (.A0(_0601_),
    .A1(_0602_),
    .S(_0186_),
    .Y(_0603_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_139 ();
 sky130_fd_sc_hd__mux4_2 _4174_ (.A0(\dp.rf.rf[2][26] ),
    .A1(\dp.rf.rf[3][26] ),
    .A2(\dp.rf.rf[6][26] ),
    .A3(\dp.rf.rf[7][26] ),
    .S0(net810),
    .S1(net806),
    .X(_0605_));
 sky130_fd_sc_hd__inv_1 _4175_ (.A(\dp.rf.rf[4][26] ),
    .Y(_0606_));
 sky130_fd_sc_hd__mux2i_1 _4176_ (.A0(\dp.rf.rf[1][26] ),
    .A1(\dp.rf.rf[5][26] ),
    .S(net806),
    .Y(_0607_));
 sky130_fd_sc_hd__a221oi_1 _4177_ (.A1(_0606_),
    .A2(net801),
    .B1(_0607_),
    .B2(net810),
    .C1(net808),
    .Y(_0608_));
 sky130_fd_sc_hd__a211oi_2 _4178_ (.A1(net808),
    .A2(_0605_),
    .B1(_0608_),
    .C1(net789),
    .Y(_0609_));
 sky130_fd_sc_hd__a211oi_4 _4179_ (.A1(_0193_),
    .A2(_0603_),
    .B1(_0609_),
    .C1(_0293_),
    .Y(_0610_));
 sky130_fd_sc_hd__inv_1 _4180_ (.A(\dp.rf.rf[28][26] ),
    .Y(_0611_));
 sky130_fd_sc_hd__mux2i_1 _4181_ (.A0(\dp.rf.rf[25][26] ),
    .A1(\dp.rf.rf[29][26] ),
    .S(net806),
    .Y(_0612_));
 sky130_fd_sc_hd__a221oi_1 _4182_ (.A1(_0611_),
    .A2(net801),
    .B1(_0612_),
    .B2(net811),
    .C1(net808),
    .Y(_0613_));
 sky130_fd_sc_hd__o21ai_2 _4183_ (.A1(\dp.rf.rf[24][26] ),
    .A2(net798),
    .B1(_0613_),
    .Y(_0614_));
 sky130_fd_sc_hd__mux4_2 _4184_ (.A0(\dp.rf.rf[26][26] ),
    .A1(\dp.rf.rf[27][26] ),
    .A2(\dp.rf.rf[30][26] ),
    .A3(\dp.rf.rf[31][26] ),
    .S0(net811),
    .S1(net806),
    .X(_0615_));
 sky130_fd_sc_hd__a21oi_2 _4185_ (.A1(net786),
    .A2(_0615_),
    .B1(_0192_),
    .Y(_0616_));
 sky130_fd_sc_hd__mux4_2 _4186_ (.A0(\dp.rf.rf[16][26] ),
    .A1(\dp.rf.rf[17][26] ),
    .A2(\dp.rf.rf[20][26] ),
    .A3(\dp.rf.rf[21][26] ),
    .S0(net811),
    .S1(net806),
    .X(_0617_));
 sky130_fd_sc_hd__mux4_2 _4187_ (.A0(\dp.rf.rf[18][26] ),
    .A1(\dp.rf.rf[19][26] ),
    .A2(\dp.rf.rf[22][26] ),
    .A3(\dp.rf.rf[23][26] ),
    .S0(net811),
    .S1(net806),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_1 _4188_ (.A0(_0617_),
    .A1(_0618_),
    .S(net808),
    .X(_0619_));
 sky130_fd_sc_hd__a21oi_4 _4189_ (.A1(_0143_),
    .A2(net802),
    .B1(_0468_),
    .Y(_0620_));
 sky130_fd_sc_hd__o21ai_2 _4190_ (.A1(net10),
    .A2(_0619_),
    .B1(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__a21oi_4 _4191_ (.A1(_0614_),
    .A2(_0616_),
    .B1(_0621_),
    .Y(_0622_));
 sky130_fd_sc_hd__nor2_4 _4192_ (.A(_0610_),
    .B(_0622_),
    .Y(_3246_[0]));
 sky130_fd_sc_hd__a21o_4 _4193_ (.A1(net18),
    .A2(net799),
    .B1(_0349_),
    .X(_3548_[0]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_138 ();
 sky130_fd_sc_hd__mux4_2 _4195_ (.A0(\dp.rf.rf[16][25] ),
    .A1(\dp.rf.rf[17][25] ),
    .A2(\dp.rf.rf[18][25] ),
    .A3(\dp.rf.rf[19][25] ),
    .S0(net825),
    .S1(net819),
    .X(_0624_));
 sky130_fd_sc_hd__mux4_2 _4196_ (.A0(\dp.rf.rf[20][25] ),
    .A1(\dp.rf.rf[21][25] ),
    .A2(\dp.rf.rf[22][25] ),
    .A3(\dp.rf.rf[23][25] ),
    .S0(net825),
    .S1(net819),
    .X(_0625_));
 sky130_fd_sc_hd__mux4_2 _4197_ (.A0(\dp.rf.rf[24][25] ),
    .A1(\dp.rf.rf[25][25] ),
    .A2(\dp.rf.rf[26][25] ),
    .A3(\dp.rf.rf[27][25] ),
    .S0(net825),
    .S1(net819),
    .X(_0626_));
 sky130_fd_sc_hd__mux4_2 _4198_ (.A0(\dp.rf.rf[28][25] ),
    .A1(\dp.rf.rf[29][25] ),
    .A2(\dp.rf.rf[30][25] ),
    .A3(\dp.rf.rf[31][25] ),
    .S0(net825),
    .S1(net819),
    .X(_0627_));
 sky130_fd_sc_hd__mux4_2 _4199_ (.A0(_0624_),
    .A1(_0625_),
    .A2(_0626_),
    .A3(_0627_),
    .S0(net15),
    .S1(net16),
    .X(_0628_));
 sky130_fd_sc_hd__mux4_2 _4200_ (.A0(\dp.rf.rf[0][25] ),
    .A1(\dp.rf.rf[1][25] ),
    .A2(\dp.rf.rf[2][25] ),
    .A3(\dp.rf.rf[3][25] ),
    .S0(net825),
    .S1(net819),
    .X(_0629_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_135 ();
 sky130_fd_sc_hd__mux4_2 _4204_ (.A0(\dp.rf.rf[4][25] ),
    .A1(\dp.rf.rf[5][25] ),
    .A2(\dp.rf.rf[6][25] ),
    .A3(\dp.rf.rf[7][25] ),
    .S0(net825),
    .S1(net819),
    .X(_0633_));
 sky130_fd_sc_hd__mux4_2 _4205_ (.A0(\dp.rf.rf[8][25] ),
    .A1(\dp.rf.rf[9][25] ),
    .A2(\dp.rf.rf[10][25] ),
    .A3(\dp.rf.rf[11][25] ),
    .S0(net825),
    .S1(net819),
    .X(_0634_));
 sky130_fd_sc_hd__mux4_2 _4206_ (.A0(\dp.rf.rf[12][25] ),
    .A1(\dp.rf.rf[13][25] ),
    .A2(\dp.rf.rf[14][25] ),
    .A3(\dp.rf.rf[15][25] ),
    .S0(net825),
    .S1(net819),
    .X(_0635_));
 sky130_fd_sc_hd__mux4_2 _4207_ (.A0(_0629_),
    .A1(_0633_),
    .A2(_0634_),
    .A3(_0635_),
    .S0(net15),
    .S1(net16),
    .X(_0636_));
 sky130_fd_sc_hd__a22o_4 _4208_ (.A1(net17),
    .A2(_0628_),
    .B1(_0636_),
    .B2(_0337_),
    .X(_0637_));
 sky130_fd_sc_hd__mux2_1 _4209_ (.A0(_3548_[0]),
    .A1(_0637_),
    .S(_0121_),
    .X(_0638_));
 sky130_fd_sc_hd__xnor2_1 _4210_ (.A(_0151_),
    .B(_0638_),
    .Y(_3251_[0]));
 sky130_fd_sc_hd__inv_1 _4211_ (.A(_3251_[0]),
    .Y(_3255_[0]));
 sky130_fd_sc_hd__mux4_2 _4212_ (.A0(\dp.rf.rf[10][25] ),
    .A1(\dp.rf.rf[11][25] ),
    .A2(\dp.rf.rf[14][25] ),
    .A3(\dp.rf.rf[15][25] ),
    .S0(net811),
    .S1(net807),
    .X(_0639_));
 sky130_fd_sc_hd__nand2_1 _4213_ (.A(net808),
    .B(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__mux4_2 _4214_ (.A0(\dp.rf.rf[8][25] ),
    .A1(\dp.rf.rf[9][25] ),
    .A2(\dp.rf.rf[12][25] ),
    .A3(\dp.rf.rf[13][25] ),
    .S0(net811),
    .S1(net807),
    .X(_0641_));
 sky130_fd_sc_hd__nand2_1 _4215_ (.A(_0186_),
    .B(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__nand3_2 _4216_ (.A(net796),
    .B(_0640_),
    .C(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__mux2_1 _4217_ (.A0(\dp.rf.rf[6][25] ),
    .A1(\dp.rf.rf[7][25] ),
    .S(net811),
    .X(_0644_));
 sky130_fd_sc_hd__o21ai_0 _4218_ (.A1(net800),
    .A2(_0644_),
    .B1(net786),
    .Y(_0645_));
 sky130_fd_sc_hd__a221oi_1 _4219_ (.A1(\dp.rf.rf[3][25] ),
    .A2(net811),
    .B1(net787),
    .B2(\dp.rf.rf[2][25] ),
    .C1(net792),
    .Y(_0646_));
 sky130_fd_sc_hd__inv_1 _4220_ (.A(\dp.rf.rf[4][25] ),
    .Y(_0647_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_134 ();
 sky130_fd_sc_hd__mux2i_1 _4222_ (.A0(\dp.rf.rf[1][25] ),
    .A1(\dp.rf.rf[5][25] ),
    .S(net807),
    .Y(_0649_));
 sky130_fd_sc_hd__a221oi_1 _4223_ (.A1(_0647_),
    .A2(net801),
    .B1(_0649_),
    .B2(net811),
    .C1(net808),
    .Y(_0650_));
 sky130_fd_sc_hd__o22ai_1 _4224_ (.A1(\dp.rf.rf[0][25] ),
    .A2(_0412_),
    .B1(_0650_),
    .B2(net789),
    .Y(_0651_));
 sky130_fd_sc_hd__o21ai_2 _4225_ (.A1(_0645_),
    .A2(_0646_),
    .B1(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__inv_1 _4226_ (.A(\dp.rf.rf[28][25] ),
    .Y(_0653_));
 sky130_fd_sc_hd__mux2i_1 _4227_ (.A0(\dp.rf.rf[25][25] ),
    .A1(\dp.rf.rf[29][25] ),
    .S(net806),
    .Y(_0654_));
 sky130_fd_sc_hd__a221oi_1 _4228_ (.A1(_0653_),
    .A2(net801),
    .B1(_0654_),
    .B2(net811),
    .C1(net808),
    .Y(_0655_));
 sky130_fd_sc_hd__o21ai_0 _4229_ (.A1(\dp.rf.rf[24][25] ),
    .A2(net798),
    .B1(_0655_),
    .Y(_0656_));
 sky130_fd_sc_hd__mux4_2 _4230_ (.A0(\dp.rf.rf[26][25] ),
    .A1(\dp.rf.rf[27][25] ),
    .A2(\dp.rf.rf[30][25] ),
    .A3(\dp.rf.rf[31][25] ),
    .S0(net811),
    .S1(net806),
    .X(_0657_));
 sky130_fd_sc_hd__a21oi_1 _4231_ (.A1(net786),
    .A2(_0657_),
    .B1(_0192_),
    .Y(_0658_));
 sky130_fd_sc_hd__mux4_2 _4232_ (.A0(\dp.rf.rf[18][25] ),
    .A1(\dp.rf.rf[19][25] ),
    .A2(\dp.rf.rf[22][25] ),
    .A3(\dp.rf.rf[23][25] ),
    .S0(net811),
    .S1(net806),
    .X(_0659_));
 sky130_fd_sc_hd__or2_0 _4233_ (.A(net811),
    .B(net806),
    .X(_0660_));
 sky130_fd_sc_hd__a211o_1 _4234_ (.A1(net808),
    .A2(_0659_),
    .B1(_0660_),
    .C1(net10),
    .X(_0661_));
 sky130_fd_sc_hd__a21oi_1 _4235_ (.A1(_0347_),
    .A2(_0661_),
    .B1(\dp.rf.rf[16][25] ),
    .Y(_0662_));
 sky130_fd_sc_hd__inv_1 _4236_ (.A(\dp.rf.rf[20][25] ),
    .Y(_0663_));
 sky130_fd_sc_hd__mux2i_1 _4237_ (.A0(\dp.rf.rf[17][25] ),
    .A1(\dp.rf.rf[21][25] ),
    .S(net806),
    .Y(_0664_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_133 ();
 sky130_fd_sc_hd__a221oi_1 _4239_ (.A1(_0663_),
    .A2(net801),
    .B1(_0664_),
    .B2(net811),
    .C1(net808),
    .Y(_0666_));
 sky130_fd_sc_hd__a211oi_1 _4240_ (.A1(net808),
    .A2(_0659_),
    .B1(_0666_),
    .C1(net10),
    .Y(_0667_));
 sky130_fd_sc_hd__a2111oi_2 _4241_ (.A1(_0656_),
    .A2(_0658_),
    .B1(net795),
    .C1(_0662_),
    .D1(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__a31oi_4 _4242_ (.A1(_0185_),
    .A2(_0643_),
    .A3(_0652_),
    .B1(_0668_),
    .Y(_3254_[0]));
 sky130_fd_sc_hd__nor2b_4 _4243_ (.A(net818),
    .B_N(net817),
    .Y(_0669_));
 sky130_fd_sc_hd__mux4_2 _4244_ (.A0(\dp.rf.rf[8][24] ),
    .A1(\dp.rf.rf[9][24] ),
    .A2(\dp.rf.rf[10][24] ),
    .A3(\dp.rf.rf[11][24] ),
    .S0(net826),
    .S1(net820),
    .X(_0670_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_131 ();
 sky130_fd_sc_hd__mux4_2 _4247_ (.A0(\dp.rf.rf[0][24] ),
    .A1(\dp.rf.rf[1][24] ),
    .A2(\dp.rf.rf[2][24] ),
    .A3(\dp.rf.rf[3][24] ),
    .S0(net826),
    .S1(net820),
    .X(_0673_));
 sky130_fd_sc_hd__nor2_4 _4248_ (.A(net818),
    .B(net817),
    .Y(_0674_));
 sky130_fd_sc_hd__a22oi_1 _4249_ (.A1(_0669_),
    .A2(_0670_),
    .B1(_0673_),
    .B2(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__and2_4 _4250_ (.A(net818),
    .B(net817),
    .X(_0676_));
 sky130_fd_sc_hd__mux4_2 _4251_ (.A0(\dp.rf.rf[12][24] ),
    .A1(\dp.rf.rf[13][24] ),
    .A2(\dp.rf.rf[14][24] ),
    .A3(\dp.rf.rf[15][24] ),
    .S0(net826),
    .S1(net820),
    .X(_0677_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_130 ();
 sky130_fd_sc_hd__mux4_2 _4253_ (.A0(\dp.rf.rf[4][24] ),
    .A1(\dp.rf.rf[5][24] ),
    .A2(\dp.rf.rf[6][24] ),
    .A3(\dp.rf.rf[7][24] ),
    .S0(net826),
    .S1(net820),
    .X(_0679_));
 sky130_fd_sc_hd__nor2b_4 _4254_ (.A(net817),
    .B_N(net818),
    .Y(_0680_));
 sky130_fd_sc_hd__a22oi_1 _4255_ (.A1(_0676_),
    .A2(_0677_),
    .B1(_0679_),
    .B2(_0680_),
    .Y(_0681_));
 sky130_fd_sc_hd__nand2_1 _4256_ (.A(_0675_),
    .B(_0681_),
    .Y(_0682_));
 sky130_fd_sc_hd__mux4_2 _4257_ (.A0(\dp.rf.rf[16][24] ),
    .A1(\dp.rf.rf[17][24] ),
    .A2(\dp.rf.rf[18][24] ),
    .A3(\dp.rf.rf[19][24] ),
    .S0(net826),
    .S1(net820),
    .X(_0683_));
 sky130_fd_sc_hd__mux4_2 _4258_ (.A0(\dp.rf.rf[24][24] ),
    .A1(\dp.rf.rf[25][24] ),
    .A2(\dp.rf.rf[26][24] ),
    .A3(\dp.rf.rf[27][24] ),
    .S0(net826),
    .S1(net820),
    .X(_0684_));
 sky130_fd_sc_hd__a22oi_1 _4259_ (.A1(_0683_),
    .A2(_0674_),
    .B1(_0669_),
    .B2(_0684_),
    .Y(_0685_));
 sky130_fd_sc_hd__mux4_2 _4260_ (.A0(\dp.rf.rf[20][24] ),
    .A1(\dp.rf.rf[21][24] ),
    .A2(\dp.rf.rf[22][24] ),
    .A3(\dp.rf.rf[23][24] ),
    .S0(net826),
    .S1(net820),
    .X(_0686_));
 sky130_fd_sc_hd__mux4_2 _4261_ (.A0(\dp.rf.rf[28][24] ),
    .A1(\dp.rf.rf[29][24] ),
    .A2(\dp.rf.rf[30][24] ),
    .A3(\dp.rf.rf[31][24] ),
    .S0(net826),
    .S1(net820),
    .X(_0687_));
 sky130_fd_sc_hd__a22oi_1 _4262_ (.A1(_0686_),
    .A2(_0680_),
    .B1(_0676_),
    .B2(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__a21oi_1 _4263_ (.A1(_0685_),
    .A2(_0688_),
    .B1(_0092_),
    .Y(_0689_));
 sky130_fd_sc_hd__a21oi_2 _4264_ (.A1(_0337_),
    .A2(_0682_),
    .B1(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__a21o_4 _4265_ (.A1(net17),
    .A2(net799),
    .B1(_0349_),
    .X(_3544_[0]));
 sky130_fd_sc_hd__nor2_1 _4266_ (.A(_0121_),
    .B(_3544_[0]),
    .Y(_0691_));
 sky130_fd_sc_hd__a21oi_1 _4267_ (.A1(_0121_),
    .A2(_0690_),
    .B1(_0691_),
    .Y(_0692_));
 sky130_fd_sc_hd__xnor2_1 _4268_ (.A(_0151_),
    .B(_0692_),
    .Y(_3259_[0]));
 sky130_fd_sc_hd__inv_1 _4269_ (.A(_3259_[0]),
    .Y(_3263_[0]));
 sky130_fd_sc_hd__nand2_1 _4270_ (.A(\dp.rf.rf[2][24] ),
    .B(net808),
    .Y(_0693_));
 sky130_fd_sc_hd__nand2_1 _4271_ (.A(_0386_),
    .B(_0693_),
    .Y(_0694_));
 sky130_fd_sc_hd__a21oi_1 _4272_ (.A1(_0347_),
    .A2(_0694_),
    .B1(\dp.rf.rf[0][24] ),
    .Y(_0695_));
 sky130_fd_sc_hd__mux4_2 _4273_ (.A0(\dp.rf.rf[10][24] ),
    .A1(\dp.rf.rf[11][24] ),
    .A2(\dp.rf.rf[14][24] ),
    .A3(\dp.rf.rf[15][24] ),
    .S0(net810),
    .S1(net806),
    .X(_0696_));
 sky130_fd_sc_hd__nand2_1 _4274_ (.A(net808),
    .B(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__mux4_2 _4275_ (.A0(\dp.rf.rf[8][24] ),
    .A1(\dp.rf.rf[9][24] ),
    .A2(\dp.rf.rf[12][24] ),
    .A3(\dp.rf.rf[13][24] ),
    .S0(net810),
    .S1(net806),
    .X(_0698_));
 sky130_fd_sc_hd__nand2_1 _4276_ (.A(_0186_),
    .B(_0698_),
    .Y(_0699_));
 sky130_fd_sc_hd__and3_4 _4277_ (.A(_0193_),
    .B(_0697_),
    .C(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__mux4_2 _4278_ (.A0(\dp.rf.rf[2][24] ),
    .A1(\dp.rf.rf[3][24] ),
    .A2(\dp.rf.rf[6][24] ),
    .A3(\dp.rf.rf[7][24] ),
    .S0(net810),
    .S1(net805),
    .X(_0701_));
 sky130_fd_sc_hd__inv_1 _4279_ (.A(\dp.rf.rf[4][24] ),
    .Y(_0702_));
 sky130_fd_sc_hd__mux2i_1 _4280_ (.A0(\dp.rf.rf[1][24] ),
    .A1(\dp.rf.rf[5][24] ),
    .S(net805),
    .Y(_0703_));
 sky130_fd_sc_hd__a221oi_1 _4281_ (.A1(_0702_),
    .A2(net801),
    .B1(_0703_),
    .B2(net810),
    .C1(net808),
    .Y(_0704_));
 sky130_fd_sc_hd__a211oi_1 _4282_ (.A1(net808),
    .A2(_0701_),
    .B1(_0704_),
    .C1(net789),
    .Y(_0705_));
 sky130_fd_sc_hd__nor4_2 _4283_ (.A(_0293_),
    .B(_0695_),
    .C(_0700_),
    .D(_0705_),
    .Y(_0706_));
 sky130_fd_sc_hd__inv_1 _4284_ (.A(\dp.rf.rf[28][24] ),
    .Y(_0707_));
 sky130_fd_sc_hd__mux2i_1 _4285_ (.A0(\dp.rf.rf[25][24] ),
    .A1(\dp.rf.rf[29][24] ),
    .S(net805),
    .Y(_0708_));
 sky130_fd_sc_hd__a221oi_1 _4286_ (.A1(_0707_),
    .A2(net801),
    .B1(_0708_),
    .B2(net810),
    .C1(net808),
    .Y(_0709_));
 sky130_fd_sc_hd__o21ai_0 _4287_ (.A1(\dp.rf.rf[24][24] ),
    .A2(net798),
    .B1(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_129 ();
 sky130_fd_sc_hd__mux4_2 _4289_ (.A0(\dp.rf.rf[26][24] ),
    .A1(\dp.rf.rf[27][24] ),
    .A2(\dp.rf.rf[30][24] ),
    .A3(\dp.rf.rf[31][24] ),
    .S0(net810),
    .S1(net805),
    .X(_0712_));
 sky130_fd_sc_hd__nand2_1 _4290_ (.A(net786),
    .B(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__nand2_1 _4291_ (.A(net808),
    .B(_0192_),
    .Y(_0714_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_128 ();
 sky130_fd_sc_hd__mux4_2 _4293_ (.A0(\dp.rf.rf[18][24] ),
    .A1(\dp.rf.rf[19][24] ),
    .A2(\dp.rf.rf[22][24] ),
    .A3(\dp.rf.rf[23][24] ),
    .S0(net810),
    .S1(net805),
    .X(_0716_));
 sky130_fd_sc_hd__mux4_2 _4294_ (.A0(\dp.rf.rf[16][24] ),
    .A1(\dp.rf.rf[17][24] ),
    .A2(\dp.rf.rf[20][24] ),
    .A3(\dp.rf.rf[21][24] ),
    .S0(net810),
    .S1(net805),
    .X(_0717_));
 sky130_fd_sc_hd__o22ai_1 _4295_ (.A1(_0714_),
    .A2(_0716_),
    .B1(_0717_),
    .B2(_0179_),
    .Y(_0718_));
 sky130_fd_sc_hd__a311oi_2 _4296_ (.A1(net10),
    .A2(_0710_),
    .A3(_0713_),
    .B1(_0718_),
    .C1(_0224_),
    .Y(_0719_));
 sky130_fd_sc_hd__nor2_4 _4297_ (.A(_0706_),
    .B(_0719_),
    .Y(_3262_[0]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_127 ();
 sky130_fd_sc_hd__mux4_2 _4299_ (.A0(\dp.rf.rf[16][23] ),
    .A1(\dp.rf.rf[17][23] ),
    .A2(\dp.rf.rf[18][23] ),
    .A3(\dp.rf.rf[19][23] ),
    .S0(net825),
    .S1(net819),
    .X(_0721_));
 sky130_fd_sc_hd__mux4_2 _4300_ (.A0(\dp.rf.rf[20][23] ),
    .A1(\dp.rf.rf[21][23] ),
    .A2(\dp.rf.rf[22][23] ),
    .A3(\dp.rf.rf[23][23] ),
    .S0(net825),
    .S1(net819),
    .X(_0722_));
 sky130_fd_sc_hd__mux4_2 _4301_ (.A0(\dp.rf.rf[24][23] ),
    .A1(\dp.rf.rf[25][23] ),
    .A2(\dp.rf.rf[26][23] ),
    .A3(\dp.rf.rf[27][23] ),
    .S0(net825),
    .S1(net819),
    .X(_0723_));
 sky130_fd_sc_hd__mux4_2 _4302_ (.A0(\dp.rf.rf[28][23] ),
    .A1(\dp.rf.rf[29][23] ),
    .A2(\dp.rf.rf[30][23] ),
    .A3(\dp.rf.rf[31][23] ),
    .S0(net825),
    .S1(net819),
    .X(_0724_));
 sky130_fd_sc_hd__mux4_2 _4303_ (.A0(_0721_),
    .A1(_0722_),
    .A2(_0723_),
    .A3(_0724_),
    .S0(net15),
    .S1(net817),
    .X(_0725_));
 sky130_fd_sc_hd__mux4_2 _4304_ (.A0(\dp.rf.rf[0][23] ),
    .A1(\dp.rf.rf[1][23] ),
    .A2(\dp.rf.rf[2][23] ),
    .A3(\dp.rf.rf[3][23] ),
    .S0(net13),
    .S1(net14),
    .X(_0726_));
 sky130_fd_sc_hd__mux4_2 _4305_ (.A0(\dp.rf.rf[4][23] ),
    .A1(\dp.rf.rf[5][23] ),
    .A2(\dp.rf.rf[6][23] ),
    .A3(\dp.rf.rf[7][23] ),
    .S0(net13),
    .S1(net14),
    .X(_0727_));
 sky130_fd_sc_hd__mux4_2 _4306_ (.A0(\dp.rf.rf[8][23] ),
    .A1(\dp.rf.rf[9][23] ),
    .A2(\dp.rf.rf[10][23] ),
    .A3(\dp.rf.rf[11][23] ),
    .S0(net13),
    .S1(net14),
    .X(_0728_));
 sky130_fd_sc_hd__mux4_2 _4307_ (.A0(\dp.rf.rf[12][23] ),
    .A1(\dp.rf.rf[13][23] ),
    .A2(\dp.rf.rf[14][23] ),
    .A3(\dp.rf.rf[15][23] ),
    .S0(net13),
    .S1(net14),
    .X(_0729_));
 sky130_fd_sc_hd__mux4_2 _4308_ (.A0(_0726_),
    .A1(_0727_),
    .A2(_0728_),
    .A3(_0729_),
    .S0(net15),
    .S1(net16),
    .X(_0730_));
 sky130_fd_sc_hd__a22o_4 _4309_ (.A1(net17),
    .A2(_0725_),
    .B1(_0730_),
    .B2(_0337_),
    .X(_0731_));
 sky130_fd_sc_hd__inv_6 _4310_ (.A(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__a21o_1 _4311_ (.A1(net817),
    .A2(net799),
    .B1(_0349_),
    .X(_3540_[0]));
 sky130_fd_sc_hd__nand2_1 _4312_ (.A(net782),
    .B(_3540_[0]),
    .Y(_0733_));
 sky130_fd_sc_hd__o21ai_0 _4313_ (.A1(net782),
    .A2(_0732_),
    .B1(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__xnor2_1 _4314_ (.A(_0151_),
    .B(_0734_),
    .Y(_3267_[0]));
 sky130_fd_sc_hd__inv_1 _4315_ (.A(_3267_[0]),
    .Y(_3271_[0]));
 sky130_fd_sc_hd__mux4_2 _4316_ (.A0(\dp.rf.rf[2][23] ),
    .A1(\dp.rf.rf[3][23] ),
    .A2(\dp.rf.rf[6][23] ),
    .A3(\dp.rf.rf[7][23] ),
    .S0(net813),
    .S1(net807),
    .X(_0735_));
 sky130_fd_sc_hd__nand2_1 _4317_ (.A(net808),
    .B(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__mux2_1 _4318_ (.A0(\dp.rf.rf[1][23] ),
    .A1(\dp.rf.rf[5][23] ),
    .S(net807),
    .X(_0737_));
 sky130_fd_sc_hd__o221ai_1 _4319_ (.A1(\dp.rf.rf[4][23] ),
    .A2(_0395_),
    .B1(_0737_),
    .B2(_0400_),
    .C1(_0186_),
    .Y(_0738_));
 sky130_fd_sc_hd__nand3_2 _4320_ (.A(net785),
    .B(_0736_),
    .C(_0738_),
    .Y(_0739_));
 sky130_fd_sc_hd__mux4_2 _4321_ (.A0(\dp.rf.rf[10][23] ),
    .A1(\dp.rf.rf[11][23] ),
    .A2(\dp.rf.rf[14][23] ),
    .A3(\dp.rf.rf[15][23] ),
    .S0(net813),
    .S1(net807),
    .X(_0740_));
 sky130_fd_sc_hd__nand2_1 _4322_ (.A(net808),
    .B(_0740_),
    .Y(_0741_));
 sky130_fd_sc_hd__mux4_2 _4323_ (.A0(\dp.rf.rf[8][23] ),
    .A1(\dp.rf.rf[9][23] ),
    .A2(\dp.rf.rf[12][23] ),
    .A3(\dp.rf.rf[13][23] ),
    .S0(net813),
    .S1(net807),
    .X(_0742_));
 sky130_fd_sc_hd__nand2_1 _4324_ (.A(_0186_),
    .B(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__nand3_2 _4325_ (.A(net796),
    .B(_0741_),
    .C(_0743_),
    .Y(_0744_));
 sky130_fd_sc_hd__nand4_1 _4326_ (.A(net1),
    .B(net12),
    .C(net23),
    .D(net297),
    .Y(_0745_));
 sky130_fd_sc_hd__o2bb2ai_4 _4327_ (.A1_N(net297),
    .A2_N(_0400_),
    .B1(_0135_),
    .B2(_0745_),
    .Y(_0746_));
 sky130_fd_sc_hd__and2_0 _4328_ (.A(\dp.rf.rf[27][23] ),
    .B(net811),
    .X(_0747_));
 sky130_fd_sc_hd__mux2i_1 _4329_ (.A0(\dp.rf.rf[30][23] ),
    .A1(\dp.rf.rf[31][23] ),
    .S(net811),
    .Y(_0748_));
 sky130_fd_sc_hd__nand2_1 _4330_ (.A(net807),
    .B(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__o311ai_0 _4331_ (.A1(net792),
    .A2(_0746_),
    .A3(_0747_),
    .B1(net786),
    .C1(_0749_),
    .Y(_0750_));
 sky130_fd_sc_hd__inv_1 _4332_ (.A(\dp.rf.rf[28][23] ),
    .Y(_0751_));
 sky130_fd_sc_hd__mux2i_1 _4333_ (.A0(\dp.rf.rf[25][23] ),
    .A1(\dp.rf.rf[29][23] ),
    .S(net807),
    .Y(_0752_));
 sky130_fd_sc_hd__a221oi_1 _4334_ (.A1(_0751_),
    .A2(net801),
    .B1(_0752_),
    .B2(net811),
    .C1(net808),
    .Y(_0753_));
 sky130_fd_sc_hd__o21ai_0 _4335_ (.A1(\dp.rf.rf[24][23] ),
    .A2(net798),
    .B1(_0753_),
    .Y(_0754_));
 sky130_fd_sc_hd__a31oi_1 _4336_ (.A1(net796),
    .A2(_0750_),
    .A3(_0754_),
    .B1(net795),
    .Y(_0755_));
 sky130_fd_sc_hd__mux2_1 _4337_ (.A0(\dp.rf.rf[22][23] ),
    .A1(\dp.rf.rf[23][23] ),
    .S(net811),
    .X(_0756_));
 sky130_fd_sc_hd__o21ai_0 _4338_ (.A1(net800),
    .A2(_0756_),
    .B1(net786),
    .Y(_0757_));
 sky130_fd_sc_hd__a221oi_1 _4339_ (.A1(\dp.rf.rf[19][23] ),
    .A2(net811),
    .B1(net787),
    .B2(\dp.rf.rf[18][23] ),
    .C1(net792),
    .Y(_0758_));
 sky130_fd_sc_hd__inv_1 _4340_ (.A(\dp.rf.rf[20][23] ),
    .Y(_0759_));
 sky130_fd_sc_hd__mux2i_1 _4341_ (.A0(\dp.rf.rf[17][23] ),
    .A1(\dp.rf.rf[21][23] ),
    .S(net806),
    .Y(_0760_));
 sky130_fd_sc_hd__a221oi_1 _4342_ (.A1(_0759_),
    .A2(net801),
    .B1(_0760_),
    .B2(net811),
    .C1(net808),
    .Y(_0761_));
 sky130_fd_sc_hd__o22ai_1 _4343_ (.A1(\dp.rf.rf[16][23] ),
    .A2(_0412_),
    .B1(_0761_),
    .B2(net789),
    .Y(_0762_));
 sky130_fd_sc_hd__o21ai_2 _4344_ (.A1(_0757_),
    .A2(_0758_),
    .B1(_0762_),
    .Y(_0763_));
 sky130_fd_sc_hd__a32oi_4 _4345_ (.A1(_0185_),
    .A2(_0739_),
    .A3(_0744_),
    .B1(_0755_),
    .B2(_0763_),
    .Y(_3270_[0]));
 sky130_fd_sc_hd__a21o_4 _4346_ (.A1(net818),
    .A2(net799),
    .B1(_0349_),
    .X(_3536_[0]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_126 ();
 sky130_fd_sc_hd__mux4_2 _4348_ (.A0(\dp.rf.rf[16][22] ),
    .A1(\dp.rf.rf[17][22] ),
    .A2(\dp.rf.rf[18][22] ),
    .A3(\dp.rf.rf[19][22] ),
    .S0(net825),
    .S1(net819),
    .X(_0765_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_124 ();
 sky130_fd_sc_hd__mux4_2 _4351_ (.A0(\dp.rf.rf[20][22] ),
    .A1(\dp.rf.rf[21][22] ),
    .A2(\dp.rf.rf[22][22] ),
    .A3(\dp.rf.rf[23][22] ),
    .S0(net825),
    .S1(net819),
    .X(_0768_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_122 ();
 sky130_fd_sc_hd__mux4_2 _4354_ (.A0(\dp.rf.rf[24][22] ),
    .A1(\dp.rf.rf[25][22] ),
    .A2(\dp.rf.rf[26][22] ),
    .A3(\dp.rf.rf[27][22] ),
    .S0(net825),
    .S1(net819),
    .X(_0771_));
 sky130_fd_sc_hd__mux4_2 _4355_ (.A0(\dp.rf.rf[28][22] ),
    .A1(\dp.rf.rf[29][22] ),
    .A2(\dp.rf.rf[30][22] ),
    .A3(\dp.rf.rf[31][22] ),
    .S0(net825),
    .S1(net819),
    .X(_0772_));
 sky130_fd_sc_hd__mux4_2 _4356_ (.A0(_0765_),
    .A1(_0768_),
    .A2(_0771_),
    .A3(_0772_),
    .S0(net15),
    .S1(net817),
    .X(_0773_));
 sky130_fd_sc_hd__nand2_2 _4357_ (.A(net17),
    .B(_0773_),
    .Y(_0774_));
 sky130_fd_sc_hd__mux4_2 _4358_ (.A0(\dp.rf.rf[0][22] ),
    .A1(\dp.rf.rf[1][22] ),
    .A2(\dp.rf.rf[2][22] ),
    .A3(\dp.rf.rf[3][22] ),
    .S0(net825),
    .S1(net819),
    .X(_0775_));
 sky130_fd_sc_hd__mux4_2 _4359_ (.A0(\dp.rf.rf[4][22] ),
    .A1(\dp.rf.rf[5][22] ),
    .A2(\dp.rf.rf[6][22] ),
    .A3(\dp.rf.rf[7][22] ),
    .S0(net825),
    .S1(net819),
    .X(_0776_));
 sky130_fd_sc_hd__mux4_2 _4360_ (.A0(\dp.rf.rf[8][22] ),
    .A1(\dp.rf.rf[9][22] ),
    .A2(\dp.rf.rf[10][22] ),
    .A3(\dp.rf.rf[11][22] ),
    .S0(net825),
    .S1(net819),
    .X(_0777_));
 sky130_fd_sc_hd__mux4_2 _4361_ (.A0(\dp.rf.rf[12][22] ),
    .A1(\dp.rf.rf[13][22] ),
    .A2(\dp.rf.rf[14][22] ),
    .A3(\dp.rf.rf[15][22] ),
    .S0(net825),
    .S1(net819),
    .X(_0778_));
 sky130_fd_sc_hd__mux4_2 _4362_ (.A0(_0775_),
    .A1(_0776_),
    .A2(_0777_),
    .A3(_0778_),
    .S0(net15),
    .S1(net16),
    .X(_0779_));
 sky130_fd_sc_hd__nand2_4 _4363_ (.A(_0092_),
    .B(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__nand2_4 _4364_ (.A(_0774_),
    .B(_0780_),
    .Y(_0781_));
 sky130_fd_sc_hd__nand2_4 _4365_ (.A(_0351_),
    .B(_0781_),
    .Y(_0782_));
 sky130_fd_sc_hd__nor2_1 _4366_ (.A(net782),
    .B(_0782_),
    .Y(_0783_));
 sky130_fd_sc_hd__a21oi_2 _4367_ (.A1(net782),
    .A2(_3536_[0]),
    .B1(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__xor2_1 _4368_ (.A(_0151_),
    .B(_0784_),
    .X(_3275_[0]));
 sky130_fd_sc_hd__inv_1 _4369_ (.A(_3275_[0]),
    .Y(_3279_[0]));
 sky130_fd_sc_hd__nor2b_1 _4370_ (.A(net812),
    .B_N(\dp.rf.rf[30][22] ),
    .Y(_0785_));
 sky130_fd_sc_hd__a211oi_1 _4371_ (.A1(\dp.rf.rf[31][22] ),
    .A2(net812),
    .B1(net800),
    .C1(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_121 ();
 sky130_fd_sc_hd__a221oi_1 _4373_ (.A1(\dp.rf.rf[27][22] ),
    .A2(net812),
    .B1(net787),
    .B2(\dp.rf.rf[26][22] ),
    .C1(net792),
    .Y(_0788_));
 sky130_fd_sc_hd__inv_1 _4374_ (.A(\dp.rf.rf[28][22] ),
    .Y(_0789_));
 sky130_fd_sc_hd__mux2i_1 _4375_ (.A0(\dp.rf.rf[25][22] ),
    .A1(\dp.rf.rf[29][22] ),
    .S(net806),
    .Y(_0790_));
 sky130_fd_sc_hd__a221oi_1 _4376_ (.A1(_0789_),
    .A2(net801),
    .B1(_0790_),
    .B2(net812),
    .C1(net808),
    .Y(_0791_));
 sky130_fd_sc_hd__o21ai_0 _4377_ (.A1(\dp.rf.rf[24][22] ),
    .A2(net798),
    .B1(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__o311ai_1 _4378_ (.A1(_0477_),
    .A2(_0786_),
    .A3(_0788_),
    .B1(_0792_),
    .C1(net796),
    .Y(_0793_));
 sky130_fd_sc_hd__mux2_1 _4379_ (.A0(\dp.rf.rf[22][22] ),
    .A1(\dp.rf.rf[23][22] ),
    .S(net812),
    .X(_0794_));
 sky130_fd_sc_hd__o21ai_0 _4380_ (.A1(net800),
    .A2(_0794_),
    .B1(net786),
    .Y(_0795_));
 sky130_fd_sc_hd__a221oi_1 _4381_ (.A1(\dp.rf.rf[19][22] ),
    .A2(net812),
    .B1(net787),
    .B2(\dp.rf.rf[18][22] ),
    .C1(net792),
    .Y(_0796_));
 sky130_fd_sc_hd__inv_1 _4382_ (.A(\dp.rf.rf[20][22] ),
    .Y(_0797_));
 sky130_fd_sc_hd__mux2i_1 _4383_ (.A0(\dp.rf.rf[17][22] ),
    .A1(\dp.rf.rf[21][22] ),
    .S(net805),
    .Y(_0798_));
 sky130_fd_sc_hd__a221oi_1 _4384_ (.A1(_0797_),
    .A2(net801),
    .B1(_0798_),
    .B2(net812),
    .C1(net808),
    .Y(_0799_));
 sky130_fd_sc_hd__o22ai_1 _4385_ (.A1(\dp.rf.rf[16][22] ),
    .A2(_0412_),
    .B1(_0799_),
    .B2(net789),
    .Y(_0800_));
 sky130_fd_sc_hd__o21ai_2 _4386_ (.A1(_0795_),
    .A2(_0796_),
    .B1(_0800_),
    .Y(_0801_));
 sky130_fd_sc_hd__mux4_2 _4387_ (.A0(\dp.rf.rf[10][22] ),
    .A1(\dp.rf.rf[11][22] ),
    .A2(\dp.rf.rf[14][22] ),
    .A3(\dp.rf.rf[15][22] ),
    .S0(net813),
    .S1(net806),
    .X(_0802_));
 sky130_fd_sc_hd__mux4_2 _4388_ (.A0(\dp.rf.rf[8][22] ),
    .A1(\dp.rf.rf[9][22] ),
    .A2(\dp.rf.rf[12][22] ),
    .A3(\dp.rf.rf[13][22] ),
    .S0(net813),
    .S1(net806),
    .X(_0803_));
 sky130_fd_sc_hd__mux2i_1 _4389_ (.A0(_0802_),
    .A1(_0803_),
    .S(_0186_),
    .Y(_0804_));
 sky130_fd_sc_hd__mux4_2 _4390_ (.A0(\dp.rf.rf[2][22] ),
    .A1(\dp.rf.rf[3][22] ),
    .A2(\dp.rf.rf[6][22] ),
    .A3(\dp.rf.rf[7][22] ),
    .S0(net813),
    .S1(net806),
    .X(_0805_));
 sky130_fd_sc_hd__inv_1 _4391_ (.A(\dp.rf.rf[4][22] ),
    .Y(_0806_));
 sky130_fd_sc_hd__mux2i_1 _4392_ (.A0(\dp.rf.rf[1][22] ),
    .A1(\dp.rf.rf[5][22] ),
    .S(net806),
    .Y(_0807_));
 sky130_fd_sc_hd__a221oi_1 _4393_ (.A1(_0806_),
    .A2(net801),
    .B1(_0807_),
    .B2(net813),
    .C1(net808),
    .Y(_0808_));
 sky130_fd_sc_hd__a211oi_1 _4394_ (.A1(net808),
    .A2(_0805_),
    .B1(_0808_),
    .C1(net789),
    .Y(_0809_));
 sky130_fd_sc_hd__a211oi_2 _4395_ (.A1(net796),
    .A2(_0804_),
    .B1(_0809_),
    .C1(_0293_),
    .Y(_0810_));
 sky130_fd_sc_hd__a31oi_4 _4396_ (.A1(net783),
    .A2(_0793_),
    .A3(_0801_),
    .B1(_0810_),
    .Y(_3278_[0]));
 sky130_fd_sc_hd__mux4_2 _4397_ (.A0(\dp.rf.rf[16][21] ),
    .A1(\dp.rf.rf[17][21] ),
    .A2(\dp.rf.rf[18][21] ),
    .A3(\dp.rf.rf[19][21] ),
    .S0(net825),
    .S1(net819),
    .X(_0811_));
 sky130_fd_sc_hd__mux4_2 _4398_ (.A0(\dp.rf.rf[20][21] ),
    .A1(\dp.rf.rf[21][21] ),
    .A2(\dp.rf.rf[22][21] ),
    .A3(\dp.rf.rf[23][21] ),
    .S0(net825),
    .S1(net819),
    .X(_0812_));
 sky130_fd_sc_hd__mux4_2 _4399_ (.A0(\dp.rf.rf[24][21] ),
    .A1(\dp.rf.rf[25][21] ),
    .A2(\dp.rf.rf[26][21] ),
    .A3(\dp.rf.rf[27][21] ),
    .S0(net825),
    .S1(net819),
    .X(_0813_));
 sky130_fd_sc_hd__mux4_2 _4400_ (.A0(\dp.rf.rf[28][21] ),
    .A1(\dp.rf.rf[29][21] ),
    .A2(\dp.rf.rf[30][21] ),
    .A3(\dp.rf.rf[31][21] ),
    .S0(net825),
    .S1(net819),
    .X(_0814_));
 sky130_fd_sc_hd__mux4_2 _4401_ (.A0(_0811_),
    .A1(_0812_),
    .A2(_0813_),
    .A3(_0814_),
    .S0(net15),
    .S1(net817),
    .X(_0815_));
 sky130_fd_sc_hd__mux4_2 _4402_ (.A0(\dp.rf.rf[0][21] ),
    .A1(\dp.rf.rf[1][21] ),
    .A2(\dp.rf.rf[2][21] ),
    .A3(\dp.rf.rf[3][21] ),
    .S0(net13),
    .S1(net14),
    .X(_0816_));
 sky130_fd_sc_hd__mux4_2 _4403_ (.A0(\dp.rf.rf[4][21] ),
    .A1(\dp.rf.rf[5][21] ),
    .A2(\dp.rf.rf[6][21] ),
    .A3(\dp.rf.rf[7][21] ),
    .S0(net13),
    .S1(net14),
    .X(_0817_));
 sky130_fd_sc_hd__mux4_2 _4404_ (.A0(\dp.rf.rf[8][21] ),
    .A1(\dp.rf.rf[9][21] ),
    .A2(\dp.rf.rf[10][21] ),
    .A3(\dp.rf.rf[11][21] ),
    .S0(net13),
    .S1(net14),
    .X(_0818_));
 sky130_fd_sc_hd__mux4_2 _4405_ (.A0(\dp.rf.rf[12][21] ),
    .A1(\dp.rf.rf[13][21] ),
    .A2(\dp.rf.rf[14][21] ),
    .A3(\dp.rf.rf[15][21] ),
    .S0(net13),
    .S1(net14),
    .X(_0819_));
 sky130_fd_sc_hd__mux4_2 _4406_ (.A0(_0816_),
    .A1(_0817_),
    .A2(_0818_),
    .A3(_0819_),
    .S0(net15),
    .S1(net16),
    .X(_0820_));
 sky130_fd_sc_hd__a22o_4 _4407_ (.A1(net17),
    .A2(_0815_),
    .B1(_0820_),
    .B2(_0337_),
    .X(_0821_));
 sky130_fd_sc_hd__nand2_1 _4408_ (.A(_0121_),
    .B(_0821_),
    .Y(_0822_));
 sky130_fd_sc_hd__a21o_1 _4409_ (.A1(net820),
    .A2(net799),
    .B1(_0349_),
    .X(_3532_[0]));
 sky130_fd_sc_hd__nand2_1 _4410_ (.A(net782),
    .B(_3532_[0]),
    .Y(_0823_));
 sky130_fd_sc_hd__nand2_1 _4411_ (.A(_0822_),
    .B(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__xnor2_1 _4412_ (.A(_0151_),
    .B(_0824_),
    .Y(_3283_[0]));
 sky130_fd_sc_hd__inv_1 _4413_ (.A(_3283_[0]),
    .Y(_3287_[0]));
 sky130_fd_sc_hd__mux2_1 _4414_ (.A0(\dp.rf.rf[22][21] ),
    .A1(\dp.rf.rf[23][21] ),
    .S(net811),
    .X(_0825_));
 sky130_fd_sc_hd__o21ai_0 _4415_ (.A1(net800),
    .A2(_0825_),
    .B1(net786),
    .Y(_0826_));
 sky130_fd_sc_hd__a221oi_1 _4416_ (.A1(\dp.rf.rf[19][21] ),
    .A2(net811),
    .B1(net787),
    .B2(\dp.rf.rf[18][21] ),
    .C1(net792),
    .Y(_0827_));
 sky130_fd_sc_hd__inv_1 _4417_ (.A(\dp.rf.rf[20][21] ),
    .Y(_0828_));
 sky130_fd_sc_hd__mux2i_1 _4418_ (.A0(\dp.rf.rf[17][21] ),
    .A1(\dp.rf.rf[21][21] ),
    .S(net806),
    .Y(_0829_));
 sky130_fd_sc_hd__a221oi_1 _4419_ (.A1(_0828_),
    .A2(net801),
    .B1(_0829_),
    .B2(net811),
    .C1(net808),
    .Y(_0830_));
 sky130_fd_sc_hd__o22ai_1 _4420_ (.A1(\dp.rf.rf[16][21] ),
    .A2(_0412_),
    .B1(_0830_),
    .B2(net789),
    .Y(_0831_));
 sky130_fd_sc_hd__o21ai_2 _4421_ (.A1(_0826_),
    .A2(_0827_),
    .B1(_0831_),
    .Y(_0832_));
 sky130_fd_sc_hd__mux2_1 _4422_ (.A0(\dp.rf.rf[30][21] ),
    .A1(\dp.rf.rf[31][21] ),
    .S(net811),
    .X(_0833_));
 sky130_fd_sc_hd__o21ai_0 _4423_ (.A1(net800),
    .A2(_0833_),
    .B1(_0469_),
    .Y(_0834_));
 sky130_fd_sc_hd__a221oi_1 _4424_ (.A1(\dp.rf.rf[27][21] ),
    .A2(net811),
    .B1(net787),
    .B2(\dp.rf.rf[26][21] ),
    .C1(net792),
    .Y(_0835_));
 sky130_fd_sc_hd__mux4_2 _4425_ (.A0(\dp.rf.rf[24][21] ),
    .A1(\dp.rf.rf[25][21] ),
    .A2(\dp.rf.rf[28][21] ),
    .A3(\dp.rf.rf[29][21] ),
    .S0(net811),
    .S1(net806),
    .X(_0836_));
 sky130_fd_sc_hd__a21oi_1 _4426_ (.A1(_0186_),
    .A2(_0836_),
    .B1(_0192_),
    .Y(_0837_));
 sky130_fd_sc_hd__o22ai_2 _4427_ (.A1(_0834_),
    .A2(_0835_),
    .B1(_0837_),
    .B2(net795),
    .Y(_0838_));
 sky130_fd_sc_hd__mux4_2 _4428_ (.A0(\dp.rf.rf[10][21] ),
    .A1(\dp.rf.rf[11][21] ),
    .A2(\dp.rf.rf[14][21] ),
    .A3(\dp.rf.rf[15][21] ),
    .S0(net813),
    .S1(net804),
    .X(_0839_));
 sky130_fd_sc_hd__mux4_2 _4429_ (.A0(\dp.rf.rf[8][21] ),
    .A1(\dp.rf.rf[9][21] ),
    .A2(\dp.rf.rf[12][21] ),
    .A3(\dp.rf.rf[13][21] ),
    .S0(net813),
    .S1(net804),
    .X(_0840_));
 sky130_fd_sc_hd__mux2i_1 _4430_ (.A0(_0839_),
    .A1(_0840_),
    .S(_0186_),
    .Y(_0841_));
 sky130_fd_sc_hd__mux4_2 _4431_ (.A0(\dp.rf.rf[2][21] ),
    .A1(\dp.rf.rf[3][21] ),
    .A2(\dp.rf.rf[6][21] ),
    .A3(\dp.rf.rf[7][21] ),
    .S0(net813),
    .S1(net804),
    .X(_0842_));
 sky130_fd_sc_hd__inv_1 _4432_ (.A(\dp.rf.rf[4][21] ),
    .Y(_0843_));
 sky130_fd_sc_hd__mux2i_1 _4433_ (.A0(\dp.rf.rf[1][21] ),
    .A1(\dp.rf.rf[5][21] ),
    .S(net804),
    .Y(_0844_));
 sky130_fd_sc_hd__a221oi_1 _4434_ (.A1(_0843_),
    .A2(net801),
    .B1(_0844_),
    .B2(net813),
    .C1(net808),
    .Y(_0845_));
 sky130_fd_sc_hd__a211oi_2 _4435_ (.A1(net808),
    .A2(_0842_),
    .B1(_0845_),
    .C1(net789),
    .Y(_0846_));
 sky130_fd_sc_hd__a211oi_4 _4436_ (.A1(net796),
    .A2(_0841_),
    .B1(_0846_),
    .C1(_0293_),
    .Y(_0847_));
 sky130_fd_sc_hd__a21oi_4 _4437_ (.A1(_0832_),
    .A2(_0838_),
    .B1(_0847_),
    .Y(_3286_[0]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_120 ();
 sky130_fd_sc_hd__a21o_1 _4439_ (.A1(net826),
    .A2(net799),
    .B1(_0349_),
    .X(_3528_[0]));
 sky130_fd_sc_hd__mux4_2 _4440_ (.A0(\dp.rf.rf[28][20] ),
    .A1(\dp.rf.rf[29][20] ),
    .A2(\dp.rf.rf[30][20] ),
    .A3(\dp.rf.rf[31][20] ),
    .S0(net826),
    .S1(net820),
    .X(_0849_));
 sky130_fd_sc_hd__mux4_2 _4441_ (.A0(\dp.rf.rf[20][20] ),
    .A1(\dp.rf.rf[21][20] ),
    .A2(\dp.rf.rf[22][20] ),
    .A3(\dp.rf.rf[23][20] ),
    .S0(net826),
    .S1(net820),
    .X(_0850_));
 sky130_fd_sc_hd__a22oi_1 _4442_ (.A1(_0676_),
    .A2(_0849_),
    .B1(_0850_),
    .B2(_0680_),
    .Y(_0851_));
 sky130_fd_sc_hd__mux4_2 _4443_ (.A0(\dp.rf.rf[16][20] ),
    .A1(\dp.rf.rf[17][20] ),
    .A2(\dp.rf.rf[18][20] ),
    .A3(\dp.rf.rf[19][20] ),
    .S0(net826),
    .S1(net820),
    .X(_0852_));
 sky130_fd_sc_hd__mux4_2 _4444_ (.A0(\dp.rf.rf[24][20] ),
    .A1(\dp.rf.rf[25][20] ),
    .A2(\dp.rf.rf[26][20] ),
    .A3(\dp.rf.rf[27][20] ),
    .S0(net826),
    .S1(net820),
    .X(_0853_));
 sky130_fd_sc_hd__a22oi_1 _4445_ (.A1(_0674_),
    .A2(_0852_),
    .B1(_0853_),
    .B2(_0669_),
    .Y(_0854_));
 sky130_fd_sc_hd__nand2_1 _4446_ (.A(_0851_),
    .B(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__nand2_1 _4447_ (.A(net826),
    .B(\dp.rf.rf[1][20] ),
    .Y(_0856_));
 sky130_fd_sc_hd__mux2i_1 _4448_ (.A0(\dp.rf.rf[2][20] ),
    .A1(\dp.rf.rf[3][20] ),
    .S(net826),
    .Y(_0857_));
 sky130_fd_sc_hd__mux2i_1 _4449_ (.A0(\dp.rf.rf[4][20] ),
    .A1(\dp.rf.rf[5][20] ),
    .S(net826),
    .Y(_0858_));
 sky130_fd_sc_hd__mux2i_1 _4450_ (.A0(\dp.rf.rf[6][20] ),
    .A1(\dp.rf.rf[7][20] ),
    .S(net826),
    .Y(_0859_));
 sky130_fd_sc_hd__mux4_2 _4451_ (.A0(_0856_),
    .A1(_0857_),
    .A2(_0858_),
    .A3(_0859_),
    .S0(net820),
    .S1(net818),
    .X(_0860_));
 sky130_fd_sc_hd__nor2b_4 _4452_ (.A(net17),
    .B_N(net817),
    .Y(_0861_));
 sky130_fd_sc_hd__mux4_2 _4453_ (.A0(\dp.rf.rf[8][20] ),
    .A1(\dp.rf.rf[9][20] ),
    .A2(\dp.rf.rf[10][20] ),
    .A3(\dp.rf.rf[11][20] ),
    .S0(net826),
    .S1(net820),
    .X(_0862_));
 sky130_fd_sc_hd__mux4_2 _4454_ (.A0(\dp.rf.rf[12][20] ),
    .A1(\dp.rf.rf[13][20] ),
    .A2(\dp.rf.rf[14][20] ),
    .A3(\dp.rf.rf[15][20] ),
    .S0(net826),
    .S1(net820),
    .X(_0863_));
 sky130_fd_sc_hd__mux2i_1 _4455_ (.A0(_0862_),
    .A1(_0863_),
    .S(net818),
    .Y(_0864_));
 sky130_fd_sc_hd__a22oi_2 _4456_ (.A1(_0109_),
    .A2(_0860_),
    .B1(_0861_),
    .B2(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__o21ai_2 _4457_ (.A1(_0092_),
    .A2(_0855_),
    .B1(_0865_),
    .Y(_0866_));
 sky130_fd_sc_hd__nor2_1 _4458_ (.A(net782),
    .B(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hd__a21oi_1 _4459_ (.A1(net782),
    .A2(_3528_[0]),
    .B1(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__xor2_1 _4460_ (.A(_0151_),
    .B(_0868_),
    .X(_3291_[0]));
 sky130_fd_sc_hd__inv_1 _4461_ (.A(_3291_[0]),
    .Y(_3295_[0]));
 sky130_fd_sc_hd__nand4_1 _4462_ (.A(net1),
    .B(net12),
    .C(net23),
    .D(\dp.rf.rf[26][20] ),
    .Y(_0869_));
 sky130_fd_sc_hd__o2bb2ai_1 _4463_ (.A1_N(\dp.rf.rf[26][20] ),
    .A2_N(_0400_),
    .B1(_0135_),
    .B2(_0869_),
    .Y(_0870_));
 sky130_fd_sc_hd__and2_0 _4464_ (.A(\dp.rf.rf[27][20] ),
    .B(net810),
    .X(_0871_));
 sky130_fd_sc_hd__mux2i_1 _4465_ (.A0(\dp.rf.rf[30][20] ),
    .A1(\dp.rf.rf[31][20] ),
    .S(net810),
    .Y(_0872_));
 sky130_fd_sc_hd__nand2_1 _4466_ (.A(net805),
    .B(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__o311ai_0 _4467_ (.A1(_0259_),
    .A2(_0870_),
    .A3(_0871_),
    .B1(_0469_),
    .C1(_0873_),
    .Y(_0874_));
 sky130_fd_sc_hd__mux2i_1 _4468_ (.A0(\dp.rf.rf[24][20] ),
    .A1(\dp.rf.rf[28][20] ),
    .S(net805),
    .Y(_0875_));
 sky130_fd_sc_hd__mux2i_1 _4469_ (.A0(\dp.rf.rf[25][20] ),
    .A1(\dp.rf.rf[29][20] ),
    .S(net805),
    .Y(_0876_));
 sky130_fd_sc_hd__o22ai_1 _4470_ (.A1(_0183_),
    .A2(_0875_),
    .B1(_0876_),
    .B2(_0211_),
    .Y(_0877_));
 sky130_fd_sc_hd__o21ai_0 _4471_ (.A1(_0192_),
    .A2(_0877_),
    .B1(_0620_),
    .Y(_0878_));
 sky130_fd_sc_hd__mux2i_1 _4472_ (.A0(\dp.rf.rf[22][20] ),
    .A1(\dp.rf.rf[23][20] ),
    .S(net810),
    .Y(_0879_));
 sky130_fd_sc_hd__mux2i_1 _4473_ (.A0(\dp.rf.rf[18][20] ),
    .A1(\dp.rf.rf[19][20] ),
    .S(net810),
    .Y(_0880_));
 sky130_fd_sc_hd__a221o_1 _4474_ (.A1(net805),
    .A2(_0879_),
    .B1(_0880_),
    .B2(_0513_),
    .C1(_0477_),
    .X(_0881_));
 sky130_fd_sc_hd__inv_1 _4475_ (.A(\dp.rf.rf[20][20] ),
    .Y(_0882_));
 sky130_fd_sc_hd__mux2i_1 _4476_ (.A0(\dp.rf.rf[17][20] ),
    .A1(\dp.rf.rf[21][20] ),
    .S(net805),
    .Y(_0883_));
 sky130_fd_sc_hd__a221oi_1 _4477_ (.A1(_0882_),
    .A2(net801),
    .B1(_0883_),
    .B2(net810),
    .C1(net808),
    .Y(_0884_));
 sky130_fd_sc_hd__o22ai_1 _4478_ (.A1(\dp.rf.rf[16][20] ),
    .A2(_0412_),
    .B1(_0884_),
    .B2(net789),
    .Y(_0885_));
 sky130_fd_sc_hd__a22oi_2 _4479_ (.A1(_0874_),
    .A2(_0878_),
    .B1(_0881_),
    .B2(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__mux4_2 _4480_ (.A0(\dp.rf.rf[10][20] ),
    .A1(\dp.rf.rf[11][20] ),
    .A2(\dp.rf.rf[14][20] ),
    .A3(\dp.rf.rf[15][20] ),
    .S0(net811),
    .S1(net806),
    .X(_0887_));
 sky130_fd_sc_hd__mux4_2 _4481_ (.A0(\dp.rf.rf[8][20] ),
    .A1(\dp.rf.rf[9][20] ),
    .A2(\dp.rf.rf[12][20] ),
    .A3(\dp.rf.rf[13][20] ),
    .S0(net811),
    .S1(net806),
    .X(_0888_));
 sky130_fd_sc_hd__mux2i_1 _4482_ (.A0(_0887_),
    .A1(_0888_),
    .S(_0186_),
    .Y(_0889_));
 sky130_fd_sc_hd__mux4_2 _4483_ (.A0(\dp.rf.rf[2][20] ),
    .A1(\dp.rf.rf[3][20] ),
    .A2(\dp.rf.rf[6][20] ),
    .A3(\dp.rf.rf[7][20] ),
    .S0(net811),
    .S1(net806),
    .X(_0890_));
 sky130_fd_sc_hd__inv_1 _4484_ (.A(\dp.rf.rf[4][20] ),
    .Y(_0891_));
 sky130_fd_sc_hd__mux2i_1 _4485_ (.A0(\dp.rf.rf[1][20] ),
    .A1(\dp.rf.rf[5][20] ),
    .S(net806),
    .Y(_0892_));
 sky130_fd_sc_hd__a221oi_1 _4486_ (.A1(_0891_),
    .A2(net801),
    .B1(_0892_),
    .B2(net811),
    .C1(net808),
    .Y(_0893_));
 sky130_fd_sc_hd__a21oi_2 _4487_ (.A1(net808),
    .A2(_0890_),
    .B1(_0893_),
    .Y(_0894_));
 sky130_fd_sc_hd__a221oi_4 _4488_ (.A1(_0193_),
    .A2(_0889_),
    .B1(_0894_),
    .B2(net785),
    .C1(_0293_),
    .Y(_0895_));
 sky130_fd_sc_hd__nor2_4 _4489_ (.A(_0886_),
    .B(_0895_),
    .Y(_3294_[0]));
 sky130_fd_sc_hd__and2_4 _4490_ (.A(_0143_),
    .B(_0118_),
    .X(_0896_));
 sky130_fd_sc_hd__nand2_8 _4491_ (.A(net26),
    .B(_0896_),
    .Y(_0897_));
 sky130_fd_sc_hd__and3_4 _4492_ (.A(net25),
    .B(_0347_),
    .C(_0897_),
    .X(_0898_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_119 ();
 sky130_fd_sc_hd__a221oi_2 _4494_ (.A1(net10),
    .A2(net799),
    .B1(_0146_),
    .B2(net11),
    .C1(_0898_),
    .Y(_0900_));
 sky130_fd_sc_hd__nand2_8 _4495_ (.A(net29),
    .B(_0042_),
    .Y(_0901_));
 sky130_fd_sc_hd__nand2_8 _4496_ (.A(_0901_),
    .B(_0897_),
    .Y(_0902_));
 sky130_fd_sc_hd__a211oi_1 _4497_ (.A1(net11),
    .A2(net799),
    .B1(_0349_),
    .C1(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__a21oi_2 _4498_ (.A1(_0900_),
    .A2(_0902_),
    .B1(_0903_),
    .Y(_3524_[0]));
 sky130_fd_sc_hd__mux4_2 _4499_ (.A0(\dp.rf.rf[16][19] ),
    .A1(\dp.rf.rf[17][19] ),
    .A2(\dp.rf.rf[18][19] ),
    .A3(\dp.rf.rf[19][19] ),
    .S0(net825),
    .S1(net819),
    .X(_0904_));
 sky130_fd_sc_hd__mux4_2 _4500_ (.A0(\dp.rf.rf[20][19] ),
    .A1(\dp.rf.rf[21][19] ),
    .A2(\dp.rf.rf[22][19] ),
    .A3(\dp.rf.rf[23][19] ),
    .S0(net825),
    .S1(net819),
    .X(_0905_));
 sky130_fd_sc_hd__mux4_2 _4501_ (.A0(\dp.rf.rf[24][19] ),
    .A1(\dp.rf.rf[25][19] ),
    .A2(\dp.rf.rf[26][19] ),
    .A3(\dp.rf.rf[27][19] ),
    .S0(net13),
    .S1(net14),
    .X(_0906_));
 sky130_fd_sc_hd__mux4_2 _4502_ (.A0(\dp.rf.rf[28][19] ),
    .A1(\dp.rf.rf[29][19] ),
    .A2(\dp.rf.rf[30][19] ),
    .A3(\dp.rf.rf[31][19] ),
    .S0(net13),
    .S1(net14),
    .X(_0907_));
 sky130_fd_sc_hd__mux4_2 _4503_ (.A0(_0904_),
    .A1(_0905_),
    .A2(_0906_),
    .A3(_0907_),
    .S0(net818),
    .S1(net16),
    .X(_0908_));
 sky130_fd_sc_hd__nand2_2 _4504_ (.A(net17),
    .B(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__mux4_2 _4505_ (.A0(\dp.rf.rf[0][19] ),
    .A1(\dp.rf.rf[1][19] ),
    .A2(\dp.rf.rf[2][19] ),
    .A3(\dp.rf.rf[3][19] ),
    .S0(net13),
    .S1(net14),
    .X(_0910_));
 sky130_fd_sc_hd__mux4_2 _4506_ (.A0(\dp.rf.rf[4][19] ),
    .A1(\dp.rf.rf[5][19] ),
    .A2(\dp.rf.rf[6][19] ),
    .A3(\dp.rf.rf[7][19] ),
    .S0(net13),
    .S1(net14),
    .X(_0911_));
 sky130_fd_sc_hd__mux4_2 _4507_ (.A0(\dp.rf.rf[8][19] ),
    .A1(\dp.rf.rf[9][19] ),
    .A2(\dp.rf.rf[10][19] ),
    .A3(\dp.rf.rf[11][19] ),
    .S0(net13),
    .S1(net14),
    .X(_0912_));
 sky130_fd_sc_hd__mux4_2 _4508_ (.A0(\dp.rf.rf[12][19] ),
    .A1(\dp.rf.rf[13][19] ),
    .A2(\dp.rf.rf[14][19] ),
    .A3(\dp.rf.rf[15][19] ),
    .S0(net13),
    .S1(net14),
    .X(_0913_));
 sky130_fd_sc_hd__mux4_2 _4509_ (.A0(_0910_),
    .A1(_0911_),
    .A2(_0912_),
    .A3(_0913_),
    .S0(net15),
    .S1(net16),
    .X(_0914_));
 sky130_fd_sc_hd__nand2_2 _4510_ (.A(_0092_),
    .B(_0914_),
    .Y(_0915_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_118 ();
 sky130_fd_sc_hd__a21oi_4 _4512_ (.A1(_0909_),
    .A2(_0915_),
    .B1(_0111_),
    .Y(_0917_));
 sky130_fd_sc_hd__mux2i_1 _4513_ (.A0(_3524_[0]),
    .A1(_0917_),
    .S(_0121_),
    .Y(_0918_));
 sky130_fd_sc_hd__xor2_1 _4514_ (.A(_0151_),
    .B(_0918_),
    .X(_3299_[0]));
 sky130_fd_sc_hd__inv_1 _4515_ (.A(_3299_[0]),
    .Y(_3303_[0]));
 sky130_fd_sc_hd__mux4_2 _4516_ (.A0(\dp.rf.rf[26][19] ),
    .A1(\dp.rf.rf[27][19] ),
    .A2(\dp.rf.rf[30][19] ),
    .A3(\dp.rf.rf[31][19] ),
    .S0(net812),
    .S1(net804),
    .X(_0919_));
 sky130_fd_sc_hd__mux4_2 _4517_ (.A0(\dp.rf.rf[24][19] ),
    .A1(\dp.rf.rf[25][19] ),
    .A2(\dp.rf.rf[28][19] ),
    .A3(\dp.rf.rf[29][19] ),
    .S0(net812),
    .S1(net804),
    .X(_0920_));
 sky130_fd_sc_hd__a221o_1 _4518_ (.A1(net786),
    .A2(_0919_),
    .B1(_0920_),
    .B2(_0186_),
    .C1(_0255_),
    .X(_0921_));
 sky130_fd_sc_hd__mux2_1 _4519_ (.A0(\dp.rf.rf[22][19] ),
    .A1(\dp.rf.rf[23][19] ),
    .S(net812),
    .X(_0922_));
 sky130_fd_sc_hd__o21ai_0 _4520_ (.A1(net800),
    .A2(_0922_),
    .B1(net786),
    .Y(_0923_));
 sky130_fd_sc_hd__a221oi_1 _4521_ (.A1(\dp.rf.rf[19][19] ),
    .A2(net812),
    .B1(_0298_),
    .B2(\dp.rf.rf[18][19] ),
    .C1(_0259_),
    .Y(_0924_));
 sky130_fd_sc_hd__inv_1 _4522_ (.A(\dp.rf.rf[20][19] ),
    .Y(_0925_));
 sky130_fd_sc_hd__mux2i_1 _4523_ (.A0(\dp.rf.rf[17][19] ),
    .A1(\dp.rf.rf[21][19] ),
    .S(net804),
    .Y(_0926_));
 sky130_fd_sc_hd__a221oi_1 _4524_ (.A1(_0925_),
    .A2(net801),
    .B1(_0926_),
    .B2(net812),
    .C1(net8),
    .Y(_0927_));
 sky130_fd_sc_hd__o22ai_1 _4525_ (.A1(\dp.rf.rf[16][19] ),
    .A2(_0412_),
    .B1(_0927_),
    .B2(_0265_),
    .Y(_0928_));
 sky130_fd_sc_hd__o21ai_2 _4526_ (.A1(_0923_),
    .A2(_0924_),
    .B1(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__mux4_2 _4527_ (.A0(\dp.rf.rf[2][19] ),
    .A1(\dp.rf.rf[3][19] ),
    .A2(\dp.rf.rf[6][19] ),
    .A3(\dp.rf.rf[7][19] ),
    .S0(net809),
    .S1(net804),
    .X(_0930_));
 sky130_fd_sc_hd__nand2_1 _4528_ (.A(net8),
    .B(_0930_),
    .Y(_0931_));
 sky130_fd_sc_hd__mux2_1 _4529_ (.A0(\dp.rf.rf[1][19] ),
    .A1(\dp.rf.rf[5][19] ),
    .S(net804),
    .X(_0932_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_117 ();
 sky130_fd_sc_hd__o221ai_1 _4531_ (.A1(\dp.rf.rf[4][19] ),
    .A2(_0395_),
    .B1(_0932_),
    .B2(_0400_),
    .C1(_0186_),
    .Y(_0934_));
 sky130_fd_sc_hd__a31oi_2 _4532_ (.A1(_0389_),
    .A2(_0931_),
    .A3(_0934_),
    .B1(_0293_),
    .Y(_0935_));
 sky130_fd_sc_hd__a221oi_1 _4533_ (.A1(\dp.rf.rf[11][19] ),
    .A2(net809),
    .B1(_0298_),
    .B2(\dp.rf.rf[10][19] ),
    .C1(_0259_),
    .Y(_0936_));
 sky130_fd_sc_hd__mux2_1 _4534_ (.A0(\dp.rf.rf[14][19] ),
    .A1(\dp.rf.rf[15][19] ),
    .S(net809),
    .X(_0937_));
 sky130_fd_sc_hd__o21ai_0 _4535_ (.A1(net800),
    .A2(_0937_),
    .B1(net786),
    .Y(_0938_));
 sky130_fd_sc_hd__mux4_2 _4536_ (.A0(\dp.rf.rf[8][19] ),
    .A1(\dp.rf.rf[9][19] ),
    .A2(\dp.rf.rf[12][19] ),
    .A3(\dp.rf.rf[13][19] ),
    .S0(net809),
    .S1(net9),
    .X(_0939_));
 sky130_fd_sc_hd__a21oi_1 _4537_ (.A1(_0186_),
    .A2(_0939_),
    .B1(_0255_),
    .Y(_0940_));
 sky130_fd_sc_hd__o21ai_2 _4538_ (.A1(_0936_),
    .A2(_0938_),
    .B1(_0940_),
    .Y(_0941_));
 sky130_fd_sc_hd__a32oi_4 _4539_ (.A1(net783),
    .A2(_0921_),
    .A3(_0929_),
    .B1(_0935_),
    .B2(_0941_),
    .Y(_3302_[0]));
 sky130_fd_sc_hd__mux4_2 _4540_ (.A0(\dp.rf.rf[16][18] ),
    .A1(\dp.rf.rf[17][18] ),
    .A2(\dp.rf.rf[18][18] ),
    .A3(\dp.rf.rf[19][18] ),
    .S0(net825),
    .S1(net819),
    .X(_0942_));
 sky130_fd_sc_hd__mux4_2 _4541_ (.A0(\dp.rf.rf[20][18] ),
    .A1(\dp.rf.rf[21][18] ),
    .A2(\dp.rf.rf[22][18] ),
    .A3(\dp.rf.rf[23][18] ),
    .S0(net825),
    .S1(net819),
    .X(_0943_));
 sky130_fd_sc_hd__mux4_2 _4542_ (.A0(\dp.rf.rf[24][18] ),
    .A1(\dp.rf.rf[25][18] ),
    .A2(\dp.rf.rf[26][18] ),
    .A3(\dp.rf.rf[27][18] ),
    .S0(net825),
    .S1(net819),
    .X(_0944_));
 sky130_fd_sc_hd__mux4_2 _4543_ (.A0(\dp.rf.rf[28][18] ),
    .A1(\dp.rf.rf[29][18] ),
    .A2(\dp.rf.rf[30][18] ),
    .A3(\dp.rf.rf[31][18] ),
    .S0(net825),
    .S1(net819),
    .X(_0945_));
 sky130_fd_sc_hd__mux4_2 _4544_ (.A0(_0942_),
    .A1(_0943_),
    .A2(_0944_),
    .A3(_0945_),
    .S0(net15),
    .S1(net817),
    .X(_0946_));
 sky130_fd_sc_hd__mux4_2 _4545_ (.A0(\dp.rf.rf[0][18] ),
    .A1(\dp.rf.rf[1][18] ),
    .A2(\dp.rf.rf[2][18] ),
    .A3(\dp.rf.rf[3][18] ),
    .S0(net13),
    .S1(net14),
    .X(_0947_));
 sky130_fd_sc_hd__mux4_2 _4546_ (.A0(\dp.rf.rf[4][18] ),
    .A1(\dp.rf.rf[5][18] ),
    .A2(\dp.rf.rf[6][18] ),
    .A3(\dp.rf.rf[7][18] ),
    .S0(net13),
    .S1(net14),
    .X(_0948_));
 sky130_fd_sc_hd__mux4_2 _4547_ (.A0(\dp.rf.rf[8][18] ),
    .A1(\dp.rf.rf[9][18] ),
    .A2(\dp.rf.rf[10][18] ),
    .A3(\dp.rf.rf[11][18] ),
    .S0(net13),
    .S1(net14),
    .X(_0949_));
 sky130_fd_sc_hd__mux4_2 _4548_ (.A0(\dp.rf.rf[12][18] ),
    .A1(\dp.rf.rf[13][18] ),
    .A2(\dp.rf.rf[14][18] ),
    .A3(\dp.rf.rf[15][18] ),
    .S0(net13),
    .S1(net14),
    .X(_0950_));
 sky130_fd_sc_hd__mux4_2 _4549_ (.A0(_0947_),
    .A1(_0948_),
    .A2(_0949_),
    .A3(_0950_),
    .S0(net15),
    .S1(net16),
    .X(_0951_));
 sky130_fd_sc_hd__a22oi_2 _4550_ (.A1(net17),
    .A2(_0946_),
    .B1(_0951_),
    .B2(_0337_),
    .Y(_0952_));
 sky130_fd_sc_hd__a221oi_1 _4551_ (.A1(net805),
    .A2(net799),
    .B1(_0146_),
    .B2(net10),
    .C1(_0898_),
    .Y(_0953_));
 sky130_fd_sc_hd__mux2i_2 _4552_ (.A0(_0900_),
    .A1(_0953_),
    .S(_0902_),
    .Y(_3520_[0]));
 sky130_fd_sc_hd__nor2_1 _4553_ (.A(_0121_),
    .B(_3520_[0]),
    .Y(_0954_));
 sky130_fd_sc_hd__a21oi_1 _4554_ (.A1(_0121_),
    .A2(_0952_),
    .B1(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__xnor2_2 _4555_ (.A(_0151_),
    .B(_0955_),
    .Y(_3307_[0]));
 sky130_fd_sc_hd__inv_1 _4556_ (.A(_3307_[0]),
    .Y(_3311_[0]));
 sky130_fd_sc_hd__mux2i_1 _4557_ (.A0(\dp.rf.rf[22][18] ),
    .A1(\dp.rf.rf[23][18] ),
    .S(net812),
    .Y(_0956_));
 sky130_fd_sc_hd__mux2i_1 _4558_ (.A0(\dp.rf.rf[18][18] ),
    .A1(\dp.rf.rf[19][18] ),
    .S(net812),
    .Y(_0957_));
 sky130_fd_sc_hd__a221o_1 _4559_ (.A1(net807),
    .A2(_0956_),
    .B1(_0957_),
    .B2(_0513_),
    .C1(_0477_),
    .X(_0958_));
 sky130_fd_sc_hd__inv_1 _4560_ (.A(\dp.rf.rf[20][18] ),
    .Y(_0959_));
 sky130_fd_sc_hd__mux2i_1 _4561_ (.A0(\dp.rf.rf[17][18] ),
    .A1(\dp.rf.rf[21][18] ),
    .S(net807),
    .Y(_0960_));
 sky130_fd_sc_hd__a221oi_1 _4562_ (.A1(_0959_),
    .A2(net801),
    .B1(_0960_),
    .B2(net812),
    .C1(net808),
    .Y(_0961_));
 sky130_fd_sc_hd__o22ai_1 _4563_ (.A1(\dp.rf.rf[16][18] ),
    .A2(_0412_),
    .B1(_0961_),
    .B2(net789),
    .Y(_0962_));
 sky130_fd_sc_hd__a21oi_2 _4564_ (.A1(_0958_),
    .A2(_0962_),
    .B1(net795),
    .Y(_0963_));
 sky130_fd_sc_hd__nor2b_1 _4565_ (.A(net813),
    .B_N(\dp.rf.rf[30][18] ),
    .Y(_0964_));
 sky130_fd_sc_hd__a211oi_1 _4566_ (.A1(\dp.rf.rf[31][18] ),
    .A2(net813),
    .B1(net800),
    .C1(_0964_),
    .Y(_0965_));
 sky130_fd_sc_hd__a221oi_1 _4567_ (.A1(\dp.rf.rf[27][18] ),
    .A2(net813),
    .B1(net787),
    .B2(\dp.rf.rf[26][18] ),
    .C1(net792),
    .Y(_0966_));
 sky130_fd_sc_hd__inv_1 _4568_ (.A(\dp.rf.rf[28][18] ),
    .Y(_0967_));
 sky130_fd_sc_hd__mux2i_1 _4569_ (.A0(\dp.rf.rf[25][18] ),
    .A1(\dp.rf.rf[29][18] ),
    .S(net807),
    .Y(_0968_));
 sky130_fd_sc_hd__a221oi_1 _4570_ (.A1(_0967_),
    .A2(net801),
    .B1(_0968_),
    .B2(net813),
    .C1(net808),
    .Y(_0969_));
 sky130_fd_sc_hd__o21ai_0 _4571_ (.A1(\dp.rf.rf[24][18] ),
    .A2(net798),
    .B1(_0969_),
    .Y(_0970_));
 sky130_fd_sc_hd__o311ai_2 _4572_ (.A1(_0477_),
    .A2(_0965_),
    .A3(_0966_),
    .B1(_0970_),
    .C1(net796),
    .Y(_0971_));
 sky130_fd_sc_hd__mux4_2 _4573_ (.A0(\dp.rf.rf[10][18] ),
    .A1(\dp.rf.rf[11][18] ),
    .A2(\dp.rf.rf[14][18] ),
    .A3(\dp.rf.rf[15][18] ),
    .S0(net813),
    .S1(net806),
    .X(_0972_));
 sky130_fd_sc_hd__mux4_2 _4574_ (.A0(\dp.rf.rf[8][18] ),
    .A1(\dp.rf.rf[9][18] ),
    .A2(\dp.rf.rf[12][18] ),
    .A3(\dp.rf.rf[13][18] ),
    .S0(net813),
    .S1(net806),
    .X(_0973_));
 sky130_fd_sc_hd__mux2i_1 _4575_ (.A0(_0972_),
    .A1(_0973_),
    .S(_0186_),
    .Y(_0974_));
 sky130_fd_sc_hd__mux4_2 _4576_ (.A0(\dp.rf.rf[2][18] ),
    .A1(\dp.rf.rf[3][18] ),
    .A2(\dp.rf.rf[6][18] ),
    .A3(\dp.rf.rf[7][18] ),
    .S0(net813),
    .S1(net806),
    .X(_0975_));
 sky130_fd_sc_hd__inv_1 _4577_ (.A(\dp.rf.rf[4][18] ),
    .Y(_0976_));
 sky130_fd_sc_hd__mux2i_1 _4578_ (.A0(\dp.rf.rf[1][18] ),
    .A1(\dp.rf.rf[5][18] ),
    .S(net806),
    .Y(_0977_));
 sky130_fd_sc_hd__a221oi_1 _4579_ (.A1(_0976_),
    .A2(net801),
    .B1(_0977_),
    .B2(net813),
    .C1(net808),
    .Y(_0978_));
 sky130_fd_sc_hd__a211oi_1 _4580_ (.A1(net808),
    .A2(_0975_),
    .B1(_0978_),
    .C1(net789),
    .Y(_0979_));
 sky130_fd_sc_hd__a211oi_2 _4581_ (.A1(net796),
    .A2(_0974_),
    .B1(_0979_),
    .C1(_0293_),
    .Y(_0980_));
 sky130_fd_sc_hd__a21oi_4 _4582_ (.A1(_0963_),
    .A2(_0971_),
    .B1(_0980_),
    .Y(_3310_[0]));
 sky130_fd_sc_hd__mux4_2 _4583_ (.A0(\dp.rf.rf[16][17] ),
    .A1(\dp.rf.rf[17][17] ),
    .A2(\dp.rf.rf[18][17] ),
    .A3(\dp.rf.rf[19][17] ),
    .S0(net825),
    .S1(net819),
    .X(_0981_));
 sky130_fd_sc_hd__mux4_2 _4584_ (.A0(\dp.rf.rf[20][17] ),
    .A1(\dp.rf.rf[21][17] ),
    .A2(\dp.rf.rf[22][17] ),
    .A3(\dp.rf.rf[23][17] ),
    .S0(net825),
    .S1(net819),
    .X(_0982_));
 sky130_fd_sc_hd__mux4_2 _4585_ (.A0(\dp.rf.rf[24][17] ),
    .A1(\dp.rf.rf[25][17] ),
    .A2(\dp.rf.rf[26][17] ),
    .A3(\dp.rf.rf[27][17] ),
    .S0(net825),
    .S1(net819),
    .X(_0983_));
 sky130_fd_sc_hd__mux4_2 _4586_ (.A0(\dp.rf.rf[28][17] ),
    .A1(\dp.rf.rf[29][17] ),
    .A2(\dp.rf.rf[30][17] ),
    .A3(\dp.rf.rf[31][17] ),
    .S0(net825),
    .S1(net819),
    .X(_0984_));
 sky130_fd_sc_hd__mux4_2 _4587_ (.A0(_0981_),
    .A1(_0982_),
    .A2(_0983_),
    .A3(_0984_),
    .S0(net15),
    .S1(net16),
    .X(_0985_));
 sky130_fd_sc_hd__nand2_2 _4588_ (.A(net17),
    .B(_0985_),
    .Y(_0986_));
 sky130_fd_sc_hd__mux4_2 _4589_ (.A0(\dp.rf.rf[0][17] ),
    .A1(\dp.rf.rf[1][17] ),
    .A2(\dp.rf.rf[2][17] ),
    .A3(\dp.rf.rf[3][17] ),
    .S0(net13),
    .S1(net14),
    .X(_0987_));
 sky130_fd_sc_hd__mux4_2 _4590_ (.A0(\dp.rf.rf[4][17] ),
    .A1(\dp.rf.rf[5][17] ),
    .A2(\dp.rf.rf[6][17] ),
    .A3(\dp.rf.rf[7][17] ),
    .S0(net13),
    .S1(net14),
    .X(_0988_));
 sky130_fd_sc_hd__mux4_2 _4591_ (.A0(\dp.rf.rf[8][17] ),
    .A1(\dp.rf.rf[9][17] ),
    .A2(\dp.rf.rf[10][17] ),
    .A3(\dp.rf.rf[11][17] ),
    .S0(net13),
    .S1(net14),
    .X(_0989_));
 sky130_fd_sc_hd__mux4_2 _4592_ (.A0(\dp.rf.rf[12][17] ),
    .A1(\dp.rf.rf[13][17] ),
    .A2(\dp.rf.rf[14][17] ),
    .A3(\dp.rf.rf[15][17] ),
    .S0(net13),
    .S1(net14),
    .X(_0990_));
 sky130_fd_sc_hd__mux4_2 _4593_ (.A0(_0987_),
    .A1(_0988_),
    .A2(_0989_),
    .A3(_0990_),
    .S0(net15),
    .S1(net16),
    .X(_0991_));
 sky130_fd_sc_hd__nand2_2 _4594_ (.A(_0092_),
    .B(_0991_),
    .Y(_0992_));
 sky130_fd_sc_hd__nand2_2 _4595_ (.A(_0986_),
    .B(_0992_),
    .Y(_0993_));
 sky130_fd_sc_hd__nand2_4 _4596_ (.A(_0351_),
    .B(_0993_),
    .Y(_0994_));
 sky130_fd_sc_hd__a221oi_1 _4597_ (.A1(net8),
    .A2(net799),
    .B1(_0146_),
    .B2(net805),
    .C1(_0898_),
    .Y(_0995_));
 sky130_fd_sc_hd__mux2i_1 _4598_ (.A0(_0953_),
    .A1(_0995_),
    .S(_0902_),
    .Y(_3516_[0]));
 sky130_fd_sc_hd__nand2_1 _4599_ (.A(net782),
    .B(_3516_[0]),
    .Y(_0996_));
 sky130_fd_sc_hd__o21ai_2 _4600_ (.A1(net782),
    .A2(_0994_),
    .B1(_0996_),
    .Y(_0997_));
 sky130_fd_sc_hd__xnor2_1 _4601_ (.A(_0151_),
    .B(_0997_),
    .Y(_3315_[0]));
 sky130_fd_sc_hd__inv_1 _4602_ (.A(_3315_[0]),
    .Y(_3319_[0]));
 sky130_fd_sc_hd__mux2_1 _4603_ (.A0(\dp.rf.rf[1][17] ),
    .A1(\dp.rf.rf[5][17] ),
    .S(net804),
    .X(_0998_));
 sky130_fd_sc_hd__o22ai_1 _4604_ (.A1(\dp.rf.rf[4][17] ),
    .A2(_0395_),
    .B1(_0998_),
    .B2(_0400_),
    .Y(_0999_));
 sky130_fd_sc_hd__mux4_2 _4605_ (.A0(\dp.rf.rf[2][17] ),
    .A1(\dp.rf.rf[3][17] ),
    .A2(\dp.rf.rf[6][17] ),
    .A3(\dp.rf.rf[7][17] ),
    .S0(net812),
    .S1(net804),
    .X(_1000_));
 sky130_fd_sc_hd__nand2_1 _4606_ (.A(net808),
    .B(_1000_),
    .Y(_1001_));
 sky130_fd_sc_hd__o211ai_1 _4607_ (.A1(net808),
    .A2(_0999_),
    .B1(_1001_),
    .C1(_0389_),
    .Y(_1002_));
 sky130_fd_sc_hd__mux4_2 _4608_ (.A0(\dp.rf.rf[10][17] ),
    .A1(\dp.rf.rf[11][17] ),
    .A2(\dp.rf.rf[14][17] ),
    .A3(\dp.rf.rf[15][17] ),
    .S0(net812),
    .S1(net804),
    .X(_1003_));
 sky130_fd_sc_hd__nand2_1 _4609_ (.A(net808),
    .B(_1003_),
    .Y(_1004_));
 sky130_fd_sc_hd__mux4_2 _4610_ (.A0(\dp.rf.rf[8][17] ),
    .A1(\dp.rf.rf[9][17] ),
    .A2(\dp.rf.rf[12][17] ),
    .A3(\dp.rf.rf[13][17] ),
    .S0(net812),
    .S1(net804),
    .X(_1005_));
 sky130_fd_sc_hd__nand2_1 _4611_ (.A(_0186_),
    .B(_1005_),
    .Y(_1006_));
 sky130_fd_sc_hd__nand3_2 _4612_ (.A(net796),
    .B(_1004_),
    .C(_1006_),
    .Y(_1007_));
 sky130_fd_sc_hd__mux2i_1 _4613_ (.A0(\dp.rf.rf[30][17] ),
    .A1(\dp.rf.rf[31][17] ),
    .S(net812),
    .Y(_1008_));
 sky130_fd_sc_hd__nand2_1 _4614_ (.A(net806),
    .B(_1008_),
    .Y(_1009_));
 sky130_fd_sc_hd__a221o_1 _4615_ (.A1(\dp.rf.rf[27][17] ),
    .A2(net812),
    .B1(_0298_),
    .B2(\dp.rf.rf[26][17] ),
    .C1(_0259_),
    .X(_1010_));
 sky130_fd_sc_hd__mux4_2 _4616_ (.A0(\dp.rf.rf[24][17] ),
    .A1(\dp.rf.rf[25][17] ),
    .A2(\dp.rf.rf[28][17] ),
    .A3(\dp.rf.rf[29][17] ),
    .S0(net812),
    .S1(net806),
    .X(_1011_));
 sky130_fd_sc_hd__nand2_1 _4617_ (.A(_0186_),
    .B(_1011_),
    .Y(_1012_));
 sky130_fd_sc_hd__a21oi_1 _4618_ (.A1(net796),
    .A2(_1012_),
    .B1(_0224_),
    .Y(_1013_));
 sky130_fd_sc_hd__a31o_4 _4619_ (.A1(_0469_),
    .A2(_1009_),
    .A3(_1010_),
    .B1(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__mux2_1 _4620_ (.A0(\dp.rf.rf[22][17] ),
    .A1(\dp.rf.rf[23][17] ),
    .S(net812),
    .X(_1015_));
 sky130_fd_sc_hd__o21ai_0 _4621_ (.A1(net800),
    .A2(_1015_),
    .B1(net786),
    .Y(_1016_));
 sky130_fd_sc_hd__a221oi_1 _4622_ (.A1(\dp.rf.rf[19][17] ),
    .A2(net812),
    .B1(_0298_),
    .B2(\dp.rf.rf[18][17] ),
    .C1(_0259_),
    .Y(_1017_));
 sky130_fd_sc_hd__inv_1 _4623_ (.A(\dp.rf.rf[20][17] ),
    .Y(_1018_));
 sky130_fd_sc_hd__mux2i_1 _4624_ (.A0(\dp.rf.rf[17][17] ),
    .A1(\dp.rf.rf[21][17] ),
    .S(net806),
    .Y(_1019_));
 sky130_fd_sc_hd__a221oi_1 _4625_ (.A1(_1018_),
    .A2(net801),
    .B1(_1019_),
    .B2(net812),
    .C1(net808),
    .Y(_1020_));
 sky130_fd_sc_hd__o22ai_1 _4626_ (.A1(\dp.rf.rf[16][17] ),
    .A2(_0412_),
    .B1(_1020_),
    .B2(_0265_),
    .Y(_1021_));
 sky130_fd_sc_hd__o21ai_2 _4627_ (.A1(_1016_),
    .A2(_1017_),
    .B1(_1021_),
    .Y(_1022_));
 sky130_fd_sc_hd__a32oi_4 _4628_ (.A1(net781),
    .A2(_1002_),
    .A3(_1007_),
    .B1(_1014_),
    .B2(_1022_),
    .Y(_3318_[0]));
 sky130_fd_sc_hd__nand2_1 _4629_ (.A(net826),
    .B(\dp.rf.rf[1][16] ),
    .Y(_1023_));
 sky130_fd_sc_hd__mux2i_1 _4630_ (.A0(\dp.rf.rf[2][16] ),
    .A1(\dp.rf.rf[3][16] ),
    .S(net826),
    .Y(_1024_));
 sky130_fd_sc_hd__mux2i_1 _4631_ (.A0(\dp.rf.rf[4][16] ),
    .A1(\dp.rf.rf[5][16] ),
    .S(net826),
    .Y(_1025_));
 sky130_fd_sc_hd__mux2i_1 _4632_ (.A0(\dp.rf.rf[6][16] ),
    .A1(\dp.rf.rf[7][16] ),
    .S(net826),
    .Y(_1026_));
 sky130_fd_sc_hd__mux4_2 _4633_ (.A0(_1023_),
    .A1(_1024_),
    .A2(_1025_),
    .A3(_1026_),
    .S0(net820),
    .S1(net818),
    .X(_1027_));
 sky130_fd_sc_hd__mux4_2 _4634_ (.A0(\dp.rf.rf[8][16] ),
    .A1(\dp.rf.rf[9][16] ),
    .A2(\dp.rf.rf[10][16] ),
    .A3(\dp.rf.rf[11][16] ),
    .S0(net826),
    .S1(net820),
    .X(_1028_));
 sky130_fd_sc_hd__mux4_2 _4635_ (.A0(\dp.rf.rf[12][16] ),
    .A1(\dp.rf.rf[13][16] ),
    .A2(\dp.rf.rf[14][16] ),
    .A3(\dp.rf.rf[15][16] ),
    .S0(net826),
    .S1(net820),
    .X(_1029_));
 sky130_fd_sc_hd__mux2i_1 _4636_ (.A0(_1028_),
    .A1(_1029_),
    .S(net818),
    .Y(_1030_));
 sky130_fd_sc_hd__a22oi_2 _4637_ (.A1(_0109_),
    .A2(_1027_),
    .B1(_1030_),
    .B2(_0861_),
    .Y(_1031_));
 sky130_fd_sc_hd__mux4_2 _4638_ (.A0(\dp.rf.rf[28][16] ),
    .A1(\dp.rf.rf[29][16] ),
    .A2(\dp.rf.rf[30][16] ),
    .A3(\dp.rf.rf[31][16] ),
    .S0(net826),
    .S1(net820),
    .X(_1032_));
 sky130_fd_sc_hd__mux4_2 _4639_ (.A0(\dp.rf.rf[20][16] ),
    .A1(\dp.rf.rf[21][16] ),
    .A2(\dp.rf.rf[22][16] ),
    .A3(\dp.rf.rf[23][16] ),
    .S0(net826),
    .S1(net820),
    .X(_1033_));
 sky130_fd_sc_hd__a22oi_1 _4640_ (.A1(_0676_),
    .A2(_1032_),
    .B1(_1033_),
    .B2(_0680_),
    .Y(_1034_));
 sky130_fd_sc_hd__mux4_2 _4641_ (.A0(\dp.rf.rf[16][16] ),
    .A1(\dp.rf.rf[17][16] ),
    .A2(\dp.rf.rf[18][16] ),
    .A3(\dp.rf.rf[19][16] ),
    .S0(net826),
    .S1(net820),
    .X(_1035_));
 sky130_fd_sc_hd__mux4_2 _4642_ (.A0(\dp.rf.rf[24][16] ),
    .A1(\dp.rf.rf[25][16] ),
    .A2(\dp.rf.rf[26][16] ),
    .A3(\dp.rf.rf[27][16] ),
    .S0(net826),
    .S1(net820),
    .X(_1036_));
 sky130_fd_sc_hd__a22oi_1 _4643_ (.A1(_0674_),
    .A2(_1035_),
    .B1(_1036_),
    .B2(_0669_),
    .Y(_1037_));
 sky130_fd_sc_hd__nand3_2 _4644_ (.A(net17),
    .B(_1034_),
    .C(_1037_),
    .Y(_1038_));
 sky130_fd_sc_hd__nand2_4 _4645_ (.A(_1031_),
    .B(_1038_),
    .Y(_1039_));
 sky130_fd_sc_hd__a221oi_1 _4646_ (.A1(net810),
    .A2(net799),
    .B1(_0146_),
    .B2(net8),
    .C1(_0898_),
    .Y(_1040_));
 sky130_fd_sc_hd__mux2i_1 _4647_ (.A0(_0995_),
    .A1(_1040_),
    .S(_0902_),
    .Y(_3512_[0]));
 sky130_fd_sc_hd__nand2_1 _4648_ (.A(net782),
    .B(_3512_[0]),
    .Y(_1041_));
 sky130_fd_sc_hd__o21ai_2 _4649_ (.A1(net782),
    .A2(_1039_),
    .B1(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__xnor2_1 _4650_ (.A(_0151_),
    .B(_1042_),
    .Y(_3323_[0]));
 sky130_fd_sc_hd__inv_1 _4651_ (.A(_3323_[0]),
    .Y(_3327_[0]));
 sky130_fd_sc_hd__nand4_1 _4652_ (.A(net1),
    .B(net12),
    .C(net23),
    .D(\dp.rf.rf[26][16] ),
    .Y(_1043_));
 sky130_fd_sc_hd__o2bb2ai_1 _4653_ (.A1_N(\dp.rf.rf[26][16] ),
    .A2_N(_0400_),
    .B1(_0135_),
    .B2(_1043_),
    .Y(_1044_));
 sky130_fd_sc_hd__and2_0 _4654_ (.A(\dp.rf.rf[27][16] ),
    .B(net810),
    .X(_1045_));
 sky130_fd_sc_hd__mux2i_1 _4655_ (.A0(\dp.rf.rf[30][16] ),
    .A1(\dp.rf.rf[31][16] ),
    .S(net810),
    .Y(_1046_));
 sky130_fd_sc_hd__nand2_1 _4656_ (.A(net805),
    .B(_1046_),
    .Y(_1047_));
 sky130_fd_sc_hd__o311ai_1 _4657_ (.A1(_0259_),
    .A2(_1044_),
    .A3(_1045_),
    .B1(_0469_),
    .C1(_1047_),
    .Y(_1048_));
 sky130_fd_sc_hd__mux2i_1 _4658_ (.A0(\dp.rf.rf[24][16] ),
    .A1(\dp.rf.rf[28][16] ),
    .S(net805),
    .Y(_1049_));
 sky130_fd_sc_hd__mux2i_1 _4659_ (.A0(\dp.rf.rf[25][16] ),
    .A1(\dp.rf.rf[29][16] ),
    .S(net805),
    .Y(_1050_));
 sky130_fd_sc_hd__o22ai_1 _4660_ (.A1(_0183_),
    .A2(_1049_),
    .B1(_1050_),
    .B2(_0211_),
    .Y(_1051_));
 sky130_fd_sc_hd__o21ai_0 _4661_ (.A1(net793),
    .A2(_1051_),
    .B1(_0620_),
    .Y(_1052_));
 sky130_fd_sc_hd__nand4_1 _4662_ (.A(net1),
    .B(net12),
    .C(net23),
    .D(\dp.rf.rf[18][16] ),
    .Y(_1053_));
 sky130_fd_sc_hd__o2bb2ai_1 _4663_ (.A1_N(\dp.rf.rf[18][16] ),
    .A2_N(_0400_),
    .B1(_0135_),
    .B2(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__and2_0 _4664_ (.A(\dp.rf.rf[19][16] ),
    .B(net810),
    .X(_1055_));
 sky130_fd_sc_hd__mux2i_1 _4665_ (.A0(\dp.rf.rf[22][16] ),
    .A1(\dp.rf.rf[23][16] ),
    .S(net810),
    .Y(_1056_));
 sky130_fd_sc_hd__nand2_1 _4666_ (.A(net805),
    .B(_1056_),
    .Y(_1057_));
 sky130_fd_sc_hd__o311ai_0 _4667_ (.A1(_0259_),
    .A2(_1054_),
    .A3(_1055_),
    .B1(net786),
    .C1(_1057_),
    .Y(_1058_));
 sky130_fd_sc_hd__inv_1 _4668_ (.A(\dp.rf.rf[20][16] ),
    .Y(_1059_));
 sky130_fd_sc_hd__mux2i_1 _4669_ (.A0(\dp.rf.rf[17][16] ),
    .A1(\dp.rf.rf[21][16] ),
    .S(net805),
    .Y(_1060_));
 sky130_fd_sc_hd__a221oi_1 _4670_ (.A1(_1059_),
    .A2(net801),
    .B1(_1060_),
    .B2(net810),
    .C1(net8),
    .Y(_1061_));
 sky130_fd_sc_hd__o22ai_1 _4671_ (.A1(\dp.rf.rf[16][16] ),
    .A2(_0412_),
    .B1(_1061_),
    .B2(net789),
    .Y(_1062_));
 sky130_fd_sc_hd__a22oi_2 _4672_ (.A1(_1048_),
    .A2(_1052_),
    .B1(_1058_),
    .B2(_1062_),
    .Y(_1063_));
 sky130_fd_sc_hd__mux4_2 _4673_ (.A0(\dp.rf.rf[10][16] ),
    .A1(\dp.rf.rf[11][16] ),
    .A2(\dp.rf.rf[14][16] ),
    .A3(\dp.rf.rf[15][16] ),
    .S0(net811),
    .S1(net806),
    .X(_1064_));
 sky130_fd_sc_hd__mux4_2 _4674_ (.A0(\dp.rf.rf[8][16] ),
    .A1(\dp.rf.rf[9][16] ),
    .A2(\dp.rf.rf[12][16] ),
    .A3(\dp.rf.rf[13][16] ),
    .S0(net811),
    .S1(net806),
    .X(_1065_));
 sky130_fd_sc_hd__mux2i_1 _4675_ (.A0(_1064_),
    .A1(_1065_),
    .S(_0186_),
    .Y(_1066_));
 sky130_fd_sc_hd__mux4_2 _4676_ (.A0(\dp.rf.rf[2][16] ),
    .A1(\dp.rf.rf[3][16] ),
    .A2(\dp.rf.rf[6][16] ),
    .A3(\dp.rf.rf[7][16] ),
    .S0(net811),
    .S1(net805),
    .X(_1067_));
 sky130_fd_sc_hd__inv_1 _4677_ (.A(\dp.rf.rf[4][16] ),
    .Y(_1068_));
 sky130_fd_sc_hd__mux2i_1 _4678_ (.A0(\dp.rf.rf[1][16] ),
    .A1(\dp.rf.rf[5][16] ),
    .S(net805),
    .Y(_1069_));
 sky130_fd_sc_hd__a221oi_1 _4679_ (.A1(_1068_),
    .A2(net801),
    .B1(_1069_),
    .B2(net811),
    .C1(net808),
    .Y(_1070_));
 sky130_fd_sc_hd__a21oi_2 _4680_ (.A1(net808),
    .A2(_1067_),
    .B1(_1070_),
    .Y(_1071_));
 sky130_fd_sc_hd__a221oi_4 _4681_ (.A1(_0193_),
    .A2(_1066_),
    .B1(_1071_),
    .B2(net785),
    .C1(_0293_),
    .Y(_1072_));
 sky130_fd_sc_hd__nor2_4 _4682_ (.A(_1063_),
    .B(_1072_),
    .Y(_3326_[0]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_116 ();
 sky130_fd_sc_hd__a221oi_1 _4684_ (.A1(net6),
    .A2(net799),
    .B1(_0146_),
    .B2(net810),
    .C1(_0898_),
    .Y(_1074_));
 sky130_fd_sc_hd__mux2i_1 _4685_ (.A0(_1040_),
    .A1(_1074_),
    .S(_0902_),
    .Y(_3508_[0]));
 sky130_fd_sc_hd__nand2_1 _4686_ (.A(net782),
    .B(_3508_[0]),
    .Y(_1075_));
 sky130_fd_sc_hd__mux4_2 _4687_ (.A0(\dp.rf.rf[16][15] ),
    .A1(\dp.rf.rf[17][15] ),
    .A2(\dp.rf.rf[18][15] ),
    .A3(\dp.rf.rf[19][15] ),
    .S0(net822),
    .S1(net14),
    .X(_1076_));
 sky130_fd_sc_hd__mux4_2 _4688_ (.A0(\dp.rf.rf[20][15] ),
    .A1(\dp.rf.rf[21][15] ),
    .A2(\dp.rf.rf[22][15] ),
    .A3(\dp.rf.rf[23][15] ),
    .S0(net822),
    .S1(net14),
    .X(_1077_));
 sky130_fd_sc_hd__mux4_2 _4689_ (.A0(\dp.rf.rf[24][15] ),
    .A1(\dp.rf.rf[25][15] ),
    .A2(\dp.rf.rf[26][15] ),
    .A3(\dp.rf.rf[27][15] ),
    .S0(net822),
    .S1(net14),
    .X(_1078_));
 sky130_fd_sc_hd__mux4_2 _4690_ (.A0(\dp.rf.rf[28][15] ),
    .A1(\dp.rf.rf[29][15] ),
    .A2(\dp.rf.rf[30][15] ),
    .A3(\dp.rf.rf[31][15] ),
    .S0(net822),
    .S1(net14),
    .X(_1079_));
 sky130_fd_sc_hd__mux4_2 _4691_ (.A0(_1076_),
    .A1(_1077_),
    .A2(_1078_),
    .A3(_1079_),
    .S0(net818),
    .S1(net16),
    .X(_1080_));
 sky130_fd_sc_hd__nand2_1 _4692_ (.A(net17),
    .B(_1080_),
    .Y(_1081_));
 sky130_fd_sc_hd__mux4_2 _4693_ (.A0(\dp.rf.rf[0][15] ),
    .A1(\dp.rf.rf[1][15] ),
    .A2(\dp.rf.rf[2][15] ),
    .A3(\dp.rf.rf[3][15] ),
    .S0(net822),
    .S1(net14),
    .X(_1082_));
 sky130_fd_sc_hd__mux4_2 _4694_ (.A0(\dp.rf.rf[4][15] ),
    .A1(\dp.rf.rf[5][15] ),
    .A2(\dp.rf.rf[6][15] ),
    .A3(\dp.rf.rf[7][15] ),
    .S0(net822),
    .S1(net14),
    .X(_1083_));
 sky130_fd_sc_hd__mux4_2 _4695_ (.A0(\dp.rf.rf[8][15] ),
    .A1(\dp.rf.rf[9][15] ),
    .A2(\dp.rf.rf[10][15] ),
    .A3(\dp.rf.rf[11][15] ),
    .S0(net822),
    .S1(net14),
    .X(_1084_));
 sky130_fd_sc_hd__mux4_2 _4696_ (.A0(\dp.rf.rf[12][15] ),
    .A1(\dp.rf.rf[13][15] ),
    .A2(\dp.rf.rf[14][15] ),
    .A3(\dp.rf.rf[15][15] ),
    .S0(net822),
    .S1(net14),
    .X(_1085_));
 sky130_fd_sc_hd__mux4_2 _4697_ (.A0(_1082_),
    .A1(_1083_),
    .A2(_1084_),
    .A3(_1085_),
    .S0(net818),
    .S1(net16),
    .X(_1086_));
 sky130_fd_sc_hd__nand2_2 _4698_ (.A(_0092_),
    .B(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__a21oi_4 _4699_ (.A1(_1081_),
    .A2(_1087_),
    .B1(_0111_),
    .Y(_1088_));
 sky130_fd_sc_hd__nand2_1 _4700_ (.A(_0121_),
    .B(_1088_),
    .Y(_1089_));
 sky130_fd_sc_hd__nand2_2 _4701_ (.A(_1075_),
    .B(_1089_),
    .Y(_1090_));
 sky130_fd_sc_hd__xnor2_1 _4702_ (.A(_0151_),
    .B(_1090_),
    .Y(_3331_[0]));
 sky130_fd_sc_hd__inv_1 _4703_ (.A(_3331_[0]),
    .Y(_3335_[0]));
 sky130_fd_sc_hd__mux4_2 _4704_ (.A0(\dp.rf.rf[26][15] ),
    .A1(\dp.rf.rf[27][15] ),
    .A2(\dp.rf.rf[30][15] ),
    .A3(\dp.rf.rf[31][15] ),
    .S0(net7),
    .S1(net9),
    .X(_1091_));
 sky130_fd_sc_hd__nand2_1 _4705_ (.A(net8),
    .B(_1091_),
    .Y(_1092_));
 sky130_fd_sc_hd__mux4_2 _4706_ (.A0(\dp.rf.rf[24][15] ),
    .A1(\dp.rf.rf[25][15] ),
    .A2(\dp.rf.rf[28][15] ),
    .A3(\dp.rf.rf[29][15] ),
    .S0(net7),
    .S1(net9),
    .X(_1093_));
 sky130_fd_sc_hd__nand2_1 _4707_ (.A(_0186_),
    .B(_1093_),
    .Y(_1094_));
 sky130_fd_sc_hd__a31oi_1 _4708_ (.A1(net10),
    .A2(_1092_),
    .A3(_1094_),
    .B1(net794),
    .Y(_1095_));
 sky130_fd_sc_hd__mux2_1 _4709_ (.A0(\dp.rf.rf[22][15] ),
    .A1(\dp.rf.rf[23][15] ),
    .S(net7),
    .X(_1096_));
 sky130_fd_sc_hd__o21ai_0 _4710_ (.A1(_0231_),
    .A2(_1096_),
    .B1(net786),
    .Y(_1097_));
 sky130_fd_sc_hd__a221oi_1 _4711_ (.A1(\dp.rf.rf[19][15] ),
    .A2(net7),
    .B1(net788),
    .B2(\dp.rf.rf[18][15] ),
    .C1(net791),
    .Y(_1098_));
 sky130_fd_sc_hd__inv_1 _4712_ (.A(\dp.rf.rf[20][15] ),
    .Y(_1099_));
 sky130_fd_sc_hd__mux2i_1 _4713_ (.A0(\dp.rf.rf[17][15] ),
    .A1(\dp.rf.rf[21][15] ),
    .S(net9),
    .Y(_1100_));
 sky130_fd_sc_hd__a221oi_1 _4714_ (.A1(_1099_),
    .A2(net801),
    .B1(_1100_),
    .B2(net7),
    .C1(net8),
    .Y(_1101_));
 sky130_fd_sc_hd__o22ai_1 _4715_ (.A1(\dp.rf.rf[16][15] ),
    .A2(net784),
    .B1(_1101_),
    .B2(_0265_),
    .Y(_1102_));
 sky130_fd_sc_hd__o21ai_0 _4716_ (.A1(_1097_),
    .A2(_1098_),
    .B1(_1102_),
    .Y(_1103_));
 sky130_fd_sc_hd__mux4_2 _4717_ (.A0(\dp.rf.rf[8][15] ),
    .A1(\dp.rf.rf[9][15] ),
    .A2(\dp.rf.rf[12][15] ),
    .A3(\dp.rf.rf[13][15] ),
    .S0(net7),
    .S1(net9),
    .X(_1104_));
 sky130_fd_sc_hd__nand2_1 _4718_ (.A(_0186_),
    .B(_1104_),
    .Y(_1105_));
 sky130_fd_sc_hd__mux4_2 _4719_ (.A0(\dp.rf.rf[10][15] ),
    .A1(\dp.rf.rf[11][15] ),
    .A2(\dp.rf.rf[14][15] ),
    .A3(\dp.rf.rf[15][15] ),
    .S0(net7),
    .S1(net9),
    .X(_1106_));
 sky130_fd_sc_hd__nand2_1 _4720_ (.A(net8),
    .B(_1106_),
    .Y(_1107_));
 sky130_fd_sc_hd__mux4_2 _4721_ (.A0(\dp.rf.rf[2][15] ),
    .A1(\dp.rf.rf[3][15] ),
    .A2(\dp.rf.rf[6][15] ),
    .A3(\dp.rf.rf[7][15] ),
    .S0(net7),
    .S1(net9),
    .X(_1108_));
 sky130_fd_sc_hd__inv_1 _4722_ (.A(\dp.rf.rf[4][15] ),
    .Y(_1109_));
 sky130_fd_sc_hd__mux2i_1 _4723_ (.A0(\dp.rf.rf[1][15] ),
    .A1(\dp.rf.rf[5][15] ),
    .S(net9),
    .Y(_1110_));
 sky130_fd_sc_hd__a221oi_1 _4724_ (.A1(_1109_),
    .A2(_0173_),
    .B1(_1110_),
    .B2(net7),
    .C1(net8),
    .Y(_1111_));
 sky130_fd_sc_hd__a211oi_1 _4725_ (.A1(net8),
    .A2(_1108_),
    .B1(_1111_),
    .C1(_0265_),
    .Y(_1112_));
 sky130_fd_sc_hd__a31oi_1 _4726_ (.A1(net797),
    .A2(_1105_),
    .A3(_1107_),
    .B1(_1112_),
    .Y(_1113_));
 sky130_fd_sc_hd__a22oi_2 _4727_ (.A1(_1095_),
    .A2(_1103_),
    .B1(_1113_),
    .B2(net780),
    .Y(_3334_[0]));
 sky130_fd_sc_hd__mux4_2 _4728_ (.A0(\dp.rf.rf[16][14] ),
    .A1(\dp.rf.rf[17][14] ),
    .A2(\dp.rf.rf[18][14] ),
    .A3(\dp.rf.rf[19][14] ),
    .S0(net822),
    .S1(net14),
    .X(_1114_));
 sky130_fd_sc_hd__mux4_2 _4729_ (.A0(\dp.rf.rf[20][14] ),
    .A1(\dp.rf.rf[21][14] ),
    .A2(\dp.rf.rf[22][14] ),
    .A3(\dp.rf.rf[23][14] ),
    .S0(net822),
    .S1(net14),
    .X(_1115_));
 sky130_fd_sc_hd__mux4_2 _4730_ (.A0(\dp.rf.rf[24][14] ),
    .A1(\dp.rf.rf[25][14] ),
    .A2(\dp.rf.rf[26][14] ),
    .A3(\dp.rf.rf[27][14] ),
    .S0(net822),
    .S1(net14),
    .X(_1116_));
 sky130_fd_sc_hd__mux4_2 _4731_ (.A0(\dp.rf.rf[28][14] ),
    .A1(\dp.rf.rf[29][14] ),
    .A2(\dp.rf.rf[30][14] ),
    .A3(\dp.rf.rf[31][14] ),
    .S0(net822),
    .S1(net14),
    .X(_1117_));
 sky130_fd_sc_hd__mux4_2 _4732_ (.A0(_1114_),
    .A1(_1115_),
    .A2(_1116_),
    .A3(_1117_),
    .S0(net15),
    .S1(net16),
    .X(_1118_));
 sky130_fd_sc_hd__mux4_2 _4733_ (.A0(\dp.rf.rf[0][14] ),
    .A1(\dp.rf.rf[1][14] ),
    .A2(\dp.rf.rf[2][14] ),
    .A3(\dp.rf.rf[3][14] ),
    .S0(net822),
    .S1(net14),
    .X(_1119_));
 sky130_fd_sc_hd__mux4_2 _4734_ (.A0(\dp.rf.rf[4][14] ),
    .A1(\dp.rf.rf[5][14] ),
    .A2(\dp.rf.rf[6][14] ),
    .A3(\dp.rf.rf[7][14] ),
    .S0(net822),
    .S1(net14),
    .X(_1120_));
 sky130_fd_sc_hd__mux4_2 _4735_ (.A0(\dp.rf.rf[8][14] ),
    .A1(\dp.rf.rf[9][14] ),
    .A2(\dp.rf.rf[10][14] ),
    .A3(\dp.rf.rf[11][14] ),
    .S0(net822),
    .S1(net14),
    .X(_1121_));
 sky130_fd_sc_hd__mux4_2 _4736_ (.A0(\dp.rf.rf[12][14] ),
    .A1(\dp.rf.rf[13][14] ),
    .A2(\dp.rf.rf[14][14] ),
    .A3(\dp.rf.rf[15][14] ),
    .S0(net822),
    .S1(net14),
    .X(_1122_));
 sky130_fd_sc_hd__mux4_2 _4737_ (.A0(_1119_),
    .A1(_1120_),
    .A2(_1121_),
    .A3(_1122_),
    .S0(net15),
    .S1(net16),
    .X(_1123_));
 sky130_fd_sc_hd__mux2_8 _4738_ (.A0(_1118_),
    .A1(_1123_),
    .S(_0092_),
    .X(_1124_));
 sky130_fd_sc_hd__nand2_8 _4739_ (.A(_1124_),
    .B(_0351_),
    .Y(_1125_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_114 ();
 sky130_fd_sc_hd__a221oi_1 _4742_ (.A1(net5),
    .A2(net799),
    .B1(_0146_),
    .B2(net6),
    .C1(_0898_),
    .Y(_1128_));
 sky130_fd_sc_hd__mux2i_1 _4743_ (.A0(_1074_),
    .A1(_1128_),
    .S(_0902_),
    .Y(_3504_[0]));
 sky130_fd_sc_hd__nand2_1 _4744_ (.A(net782),
    .B(_3504_[0]),
    .Y(_1129_));
 sky130_fd_sc_hd__o21ai_4 _4745_ (.A1(_0148_),
    .A2(_1125_),
    .B1(_1129_),
    .Y(_1130_));
 sky130_fd_sc_hd__xnor2_1 _4746_ (.A(_1130_),
    .B(_0151_),
    .Y(_3339_[0]));
 sky130_fd_sc_hd__inv_1 _4747_ (.A(net263),
    .Y(_3343_[0]));
 sky130_fd_sc_hd__mux4_2 _4748_ (.A0(\dp.rf.rf[10][14] ),
    .A1(\dp.rf.rf[11][14] ),
    .A2(\dp.rf.rf[14][14] ),
    .A3(\dp.rf.rf[15][14] ),
    .S0(net809),
    .S1(net9),
    .X(_1131_));
 sky130_fd_sc_hd__nand2_1 _4749_ (.A(net8),
    .B(_1131_),
    .Y(_1132_));
 sky130_fd_sc_hd__mux4_2 _4750_ (.A0(net265),
    .A1(net266),
    .A2(net283),
    .A3(net284),
    .S0(net809),
    .S1(net9),
    .X(_1133_));
 sky130_fd_sc_hd__nand2_1 _4751_ (.A(_0186_),
    .B(_1133_),
    .Y(_1134_));
 sky130_fd_sc_hd__nand3_2 _4752_ (.A(net797),
    .B(_1132_),
    .C(_1134_),
    .Y(_1135_));
 sky130_fd_sc_hd__mux2_1 _4753_ (.A0(\dp.rf.rf[6][14] ),
    .A1(\dp.rf.rf[7][14] ),
    .S(net7),
    .X(_1136_));
 sky130_fd_sc_hd__o21ai_0 _4754_ (.A1(_0231_),
    .A2(_1136_),
    .B1(_0304_),
    .Y(_1137_));
 sky130_fd_sc_hd__a221oi_1 _4755_ (.A1(\dp.rf.rf[3][14] ),
    .A2(net7),
    .B1(net788),
    .B2(\dp.rf.rf[2][14] ),
    .C1(net791),
    .Y(_1138_));
 sky130_fd_sc_hd__inv_1 _4756_ (.A(\dp.rf.rf[4][14] ),
    .Y(_1139_));
 sky130_fd_sc_hd__mux2i_1 _4757_ (.A0(\dp.rf.rf[1][14] ),
    .A1(\dp.rf.rf[5][14] ),
    .S(net9),
    .Y(_1140_));
 sky130_fd_sc_hd__a221oi_1 _4758_ (.A1(_1139_),
    .A2(_0173_),
    .B1(_1140_),
    .B2(net7),
    .C1(net8),
    .Y(_1141_));
 sky130_fd_sc_hd__o22ai_1 _4759_ (.A1(\dp.rf.rf[0][14] ),
    .A2(net784),
    .B1(_1141_),
    .B2(_0265_),
    .Y(_1142_));
 sky130_fd_sc_hd__o21ai_2 _4760_ (.A1(_1137_),
    .A2(_1138_),
    .B1(_1142_),
    .Y(_1143_));
 sky130_fd_sc_hd__mux4_2 _4761_ (.A0(\dp.rf.rf[26][14] ),
    .A1(\dp.rf.rf[27][14] ),
    .A2(\dp.rf.rf[30][14] ),
    .A3(\dp.rf.rf[31][14] ),
    .S0(net809),
    .S1(net9),
    .X(_1144_));
 sky130_fd_sc_hd__nand2_1 _4762_ (.A(net8),
    .B(_1144_),
    .Y(_1145_));
 sky130_fd_sc_hd__mux4_2 _4763_ (.A0(\dp.rf.rf[24][14] ),
    .A1(\dp.rf.rf[25][14] ),
    .A2(\dp.rf.rf[28][14] ),
    .A3(\dp.rf.rf[29][14] ),
    .S0(net809),
    .S1(net9),
    .X(_1146_));
 sky130_fd_sc_hd__nand2_1 _4764_ (.A(_0186_),
    .B(_1146_),
    .Y(_1147_));
 sky130_fd_sc_hd__a31oi_2 _4765_ (.A1(net10),
    .A2(_1145_),
    .A3(_1147_),
    .B1(net794),
    .Y(_1148_));
 sky130_fd_sc_hd__mux2_1 _4766_ (.A0(\dp.rf.rf[22][14] ),
    .A1(\dp.rf.rf[23][14] ),
    .S(net809),
    .X(_1149_));
 sky130_fd_sc_hd__o21ai_0 _4767_ (.A1(_0231_),
    .A2(_1149_),
    .B1(_0304_),
    .Y(_1150_));
 sky130_fd_sc_hd__a221oi_1 _4768_ (.A1(\dp.rf.rf[19][14] ),
    .A2(net809),
    .B1(net788),
    .B2(\dp.rf.rf[18][14] ),
    .C1(net791),
    .Y(_1151_));
 sky130_fd_sc_hd__inv_1 _4769_ (.A(\dp.rf.rf[20][14] ),
    .Y(_1152_));
 sky130_fd_sc_hd__mux2i_1 _4770_ (.A0(\dp.rf.rf[17][14] ),
    .A1(\dp.rf.rf[21][14] ),
    .S(net9),
    .Y(_1153_));
 sky130_fd_sc_hd__a221oi_1 _4771_ (.A1(_1152_),
    .A2(_0173_),
    .B1(_1153_),
    .B2(net809),
    .C1(net8),
    .Y(_1154_));
 sky130_fd_sc_hd__o22ai_1 _4772_ (.A1(\dp.rf.rf[16][14] ),
    .A2(net784),
    .B1(_1154_),
    .B2(_0265_),
    .Y(_1155_));
 sky130_fd_sc_hd__o21ai_2 _4773_ (.A1(_1150_),
    .A2(_1151_),
    .B1(_1155_),
    .Y(_1156_));
 sky130_fd_sc_hd__a32oi_4 _4774_ (.A1(net780),
    .A2(_1135_),
    .A3(_1143_),
    .B1(_1148_),
    .B2(_1156_),
    .Y(_3342_[0]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_112 ();
 sky130_fd_sc_hd__a221oi_1 _4777_ (.A1(net815),
    .A2(net799),
    .B1(_0146_),
    .B2(net5),
    .C1(_0898_),
    .Y(_1159_));
 sky130_fd_sc_hd__mux2i_2 _4778_ (.A0(_1128_),
    .A1(_1159_),
    .S(_0902_),
    .Y(_3500_[0]));
 sky130_fd_sc_hd__nand2_1 _4779_ (.A(net782),
    .B(_3500_[0]),
    .Y(_1160_));
 sky130_fd_sc_hd__mux4_2 _4780_ (.A0(\dp.rf.rf[16][13] ),
    .A1(\dp.rf.rf[17][13] ),
    .A2(\dp.rf.rf[18][13] ),
    .A3(\dp.rf.rf[19][13] ),
    .S0(net13),
    .S1(net14),
    .X(_1161_));
 sky130_fd_sc_hd__mux4_2 _4781_ (.A0(\dp.rf.rf[20][13] ),
    .A1(\dp.rf.rf[21][13] ),
    .A2(\dp.rf.rf[22][13] ),
    .A3(\dp.rf.rf[23][13] ),
    .S0(net13),
    .S1(net14),
    .X(_1162_));
 sky130_fd_sc_hd__mux4_2 _4782_ (.A0(\dp.rf.rf[24][13] ),
    .A1(\dp.rf.rf[25][13] ),
    .A2(\dp.rf.rf[26][13] ),
    .A3(\dp.rf.rf[27][13] ),
    .S0(net13),
    .S1(net14),
    .X(_1163_));
 sky130_fd_sc_hd__mux4_2 _4783_ (.A0(\dp.rf.rf[28][13] ),
    .A1(\dp.rf.rf[29][13] ),
    .A2(\dp.rf.rf[30][13] ),
    .A3(\dp.rf.rf[31][13] ),
    .S0(net13),
    .S1(net14),
    .X(_1164_));
 sky130_fd_sc_hd__mux4_2 _4784_ (.A0(_1161_),
    .A1(_1162_),
    .A2(_1163_),
    .A3(_1164_),
    .S0(net818),
    .S1(net16),
    .X(_1165_));
 sky130_fd_sc_hd__nand2_2 _4785_ (.A(net17),
    .B(_1165_),
    .Y(_1166_));
 sky130_fd_sc_hd__mux4_2 _4786_ (.A0(\dp.rf.rf[0][13] ),
    .A1(\dp.rf.rf[1][13] ),
    .A2(\dp.rf.rf[2][13] ),
    .A3(\dp.rf.rf[3][13] ),
    .S0(net13),
    .S1(net819),
    .X(_1167_));
 sky130_fd_sc_hd__mux4_2 _4787_ (.A0(\dp.rf.rf[4][13] ),
    .A1(\dp.rf.rf[5][13] ),
    .A2(\dp.rf.rf[6][13] ),
    .A3(\dp.rf.rf[7][13] ),
    .S0(net13),
    .S1(net819),
    .X(_1168_));
 sky130_fd_sc_hd__mux4_2 _4788_ (.A0(\dp.rf.rf[8][13] ),
    .A1(\dp.rf.rf[9][13] ),
    .A2(\dp.rf.rf[10][13] ),
    .A3(\dp.rf.rf[11][13] ),
    .S0(net13),
    .S1(net14),
    .X(_1169_));
 sky130_fd_sc_hd__mux4_2 _4789_ (.A0(\dp.rf.rf[12][13] ),
    .A1(\dp.rf.rf[13][13] ),
    .A2(\dp.rf.rf[14][13] ),
    .A3(\dp.rf.rf[15][13] ),
    .S0(net13),
    .S1(net14),
    .X(_1170_));
 sky130_fd_sc_hd__mux4_2 _4790_ (.A0(_1167_),
    .A1(_1168_),
    .A2(_1169_),
    .A3(_1170_),
    .S0(net818),
    .S1(net16),
    .X(_1171_));
 sky130_fd_sc_hd__nand2_2 _4791_ (.A(_0092_),
    .B(_1171_),
    .Y(_1172_));
 sky130_fd_sc_hd__a21oi_4 _4792_ (.A1(_1166_),
    .A2(_1172_),
    .B1(_0111_),
    .Y(_1173_));
 sky130_fd_sc_hd__nand2_1 _4793_ (.A(_0121_),
    .B(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__nand2_2 _4794_ (.A(_1160_),
    .B(_1174_),
    .Y(_1175_));
 sky130_fd_sc_hd__xnor2_1 _4795_ (.A(_0151_),
    .B(_1175_),
    .Y(_3347_[0]));
 sky130_fd_sc_hd__inv_1 _4796_ (.A(_3347_[0]),
    .Y(_3351_[0]));
 sky130_fd_sc_hd__a221oi_1 _4797_ (.A1(\dp.rf.rf[11][13] ),
    .A2(net809),
    .B1(_0298_),
    .B2(\dp.rf.rf[10][13] ),
    .C1(_0259_),
    .Y(_1176_));
 sky130_fd_sc_hd__mux2_1 _4798_ (.A0(\dp.rf.rf[14][13] ),
    .A1(\dp.rf.rf[15][13] ),
    .S(net809),
    .X(_1177_));
 sky130_fd_sc_hd__o21ai_0 _4799_ (.A1(net800),
    .A2(_1177_),
    .B1(net786),
    .Y(_1178_));
 sky130_fd_sc_hd__mux4_2 _4800_ (.A0(\dp.rf.rf[8][13] ),
    .A1(\dp.rf.rf[9][13] ),
    .A2(\dp.rf.rf[12][13] ),
    .A3(\dp.rf.rf[13][13] ),
    .S0(net809),
    .S1(net9),
    .X(_1179_));
 sky130_fd_sc_hd__a21oi_1 _4801_ (.A1(_0186_),
    .A2(_1179_),
    .B1(_0255_),
    .Y(_1180_));
 sky130_fd_sc_hd__o21ai_2 _4802_ (.A1(_1176_),
    .A2(_1178_),
    .B1(_1180_),
    .Y(_1181_));
 sky130_fd_sc_hd__mux2i_1 _4803_ (.A0(\dp.rf.rf[6][13] ),
    .A1(\dp.rf.rf[7][13] ),
    .S(net812),
    .Y(_1182_));
 sky130_fd_sc_hd__mux2i_1 _4804_ (.A0(\dp.rf.rf[2][13] ),
    .A1(\dp.rf.rf[3][13] ),
    .S(net812),
    .Y(_1183_));
 sky130_fd_sc_hd__a221o_1 _4805_ (.A1(net9),
    .A2(_1182_),
    .B1(_1183_),
    .B2(_0513_),
    .C1(_0186_),
    .X(_1184_));
 sky130_fd_sc_hd__inv_1 _4806_ (.A(\dp.rf.rf[4][13] ),
    .Y(_1185_));
 sky130_fd_sc_hd__mux2i_1 _4807_ (.A0(\dp.rf.rf[1][13] ),
    .A1(\dp.rf.rf[5][13] ),
    .S(net9),
    .Y(_1186_));
 sky130_fd_sc_hd__a221oi_1 _4808_ (.A1(_1185_),
    .A2(_0173_),
    .B1(_1186_),
    .B2(net812),
    .C1(net8),
    .Y(_1187_));
 sky130_fd_sc_hd__o22ai_1 _4809_ (.A1(\dp.rf.rf[0][13] ),
    .A2(_0166_),
    .B1(_1187_),
    .B2(_0137_),
    .Y(_1188_));
 sky130_fd_sc_hd__nand3_2 _4810_ (.A(_0192_),
    .B(_1184_),
    .C(_1188_),
    .Y(_1189_));
 sky130_fd_sc_hd__mux4_2 _4811_ (.A0(\dp.rf.rf[26][13] ),
    .A1(\dp.rf.rf[27][13] ),
    .A2(\dp.rf.rf[30][13] ),
    .A3(\dp.rf.rf[31][13] ),
    .S0(net809),
    .S1(net9),
    .X(_1190_));
 sky130_fd_sc_hd__nand2_1 _4812_ (.A(net8),
    .B(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__mux4_2 _4813_ (.A0(\dp.rf.rf[24][13] ),
    .A1(\dp.rf.rf[25][13] ),
    .A2(\dp.rf.rf[28][13] ),
    .A3(\dp.rf.rf[29][13] ),
    .S0(net809),
    .S1(net9),
    .X(_1192_));
 sky130_fd_sc_hd__nand2_1 _4814_ (.A(_0186_),
    .B(_1192_),
    .Y(_1193_));
 sky130_fd_sc_hd__a31oi_2 _4815_ (.A1(net10),
    .A2(_1191_),
    .A3(_1193_),
    .B1(net794),
    .Y(_1194_));
 sky130_fd_sc_hd__mux2_1 _4816_ (.A0(\dp.rf.rf[22][13] ),
    .A1(\dp.rf.rf[23][13] ),
    .S(net809),
    .X(_1195_));
 sky130_fd_sc_hd__o21ai_0 _4817_ (.A1(net800),
    .A2(_1195_),
    .B1(net786),
    .Y(_1196_));
 sky130_fd_sc_hd__a221oi_1 _4818_ (.A1(\dp.rf.rf[19][13] ),
    .A2(net809),
    .B1(net788),
    .B2(\dp.rf.rf[18][13] ),
    .C1(net791),
    .Y(_1197_));
 sky130_fd_sc_hd__inv_1 _4819_ (.A(\dp.rf.rf[20][13] ),
    .Y(_1198_));
 sky130_fd_sc_hd__mux2i_1 _4820_ (.A0(\dp.rf.rf[17][13] ),
    .A1(\dp.rf.rf[21][13] ),
    .S(net9),
    .Y(_1199_));
 sky130_fd_sc_hd__a221oi_1 _4821_ (.A1(_1198_),
    .A2(_0173_),
    .B1(_1199_),
    .B2(net809),
    .C1(net8),
    .Y(_1200_));
 sky130_fd_sc_hd__o22ai_1 _4822_ (.A1(\dp.rf.rf[16][13] ),
    .A2(net784),
    .B1(_1200_),
    .B2(_0265_),
    .Y(_1201_));
 sky130_fd_sc_hd__o21ai_2 _4823_ (.A1(_1196_),
    .A2(_1197_),
    .B1(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__a32oi_4 _4824_ (.A1(net781),
    .A2(_1181_),
    .A3(_1189_),
    .B1(_1194_),
    .B2(_1202_),
    .Y(_1203_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_111 ();
 sky130_fd_sc_hd__mux4_2 _4826_ (.A0(\dp.rf.rf[16][12] ),
    .A1(\dp.rf.rf[17][12] ),
    .A2(\dp.rf.rf[18][12] ),
    .A3(\dp.rf.rf[19][12] ),
    .S0(net823),
    .S1(net821),
    .X(_1204_));
 sky130_fd_sc_hd__mux4_2 _4827_ (.A0(\dp.rf.rf[20][12] ),
    .A1(\dp.rf.rf[21][12] ),
    .A2(\dp.rf.rf[22][12] ),
    .A3(\dp.rf.rf[23][12] ),
    .S0(net823),
    .S1(net821),
    .X(_1205_));
 sky130_fd_sc_hd__mux4_2 _4828_ (.A0(\dp.rf.rf[24][12] ),
    .A1(\dp.rf.rf[25][12] ),
    .A2(\dp.rf.rf[26][12] ),
    .A3(\dp.rf.rf[27][12] ),
    .S0(net823),
    .S1(net821),
    .X(_1206_));
 sky130_fd_sc_hd__mux4_2 _4829_ (.A0(\dp.rf.rf[28][12] ),
    .A1(\dp.rf.rf[29][12] ),
    .A2(\dp.rf.rf[30][12] ),
    .A3(\dp.rf.rf[31][12] ),
    .S0(net823),
    .S1(net821),
    .X(_1207_));
 sky130_fd_sc_hd__mux4_2 _4830_ (.A0(_1204_),
    .A1(_1205_),
    .A2(_1206_),
    .A3(_1207_),
    .S0(net15),
    .S1(net16),
    .X(_1208_));
 sky130_fd_sc_hd__mux4_2 _4831_ (.A0(\dp.rf.rf[0][12] ),
    .A1(\dp.rf.rf[1][12] ),
    .A2(\dp.rf.rf[2][12] ),
    .A3(\dp.rf.rf[3][12] ),
    .S0(net823),
    .S1(net821),
    .X(_1209_));
 sky130_fd_sc_hd__mux4_2 _4832_ (.A0(\dp.rf.rf[4][12] ),
    .A1(\dp.rf.rf[5][12] ),
    .A2(\dp.rf.rf[6][12] ),
    .A3(\dp.rf.rf[7][12] ),
    .S0(net823),
    .S1(net821),
    .X(_1210_));
 sky130_fd_sc_hd__mux4_2 _4833_ (.A0(\dp.rf.rf[8][12] ),
    .A1(\dp.rf.rf[9][12] ),
    .A2(\dp.rf.rf[10][12] ),
    .A3(\dp.rf.rf[11][12] ),
    .S0(net823),
    .S1(net821),
    .X(_1211_));
 sky130_fd_sc_hd__mux4_2 _4834_ (.A0(\dp.rf.rf[12][12] ),
    .A1(\dp.rf.rf[13][12] ),
    .A2(\dp.rf.rf[14][12] ),
    .A3(\dp.rf.rf[15][12] ),
    .S0(net823),
    .S1(net821),
    .X(_1212_));
 sky130_fd_sc_hd__mux4_2 _4835_ (.A0(_1209_),
    .A1(_1210_),
    .A2(_1211_),
    .A3(_1212_),
    .S0(net15),
    .S1(net16),
    .X(_1213_));
 sky130_fd_sc_hd__mux2i_4 _4836_ (.A0(_1208_),
    .A1(_1213_),
    .S(_0092_),
    .Y(_1214_));
 sky130_fd_sc_hd__nor2_4 _4837_ (.A(_0111_),
    .B(_1214_),
    .Y(_1215_));
 sky130_fd_sc_hd__nand3_1 _4838_ (.A(net25),
    .B(_0347_),
    .C(_0897_),
    .Y(_1216_));
 sky130_fd_sc_hd__o21ai_0 _4839_ (.A1(net799),
    .A2(_0146_),
    .B1(net4),
    .Y(_1217_));
 sky130_fd_sc_hd__a21oi_1 _4840_ (.A1(_1216_),
    .A2(_1217_),
    .B1(_0121_),
    .Y(_1218_));
 sky130_fd_sc_hd__a21oi_2 _4841_ (.A1(_0121_),
    .A2(_1215_),
    .B1(_1218_),
    .Y(_1219_));
 sky130_fd_sc_hd__xor2_1 _4842_ (.A(_0151_),
    .B(_1219_),
    .X(_3355_[0]));
 sky130_fd_sc_hd__inv_1 _4843_ (.A(_3355_[0]),
    .Y(_3359_[0]));
 sky130_fd_sc_hd__mux4_2 _4844_ (.A0(\dp.rf.rf[2][12] ),
    .A1(\dp.rf.rf[3][12] ),
    .A2(\dp.rf.rf[6][12] ),
    .A3(\dp.rf.rf[7][12] ),
    .S0(net7),
    .S1(net9),
    .X(_1220_));
 sky130_fd_sc_hd__nand2_1 _4845_ (.A(_0304_),
    .B(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hd__inv_1 _4846_ (.A(\dp.rf.rf[4][12] ),
    .Y(_1222_));
 sky130_fd_sc_hd__mux2i_1 _4847_ (.A0(\dp.rf.rf[1][12] ),
    .A1(\dp.rf.rf[5][12] ),
    .S(net9),
    .Y(_1223_));
 sky130_fd_sc_hd__a221oi_1 _4848_ (.A1(_1222_),
    .A2(_0173_),
    .B1(_1223_),
    .B2(net7),
    .C1(net8),
    .Y(_1224_));
 sky130_fd_sc_hd__o22ai_1 _4849_ (.A1(\dp.rf.rf[0][12] ),
    .A2(net784),
    .B1(_1224_),
    .B2(net790),
    .Y(_1225_));
 sky130_fd_sc_hd__mux4_2 _4850_ (.A0(\dp.rf.rf[8][12] ),
    .A1(\dp.rf.rf[9][12] ),
    .A2(\dp.rf.rf[12][12] ),
    .A3(\dp.rf.rf[13][12] ),
    .S0(net7),
    .S1(net9),
    .X(_1226_));
 sky130_fd_sc_hd__mux4_2 _4851_ (.A0(\dp.rf.rf[10][12] ),
    .A1(\dp.rf.rf[11][12] ),
    .A2(\dp.rf.rf[14][12] ),
    .A3(\dp.rf.rf[15][12] ),
    .S0(net7),
    .S1(net9),
    .X(_1227_));
 sky130_fd_sc_hd__mux2i_1 _4852_ (.A0(_1226_),
    .A1(_1227_),
    .S(net8),
    .Y(_1228_));
 sky130_fd_sc_hd__a22oi_2 _4853_ (.A1(_1221_),
    .A2(_1225_),
    .B1(_1228_),
    .B2(net797),
    .Y(_1229_));
 sky130_fd_sc_hd__mux4_2 _4854_ (.A0(\dp.rf.rf[26][12] ),
    .A1(\dp.rf.rf[27][12] ),
    .A2(\dp.rf.rf[30][12] ),
    .A3(\dp.rf.rf[31][12] ),
    .S0(net809),
    .S1(net9),
    .X(_1230_));
 sky130_fd_sc_hd__nand2_1 _4855_ (.A(net8),
    .B(_1230_),
    .Y(_1231_));
 sky130_fd_sc_hd__mux4_2 _4856_ (.A0(\dp.rf.rf[24][12] ),
    .A1(\dp.rf.rf[25][12] ),
    .A2(\dp.rf.rf[28][12] ),
    .A3(\dp.rf.rf[29][12] ),
    .S0(net7),
    .S1(net9),
    .X(_1232_));
 sky130_fd_sc_hd__a21oi_1 _4857_ (.A1(_0186_),
    .A2(_1232_),
    .B1(_0255_),
    .Y(_1233_));
 sky130_fd_sc_hd__a21oi_1 _4858_ (.A1(_1231_),
    .A2(_1233_),
    .B1(net794),
    .Y(_1234_));
 sky130_fd_sc_hd__mux2_1 _4859_ (.A0(\dp.rf.rf[22][12] ),
    .A1(\dp.rf.rf[23][12] ),
    .S(net7),
    .X(_1235_));
 sky130_fd_sc_hd__o21ai_0 _4860_ (.A1(_0231_),
    .A2(_1235_),
    .B1(_0304_),
    .Y(_1236_));
 sky130_fd_sc_hd__a221oi_1 _4861_ (.A1(\dp.rf.rf[19][12] ),
    .A2(net7),
    .B1(net788),
    .B2(\dp.rf.rf[18][12] ),
    .C1(net791),
    .Y(_1237_));
 sky130_fd_sc_hd__inv_1 _4862_ (.A(\dp.rf.rf[20][12] ),
    .Y(_1238_));
 sky130_fd_sc_hd__mux2i_1 _4863_ (.A0(\dp.rf.rf[17][12] ),
    .A1(\dp.rf.rf[21][12] ),
    .S(net9),
    .Y(_1239_));
 sky130_fd_sc_hd__a221oi_1 _4864_ (.A1(_1238_),
    .A2(_0173_),
    .B1(_1239_),
    .B2(net7),
    .C1(net8),
    .Y(_1240_));
 sky130_fd_sc_hd__o22ai_1 _4865_ (.A1(\dp.rf.rf[16][12] ),
    .A2(net784),
    .B1(_1240_),
    .B2(net790),
    .Y(_1241_));
 sky130_fd_sc_hd__o21ai_0 _4866_ (.A1(_1236_),
    .A2(_1237_),
    .B1(_1241_),
    .Y(_1242_));
 sky130_fd_sc_hd__a22oi_2 _4867_ (.A1(net780),
    .A2(_1229_),
    .B1(_1234_),
    .B2(_1242_),
    .Y(_3358_[0]));
 sky130_fd_sc_hd__mux4_2 _4868_ (.A0(\dp.rf.rf[16][11] ),
    .A1(\dp.rf.rf[17][11] ),
    .A2(\dp.rf.rf[18][11] ),
    .A3(\dp.rf.rf[19][11] ),
    .S0(net823),
    .S1(net14),
    .X(_1243_));
 sky130_fd_sc_hd__mux4_2 _4869_ (.A0(\dp.rf.rf[20][11] ),
    .A1(\dp.rf.rf[21][11] ),
    .A2(\dp.rf.rf[22][11] ),
    .A3(\dp.rf.rf[23][11] ),
    .S0(net823),
    .S1(net14),
    .X(_1244_));
 sky130_fd_sc_hd__mux4_2 _4870_ (.A0(\dp.rf.rf[24][11] ),
    .A1(\dp.rf.rf[25][11] ),
    .A2(\dp.rf.rf[26][11] ),
    .A3(\dp.rf.rf[27][11] ),
    .S0(net823),
    .S1(net14),
    .X(_1245_));
 sky130_fd_sc_hd__mux4_2 _4871_ (.A0(\dp.rf.rf[28][11] ),
    .A1(\dp.rf.rf[29][11] ),
    .A2(\dp.rf.rf[30][11] ),
    .A3(\dp.rf.rf[31][11] ),
    .S0(net823),
    .S1(net14),
    .X(_1246_));
 sky130_fd_sc_hd__mux4_2 _4872_ (.A0(_1243_),
    .A1(_1244_),
    .A2(_1245_),
    .A3(_1246_),
    .S0(net15),
    .S1(net16),
    .X(_1247_));
 sky130_fd_sc_hd__mux4_2 _4873_ (.A0(\dp.rf.rf[0][11] ),
    .A1(\dp.rf.rf[1][11] ),
    .A2(\dp.rf.rf[2][11] ),
    .A3(\dp.rf.rf[3][11] ),
    .S0(net824),
    .S1(net821),
    .X(_1248_));
 sky130_fd_sc_hd__mux4_2 _4874_ (.A0(\dp.rf.rf[4][11] ),
    .A1(\dp.rf.rf[5][11] ),
    .A2(\dp.rf.rf[6][11] ),
    .A3(\dp.rf.rf[7][11] ),
    .S0(net824),
    .S1(net821),
    .X(_1249_));
 sky130_fd_sc_hd__mux4_2 _4875_ (.A0(\dp.rf.rf[8][11] ),
    .A1(\dp.rf.rf[9][11] ),
    .A2(\dp.rf.rf[10][11] ),
    .A3(\dp.rf.rf[11][11] ),
    .S0(net824),
    .S1(net821),
    .X(_1250_));
 sky130_fd_sc_hd__mux4_2 _4876_ (.A0(\dp.rf.rf[12][11] ),
    .A1(\dp.rf.rf[13][11] ),
    .A2(\dp.rf.rf[14][11] ),
    .A3(\dp.rf.rf[15][11] ),
    .S0(net824),
    .S1(net821),
    .X(_1251_));
 sky130_fd_sc_hd__mux4_2 _4877_ (.A0(_1248_),
    .A1(_1249_),
    .A2(_1250_),
    .A3(_1251_),
    .S0(net15),
    .S1(net16),
    .X(_1252_));
 sky130_fd_sc_hd__a22o_4 _4878_ (.A1(net17),
    .A2(_1247_),
    .B1(_1252_),
    .B2(_0337_),
    .X(_1253_));
 sky130_fd_sc_hd__nand2_1 _4879_ (.A(_0121_),
    .B(_1253_),
    .Y(_1254_));
 sky130_fd_sc_hd__and3_4 _4880_ (.A(_0901_),
    .B(_0897_),
    .C(_0349_),
    .X(_1255_));
 sky130_fd_sc_hd__a221o_4 _4881_ (.A1(net30),
    .A2(_0139_),
    .B1(_0146_),
    .B2(net13),
    .C1(_1255_),
    .X(_3492_[0]));
 sky130_fd_sc_hd__nand2_1 _4882_ (.A(_0148_),
    .B(_3492_[0]),
    .Y(_1256_));
 sky130_fd_sc_hd__nand2_1 _4883_ (.A(_1254_),
    .B(_1256_),
    .Y(_1257_));
 sky130_fd_sc_hd__xnor2_1 _4884_ (.A(_0151_),
    .B(_1257_),
    .Y(_3363_[0]));
 sky130_fd_sc_hd__inv_1 _4885_ (.A(_3363_[0]),
    .Y(_3367_[0]));
 sky130_fd_sc_hd__a221oi_1 _4886_ (.A1(\dp.rf.rf[27][11] ),
    .A2(net7),
    .B1(net788),
    .B2(\dp.rf.rf[26][11] ),
    .C1(net791),
    .Y(_1258_));
 sky130_fd_sc_hd__nor2b_1 _4887_ (.A(net7),
    .B_N(\dp.rf.rf[30][11] ),
    .Y(_1259_));
 sky130_fd_sc_hd__a211oi_1 _4888_ (.A1(\dp.rf.rf[31][11] ),
    .A2(net7),
    .B1(_0231_),
    .C1(_1259_),
    .Y(_1260_));
 sky130_fd_sc_hd__mux4_2 _4889_ (.A0(\dp.rf.rf[24][11] ),
    .A1(\dp.rf.rf[25][11] ),
    .A2(\dp.rf.rf[28][11] ),
    .A3(\dp.rf.rf[29][11] ),
    .S0(net7),
    .S1(net9),
    .X(_1261_));
 sky130_fd_sc_hd__a21oi_1 _4890_ (.A1(_0186_),
    .A2(_1261_),
    .B1(_0255_),
    .Y(_1262_));
 sky130_fd_sc_hd__o31ai_1 _4891_ (.A1(_0477_),
    .A2(_1258_),
    .A3(_1260_),
    .B1(_1262_),
    .Y(_1263_));
 sky130_fd_sc_hd__mux2_1 _4892_ (.A0(\dp.rf.rf[22][11] ),
    .A1(\dp.rf.rf[23][11] ),
    .S(net7),
    .X(_1264_));
 sky130_fd_sc_hd__o21ai_0 _4893_ (.A1(_0231_),
    .A2(_1264_),
    .B1(_0304_),
    .Y(_1265_));
 sky130_fd_sc_hd__a221oi_1 _4894_ (.A1(\dp.rf.rf[19][11] ),
    .A2(net7),
    .B1(net788),
    .B2(\dp.rf.rf[18][11] ),
    .C1(net791),
    .Y(_1266_));
 sky130_fd_sc_hd__inv_1 _4895_ (.A(\dp.rf.rf[20][11] ),
    .Y(_1267_));
 sky130_fd_sc_hd__mux2i_1 _4896_ (.A0(\dp.rf.rf[17][11] ),
    .A1(\dp.rf.rf[21][11] ),
    .S(net9),
    .Y(_1268_));
 sky130_fd_sc_hd__a221oi_1 _4897_ (.A1(_1267_),
    .A2(_0173_),
    .B1(_1268_),
    .B2(net7),
    .C1(net8),
    .Y(_1269_));
 sky130_fd_sc_hd__o22ai_1 _4898_ (.A1(\dp.rf.rf[16][11] ),
    .A2(net784),
    .B1(_1269_),
    .B2(net790),
    .Y(_1270_));
 sky130_fd_sc_hd__o21ai_2 _4899_ (.A1(_1265_),
    .A2(_1266_),
    .B1(_1270_),
    .Y(_1271_));
 sky130_fd_sc_hd__mux4_2 _4900_ (.A0(\dp.rf.rf[8][11] ),
    .A1(\dp.rf.rf[9][11] ),
    .A2(\dp.rf.rf[12][11] ),
    .A3(\dp.rf.rf[13][11] ),
    .S0(net7),
    .S1(net9),
    .X(_1272_));
 sky130_fd_sc_hd__nand2_1 _4901_ (.A(_0186_),
    .B(_1272_),
    .Y(_1273_));
 sky130_fd_sc_hd__mux4_2 _4902_ (.A0(\dp.rf.rf[10][11] ),
    .A1(\dp.rf.rf[11][11] ),
    .A2(\dp.rf.rf[14][11] ),
    .A3(\dp.rf.rf[15][11] ),
    .S0(net7),
    .S1(net9),
    .X(_1274_));
 sky130_fd_sc_hd__nand2_1 _4903_ (.A(net8),
    .B(_1274_),
    .Y(_1275_));
 sky130_fd_sc_hd__mux4_2 _4904_ (.A0(\dp.rf.rf[2][11] ),
    .A1(\dp.rf.rf[3][11] ),
    .A2(\dp.rf.rf[6][11] ),
    .A3(\dp.rf.rf[7][11] ),
    .S0(net7),
    .S1(net9),
    .X(_1276_));
 sky130_fd_sc_hd__inv_1 _4905_ (.A(\dp.rf.rf[4][11] ),
    .Y(_1277_));
 sky130_fd_sc_hd__mux2i_1 _4906_ (.A0(\dp.rf.rf[1][11] ),
    .A1(\dp.rf.rf[5][11] ),
    .S(net9),
    .Y(_1278_));
 sky130_fd_sc_hd__a221oi_1 _4907_ (.A1(_1277_),
    .A2(_0173_),
    .B1(_1278_),
    .B2(net7),
    .C1(net8),
    .Y(_1279_));
 sky130_fd_sc_hd__a211oi_2 _4908_ (.A1(net8),
    .A2(_1276_),
    .B1(_1279_),
    .C1(net790),
    .Y(_1280_));
 sky130_fd_sc_hd__a31oi_4 _4909_ (.A1(net797),
    .A2(_1273_),
    .A3(_1275_),
    .B1(_1280_),
    .Y(_1281_));
 sky130_fd_sc_hd__a32oi_4 _4910_ (.A1(_0620_),
    .A2(_1263_),
    .A3(_1271_),
    .B1(_1281_),
    .B2(net780),
    .Y(_3366_[0]));
 sky130_fd_sc_hd__and2_4 _4911_ (.A(net816),
    .B(_0347_),
    .X(_3488_[0]));
 sky130_fd_sc_hd__mux4_2 _4912_ (.A0(\dp.rf.rf[16][10] ),
    .A1(\dp.rf.rf[17][10] ),
    .A2(\dp.rf.rf[18][10] ),
    .A3(\dp.rf.rf[19][10] ),
    .S0(net13),
    .S1(net14),
    .X(_1282_));
 sky130_fd_sc_hd__mux4_2 _4913_ (.A0(\dp.rf.rf[20][10] ),
    .A1(\dp.rf.rf[21][10] ),
    .A2(\dp.rf.rf[22][10] ),
    .A3(\dp.rf.rf[23][10] ),
    .S0(net13),
    .S1(net14),
    .X(_1283_));
 sky130_fd_sc_hd__mux4_2 _4914_ (.A0(\dp.rf.rf[24][10] ),
    .A1(\dp.rf.rf[25][10] ),
    .A2(\dp.rf.rf[26][10] ),
    .A3(\dp.rf.rf[27][10] ),
    .S0(net13),
    .S1(net14),
    .X(_1284_));
 sky130_fd_sc_hd__mux4_2 _4915_ (.A0(\dp.rf.rf[28][10] ),
    .A1(\dp.rf.rf[29][10] ),
    .A2(\dp.rf.rf[30][10] ),
    .A3(\dp.rf.rf[31][10] ),
    .S0(net13),
    .S1(net14),
    .X(_1285_));
 sky130_fd_sc_hd__mux4_2 _4916_ (.A0(_1282_),
    .A1(_1283_),
    .A2(_1284_),
    .A3(_1285_),
    .S0(net15),
    .S1(net16),
    .X(_1286_));
 sky130_fd_sc_hd__nand2_2 _4917_ (.A(net17),
    .B(_1286_),
    .Y(_1287_));
 sky130_fd_sc_hd__mux4_2 _4918_ (.A0(\dp.rf.rf[0][10] ),
    .A1(\dp.rf.rf[1][10] ),
    .A2(\dp.rf.rf[2][10] ),
    .A3(\dp.rf.rf[3][10] ),
    .S0(net13),
    .S1(net14),
    .X(_1288_));
 sky130_fd_sc_hd__mux4_2 _4919_ (.A0(\dp.rf.rf[4][10] ),
    .A1(\dp.rf.rf[5][10] ),
    .A2(\dp.rf.rf[6][10] ),
    .A3(\dp.rf.rf[7][10] ),
    .S0(net13),
    .S1(net14),
    .X(_1289_));
 sky130_fd_sc_hd__mux4_2 _4920_ (.A0(\dp.rf.rf[8][10] ),
    .A1(\dp.rf.rf[9][10] ),
    .A2(\dp.rf.rf[10][10] ),
    .A3(\dp.rf.rf[11][10] ),
    .S0(net13),
    .S1(net14),
    .X(_1290_));
 sky130_fd_sc_hd__mux4_2 _4921_ (.A0(\dp.rf.rf[12][10] ),
    .A1(\dp.rf.rf[13][10] ),
    .A2(\dp.rf.rf[14][10] ),
    .A3(\dp.rf.rf[15][10] ),
    .S0(net13),
    .S1(net14),
    .X(_1291_));
 sky130_fd_sc_hd__mux4_2 _4922_ (.A0(_1288_),
    .A1(_1289_),
    .A2(_1290_),
    .A3(_1291_),
    .S0(net818),
    .S1(net16),
    .X(_1292_));
 sky130_fd_sc_hd__nand2_2 _4923_ (.A(_0092_),
    .B(_1292_),
    .Y(_1293_));
 sky130_fd_sc_hd__nand2_4 _4924_ (.A(_1287_),
    .B(_1293_),
    .Y(_1294_));
 sky130_fd_sc_hd__nand2_4 _4925_ (.A(_0351_),
    .B(_1294_),
    .Y(_1295_));
 sky130_fd_sc_hd__nor2_1 _4926_ (.A(_0148_),
    .B(_1295_),
    .Y(_1296_));
 sky130_fd_sc_hd__a21oi_2 _4927_ (.A1(_0148_),
    .A2(_3488_[0]),
    .B1(_1296_),
    .Y(_1297_));
 sky130_fd_sc_hd__xor2_1 _4928_ (.A(_0151_),
    .B(_1297_),
    .X(_3371_[0]));
 sky130_fd_sc_hd__inv_1 _4929_ (.A(_3371_[0]),
    .Y(_3375_[0]));
 sky130_fd_sc_hd__mux4_2 _4930_ (.A0(\dp.rf.rf[26][10] ),
    .A1(\dp.rf.rf[27][10] ),
    .A2(\dp.rf.rf[30][10] ),
    .A3(\dp.rf.rf[31][10] ),
    .S0(net809),
    .S1(net9),
    .X(_1298_));
 sky130_fd_sc_hd__mux4_2 _4931_ (.A0(\dp.rf.rf[24][10] ),
    .A1(\dp.rf.rf[25][10] ),
    .A2(\dp.rf.rf[28][10] ),
    .A3(\dp.rf.rf[29][10] ),
    .S0(net809),
    .S1(net9),
    .X(_1299_));
 sky130_fd_sc_hd__a221o_4 _4932_ (.A1(net786),
    .A2(_1298_),
    .B1(_1299_),
    .B2(_0186_),
    .C1(_0255_),
    .X(_1300_));
 sky130_fd_sc_hd__mux2_1 _4933_ (.A0(\dp.rf.rf[22][10] ),
    .A1(\dp.rf.rf[23][10] ),
    .S(net809),
    .X(_1301_));
 sky130_fd_sc_hd__o21ai_0 _4934_ (.A1(_0231_),
    .A2(_1301_),
    .B1(net786),
    .Y(_1302_));
 sky130_fd_sc_hd__a221oi_1 _4935_ (.A1(\dp.rf.rf[19][10] ),
    .A2(net809),
    .B1(net788),
    .B2(\dp.rf.rf[18][10] ),
    .C1(net791),
    .Y(_1303_));
 sky130_fd_sc_hd__inv_1 _4936_ (.A(\dp.rf.rf[20][10] ),
    .Y(_1304_));
 sky130_fd_sc_hd__mux2i_1 _4937_ (.A0(\dp.rf.rf[17][10] ),
    .A1(\dp.rf.rf[21][10] ),
    .S(net9),
    .Y(_1305_));
 sky130_fd_sc_hd__a221oi_1 _4938_ (.A1(_1304_),
    .A2(_0173_),
    .B1(_1305_),
    .B2(net809),
    .C1(net8),
    .Y(_1306_));
 sky130_fd_sc_hd__o22ai_1 _4939_ (.A1(\dp.rf.rf[16][10] ),
    .A2(net784),
    .B1(_1306_),
    .B2(_0265_),
    .Y(_1307_));
 sky130_fd_sc_hd__o21ai_2 _4940_ (.A1(_1302_),
    .A2(_1303_),
    .B1(_1307_),
    .Y(_1308_));
 sky130_fd_sc_hd__mux4_2 _4941_ (.A0(\dp.rf.rf[10][10] ),
    .A1(\dp.rf.rf[11][10] ),
    .A2(\dp.rf.rf[14][10] ),
    .A3(\dp.rf.rf[15][10] ),
    .S0(net812),
    .S1(net9),
    .X(_1309_));
 sky130_fd_sc_hd__nand2_1 _4942_ (.A(net786),
    .B(_1309_),
    .Y(_1310_));
 sky130_fd_sc_hd__mux4_2 _4943_ (.A0(\dp.rf.rf[8][10] ),
    .A1(\dp.rf.rf[9][10] ),
    .A2(\dp.rf.rf[12][10] ),
    .A3(\dp.rf.rf[13][10] ),
    .S0(net812),
    .S1(net9),
    .X(_1311_));
 sky130_fd_sc_hd__a21oi_1 _4944_ (.A1(_0186_),
    .A2(_1311_),
    .B1(_0255_),
    .Y(_1312_));
 sky130_fd_sc_hd__a21oi_1 _4945_ (.A1(_1310_),
    .A2(_1312_),
    .B1(_0293_),
    .Y(_1313_));
 sky130_fd_sc_hd__mux2_1 _4946_ (.A0(\dp.rf.rf[6][10] ),
    .A1(\dp.rf.rf[7][10] ),
    .S(net7),
    .X(_1314_));
 sky130_fd_sc_hd__o21ai_0 _4947_ (.A1(net800),
    .A2(_1314_),
    .B1(net786),
    .Y(_1315_));
 sky130_fd_sc_hd__a221oi_1 _4948_ (.A1(\dp.rf.rf[3][10] ),
    .A2(net812),
    .B1(_0298_),
    .B2(\dp.rf.rf[2][10] ),
    .C1(net791),
    .Y(_1316_));
 sky130_fd_sc_hd__inv_1 _4949_ (.A(\dp.rf.rf[4][10] ),
    .Y(_1317_));
 sky130_fd_sc_hd__mux2i_1 _4950_ (.A0(\dp.rf.rf[1][10] ),
    .A1(\dp.rf.rf[5][10] ),
    .S(net9),
    .Y(_1318_));
 sky130_fd_sc_hd__a221oi_1 _4951_ (.A1(_1317_),
    .A2(_0173_),
    .B1(_1318_),
    .B2(net7),
    .C1(net8),
    .Y(_1319_));
 sky130_fd_sc_hd__o22ai_1 _4952_ (.A1(\dp.rf.rf[0][10] ),
    .A2(net784),
    .B1(_1319_),
    .B2(_0265_),
    .Y(_1320_));
 sky130_fd_sc_hd__o21ai_2 _4953_ (.A1(_1315_),
    .A2(_1316_),
    .B1(_1320_),
    .Y(_1321_));
 sky130_fd_sc_hd__a32oi_4 _4954_ (.A1(net783),
    .A2(_1300_),
    .A3(_1308_),
    .B1(_1313_),
    .B2(_1321_),
    .Y(_3374_[0]));
 sky130_fd_sc_hd__mux4_2 _4955_ (.A0(\dp.rf.rf[4][9] ),
    .A1(\dp.rf.rf[5][9] ),
    .A2(\dp.rf.rf[6][9] ),
    .A3(\dp.rf.rf[7][9] ),
    .S0(net13),
    .S1(net14),
    .X(_1322_));
 sky130_fd_sc_hd__mux4_2 _4956_ (.A0(\dp.rf.rf[12][9] ),
    .A1(\dp.rf.rf[13][9] ),
    .A2(\dp.rf.rf[14][9] ),
    .A3(\dp.rf.rf[15][9] ),
    .S0(net13),
    .S1(net14),
    .X(_1323_));
 sky130_fd_sc_hd__mux2_4 _4957_ (.A0(_1322_),
    .A1(_1323_),
    .S(net16),
    .X(_1324_));
 sky130_fd_sc_hd__mux4_2 _4958_ (.A0(\dp.rf.rf[0][9] ),
    .A1(\dp.rf.rf[1][9] ),
    .A2(\dp.rf.rf[2][9] ),
    .A3(\dp.rf.rf[3][9] ),
    .S0(net13),
    .S1(net14),
    .X(_1325_));
 sky130_fd_sc_hd__mux4_2 _4959_ (.A0(\dp.rf.rf[8][9] ),
    .A1(\dp.rf.rf[9][9] ),
    .A2(\dp.rf.rf[10][9] ),
    .A3(\dp.rf.rf[11][9] ),
    .S0(net13),
    .S1(net14),
    .X(_1326_));
 sky130_fd_sc_hd__mux2i_1 _4960_ (.A0(_1325_),
    .A1(_1326_),
    .S(net16),
    .Y(_1327_));
 sky130_fd_sc_hd__nor2_1 _4961_ (.A(net818),
    .B(_1327_),
    .Y(_1328_));
 sky130_fd_sc_hd__a21oi_4 _4962_ (.A1(net818),
    .A2(_1324_),
    .B1(_1328_),
    .Y(_1329_));
 sky130_fd_sc_hd__mux4_2 _4963_ (.A0(\dp.rf.rf[16][9] ),
    .A1(\dp.rf.rf[17][9] ),
    .A2(\dp.rf.rf[18][9] ),
    .A3(\dp.rf.rf[19][9] ),
    .S0(net13),
    .S1(net14),
    .X(_1330_));
 sky130_fd_sc_hd__mux4_2 _4964_ (.A0(\dp.rf.rf[20][9] ),
    .A1(\dp.rf.rf[21][9] ),
    .A2(\dp.rf.rf[22][9] ),
    .A3(\dp.rf.rf[23][9] ),
    .S0(net13),
    .S1(net14),
    .X(_1331_));
 sky130_fd_sc_hd__mux4_2 _4965_ (.A0(\dp.rf.rf[24][9] ),
    .A1(\dp.rf.rf[25][9] ),
    .A2(\dp.rf.rf[26][9] ),
    .A3(\dp.rf.rf[27][9] ),
    .S0(net13),
    .S1(net820),
    .X(_1332_));
 sky130_fd_sc_hd__mux4_2 _4966_ (.A0(\dp.rf.rf[28][9] ),
    .A1(\dp.rf.rf[29][9] ),
    .A2(\dp.rf.rf[30][9] ),
    .A3(\dp.rf.rf[31][9] ),
    .S0(net13),
    .S1(net820),
    .X(_1333_));
 sky130_fd_sc_hd__mux4_2 _4967_ (.A0(_1330_),
    .A1(_1331_),
    .A2(_1332_),
    .A3(_1333_),
    .S0(net818),
    .S1(net16),
    .X(_1334_));
 sky130_fd_sc_hd__nand2_2 _4968_ (.A(net17),
    .B(_1334_),
    .Y(_1335_));
 sky130_fd_sc_hd__o21a_4 _4969_ (.A1(_0492_),
    .A2(_1329_),
    .B1(_1335_),
    .X(_1336_));
 sky130_fd_sc_hd__and2_4 _4970_ (.A(net22),
    .B(_0347_),
    .X(_3484_[0]));
 sky130_fd_sc_hd__nand2_1 _4971_ (.A(_0148_),
    .B(_3484_[0]),
    .Y(_1337_));
 sky130_fd_sc_hd__o21ai_2 _4972_ (.A1(_0148_),
    .A2(_1336_),
    .B1(_1337_),
    .Y(_1338_));
 sky130_fd_sc_hd__xnor2_1 _4973_ (.A(_0151_),
    .B(_1338_),
    .Y(_3379_[0]));
 sky130_fd_sc_hd__inv_1 _4974_ (.A(_3379_[0]),
    .Y(_3383_[0]));
 sky130_fd_sc_hd__nor2b_1 _4975_ (.A(net810),
    .B_N(\dp.rf.rf[22][9] ),
    .Y(_1339_));
 sky130_fd_sc_hd__a211oi_1 _4976_ (.A1(\dp.rf.rf[23][9] ),
    .A2(net810),
    .B1(_0231_),
    .C1(_1339_),
    .Y(_1340_));
 sky130_fd_sc_hd__a221oi_1 _4977_ (.A1(\dp.rf.rf[19][9] ),
    .A2(net810),
    .B1(_0298_),
    .B2(\dp.rf.rf[18][9] ),
    .C1(_0259_),
    .Y(_1341_));
 sky130_fd_sc_hd__inv_1 _4978_ (.A(\dp.rf.rf[20][9] ),
    .Y(_1342_));
 sky130_fd_sc_hd__mux2i_1 _4979_ (.A0(\dp.rf.rf[17][9] ),
    .A1(\dp.rf.rf[21][9] ),
    .S(net804),
    .Y(_1343_));
 sky130_fd_sc_hd__a221oi_1 _4980_ (.A1(_1342_),
    .A2(net801),
    .B1(_1343_),
    .B2(net810),
    .C1(net8),
    .Y(_1344_));
 sky130_fd_sc_hd__o22ai_1 _4981_ (.A1(\dp.rf.rf[16][9] ),
    .A2(net784),
    .B1(_1344_),
    .B2(_0265_),
    .Y(_1345_));
 sky130_fd_sc_hd__o31ai_2 _4982_ (.A1(_0477_),
    .A2(_1340_),
    .A3(_1341_),
    .B1(_1345_),
    .Y(_1346_));
 sky130_fd_sc_hd__a221oi_1 _4983_ (.A1(\dp.rf.rf[27][9] ),
    .A2(net810),
    .B1(_0298_),
    .B2(\dp.rf.rf[26][9] ),
    .C1(_0259_),
    .Y(_1347_));
 sky130_fd_sc_hd__mux2_1 _4984_ (.A0(\dp.rf.rf[30][9] ),
    .A1(\dp.rf.rf[31][9] ),
    .S(net810),
    .X(_1348_));
 sky130_fd_sc_hd__o21ai_0 _4985_ (.A1(_0231_),
    .A2(_1348_),
    .B1(net8),
    .Y(_1349_));
 sky130_fd_sc_hd__mux4_2 _4986_ (.A0(\dp.rf.rf[24][9] ),
    .A1(\dp.rf.rf[25][9] ),
    .A2(\dp.rf.rf[28][9] ),
    .A3(\dp.rf.rf[29][9] ),
    .S0(net810),
    .S1(net805),
    .X(_1350_));
 sky130_fd_sc_hd__a21oi_1 _4987_ (.A1(_0186_),
    .A2(_1350_),
    .B1(_0192_),
    .Y(_1351_));
 sky130_fd_sc_hd__o21ai_2 _4988_ (.A1(_1347_),
    .A2(_1349_),
    .B1(_1351_),
    .Y(_1352_));
 sky130_fd_sc_hd__mux4_2 _4989_ (.A0(\dp.rf.rf[2][9] ),
    .A1(\dp.rf.rf[3][9] ),
    .A2(\dp.rf.rf[6][9] ),
    .A3(\dp.rf.rf[7][9] ),
    .S0(net812),
    .S1(net805),
    .X(_1353_));
 sky130_fd_sc_hd__nand2_1 _4990_ (.A(net8),
    .B(_1353_),
    .Y(_1354_));
 sky130_fd_sc_hd__mux2_1 _4991_ (.A0(\dp.rf.rf[1][9] ),
    .A1(\dp.rf.rf[5][9] ),
    .S(net805),
    .X(_1355_));
 sky130_fd_sc_hd__o221ai_1 _4992_ (.A1(\dp.rf.rf[4][9] ),
    .A2(_0395_),
    .B1(_1355_),
    .B2(_0400_),
    .C1(_0186_),
    .Y(_1356_));
 sky130_fd_sc_hd__a31oi_2 _4993_ (.A1(_0389_),
    .A2(_1354_),
    .A3(_1356_),
    .B1(_0293_),
    .Y(_1357_));
 sky130_fd_sc_hd__a221oi_1 _4994_ (.A1(\dp.rf.rf[11][9] ),
    .A2(net812),
    .B1(_0298_),
    .B2(\dp.rf.rf[10][9] ),
    .C1(_0259_),
    .Y(_1358_));
 sky130_fd_sc_hd__mux2_1 _4995_ (.A0(\dp.rf.rf[14][9] ),
    .A1(\dp.rf.rf[15][9] ),
    .S(net812),
    .X(_1359_));
 sky130_fd_sc_hd__o21ai_0 _4996_ (.A1(net800),
    .A2(_1359_),
    .B1(net786),
    .Y(_1360_));
 sky130_fd_sc_hd__mux4_2 _4997_ (.A0(\dp.rf.rf[8][9] ),
    .A1(\dp.rf.rf[9][9] ),
    .A2(\dp.rf.rf[12][9] ),
    .A3(\dp.rf.rf[13][9] ),
    .S0(net812),
    .S1(net805),
    .X(_1361_));
 sky130_fd_sc_hd__a21oi_1 _4998_ (.A1(_0186_),
    .A2(_1361_),
    .B1(net793),
    .Y(_1362_));
 sky130_fd_sc_hd__o21ai_2 _4999_ (.A1(_1358_),
    .A2(_1360_),
    .B1(_1362_),
    .Y(_1363_));
 sky130_fd_sc_hd__a32oi_4 _5000_ (.A1(_0620_),
    .A2(_1346_),
    .A3(_1352_),
    .B1(_1357_),
    .B2(_1363_),
    .Y(_1364_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_110 ();
 sky130_fd_sc_hd__and2_4 _5002_ (.A(net21),
    .B(_0347_),
    .X(_3480_[0]));
 sky130_fd_sc_hd__mux4_2 _5003_ (.A0(\dp.rf.rf[16][8] ),
    .A1(\dp.rf.rf[17][8] ),
    .A2(\dp.rf.rf[18][8] ),
    .A3(\dp.rf.rf[19][8] ),
    .S0(net13),
    .S1(net14),
    .X(_1365_));
 sky130_fd_sc_hd__mux4_2 _5004_ (.A0(\dp.rf.rf[20][8] ),
    .A1(\dp.rf.rf[21][8] ),
    .A2(\dp.rf.rf[22][8] ),
    .A3(\dp.rf.rf[23][8] ),
    .S0(net13),
    .S1(net14),
    .X(_1366_));
 sky130_fd_sc_hd__mux4_2 _5005_ (.A0(\dp.rf.rf[24][8] ),
    .A1(\dp.rf.rf[25][8] ),
    .A2(\dp.rf.rf[26][8] ),
    .A3(\dp.rf.rf[27][8] ),
    .S0(net13),
    .S1(net14),
    .X(_1367_));
 sky130_fd_sc_hd__mux4_2 _5006_ (.A0(\dp.rf.rf[28][8] ),
    .A1(\dp.rf.rf[29][8] ),
    .A2(\dp.rf.rf[30][8] ),
    .A3(\dp.rf.rf[31][8] ),
    .S0(net13),
    .S1(net14),
    .X(_1368_));
 sky130_fd_sc_hd__mux4_2 _5007_ (.A0(_1365_),
    .A1(_1366_),
    .A2(_1367_),
    .A3(_1368_),
    .S0(net818),
    .S1(net16),
    .X(_1369_));
 sky130_fd_sc_hd__mux4_2 _5008_ (.A0(\dp.rf.rf[0][8] ),
    .A1(\dp.rf.rf[1][8] ),
    .A2(\dp.rf.rf[2][8] ),
    .A3(\dp.rf.rf[3][8] ),
    .S0(net825),
    .S1(net819),
    .X(_1370_));
 sky130_fd_sc_hd__mux4_2 _5009_ (.A0(\dp.rf.rf[4][8] ),
    .A1(\dp.rf.rf[5][8] ),
    .A2(\dp.rf.rf[6][8] ),
    .A3(\dp.rf.rf[7][8] ),
    .S0(net825),
    .S1(net819),
    .X(_1371_));
 sky130_fd_sc_hd__mux2i_1 _5010_ (.A0(_1370_),
    .A1(_1371_),
    .S(net818),
    .Y(_1372_));
 sky130_fd_sc_hd__mux4_2 _5011_ (.A0(\dp.rf.rf[8][8] ),
    .A1(\dp.rf.rf[9][8] ),
    .A2(\dp.rf.rf[10][8] ),
    .A3(\dp.rf.rf[11][8] ),
    .S0(net13),
    .S1(net14),
    .X(_1373_));
 sky130_fd_sc_hd__mux4_2 _5012_ (.A0(\dp.rf.rf[12][8] ),
    .A1(\dp.rf.rf[13][8] ),
    .A2(\dp.rf.rf[14][8] ),
    .A3(\dp.rf.rf[15][8] ),
    .S0(net13),
    .S1(net14),
    .X(_1374_));
 sky130_fd_sc_hd__mux2i_1 _5013_ (.A0(_1373_),
    .A1(_1374_),
    .S(net818),
    .Y(_1375_));
 sky130_fd_sc_hd__a221oi_1 _5014_ (.A1(_0109_),
    .A2(_1372_),
    .B1(_1375_),
    .B2(_0861_),
    .C1(_0111_),
    .Y(_1376_));
 sky130_fd_sc_hd__o21ai_4 _5015_ (.A1(_0092_),
    .A2(_1369_),
    .B1(_1376_),
    .Y(_1377_));
 sky130_fd_sc_hd__nor2_1 _5016_ (.A(_0148_),
    .B(_1377_),
    .Y(_1378_));
 sky130_fd_sc_hd__a21oi_2 _5017_ (.A1(_0148_),
    .A2(_3480_[0]),
    .B1(_1378_),
    .Y(_1379_));
 sky130_fd_sc_hd__xor2_1 _5018_ (.A(_0151_),
    .B(_1379_),
    .X(_3387_[0]));
 sky130_fd_sc_hd__inv_1 _5019_ (.A(_3387_[0]),
    .Y(_3391_[0]));
 sky130_fd_sc_hd__mux4_2 _5020_ (.A0(\dp.rf.rf[18][8] ),
    .A1(\dp.rf.rf[19][8] ),
    .A2(\dp.rf.rf[22][8] ),
    .A3(\dp.rf.rf[23][8] ),
    .S0(net812),
    .S1(net805),
    .X(_1380_));
 sky130_fd_sc_hd__nand2_1 _5021_ (.A(net786),
    .B(_1380_),
    .Y(_1381_));
 sky130_fd_sc_hd__inv_1 _5022_ (.A(\dp.rf.rf[20][8] ),
    .Y(_1382_));
 sky130_fd_sc_hd__mux2i_1 _5023_ (.A0(\dp.rf.rf[17][8] ),
    .A1(\dp.rf.rf[21][8] ),
    .S(net805),
    .Y(_1383_));
 sky130_fd_sc_hd__a221oi_1 _5024_ (.A1(_1382_),
    .A2(net801),
    .B1(_1383_),
    .B2(net812),
    .C1(net8),
    .Y(_1384_));
 sky130_fd_sc_hd__o22ai_1 _5025_ (.A1(\dp.rf.rf[16][8] ),
    .A2(net784),
    .B1(_1384_),
    .B2(_0265_),
    .Y(_1385_));
 sky130_fd_sc_hd__nand2_2 _5026_ (.A(_1381_),
    .B(_1385_),
    .Y(_1386_));
 sky130_fd_sc_hd__mux4_2 _5027_ (.A0(\dp.rf.rf[26][8] ),
    .A1(\dp.rf.rf[27][8] ),
    .A2(\dp.rf.rf[30][8] ),
    .A3(\dp.rf.rf[31][8] ),
    .S0(net812),
    .S1(net805),
    .X(_1387_));
 sky130_fd_sc_hd__nand2_1 _5028_ (.A(net8),
    .B(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__mux4_2 _5029_ (.A0(\dp.rf.rf[24][8] ),
    .A1(\dp.rf.rf[25][8] ),
    .A2(\dp.rf.rf[28][8] ),
    .A3(\dp.rf.rf[29][8] ),
    .S0(net812),
    .S1(net804),
    .X(_1389_));
 sky130_fd_sc_hd__nand2_1 _5030_ (.A(_0186_),
    .B(_1389_),
    .Y(_1390_));
 sky130_fd_sc_hd__nand3_2 _5031_ (.A(net10),
    .B(_1388_),
    .C(_1390_),
    .Y(_1391_));
 sky130_fd_sc_hd__mux4_2 _5032_ (.A0(\dp.rf.rf[8][8] ),
    .A1(\dp.rf.rf[9][8] ),
    .A2(\dp.rf.rf[12][8] ),
    .A3(\dp.rf.rf[13][8] ),
    .S0(net7),
    .S1(net804),
    .X(_1392_));
 sky130_fd_sc_hd__nand2_1 _5033_ (.A(_0186_),
    .B(_1392_),
    .Y(_1393_));
 sky130_fd_sc_hd__mux4_2 _5034_ (.A0(\dp.rf.rf[10][8] ),
    .A1(\dp.rf.rf[11][8] ),
    .A2(\dp.rf.rf[14][8] ),
    .A3(\dp.rf.rf[15][8] ),
    .S0(net7),
    .S1(net804),
    .X(_1394_));
 sky130_fd_sc_hd__a21oi_1 _5035_ (.A1(net8),
    .A2(_1394_),
    .B1(net793),
    .Y(_1395_));
 sky130_fd_sc_hd__a21oi_2 _5036_ (.A1(_1393_),
    .A2(_1395_),
    .B1(_0293_),
    .Y(_1396_));
 sky130_fd_sc_hd__mux2_1 _5037_ (.A0(\dp.rf.rf[6][8] ),
    .A1(\dp.rf.rf[7][8] ),
    .S(net812),
    .X(_1397_));
 sky130_fd_sc_hd__o21ai_0 _5038_ (.A1(net800),
    .A2(_1397_),
    .B1(net786),
    .Y(_1398_));
 sky130_fd_sc_hd__a221oi_1 _5039_ (.A1(\dp.rf.rf[3][8] ),
    .A2(net812),
    .B1(_0298_),
    .B2(\dp.rf.rf[2][8] ),
    .C1(_0259_),
    .Y(_1399_));
 sky130_fd_sc_hd__inv_1 _5040_ (.A(\dp.rf.rf[4][8] ),
    .Y(_1400_));
 sky130_fd_sc_hd__mux2i_1 _5041_ (.A0(\dp.rf.rf[1][8] ),
    .A1(\dp.rf.rf[5][8] ),
    .S(net804),
    .Y(_1401_));
 sky130_fd_sc_hd__a221oi_1 _5042_ (.A1(_1400_),
    .A2(_0173_),
    .B1(_1401_),
    .B2(net812),
    .C1(net8),
    .Y(_1402_));
 sky130_fd_sc_hd__o22ai_1 _5043_ (.A1(\dp.rf.rf[0][8] ),
    .A2(net784),
    .B1(_1402_),
    .B2(_0265_),
    .Y(_1403_));
 sky130_fd_sc_hd__o21ai_2 _5044_ (.A1(_1398_),
    .A2(_1399_),
    .B1(_1403_),
    .Y(_1404_));
 sky130_fd_sc_hd__a32oi_4 _5045_ (.A1(net783),
    .A2(_1386_),
    .A3(_1391_),
    .B1(_1396_),
    .B2(_1404_),
    .Y(_1405_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_109 ();
 sky130_fd_sc_hd__mux4_2 _5047_ (.A0(\dp.rf.rf[16][7] ),
    .A1(\dp.rf.rf[17][7] ),
    .A2(\dp.rf.rf[18][7] ),
    .A3(\dp.rf.rf[19][7] ),
    .S0(net822),
    .S1(net14),
    .X(_1406_));
 sky130_fd_sc_hd__mux4_2 _5048_ (.A0(\dp.rf.rf[20][7] ),
    .A1(\dp.rf.rf[21][7] ),
    .A2(\dp.rf.rf[22][7] ),
    .A3(\dp.rf.rf[23][7] ),
    .S0(net822),
    .S1(net14),
    .X(_1407_));
 sky130_fd_sc_hd__mux4_2 _5049_ (.A0(\dp.rf.rf[24][7] ),
    .A1(\dp.rf.rf[25][7] ),
    .A2(\dp.rf.rf[26][7] ),
    .A3(\dp.rf.rf[27][7] ),
    .S0(net822),
    .S1(net14),
    .X(_1408_));
 sky130_fd_sc_hd__mux4_2 _5050_ (.A0(\dp.rf.rf[28][7] ),
    .A1(\dp.rf.rf[29][7] ),
    .A2(\dp.rf.rf[30][7] ),
    .A3(\dp.rf.rf[31][7] ),
    .S0(net822),
    .S1(net14),
    .X(_1409_));
 sky130_fd_sc_hd__mux4_2 _5051_ (.A0(_1406_),
    .A1(_1407_),
    .A2(_1408_),
    .A3(_1409_),
    .S0(net15),
    .S1(net16),
    .X(_1410_));
 sky130_fd_sc_hd__nand2_2 _5052_ (.A(net17),
    .B(_1410_),
    .Y(_1411_));
 sky130_fd_sc_hd__mux4_2 _5053_ (.A0(\dp.rf.rf[0][7] ),
    .A1(\dp.rf.rf[1][7] ),
    .A2(\dp.rf.rf[2][7] ),
    .A3(\dp.rf.rf[3][7] ),
    .S0(net822),
    .S1(net14),
    .X(_1412_));
 sky130_fd_sc_hd__mux4_2 _5054_ (.A0(\dp.rf.rf[4][7] ),
    .A1(\dp.rf.rf[5][7] ),
    .A2(\dp.rf.rf[6][7] ),
    .A3(\dp.rf.rf[7][7] ),
    .S0(net822),
    .S1(net14),
    .X(_1413_));
 sky130_fd_sc_hd__mux4_2 _5055_ (.A0(\dp.rf.rf[8][7] ),
    .A1(\dp.rf.rf[9][7] ),
    .A2(\dp.rf.rf[10][7] ),
    .A3(\dp.rf.rf[11][7] ),
    .S0(net822),
    .S1(net14),
    .X(_1414_));
 sky130_fd_sc_hd__mux4_2 _5056_ (.A0(\dp.rf.rf[12][7] ),
    .A1(\dp.rf.rf[13][7] ),
    .A2(\dp.rf.rf[14][7] ),
    .A3(\dp.rf.rf[15][7] ),
    .S0(net822),
    .S1(net14),
    .X(_1415_));
 sky130_fd_sc_hd__mux4_2 _5057_ (.A0(_1412_),
    .A1(_1413_),
    .A2(_1414_),
    .A3(_1415_),
    .S0(net15),
    .S1(net16),
    .X(_1416_));
 sky130_fd_sc_hd__nand2_2 _5058_ (.A(_0092_),
    .B(_1416_),
    .Y(_1417_));
 sky130_fd_sc_hd__a21oi_4 _5059_ (.A1(_1411_),
    .A2(_1417_),
    .B1(_0111_),
    .Y(net162));
 sky130_fd_sc_hd__and2_4 _5060_ (.A(net20),
    .B(_0347_),
    .X(_3476_[0]));
 sky130_fd_sc_hd__mux2i_1 _5061_ (.A0(net162),
    .A1(_3476_[0]),
    .S(_0148_),
    .Y(_1418_));
 sky130_fd_sc_hd__xor2_2 _5062_ (.A(_0151_),
    .B(_1418_),
    .X(_3395_[0]));
 sky130_fd_sc_hd__inv_1 _5063_ (.A(_3395_[0]),
    .Y(_3399_[0]));
 sky130_fd_sc_hd__mux4_2 _5064_ (.A0(\dp.rf.rf[10][7] ),
    .A1(\dp.rf.rf[11][7] ),
    .A2(\dp.rf.rf[14][7] ),
    .A3(\dp.rf.rf[15][7] ),
    .S0(net7),
    .S1(net9),
    .X(_1419_));
 sky130_fd_sc_hd__nand2_1 _5065_ (.A(net8),
    .B(_1419_),
    .Y(_1420_));
 sky130_fd_sc_hd__mux4_2 _5066_ (.A0(\dp.rf.rf[8][7] ),
    .A1(\dp.rf.rf[9][7] ),
    .A2(\dp.rf.rf[12][7] ),
    .A3(\dp.rf.rf[13][7] ),
    .S0(net7),
    .S1(net9),
    .X(_1421_));
 sky130_fd_sc_hd__nand2_1 _5067_ (.A(_0186_),
    .B(_1421_),
    .Y(_1422_));
 sky130_fd_sc_hd__nand3_2 _5068_ (.A(net797),
    .B(_1420_),
    .C(_1422_),
    .Y(_1423_));
 sky130_fd_sc_hd__mux2_1 _5069_ (.A0(\dp.rf.rf[1][7] ),
    .A1(\dp.rf.rf[5][7] ),
    .S(net9),
    .X(_1424_));
 sky130_fd_sc_hd__o22ai_1 _5070_ (.A1(\dp.rf.rf[4][7] ),
    .A2(_0395_),
    .B1(_1424_),
    .B2(_0400_),
    .Y(_1425_));
 sky130_fd_sc_hd__mux4_2 _5071_ (.A0(\dp.rf.rf[2][7] ),
    .A1(\dp.rf.rf[3][7] ),
    .A2(\dp.rf.rf[6][7] ),
    .A3(\dp.rf.rf[7][7] ),
    .S0(net7),
    .S1(net9),
    .X(_1426_));
 sky130_fd_sc_hd__nand2_1 _5072_ (.A(net8),
    .B(_1426_),
    .Y(_1427_));
 sky130_fd_sc_hd__o211ai_1 _5073_ (.A1(net8),
    .A2(_1425_),
    .B1(_1427_),
    .C1(_0389_),
    .Y(_1428_));
 sky130_fd_sc_hd__mux4_2 _5074_ (.A0(\dp.rf.rf[26][7] ),
    .A1(\dp.rf.rf[27][7] ),
    .A2(\dp.rf.rf[30][7] ),
    .A3(\dp.rf.rf[31][7] ),
    .S0(net809),
    .S1(net9),
    .X(_1429_));
 sky130_fd_sc_hd__nand2_1 _5075_ (.A(net8),
    .B(_1429_),
    .Y(_1430_));
 sky130_fd_sc_hd__mux4_2 _5076_ (.A0(\dp.rf.rf[24][7] ),
    .A1(\dp.rf.rf[25][7] ),
    .A2(\dp.rf.rf[28][7] ),
    .A3(\dp.rf.rf[29][7] ),
    .S0(net809),
    .S1(net9),
    .X(_1431_));
 sky130_fd_sc_hd__nand2_1 _5077_ (.A(_0186_),
    .B(_1431_),
    .Y(_1432_));
 sky130_fd_sc_hd__a31oi_2 _5078_ (.A1(net10),
    .A2(_1430_),
    .A3(_1432_),
    .B1(net794),
    .Y(_1433_));
 sky130_fd_sc_hd__mux2_1 _5079_ (.A0(\dp.rf.rf[22][7] ),
    .A1(\dp.rf.rf[23][7] ),
    .S(net809),
    .X(_1434_));
 sky130_fd_sc_hd__o21ai_0 _5080_ (.A1(_0231_),
    .A2(_1434_),
    .B1(net786),
    .Y(_1435_));
 sky130_fd_sc_hd__a221oi_1 _5081_ (.A1(\dp.rf.rf[19][7] ),
    .A2(net809),
    .B1(net788),
    .B2(\dp.rf.rf[18][7] ),
    .C1(net791),
    .Y(_1436_));
 sky130_fd_sc_hd__inv_1 _5082_ (.A(\dp.rf.rf[20][7] ),
    .Y(_1437_));
 sky130_fd_sc_hd__mux2i_1 _5083_ (.A0(\dp.rf.rf[17][7] ),
    .A1(\dp.rf.rf[21][7] ),
    .S(net9),
    .Y(_1438_));
 sky130_fd_sc_hd__a221oi_1 _5084_ (.A1(_1437_),
    .A2(_0173_),
    .B1(_1438_),
    .B2(net809),
    .C1(net8),
    .Y(_1439_));
 sky130_fd_sc_hd__o22ai_1 _5085_ (.A1(\dp.rf.rf[16][7] ),
    .A2(net784),
    .B1(_1439_),
    .B2(_0265_),
    .Y(_1440_));
 sky130_fd_sc_hd__o21ai_2 _5086_ (.A1(_1435_),
    .A2(_1436_),
    .B1(_1440_),
    .Y(_1441_));
 sky130_fd_sc_hd__a32oi_4 _5087_ (.A1(net780),
    .A2(_1423_),
    .A3(_1428_),
    .B1(_1433_),
    .B2(_1441_),
    .Y(_3398_[0]));
 sky130_fd_sc_hd__mux4_2 _5088_ (.A0(\dp.rf.rf[16][6] ),
    .A1(\dp.rf.rf[17][6] ),
    .A2(\dp.rf.rf[18][6] ),
    .A3(\dp.rf.rf[19][6] ),
    .S0(net823),
    .S1(net821),
    .X(_1442_));
 sky130_fd_sc_hd__mux4_2 _5089_ (.A0(\dp.rf.rf[20][6] ),
    .A1(\dp.rf.rf[21][6] ),
    .A2(\dp.rf.rf[22][6] ),
    .A3(\dp.rf.rf[23][6] ),
    .S0(net823),
    .S1(net821),
    .X(_1443_));
 sky130_fd_sc_hd__mux4_2 _5090_ (.A0(\dp.rf.rf[24][6] ),
    .A1(\dp.rf.rf[25][6] ),
    .A2(\dp.rf.rf[26][6] ),
    .A3(\dp.rf.rf[27][6] ),
    .S0(net823),
    .S1(net821),
    .X(_1444_));
 sky130_fd_sc_hd__mux4_2 _5091_ (.A0(\dp.rf.rf[28][6] ),
    .A1(\dp.rf.rf[29][6] ),
    .A2(\dp.rf.rf[30][6] ),
    .A3(\dp.rf.rf[31][6] ),
    .S0(net823),
    .S1(net821),
    .X(_1445_));
 sky130_fd_sc_hd__mux4_2 _5092_ (.A0(_1442_),
    .A1(_1443_),
    .A2(_1444_),
    .A3(_1445_),
    .S0(net15),
    .S1(net16),
    .X(_1446_));
 sky130_fd_sc_hd__nand2_1 _5093_ (.A(net17),
    .B(_1446_),
    .Y(_1447_));
 sky130_fd_sc_hd__mux4_2 _5094_ (.A0(\dp.rf.rf[0][6] ),
    .A1(\dp.rf.rf[1][6] ),
    .A2(\dp.rf.rf[2][6] ),
    .A3(\dp.rf.rf[3][6] ),
    .S0(net823),
    .S1(net821),
    .X(_1448_));
 sky130_fd_sc_hd__mux4_2 _5095_ (.A0(\dp.rf.rf[4][6] ),
    .A1(\dp.rf.rf[5][6] ),
    .A2(\dp.rf.rf[6][6] ),
    .A3(\dp.rf.rf[7][6] ),
    .S0(net823),
    .S1(net821),
    .X(_1449_));
 sky130_fd_sc_hd__mux4_2 _5096_ (.A0(\dp.rf.rf[8][6] ),
    .A1(\dp.rf.rf[9][6] ),
    .A2(\dp.rf.rf[10][6] ),
    .A3(\dp.rf.rf[11][6] ),
    .S0(net823),
    .S1(net821),
    .X(_1450_));
 sky130_fd_sc_hd__mux4_2 _5097_ (.A0(\dp.rf.rf[12][6] ),
    .A1(\dp.rf.rf[13][6] ),
    .A2(\dp.rf.rf[14][6] ),
    .A3(\dp.rf.rf[15][6] ),
    .S0(net823),
    .S1(net821),
    .X(_1451_));
 sky130_fd_sc_hd__mux4_2 _5098_ (.A0(_1448_),
    .A1(_1449_),
    .A2(_1450_),
    .A3(_1451_),
    .S0(net15),
    .S1(net16),
    .X(_1452_));
 sky130_fd_sc_hd__nand2_2 _5099_ (.A(_0092_),
    .B(_1452_),
    .Y(_1453_));
 sky130_fd_sc_hd__a21oi_4 _5100_ (.A1(_1447_),
    .A2(_1453_),
    .B1(_0111_),
    .Y(net161));
 sky130_fd_sc_hd__and2_4 _5101_ (.A(net19),
    .B(_0347_),
    .X(_3472_[0]));
 sky130_fd_sc_hd__mux2i_1 _5102_ (.A0(net161),
    .A1(_3472_[0]),
    .S(_0148_),
    .Y(_1454_));
 sky130_fd_sc_hd__xor2_1 _5103_ (.A(_0151_),
    .B(_1454_),
    .X(_3403_[0]));
 sky130_fd_sc_hd__inv_1 _5104_ (.A(_3403_[0]),
    .Y(_3407_[0]));
 sky130_fd_sc_hd__mux4_2 _5105_ (.A0(\dp.rf.rf[10][6] ),
    .A1(\dp.rf.rf[11][6] ),
    .A2(\dp.rf.rf[14][6] ),
    .A3(\dp.rf.rf[15][6] ),
    .S0(net7),
    .S1(net9),
    .X(_1455_));
 sky130_fd_sc_hd__nand2_1 _5106_ (.A(net8),
    .B(_1455_),
    .Y(_1456_));
 sky130_fd_sc_hd__mux4_2 _5107_ (.A0(\dp.rf.rf[8][6] ),
    .A1(\dp.rf.rf[9][6] ),
    .A2(\dp.rf.rf[12][6] ),
    .A3(\dp.rf.rf[13][6] ),
    .S0(net7),
    .S1(net9),
    .X(_1457_));
 sky130_fd_sc_hd__nand2_1 _5108_ (.A(_0186_),
    .B(_1457_),
    .Y(_1458_));
 sky130_fd_sc_hd__nand3_2 _5109_ (.A(net797),
    .B(_1456_),
    .C(_1458_),
    .Y(_1459_));
 sky130_fd_sc_hd__mux2_1 _5110_ (.A0(\dp.rf.rf[6][6] ),
    .A1(\dp.rf.rf[7][6] ),
    .S(net7),
    .X(_1460_));
 sky130_fd_sc_hd__o21ai_0 _5111_ (.A1(_0231_),
    .A2(_1460_),
    .B1(_0304_),
    .Y(_1461_));
 sky130_fd_sc_hd__a221oi_1 _5112_ (.A1(\dp.rf.rf[3][6] ),
    .A2(net7),
    .B1(net788),
    .B2(\dp.rf.rf[2][6] ),
    .C1(net791),
    .Y(_1462_));
 sky130_fd_sc_hd__inv_1 _5113_ (.A(\dp.rf.rf[4][6] ),
    .Y(_1463_));
 sky130_fd_sc_hd__mux2i_1 _5114_ (.A0(\dp.rf.rf[1][6] ),
    .A1(\dp.rf.rf[5][6] ),
    .S(net9),
    .Y(_1464_));
 sky130_fd_sc_hd__a221oi_1 _5115_ (.A1(_1463_),
    .A2(_0173_),
    .B1(_1464_),
    .B2(net7),
    .C1(net8),
    .Y(_1465_));
 sky130_fd_sc_hd__o22ai_1 _5116_ (.A1(\dp.rf.rf[0][6] ),
    .A2(net784),
    .B1(_1465_),
    .B2(net790),
    .Y(_1466_));
 sky130_fd_sc_hd__o21ai_2 _5117_ (.A1(_1461_),
    .A2(_1462_),
    .B1(_1466_),
    .Y(_1467_));
 sky130_fd_sc_hd__mux4_2 _5118_ (.A0(\dp.rf.rf[26][6] ),
    .A1(\dp.rf.rf[27][6] ),
    .A2(\dp.rf.rf[30][6] ),
    .A3(\dp.rf.rf[31][6] ),
    .S0(net7),
    .S1(net9),
    .X(_1468_));
 sky130_fd_sc_hd__nand2_1 _5119_ (.A(net8),
    .B(_1468_),
    .Y(_1469_));
 sky130_fd_sc_hd__mux4_2 _5120_ (.A0(\dp.rf.rf[24][6] ),
    .A1(\dp.rf.rf[25][6] ),
    .A2(\dp.rf.rf[28][6] ),
    .A3(\dp.rf.rf[29][6] ),
    .S0(net7),
    .S1(net9),
    .X(_1470_));
 sky130_fd_sc_hd__nand2_1 _5121_ (.A(_0186_),
    .B(_1470_),
    .Y(_1471_));
 sky130_fd_sc_hd__a31oi_2 _5122_ (.A1(net797),
    .A2(_1469_),
    .A3(_1471_),
    .B1(net794),
    .Y(_1472_));
 sky130_fd_sc_hd__mux2_1 _5123_ (.A0(\dp.rf.rf[22][6] ),
    .A1(\dp.rf.rf[23][6] ),
    .S(net7),
    .X(_1473_));
 sky130_fd_sc_hd__o21ai_0 _5124_ (.A1(_0231_),
    .A2(_1473_),
    .B1(_0304_),
    .Y(_1474_));
 sky130_fd_sc_hd__a221oi_1 _5125_ (.A1(\dp.rf.rf[19][6] ),
    .A2(net7),
    .B1(net788),
    .B2(\dp.rf.rf[18][6] ),
    .C1(net791),
    .Y(_1475_));
 sky130_fd_sc_hd__inv_1 _5126_ (.A(\dp.rf.rf[20][6] ),
    .Y(_1476_));
 sky130_fd_sc_hd__mux2i_1 _5127_ (.A0(\dp.rf.rf[17][6] ),
    .A1(\dp.rf.rf[21][6] ),
    .S(net9),
    .Y(_1477_));
 sky130_fd_sc_hd__a221oi_1 _5128_ (.A1(_1476_),
    .A2(_0173_),
    .B1(_1477_),
    .B2(net7),
    .C1(net8),
    .Y(_1478_));
 sky130_fd_sc_hd__o22ai_1 _5129_ (.A1(\dp.rf.rf[16][6] ),
    .A2(net784),
    .B1(_1478_),
    .B2(net790),
    .Y(_1479_));
 sky130_fd_sc_hd__o21ai_1 _5130_ (.A1(_1474_),
    .A2(_1475_),
    .B1(_1479_),
    .Y(_1480_));
 sky130_fd_sc_hd__a32oi_4 _5131_ (.A1(net780),
    .A2(_1459_),
    .A3(_1467_),
    .B1(_1472_),
    .B2(_1480_),
    .Y(_3406_[0]));
 sky130_fd_sc_hd__mux4_2 _5132_ (.A0(\dp.rf.rf[16][5] ),
    .A1(\dp.rf.rf[17][5] ),
    .A2(\dp.rf.rf[18][5] ),
    .A3(\dp.rf.rf[19][5] ),
    .S0(net824),
    .S1(net821),
    .X(_1481_));
 sky130_fd_sc_hd__mux4_2 _5133_ (.A0(\dp.rf.rf[20][5] ),
    .A1(\dp.rf.rf[21][5] ),
    .A2(\dp.rf.rf[22][5] ),
    .A3(\dp.rf.rf[23][5] ),
    .S0(net824),
    .S1(net821),
    .X(_1482_));
 sky130_fd_sc_hd__mux4_2 _5134_ (.A0(\dp.rf.rf[24][5] ),
    .A1(\dp.rf.rf[25][5] ),
    .A2(\dp.rf.rf[26][5] ),
    .A3(\dp.rf.rf[27][5] ),
    .S0(net824),
    .S1(net821),
    .X(_1483_));
 sky130_fd_sc_hd__mux4_2 _5135_ (.A0(\dp.rf.rf[28][5] ),
    .A1(\dp.rf.rf[29][5] ),
    .A2(\dp.rf.rf[30][5] ),
    .A3(\dp.rf.rf[31][5] ),
    .S0(net824),
    .S1(net821),
    .X(_1484_));
 sky130_fd_sc_hd__mux4_2 _5136_ (.A0(_1481_),
    .A1(_1482_),
    .A2(_1483_),
    .A3(_1484_),
    .S0(net15),
    .S1(net16),
    .X(_1485_));
 sky130_fd_sc_hd__nand2_2 _5137_ (.A(net17),
    .B(_1485_),
    .Y(_1486_));
 sky130_fd_sc_hd__mux4_2 _5138_ (.A0(\dp.rf.rf[0][5] ),
    .A1(\dp.rf.rf[1][5] ),
    .A2(\dp.rf.rf[2][5] ),
    .A3(\dp.rf.rf[3][5] ),
    .S0(net824),
    .S1(net821),
    .X(_1487_));
 sky130_fd_sc_hd__mux4_2 _5139_ (.A0(\dp.rf.rf[4][5] ),
    .A1(\dp.rf.rf[5][5] ),
    .A2(\dp.rf.rf[6][5] ),
    .A3(\dp.rf.rf[7][5] ),
    .S0(net824),
    .S1(net821),
    .X(_1488_));
 sky130_fd_sc_hd__mux4_2 _5140_ (.A0(\dp.rf.rf[8][5] ),
    .A1(\dp.rf.rf[9][5] ),
    .A2(\dp.rf.rf[10][5] ),
    .A3(\dp.rf.rf[11][5] ),
    .S0(net824),
    .S1(net821),
    .X(_1489_));
 sky130_fd_sc_hd__mux4_2 _5141_ (.A0(\dp.rf.rf[12][5] ),
    .A1(\dp.rf.rf[13][5] ),
    .A2(\dp.rf.rf[14][5] ),
    .A3(\dp.rf.rf[15][5] ),
    .S0(net824),
    .S1(net821),
    .X(_1490_));
 sky130_fd_sc_hd__mux4_2 _5142_ (.A0(_1487_),
    .A1(_1488_),
    .A2(_1489_),
    .A3(_1490_),
    .S0(net15),
    .S1(net16),
    .X(_1491_));
 sky130_fd_sc_hd__nand2_2 _5143_ (.A(_0092_),
    .B(_1491_),
    .Y(_1492_));
 sky130_fd_sc_hd__a21oi_4 _5144_ (.A1(_1486_),
    .A2(_1492_),
    .B1(_0111_),
    .Y(net160));
 sky130_fd_sc_hd__and2_4 _5145_ (.A(net18),
    .B(_0347_),
    .X(_3468_[0]));
 sky130_fd_sc_hd__mux2i_1 _5146_ (.A0(net160),
    .A1(_3468_[0]),
    .S(_0148_),
    .Y(_1493_));
 sky130_fd_sc_hd__xor2_1 _5147_ (.A(_0151_),
    .B(_1493_),
    .X(_3411_[0]));
 sky130_fd_sc_hd__inv_1 _5148_ (.A(_3411_[0]),
    .Y(_3415_[0]));
 sky130_fd_sc_hd__mux4_2 _5149_ (.A0(\dp.rf.rf[2][5] ),
    .A1(\dp.rf.rf[3][5] ),
    .A2(\dp.rf.rf[6][5] ),
    .A3(\dp.rf.rf[7][5] ),
    .S0(net7),
    .S1(net9),
    .X(_1494_));
 sky130_fd_sc_hd__nand2_1 _5150_ (.A(net8),
    .B(_1494_),
    .Y(_1495_));
 sky130_fd_sc_hd__mux2_1 _5151_ (.A0(\dp.rf.rf[1][5] ),
    .A1(\dp.rf.rf[5][5] ),
    .S(net9),
    .X(_1496_));
 sky130_fd_sc_hd__o221ai_1 _5152_ (.A1(\dp.rf.rf[4][5] ),
    .A2(_0395_),
    .B1(_1496_),
    .B2(_0400_),
    .C1(_0186_),
    .Y(_1497_));
 sky130_fd_sc_hd__nand3_2 _5153_ (.A(_0389_),
    .B(_1495_),
    .C(_1497_),
    .Y(_1498_));
 sky130_fd_sc_hd__a221oi_1 _5154_ (.A1(\dp.rf.rf[11][5] ),
    .A2(net7),
    .B1(net788),
    .B2(\dp.rf.rf[10][5] ),
    .C1(net791),
    .Y(_1499_));
 sky130_fd_sc_hd__mux2_1 _5155_ (.A0(\dp.rf.rf[14][5] ),
    .A1(\dp.rf.rf[15][5] ),
    .S(net7),
    .X(_1500_));
 sky130_fd_sc_hd__o21ai_0 _5156_ (.A1(_0231_),
    .A2(_1500_),
    .B1(_0347_),
    .Y(_1501_));
 sky130_fd_sc_hd__mux4_2 _5157_ (.A0(\dp.rf.rf[8][5] ),
    .A1(\dp.rf.rf[9][5] ),
    .A2(\dp.rf.rf[12][5] ),
    .A3(\dp.rf.rf[13][5] ),
    .S0(net7),
    .S1(net9),
    .X(_1502_));
 sky130_fd_sc_hd__nand2_1 _5158_ (.A(_0186_),
    .B(_1502_),
    .Y(_1503_));
 sky130_fd_sc_hd__o311ai_2 _5159_ (.A1(_0186_),
    .A2(_1499_),
    .A3(_1501_),
    .B1(_1503_),
    .C1(net797),
    .Y(_1504_));
 sky130_fd_sc_hd__mux4_2 _5160_ (.A0(\dp.rf.rf[26][5] ),
    .A1(\dp.rf.rf[27][5] ),
    .A2(\dp.rf.rf[30][5] ),
    .A3(\dp.rf.rf[31][5] ),
    .S0(net7),
    .S1(net9),
    .X(_1505_));
 sky130_fd_sc_hd__mux4_2 _5161_ (.A0(\dp.rf.rf[24][5] ),
    .A1(\dp.rf.rf[25][5] ),
    .A2(\dp.rf.rf[28][5] ),
    .A3(\dp.rf.rf[29][5] ),
    .S0(net7),
    .S1(net9),
    .X(_1506_));
 sky130_fd_sc_hd__a221oi_1 _5162_ (.A1(_0304_),
    .A2(_1505_),
    .B1(_1506_),
    .B2(_0186_),
    .C1(_0255_),
    .Y(_1507_));
 sky130_fd_sc_hd__nor2_2 _5163_ (.A(net794),
    .B(_1507_),
    .Y(_1508_));
 sky130_fd_sc_hd__mux2_1 _5164_ (.A0(\dp.rf.rf[22][5] ),
    .A1(\dp.rf.rf[23][5] ),
    .S(net7),
    .X(_1509_));
 sky130_fd_sc_hd__o21ai_0 _5165_ (.A1(_0231_),
    .A2(_1509_),
    .B1(_0304_),
    .Y(_1510_));
 sky130_fd_sc_hd__a221oi_1 _5166_ (.A1(\dp.rf.rf[19][5] ),
    .A2(net7),
    .B1(net788),
    .B2(\dp.rf.rf[18][5] ),
    .C1(net791),
    .Y(_1511_));
 sky130_fd_sc_hd__inv_1 _5167_ (.A(\dp.rf.rf[20][5] ),
    .Y(_1512_));
 sky130_fd_sc_hd__mux2i_1 _5168_ (.A0(\dp.rf.rf[17][5] ),
    .A1(\dp.rf.rf[21][5] ),
    .S(net9),
    .Y(_1513_));
 sky130_fd_sc_hd__a221oi_1 _5169_ (.A1(_1512_),
    .A2(_0173_),
    .B1(_1513_),
    .B2(net7),
    .C1(net8),
    .Y(_1514_));
 sky130_fd_sc_hd__o22ai_1 _5170_ (.A1(\dp.rf.rf[16][5] ),
    .A2(net784),
    .B1(_1514_),
    .B2(net790),
    .Y(_1515_));
 sky130_fd_sc_hd__o21ai_2 _5171_ (.A1(_1510_),
    .A2(_1511_),
    .B1(_1515_),
    .Y(_1516_));
 sky130_fd_sc_hd__a32oi_4 _5172_ (.A1(net780),
    .A2(_1498_),
    .A3(_1504_),
    .B1(_1508_),
    .B2(_1516_),
    .Y(_3414_[0]));
 sky130_fd_sc_hd__a22oi_2 _5173_ (.A1(_0036_),
    .A2(net803),
    .B1(_0143_),
    .B2(net802),
    .Y(_1517_));
 sky130_fd_sc_hd__a22o_4 _5174_ (.A1(net3),
    .A2(_0042_),
    .B1(_1517_),
    .B2(net17),
    .X(_3464_[0]));
 sky130_fd_sc_hd__mux4_2 _5175_ (.A0(\dp.rf.rf[16][4] ),
    .A1(\dp.rf.rf[17][4] ),
    .A2(\dp.rf.rf[18][4] ),
    .A3(\dp.rf.rf[19][4] ),
    .S0(net822),
    .S1(net14),
    .X(_1518_));
 sky130_fd_sc_hd__mux4_2 _5176_ (.A0(\dp.rf.rf[20][4] ),
    .A1(\dp.rf.rf[21][4] ),
    .A2(\dp.rf.rf[22][4] ),
    .A3(\dp.rf.rf[23][4] ),
    .S0(net822),
    .S1(net14),
    .X(_1519_));
 sky130_fd_sc_hd__mux4_2 _5177_ (.A0(\dp.rf.rf[24][4] ),
    .A1(\dp.rf.rf[25][4] ),
    .A2(\dp.rf.rf[26][4] ),
    .A3(\dp.rf.rf[27][4] ),
    .S0(net822),
    .S1(net14),
    .X(_1520_));
 sky130_fd_sc_hd__mux4_2 _5178_ (.A0(\dp.rf.rf[28][4] ),
    .A1(\dp.rf.rf[29][4] ),
    .A2(\dp.rf.rf[30][4] ),
    .A3(\dp.rf.rf[31][4] ),
    .S0(net822),
    .S1(net14),
    .X(_1521_));
 sky130_fd_sc_hd__mux4_2 _5179_ (.A0(_1518_),
    .A1(_1519_),
    .A2(_1520_),
    .A3(_1521_),
    .S0(net15),
    .S1(net16),
    .X(_1522_));
 sky130_fd_sc_hd__nand2_1 _5180_ (.A(net17),
    .B(_1522_),
    .Y(_1523_));
 sky130_fd_sc_hd__mux4_2 _5181_ (.A0(\dp.rf.rf[0][4] ),
    .A1(\dp.rf.rf[1][4] ),
    .A2(\dp.rf.rf[2][4] ),
    .A3(\dp.rf.rf[3][4] ),
    .S0(net823),
    .S1(net821),
    .X(_1524_));
 sky130_fd_sc_hd__mux4_2 _5182_ (.A0(\dp.rf.rf[4][4] ),
    .A1(\dp.rf.rf[5][4] ),
    .A2(\dp.rf.rf[6][4] ),
    .A3(\dp.rf.rf[7][4] ),
    .S0(net823),
    .S1(net14),
    .X(_1525_));
 sky130_fd_sc_hd__mux4_2 _5183_ (.A0(\dp.rf.rf[8][4] ),
    .A1(\dp.rf.rf[9][4] ),
    .A2(\dp.rf.rf[10][4] ),
    .A3(\dp.rf.rf[11][4] ),
    .S0(net823),
    .S1(net14),
    .X(_1526_));
 sky130_fd_sc_hd__mux4_2 _5184_ (.A0(\dp.rf.rf[12][4] ),
    .A1(\dp.rf.rf[13][4] ),
    .A2(\dp.rf.rf[14][4] ),
    .A3(\dp.rf.rf[15][4] ),
    .S0(net823),
    .S1(net14),
    .X(_1527_));
 sky130_fd_sc_hd__mux4_2 _5185_ (.A0(_1524_),
    .A1(_1525_),
    .A2(_1526_),
    .A3(_1527_),
    .S0(net15),
    .S1(net16),
    .X(_1528_));
 sky130_fd_sc_hd__nand2_2 _5186_ (.A(_0092_),
    .B(_1528_),
    .Y(_1529_));
 sky130_fd_sc_hd__a21oi_4 _5187_ (.A1(_1523_),
    .A2(_1529_),
    .B1(_0111_),
    .Y(net159));
 sky130_fd_sc_hd__nand2_4 _5188_ (.A(_0148_),
    .B(_3464_[0]),
    .Y(_1530_));
 sky130_fd_sc_hd__nand2_2 _5189_ (.A(_0121_),
    .B(net159),
    .Y(_1531_));
 sky130_fd_sc_hd__nand2_8 _5190_ (.A(_1531_),
    .B(_1530_),
    .Y(_1532_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_106 ();
 sky130_fd_sc_hd__xnor2_4 _5194_ (.A(_0151_),
    .B(_1532_),
    .Y(_3419_[0]));
 sky130_fd_sc_hd__inv_1 _5195_ (.A(_3419_[0]),
    .Y(_3423_[0]));
 sky130_fd_sc_hd__mux4_2 _5196_ (.A0(\dp.rf.rf[10][4] ),
    .A1(\dp.rf.rf[11][4] ),
    .A2(\dp.rf.rf[14][4] ),
    .A3(\dp.rf.rf[15][4] ),
    .S0(net809),
    .S1(net9),
    .X(_1536_));
 sky130_fd_sc_hd__nand2_1 _5197_ (.A(net8),
    .B(_1536_),
    .Y(_1537_));
 sky130_fd_sc_hd__mux4_2 _5198_ (.A0(\dp.rf.rf[8][4] ),
    .A1(\dp.rf.rf[9][4] ),
    .A2(\dp.rf.rf[12][4] ),
    .A3(\dp.rf.rf[13][4] ),
    .S0(net809),
    .S1(net9),
    .X(_1538_));
 sky130_fd_sc_hd__nand2_1 _5199_ (.A(_0186_),
    .B(_1538_),
    .Y(_1539_));
 sky130_fd_sc_hd__nand3_2 _5200_ (.A(net797),
    .B(_1537_),
    .C(_1539_),
    .Y(_1540_));
 sky130_fd_sc_hd__mux2_1 _5201_ (.A0(\dp.rf.rf[6][4] ),
    .A1(\dp.rf.rf[7][4] ),
    .S(net7),
    .X(_1541_));
 sky130_fd_sc_hd__o21ai_0 _5202_ (.A1(_0231_),
    .A2(_1541_),
    .B1(_0304_),
    .Y(_1542_));
 sky130_fd_sc_hd__a221oi_1 _5203_ (.A1(\dp.rf.rf[3][4] ),
    .A2(net7),
    .B1(net788),
    .B2(\dp.rf.rf[2][4] ),
    .C1(net791),
    .Y(_1543_));
 sky130_fd_sc_hd__inv_1 _5204_ (.A(\dp.rf.rf[4][4] ),
    .Y(_1544_));
 sky130_fd_sc_hd__mux2i_1 _5205_ (.A0(\dp.rf.rf[1][4] ),
    .A1(\dp.rf.rf[5][4] ),
    .S(net9),
    .Y(_1545_));
 sky130_fd_sc_hd__a221oi_1 _5206_ (.A1(_1544_),
    .A2(_0173_),
    .B1(_1545_),
    .B2(net7),
    .C1(net8),
    .Y(_1546_));
 sky130_fd_sc_hd__o22ai_1 _5207_ (.A1(\dp.rf.rf[0][4] ),
    .A2(net784),
    .B1(_1546_),
    .B2(net790),
    .Y(_1547_));
 sky130_fd_sc_hd__o21ai_2 _5208_ (.A1(_1542_),
    .A2(_1543_),
    .B1(_1547_),
    .Y(_1548_));
 sky130_fd_sc_hd__mux4_2 _5209_ (.A0(\dp.rf.rf[26][4] ),
    .A1(\dp.rf.rf[27][4] ),
    .A2(\dp.rf.rf[30][4] ),
    .A3(\dp.rf.rf[31][4] ),
    .S0(net809),
    .S1(net9),
    .X(_1549_));
 sky130_fd_sc_hd__nand2_1 _5210_ (.A(net8),
    .B(_1549_),
    .Y(_1550_));
 sky130_fd_sc_hd__mux4_2 _5211_ (.A0(\dp.rf.rf[24][4] ),
    .A1(\dp.rf.rf[25][4] ),
    .A2(\dp.rf.rf[28][4] ),
    .A3(\dp.rf.rf[29][4] ),
    .S0(net809),
    .S1(net9),
    .X(_1551_));
 sky130_fd_sc_hd__nand2_1 _5212_ (.A(_0186_),
    .B(_1551_),
    .Y(_1552_));
 sky130_fd_sc_hd__a31oi_2 _5213_ (.A1(net10),
    .A2(_1550_),
    .A3(_1552_),
    .B1(net794),
    .Y(_1553_));
 sky130_fd_sc_hd__mux2_1 _5214_ (.A0(\dp.rf.rf[22][4] ),
    .A1(\dp.rf.rf[23][4] ),
    .S(net7),
    .X(_1554_));
 sky130_fd_sc_hd__o21ai_0 _5215_ (.A1(_0231_),
    .A2(_1554_),
    .B1(_0304_),
    .Y(_1555_));
 sky130_fd_sc_hd__a221oi_1 _5216_ (.A1(\dp.rf.rf[19][4] ),
    .A2(net7),
    .B1(net788),
    .B2(\dp.rf.rf[18][4] ),
    .C1(net791),
    .Y(_1556_));
 sky130_fd_sc_hd__inv_1 _5217_ (.A(\dp.rf.rf[20][4] ),
    .Y(_1557_));
 sky130_fd_sc_hd__mux2i_1 _5218_ (.A0(\dp.rf.rf[17][4] ),
    .A1(\dp.rf.rf[21][4] ),
    .S(net9),
    .Y(_1558_));
 sky130_fd_sc_hd__a221oi_1 _5219_ (.A1(_1557_),
    .A2(_0173_),
    .B1(_1558_),
    .B2(net7),
    .C1(net8),
    .Y(_1559_));
 sky130_fd_sc_hd__o22ai_1 _5220_ (.A1(\dp.rf.rf[16][4] ),
    .A2(net784),
    .B1(_1559_),
    .B2(net790),
    .Y(_1560_));
 sky130_fd_sc_hd__o21ai_2 _5221_ (.A1(_1555_),
    .A2(_1556_),
    .B1(_1560_),
    .Y(_1561_));
 sky130_fd_sc_hd__a32oi_4 _5222_ (.A1(net780),
    .A2(_1540_),
    .A3(_1548_),
    .B1(_1553_),
    .B2(_1561_),
    .Y(_3422_[0]));
 sky130_fd_sc_hd__a22o_4 _5223_ (.A1(net2),
    .A2(_0042_),
    .B1(_1517_),
    .B2(net16),
    .X(_3458_[0]));
 sky130_fd_sc_hd__mux4_2 _5224_ (.A0(\dp.rf.rf[16][3] ),
    .A1(\dp.rf.rf[17][3] ),
    .A2(\dp.rf.rf[18][3] ),
    .A3(\dp.rf.rf[19][3] ),
    .S0(net822),
    .S1(net14),
    .X(_1562_));
 sky130_fd_sc_hd__mux4_2 _5225_ (.A0(\dp.rf.rf[20][3] ),
    .A1(\dp.rf.rf[21][3] ),
    .A2(\dp.rf.rf[22][3] ),
    .A3(\dp.rf.rf[23][3] ),
    .S0(net822),
    .S1(net14),
    .X(_1563_));
 sky130_fd_sc_hd__mux4_2 _5226_ (.A0(\dp.rf.rf[24][3] ),
    .A1(\dp.rf.rf[25][3] ),
    .A2(\dp.rf.rf[26][3] ),
    .A3(\dp.rf.rf[27][3] ),
    .S0(net822),
    .S1(net14),
    .X(_1564_));
 sky130_fd_sc_hd__mux4_2 _5227_ (.A0(\dp.rf.rf[28][3] ),
    .A1(\dp.rf.rf[29][3] ),
    .A2(\dp.rf.rf[30][3] ),
    .A3(\dp.rf.rf[31][3] ),
    .S0(net822),
    .S1(net14),
    .X(_1565_));
 sky130_fd_sc_hd__mux4_2 _5228_ (.A0(_1562_),
    .A1(_1563_),
    .A2(_1564_),
    .A3(_1565_),
    .S0(net818),
    .S1(net16),
    .X(_1566_));
 sky130_fd_sc_hd__mux4_2 _5229_ (.A0(\dp.rf.rf[0][3] ),
    .A1(\dp.rf.rf[1][3] ),
    .A2(\dp.rf.rf[2][3] ),
    .A3(\dp.rf.rf[3][3] ),
    .S0(net822),
    .S1(net14),
    .X(_1567_));
 sky130_fd_sc_hd__mux4_2 _5230_ (.A0(\dp.rf.rf[4][3] ),
    .A1(\dp.rf.rf[5][3] ),
    .A2(\dp.rf.rf[6][3] ),
    .A3(\dp.rf.rf[7][3] ),
    .S0(net822),
    .S1(net14),
    .X(_1568_));
 sky130_fd_sc_hd__mux4_2 _5231_ (.A0(\dp.rf.rf[8][3] ),
    .A1(\dp.rf.rf[9][3] ),
    .A2(\dp.rf.rf[10][3] ),
    .A3(\dp.rf.rf[11][3] ),
    .S0(net822),
    .S1(net14),
    .X(_1569_));
 sky130_fd_sc_hd__mux4_2 _5232_ (.A0(\dp.rf.rf[12][3] ),
    .A1(\dp.rf.rf[13][3] ),
    .A2(\dp.rf.rf[14][3] ),
    .A3(\dp.rf.rf[15][3] ),
    .S0(net822),
    .S1(net14),
    .X(_1570_));
 sky130_fd_sc_hd__mux4_2 _5233_ (.A0(_1567_),
    .A1(_1568_),
    .A2(_1569_),
    .A3(_1570_),
    .S0(net818),
    .S1(net16),
    .X(_1571_));
 sky130_fd_sc_hd__a22oi_2 _5234_ (.A1(net17),
    .A2(_1566_),
    .B1(_1571_),
    .B2(_0337_),
    .Y(_1572_));
 sky130_fd_sc_hd__clkinvlp_4 _5235_ (.A(net209),
    .Y(net158));
 sky130_fd_sc_hd__nand2_4 _5236_ (.A(_0121_),
    .B(net218),
    .Y(_1573_));
 sky130_fd_sc_hd__o21a_4 _5237_ (.A1(_0121_),
    .A2(_3458_[0]),
    .B1(_1573_),
    .X(_1574_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_104 ();
 sky130_fd_sc_hd__xnor2_4 _5240_ (.A(_0151_),
    .B(_1574_),
    .Y(_3427_[0]));
 sky130_fd_sc_hd__inv_1 _5241_ (.A(_3427_[0]),
    .Y(_3431_[0]));
 sky130_fd_sc_hd__mux2_1 _5242_ (.A0(\dp.rf.rf[14][3] ),
    .A1(\dp.rf.rf[15][3] ),
    .S(net7),
    .X(_1577_));
 sky130_fd_sc_hd__o21ai_0 _5243_ (.A1(_0231_),
    .A2(_1577_),
    .B1(net786),
    .Y(_1578_));
 sky130_fd_sc_hd__a221oi_1 _5244_ (.A1(\dp.rf.rf[11][3] ),
    .A2(net7),
    .B1(net788),
    .B2(\dp.rf.rf[10][3] ),
    .C1(net791),
    .Y(_1579_));
 sky130_fd_sc_hd__inv_1 _5245_ (.A(\dp.rf.rf[12][3] ),
    .Y(_1580_));
 sky130_fd_sc_hd__mux2i_1 _5246_ (.A0(\dp.rf.rf[9][3] ),
    .A1(\dp.rf.rf[13][3] ),
    .S(net9),
    .Y(_1581_));
 sky130_fd_sc_hd__a221oi_1 _5247_ (.A1(_1580_),
    .A2(net801),
    .B1(_1581_),
    .B2(net7),
    .C1(net8),
    .Y(_1582_));
 sky130_fd_sc_hd__a22oi_2 _5248_ (.A1(_0143_),
    .A2(net802),
    .B1(_0165_),
    .B2(_0468_),
    .Y(_1583_));
 sky130_fd_sc_hd__o32ai_1 _5249_ (.A1(net11),
    .A2(_0137_),
    .A3(_1582_),
    .B1(_1583_),
    .B2(\dp.rf.rf[8][3] ),
    .Y(_1584_));
 sky130_fd_sc_hd__o21ai_2 _5250_ (.A1(_1578_),
    .A2(_1579_),
    .B1(_1584_),
    .Y(_1585_));
 sky130_fd_sc_hd__a221oi_1 _5251_ (.A1(\dp.rf.rf[27][3] ),
    .A2(net810),
    .B1(net788),
    .B2(\dp.rf.rf[26][3] ),
    .C1(net791),
    .Y(_1586_));
 sky130_fd_sc_hd__mux2_1 _5252_ (.A0(\dp.rf.rf[30][3] ),
    .A1(\dp.rf.rf[31][3] ),
    .S(net810),
    .X(_1587_));
 sky130_fd_sc_hd__o21ai_0 _5253_ (.A1(_0231_),
    .A2(_1587_),
    .B1(net8),
    .Y(_1588_));
 sky130_fd_sc_hd__mux4_2 _5254_ (.A0(\dp.rf.rf[24][3] ),
    .A1(\dp.rf.rf[25][3] ),
    .A2(\dp.rf.rf[28][3] ),
    .A3(\dp.rf.rf[29][3] ),
    .S0(net810),
    .S1(net804),
    .X(_1589_));
 sky130_fd_sc_hd__a21oi_1 _5255_ (.A1(_0186_),
    .A2(_1589_),
    .B1(net794),
    .Y(_1590_));
 sky130_fd_sc_hd__o21ai_2 _5256_ (.A1(_1586_),
    .A2(_1588_),
    .B1(_1590_),
    .Y(_1591_));
 sky130_fd_sc_hd__nand3_4 _5257_ (.A(net797),
    .B(_1585_),
    .C(_1591_),
    .Y(_1592_));
 sky130_fd_sc_hd__a221oi_1 _5258_ (.A1(\dp.rf.rf[19][3] ),
    .A2(net7),
    .B1(net788),
    .B2(\dp.rf.rf[18][3] ),
    .C1(net791),
    .Y(_1593_));
 sky130_fd_sc_hd__mux2i_1 _5259_ (.A0(\dp.rf.rf[22][3] ),
    .A1(\dp.rf.rf[23][3] ),
    .S(net7),
    .Y(_1594_));
 sky130_fd_sc_hd__nand2_1 _5260_ (.A(net9),
    .B(_1594_),
    .Y(_1595_));
 sky130_fd_sc_hd__nand3_1 _5261_ (.A(net8),
    .B(_0347_),
    .C(_1595_),
    .Y(_1596_));
 sky130_fd_sc_hd__mux4_2 _5262_ (.A0(\dp.rf.rf[16][3] ),
    .A1(\dp.rf.rf[17][3] ),
    .A2(\dp.rf.rf[20][3] ),
    .A3(\dp.rf.rf[21][3] ),
    .S0(net7),
    .S1(net9),
    .X(_1597_));
 sky130_fd_sc_hd__nand2_1 _5263_ (.A(_0186_),
    .B(_1597_),
    .Y(_1598_));
 sky130_fd_sc_hd__o21ai_2 _5264_ (.A1(_1593_),
    .A2(_1596_),
    .B1(_1598_),
    .Y(_1599_));
 sky130_fd_sc_hd__nand3_2 _5265_ (.A(_0231_),
    .B(_0468_),
    .C(_0207_),
    .Y(_1600_));
 sky130_fd_sc_hd__mux2_1 _5266_ (.A0(\dp.rf.rf[6][3] ),
    .A1(\dp.rf.rf[7][3] ),
    .S(net7),
    .X(_1601_));
 sky130_fd_sc_hd__o21ai_0 _5267_ (.A1(_0231_),
    .A2(_1601_),
    .B1(net786),
    .Y(_1602_));
 sky130_fd_sc_hd__a221oi_1 _5268_ (.A1(\dp.rf.rf[3][3] ),
    .A2(net7),
    .B1(_0298_),
    .B2(\dp.rf.rf[2][3] ),
    .C1(net791),
    .Y(_1603_));
 sky130_fd_sc_hd__inv_1 _5269_ (.A(\dp.rf.rf[4][3] ),
    .Y(_1604_));
 sky130_fd_sc_hd__mux2i_1 _5270_ (.A0(\dp.rf.rf[1][3] ),
    .A1(\dp.rf.rf[5][3] ),
    .S(net9),
    .Y(_1605_));
 sky130_fd_sc_hd__a221oi_1 _5271_ (.A1(_1604_),
    .A2(net801),
    .B1(_1605_),
    .B2(net7),
    .C1(net8),
    .Y(_1606_));
 sky130_fd_sc_hd__o32ai_1 _5272_ (.A1(net11),
    .A2(_0137_),
    .A3(_1606_),
    .B1(_1583_),
    .B2(\dp.rf.rf[0][3] ),
    .Y(_1607_));
 sky130_fd_sc_hd__o21ai_2 _5273_ (.A1(_1602_),
    .A2(_1603_),
    .B1(_1607_),
    .Y(_1608_));
 sky130_fd_sc_hd__o2111ai_4 _5274_ (.A1(net794),
    .A2(_1599_),
    .B1(_1600_),
    .C1(_1608_),
    .D1(_0389_),
    .Y(_1609_));
 sky130_fd_sc_hd__nand2_8 _5275_ (.A(_1592_),
    .B(_1609_),
    .Y(_3426_[0]));
 sky130_fd_sc_hd__clkinvlp_4 _5276_ (.A(_3426_[0]),
    .Y(_3430_[0]));
 sky130_fd_sc_hd__a22o_4 _5277_ (.A1(net32),
    .A2(_0042_),
    .B1(_1517_),
    .B2(net818),
    .X(_3454_[0]));
 sky130_fd_sc_hd__nand2_2 _5278_ (.A(net17),
    .B(net15),
    .Y(_1610_));
 sky130_fd_sc_hd__mux4_2 _5279_ (.A0(\dp.rf.rf[20][2] ),
    .A1(\dp.rf.rf[21][2] ),
    .A2(\dp.rf.rf[22][2] ),
    .A3(\dp.rf.rf[23][2] ),
    .S0(net824),
    .S1(net821),
    .X(_1611_));
 sky130_fd_sc_hd__mux4_2 _5280_ (.A0(\dp.rf.rf[28][2] ),
    .A1(\dp.rf.rf[29][2] ),
    .A2(\dp.rf.rf[30][2] ),
    .A3(\dp.rf.rf[31][2] ),
    .S0(net823),
    .S1(net821),
    .X(_1612_));
 sky130_fd_sc_hd__mux2i_4 _5281_ (.A0(_1611_),
    .A1(_1612_),
    .S(net16),
    .Y(_1613_));
 sky130_fd_sc_hd__mux2i_1 _5282_ (.A0(\dp.rf.rf[1][2] ),
    .A1(\dp.rf.rf[9][2] ),
    .S(net16),
    .Y(_1614_));
 sky130_fd_sc_hd__a21oi_1 _5283_ (.A1(net16),
    .A2(\dp.rf.rf[8][2] ),
    .B1(net824),
    .Y(_1615_));
 sky130_fd_sc_hd__a21oi_1 _5284_ (.A1(net824),
    .A2(_1614_),
    .B1(_1615_),
    .Y(_1616_));
 sky130_fd_sc_hd__mux4_2 _5285_ (.A0(\dp.rf.rf[4][2] ),
    .A1(\dp.rf.rf[5][2] ),
    .A2(\dp.rf.rf[12][2] ),
    .A3(\dp.rf.rf[13][2] ),
    .S0(net824),
    .S1(net16),
    .X(_1617_));
 sky130_fd_sc_hd__mux4_2 _5286_ (.A0(\dp.rf.rf[2][2] ),
    .A1(\dp.rf.rf[3][2] ),
    .A2(\dp.rf.rf[10][2] ),
    .A3(\dp.rf.rf[11][2] ),
    .S0(net824),
    .S1(net16),
    .X(_1618_));
 sky130_fd_sc_hd__mux4_2 _5287_ (.A0(\dp.rf.rf[6][2] ),
    .A1(\dp.rf.rf[7][2] ),
    .A2(\dp.rf.rf[14][2] ),
    .A3(\dp.rf.rf[15][2] ),
    .S0(net824),
    .S1(net16),
    .X(_1619_));
 sky130_fd_sc_hd__mux4_2 _5288_ (.A0(_1616_),
    .A1(_1617_),
    .A2(_1618_),
    .A3(_1619_),
    .S0(net15),
    .S1(net821),
    .X(_1620_));
 sky130_fd_sc_hd__nand2_2 _5289_ (.A(_1620_),
    .B(_0092_),
    .Y(_1621_));
 sky130_fd_sc_hd__mux4_2 _5290_ (.A0(\dp.rf.rf[16][2] ),
    .A1(\dp.rf.rf[17][2] ),
    .A2(\dp.rf.rf[24][2] ),
    .A3(\dp.rf.rf[25][2] ),
    .S0(net824),
    .S1(net16),
    .X(_1622_));
 sky130_fd_sc_hd__mux2i_1 _5291_ (.A0(\dp.rf.rf[18][2] ),
    .A1(\dp.rf.rf[19][2] ),
    .S(net824),
    .Y(_1623_));
 sky130_fd_sc_hd__nand2_1 _5292_ (.A(_0079_),
    .B(_1623_),
    .Y(_1624_));
 sky130_fd_sc_hd__mux2i_1 _5293_ (.A0(\dp.rf.rf[26][2] ),
    .A1(\dp.rf.rf[27][2] ),
    .S(net823),
    .Y(_1625_));
 sky130_fd_sc_hd__nand3_1 _5294_ (.A(net821),
    .B(net16),
    .C(_1625_),
    .Y(_1626_));
 sky130_fd_sc_hd__o2111ai_4 _5295_ (.A1(net821),
    .A2(_1622_),
    .B1(_1624_),
    .C1(_1626_),
    .D1(_0094_),
    .Y(_1627_));
 sky130_fd_sc_hd__o211ai_4 _5296_ (.A1(_1610_),
    .A2(_1613_),
    .B1(_1621_),
    .C1(_1627_),
    .Y(net155));
 sky130_fd_sc_hd__mux2_8 _5297_ (.A0(_3454_[0]),
    .A1(net155),
    .S(_0121_),
    .X(_1628_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_102 ();
 sky130_fd_sc_hd__xnor2_4 _5300_ (.A(_0151_),
    .B(_1628_),
    .Y(_3435_[0]));
 sky130_fd_sc_hd__inv_1 _5301_ (.A(_3435_[0]),
    .Y(_3439_[0]));
 sky130_fd_sc_hd__mux4_2 _5302_ (.A0(\dp.rf.rf[2][2] ),
    .A1(\dp.rf.rf[3][2] ),
    .A2(\dp.rf.rf[6][2] ),
    .A3(\dp.rf.rf[7][2] ),
    .S0(net7),
    .S1(net9),
    .X(_1631_));
 sky130_fd_sc_hd__nand2_1 _5303_ (.A(net8),
    .B(_1631_),
    .Y(_1632_));
 sky130_fd_sc_hd__mux2_1 _5304_ (.A0(\dp.rf.rf[1][2] ),
    .A1(\dp.rf.rf[5][2] ),
    .S(net9),
    .X(_1633_));
 sky130_fd_sc_hd__o221ai_1 _5305_ (.A1(\dp.rf.rf[4][2] ),
    .A2(_0395_),
    .B1(_1633_),
    .B2(_0400_),
    .C1(_0186_),
    .Y(_1634_));
 sky130_fd_sc_hd__mux4_2 _5306_ (.A0(\dp.rf.rf[10][2] ),
    .A1(\dp.rf.rf[11][2] ),
    .A2(\dp.rf.rf[14][2] ),
    .A3(\dp.rf.rf[15][2] ),
    .S0(net7),
    .S1(net9),
    .X(_1635_));
 sky130_fd_sc_hd__mux4_2 _5307_ (.A0(\dp.rf.rf[8][2] ),
    .A1(\dp.rf.rf[9][2] ),
    .A2(\dp.rf.rf[12][2] ),
    .A3(\dp.rf.rf[13][2] ),
    .S0(net7),
    .S1(net9),
    .X(_1636_));
 sky130_fd_sc_hd__mux2i_1 _5308_ (.A0(_1635_),
    .A1(_1636_),
    .S(_0186_),
    .Y(_1637_));
 sky130_fd_sc_hd__a32oi_2 _5309_ (.A1(_0389_),
    .A2(_1632_),
    .A3(_1634_),
    .B1(_1637_),
    .B2(net797),
    .Y(_1638_));
 sky130_fd_sc_hd__mux4_2 _5310_ (.A0(\dp.rf.rf[26][2] ),
    .A1(\dp.rf.rf[27][2] ),
    .A2(\dp.rf.rf[30][2] ),
    .A3(\dp.rf.rf[31][2] ),
    .S0(net7),
    .S1(net9),
    .X(_1639_));
 sky130_fd_sc_hd__mux4_2 _5311_ (.A0(\dp.rf.rf[24][2] ),
    .A1(\dp.rf.rf[25][2] ),
    .A2(\dp.rf.rf[28][2] ),
    .A3(\dp.rf.rf[29][2] ),
    .S0(net7),
    .S1(net9),
    .X(_1640_));
 sky130_fd_sc_hd__o311a_1 _5312_ (.A1(\dp.rf.rf[24][2] ),
    .A2(_0134_),
    .A3(_0135_),
    .B1(_1640_),
    .C1(_0186_),
    .X(_1641_));
 sky130_fd_sc_hd__a211o_4 _5313_ (.A1(_0304_),
    .A2(_1639_),
    .B1(_1641_),
    .C1(_0192_),
    .X(_1642_));
 sky130_fd_sc_hd__mux4_2 _5314_ (.A0(\dp.rf.rf[18][2] ),
    .A1(\dp.rf.rf[19][2] ),
    .A2(\dp.rf.rf[22][2] ),
    .A3(\dp.rf.rf[23][2] ),
    .S0(net7),
    .S1(net9),
    .X(_1643_));
 sky130_fd_sc_hd__o211ai_1 _5315_ (.A1(_0134_),
    .A2(_0135_),
    .B1(_1643_),
    .C1(net8),
    .Y(_1644_));
 sky130_fd_sc_hd__mux4_2 _5316_ (.A0(\dp.rf.rf[16][2] ),
    .A1(\dp.rf.rf[17][2] ),
    .A2(\dp.rf.rf[20][2] ),
    .A3(\dp.rf.rf[21][2] ),
    .S0(net7),
    .S1(net9),
    .X(_1645_));
 sky130_fd_sc_hd__a21oi_1 _5317_ (.A1(_0186_),
    .A2(_1645_),
    .B1(net10),
    .Y(_1646_));
 sky130_fd_sc_hd__a21oi_2 _5318_ (.A1(_1644_),
    .A2(_1646_),
    .B1(net794),
    .Y(_1647_));
 sky130_fd_sc_hd__a22o_4 _5319_ (.A1(net780),
    .A2(_1638_),
    .B1(_1642_),
    .B2(_1647_),
    .X(_3434_[0]));
 sky130_fd_sc_hd__inv_6 _5320_ (.A(_3434_[0]),
    .Y(_3438_[0]));
 sky130_fd_sc_hd__a22o_4 _5321_ (.A1(net31),
    .A2(_0042_),
    .B1(_1517_),
    .B2(net14),
    .X(_3191_[0]));
 sky130_fd_sc_hd__mux2_1 _5322_ (.A0(\dp.rf.rf[26][1] ),
    .A1(\dp.rf.rf[27][1] ),
    .S(net824),
    .X(_1648_));
 sky130_fd_sc_hd__mux2i_1 _5323_ (.A0(\dp.rf.rf[18][1] ),
    .A1(\dp.rf.rf[19][1] ),
    .S(net824),
    .Y(_1649_));
 sky130_fd_sc_hd__a2bb2oi_1 _5324_ (.A1_N(_0073_),
    .A2_N(_1648_),
    .B1(_0079_),
    .B2(_1649_),
    .Y(_1650_));
 sky130_fd_sc_hd__mux2i_1 _5325_ (.A0(\dp.rf.rf[16][1] ),
    .A1(\dp.rf.rf[17][1] ),
    .S(net824),
    .Y(_1651_));
 sky130_fd_sc_hd__mux2i_1 _5326_ (.A0(\dp.rf.rf[24][1] ),
    .A1(\dp.rf.rf[25][1] ),
    .S(net824),
    .Y(_1652_));
 sky130_fd_sc_hd__a22oi_1 _5327_ (.A1(_0086_),
    .A2(_1651_),
    .B1(_1652_),
    .B2(_0064_),
    .Y(_1653_));
 sky130_fd_sc_hd__nand3_1 _5328_ (.A(_0094_),
    .B(_1650_),
    .C(_1653_),
    .Y(_1654_));
 sky130_fd_sc_hd__mux2_1 _5329_ (.A0(\dp.rf.rf[10][1] ),
    .A1(\dp.rf.rf[11][1] ),
    .S(net824),
    .X(_1655_));
 sky130_fd_sc_hd__mux2i_1 _5330_ (.A0(\dp.rf.rf[0][1] ),
    .A1(\dp.rf.rf[1][1] ),
    .S(net824),
    .Y(_1656_));
 sky130_fd_sc_hd__nand2_1 _5331_ (.A(_0086_),
    .B(_1656_),
    .Y(_1657_));
 sky130_fd_sc_hd__mux2i_1 _5332_ (.A0(\dp.rf.rf[2][1] ),
    .A1(\dp.rf.rf[3][1] ),
    .S(net824),
    .Y(_1658_));
 sky130_fd_sc_hd__mux2i_1 _5333_ (.A0(\dp.rf.rf[8][1] ),
    .A1(\dp.rf.rf[9][1] ),
    .S(net824),
    .Y(_1659_));
 sky130_fd_sc_hd__a221oi_1 _5334_ (.A1(_0079_),
    .A2(_1658_),
    .B1(_1659_),
    .B2(_0064_),
    .C1(_0089_),
    .Y(_1660_));
 sky130_fd_sc_hd__o211ai_1 _5335_ (.A1(_0073_),
    .A2(_1655_),
    .B1(_1657_),
    .C1(_1660_),
    .Y(_1661_));
 sky130_fd_sc_hd__mux4_2 _5336_ (.A0(\dp.rf.rf[4][1] ),
    .A1(\dp.rf.rf[5][1] ),
    .A2(\dp.rf.rf[6][1] ),
    .A3(\dp.rf.rf[7][1] ),
    .S0(net824),
    .S1(net821),
    .X(_1662_));
 sky130_fd_sc_hd__mux4_2 _5337_ (.A0(\dp.rf.rf[12][1] ),
    .A1(\dp.rf.rf[13][1] ),
    .A2(\dp.rf.rf[14][1] ),
    .A3(\dp.rf.rf[15][1] ),
    .S0(net824),
    .S1(net821),
    .X(_1663_));
 sky130_fd_sc_hd__mux2_1 _5338_ (.A0(_1662_),
    .A1(_1663_),
    .S(net16),
    .X(_1664_));
 sky130_fd_sc_hd__nand3_1 _5339_ (.A(_0092_),
    .B(net15),
    .C(_1664_),
    .Y(_1665_));
 sky130_fd_sc_hd__mux4_2 _5340_ (.A0(\dp.rf.rf[20][1] ),
    .A1(\dp.rf.rf[21][1] ),
    .A2(\dp.rf.rf[22][1] ),
    .A3(\dp.rf.rf[23][1] ),
    .S0(net824),
    .S1(net821),
    .X(_1666_));
 sky130_fd_sc_hd__mux4_2 _5341_ (.A0(\dp.rf.rf[28][1] ),
    .A1(\dp.rf.rf[29][1] ),
    .A2(\dp.rf.rf[30][1] ),
    .A3(\dp.rf.rf[31][1] ),
    .S0(net824),
    .S1(net821),
    .X(_1667_));
 sky130_fd_sc_hd__mux2_1 _5342_ (.A0(_1666_),
    .A1(_1667_),
    .S(net16),
    .X(_1668_));
 sky130_fd_sc_hd__nand3_1 _5343_ (.A(net17),
    .B(net15),
    .C(_1668_),
    .Y(_1669_));
 sky130_fd_sc_hd__nand4_1 _5344_ (.A(_1665_),
    .B(_1661_),
    .C(_1669_),
    .D(_1654_),
    .Y(_1670_));
 sky130_fd_sc_hd__and2_4 _5345_ (.A(_0351_),
    .B(net775),
    .X(net144));
 sky130_fd_sc_hd__and2_4 _5346_ (.A(_0148_),
    .B(_3191_[0]),
    .X(_1671_));
 sky130_fd_sc_hd__a31o_4 _5347_ (.A1(_1670_),
    .A2(_0121_),
    .A3(_0351_),
    .B1(_1671_),
    .X(_1672_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_100 ();
 sky130_fd_sc_hd__xnor2_4 _5350_ (.A(_0151_),
    .B(_1672_),
    .Y(_3186_[0]));
 sky130_fd_sc_hd__inv_1 _5351_ (.A(_3186_[0]),
    .Y(_3445_[0]));
 sky130_fd_sc_hd__a221oi_1 _5352_ (.A1(\dp.rf.rf[11][1] ),
    .A2(net7),
    .B1(net788),
    .B2(\dp.rf.rf[10][1] ),
    .C1(net791),
    .Y(_1675_));
 sky130_fd_sc_hd__mux2_1 _5353_ (.A0(\dp.rf.rf[14][1] ),
    .A1(\dp.rf.rf[15][1] ),
    .S(net7),
    .X(_1676_));
 sky130_fd_sc_hd__o21ai_0 _5354_ (.A1(_0231_),
    .A2(_1676_),
    .B1(_0304_),
    .Y(_1677_));
 sky130_fd_sc_hd__mux4_2 _5355_ (.A0(\dp.rf.rf[8][1] ),
    .A1(\dp.rf.rf[9][1] ),
    .A2(\dp.rf.rf[12][1] ),
    .A3(\dp.rf.rf[13][1] ),
    .S0(net7),
    .S1(net9),
    .X(_1678_));
 sky130_fd_sc_hd__a21oi_1 _5356_ (.A1(_0186_),
    .A2(_1678_),
    .B1(_0255_),
    .Y(_1679_));
 sky130_fd_sc_hd__o21ai_0 _5357_ (.A1(_1675_),
    .A2(_1677_),
    .B1(_1679_),
    .Y(_1680_));
 sky130_fd_sc_hd__mux4_2 _5358_ (.A0(\dp.rf.rf[0][1] ),
    .A1(\dp.rf.rf[1][1] ),
    .A2(\dp.rf.rf[4][1] ),
    .A3(\dp.rf.rf[5][1] ),
    .S0(net7),
    .S1(net9),
    .X(_1681_));
 sky130_fd_sc_hd__o211ai_1 _5359_ (.A1(\dp.rf.rf[0][1] ),
    .A2(_0347_),
    .B1(_1681_),
    .C1(_0186_),
    .Y(_1682_));
 sky130_fd_sc_hd__mux4_2 _5360_ (.A0(\dp.rf.rf[2][1] ),
    .A1(\dp.rf.rf[3][1] ),
    .A2(\dp.rf.rf[6][1] ),
    .A3(\dp.rf.rf[7][1] ),
    .S0(net7),
    .S1(net9),
    .X(_1683_));
 sky130_fd_sc_hd__a21oi_1 _5361_ (.A1(net8),
    .A2(_1683_),
    .B1(net10),
    .Y(_1684_));
 sky130_fd_sc_hd__nand2_1 _5362_ (.A(_1682_),
    .B(_1684_),
    .Y(_1685_));
 sky130_fd_sc_hd__mux4_2 _5363_ (.A0(\dp.rf.rf[18][1] ),
    .A1(\dp.rf.rf[19][1] ),
    .A2(\dp.rf.rf[22][1] ),
    .A3(\dp.rf.rf[23][1] ),
    .S0(net7),
    .S1(net9),
    .X(_1686_));
 sky130_fd_sc_hd__nand2_1 _5364_ (.A(_0304_),
    .B(_1686_),
    .Y(_1687_));
 sky130_fd_sc_hd__inv_1 _5365_ (.A(\dp.rf.rf[20][1] ),
    .Y(_1688_));
 sky130_fd_sc_hd__mux2i_1 _5366_ (.A0(\dp.rf.rf[17][1] ),
    .A1(\dp.rf.rf[21][1] ),
    .S(net9),
    .Y(_1689_));
 sky130_fd_sc_hd__a221oi_1 _5367_ (.A1(_1688_),
    .A2(_0173_),
    .B1(_1689_),
    .B2(net7),
    .C1(net8),
    .Y(_1690_));
 sky130_fd_sc_hd__o22ai_1 _5368_ (.A1(\dp.rf.rf[16][1] ),
    .A2(net784),
    .B1(_1690_),
    .B2(net790),
    .Y(_1691_));
 sky130_fd_sc_hd__a21oi_1 _5369_ (.A1(_1687_),
    .A2(_1691_),
    .B1(net794),
    .Y(_1692_));
 sky130_fd_sc_hd__a221oi_1 _5370_ (.A1(\dp.rf.rf[27][1] ),
    .A2(net7),
    .B1(net788),
    .B2(\dp.rf.rf[26][1] ),
    .C1(net791),
    .Y(_1693_));
 sky130_fd_sc_hd__mux2_1 _5371_ (.A0(\dp.rf.rf[30][1] ),
    .A1(\dp.rf.rf[31][1] ),
    .S(net7),
    .X(_1694_));
 sky130_fd_sc_hd__o21ai_0 _5372_ (.A1(_0231_),
    .A2(_1694_),
    .B1(_0304_),
    .Y(_1695_));
 sky130_fd_sc_hd__mux4_2 _5373_ (.A0(\dp.rf.rf[24][1] ),
    .A1(\dp.rf.rf[25][1] ),
    .A2(net251),
    .A3(net250),
    .S0(net7),
    .S1(net9),
    .X(_1696_));
 sky130_fd_sc_hd__a21oi_1 _5374_ (.A1(_0186_),
    .A2(_1696_),
    .B1(_0255_),
    .Y(_1697_));
 sky130_fd_sc_hd__o21ai_1 _5375_ (.A1(_1693_),
    .A2(_1695_),
    .B1(_1697_),
    .Y(_1698_));
 sky130_fd_sc_hd__a32o_4 _5376_ (.A1(net780),
    .A2(_1680_),
    .A3(_1685_),
    .B1(_1692_),
    .B2(_1698_),
    .X(_3185_[0]));
 sky130_fd_sc_hd__inv_8 _5377_ (.A(_3185_[0]),
    .Y(_1699_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_99 ();
 sky130_fd_sc_hd__nand3_2 _5379_ (.A(_0123_),
    .B(_0035_),
    .C(net803),
    .Y(_1700_));
 sky130_fd_sc_hd__nand2_2 _5380_ (.A(net5),
    .B(_1700_),
    .Y(_1701_));
 sky130_fd_sc_hd__nor2_1 _5381_ (.A(net814),
    .B(net815),
    .Y(_1702_));
 sky130_fd_sc_hd__nand2_4 _5382_ (.A(_0347_),
    .B(_0901_),
    .Y(_1703_));
 sky130_fd_sc_hd__a21oi_2 _5383_ (.A1(net27),
    .A2(_0127_),
    .B1(_0130_),
    .Y(_1704_));
 sky130_fd_sc_hd__a21oi_1 _5384_ (.A1(net814),
    .A2(net815),
    .B1(_1704_),
    .Y(_1705_));
 sky130_fd_sc_hd__nand2_4 _5385_ (.A(net814),
    .B(net815),
    .Y(_1706_));
 sky130_fd_sc_hd__a21oi_1 _5386_ (.A1(_1706_),
    .A2(_1700_),
    .B1(net5),
    .Y(_1707_));
 sky130_fd_sc_hd__a2111oi_1 _5387_ (.A1(_1701_),
    .A2(_1702_),
    .B1(_1703_),
    .C1(_1705_),
    .D1(_1707_),
    .Y(_1708_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_97 ();
 sky130_fd_sc_hd__nor4b_2 _5390_ (.A(net815),
    .B(_1703_),
    .C(_1704_),
    .D_N(net814),
    .Y(_1711_));
 sky130_fd_sc_hd__nand2_4 _5391_ (.A(net5),
    .B(net773),
    .Y(_1712_));
 sky130_fd_sc_hd__nor2_4 _5392_ (.A(net27),
    .B(_0130_),
    .Y(_1713_));
 sky130_fd_sc_hd__nor2b_1 _5393_ (.A(net814),
    .B_N(net816),
    .Y(_1714_));
 sky130_fd_sc_hd__nand2b_2 _5394_ (.A_N(net5),
    .B(net815),
    .Y(_1715_));
 sky130_fd_sc_hd__or4_4 _5395_ (.A(net799),
    .B(_1713_),
    .C(_1714_),
    .D(_1715_),
    .X(_1716_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_96 ();
 sky130_fd_sc_hd__o21ai_0 _5397_ (.A1(_3200_[0]),
    .A2(_1712_),
    .B1(_1716_),
    .Y(_1718_));
 sky130_fd_sc_hd__a21oi_1 _5398_ (.A1(_3196_[0]),
    .A2(net774),
    .B1(_1718_),
    .Y(_1719_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_95 ();
 sky130_fd_sc_hd__or4b_4 _5400_ (.A(net815),
    .B(_1703_),
    .C(_1704_),
    .D_N(net814),
    .X(_1721_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_94 ();
 sky130_fd_sc_hd__nor4_1 _5402_ (.A(_0123_),
    .B(net814),
    .C(_0127_),
    .D(_0130_),
    .Y(_1723_));
 sky130_fd_sc_hd__o21ai_2 _5403_ (.A1(net5),
    .A2(_1723_),
    .B1(net815),
    .Y(_1724_));
 sky130_fd_sc_hd__nor2_1 _5404_ (.A(net815),
    .B(_1713_),
    .Y(_1725_));
 sky130_fd_sc_hd__o21ai_2 _5405_ (.A1(net5),
    .A2(_1725_),
    .B1(net814),
    .Y(_1726_));
 sky130_fd_sc_hd__a31o_4 _5406_ (.A1(_1701_),
    .A2(_1724_),
    .A3(_1726_),
    .B1(_1703_),
    .X(_1727_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_93 ();
 sky130_fd_sc_hd__nand2_1 _5408_ (.A(_0151_),
    .B(_1727_),
    .Y(_1729_));
 sky130_fd_sc_hd__o21ai_0 _5409_ (.A1(net5),
    .A2(_1721_),
    .B1(_1729_),
    .Y(_1730_));
 sky130_fd_sc_hd__a31oi_4 _5410_ (.A1(_1701_),
    .A2(_1724_),
    .A3(_1726_),
    .B1(_1703_),
    .Y(_1731_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_92 ();
 sky130_fd_sc_hd__nor3_1 _5412_ (.A(_3197_[0]),
    .B(_0151_),
    .C(_1731_),
    .Y(_1733_));
 sky130_fd_sc_hd__a21oi_1 _5413_ (.A1(_3197_[0]),
    .A2(_1730_),
    .B1(_1733_),
    .Y(_1734_));
 sky130_fd_sc_hd__nor4b_1 _5414_ (.A(net814),
    .B(_1704_),
    .C(_1703_),
    .D_N(net5),
    .Y(_1735_));
 sky130_fd_sc_hd__clkinv_1 _5415_ (.A(_3309_[0]),
    .Y(_1736_));
 sky130_fd_sc_hd__nor2_1 _5416_ (.A(_3317_[0]),
    .B(_3316_[0]),
    .Y(_1737_));
 sky130_fd_sc_hd__nor2_1 _5417_ (.A(_1736_),
    .B(_1737_),
    .Y(_1738_));
 sky130_fd_sc_hd__o21ai_2 _5418_ (.A1(_3308_[0]),
    .A2(_1738_),
    .B1(_3301_[0]),
    .Y(_1739_));
 sky130_fd_sc_hd__nand2b_4 _5419_ (.A_N(_3300_[0]),
    .B(_1739_),
    .Y(_1740_));
 sky130_fd_sc_hd__clkinv_2 _5420_ (.A(_3413_[0]),
    .Y(_1741_));
 sky130_fd_sc_hd__clkinv_4 _5421_ (.A(_3429_[0]),
    .Y(_1742_));
 sky130_fd_sc_hd__a21oi_4 _5422_ (.A1(_3437_[0]),
    .A2(_3187_[0]),
    .B1(_3436_[0]),
    .Y(_1743_));
 sky130_fd_sc_hd__o21bai_4 _5423_ (.A1(_1743_),
    .A2(_1742_),
    .B1_N(_3428_[0]),
    .Y(_1744_));
 sky130_fd_sc_hd__a21oi_2 _5424_ (.A1(_1744_),
    .A2(_3421_[0]),
    .B1(_3420_[0]),
    .Y(_1745_));
 sky130_fd_sc_hd__o21bai_2 _5425_ (.A1(_1745_),
    .A2(_1741_),
    .B1_N(_3412_[0]),
    .Y(_1746_));
 sky130_fd_sc_hd__a21oi_2 _5426_ (.A1(_1746_),
    .A2(_3405_[0]),
    .B1(_3404_[0]),
    .Y(_1747_));
 sky130_fd_sc_hd__nand3_1 _5427_ (.A(_3381_[0]),
    .B(_3389_[0]),
    .C(_3397_[0]),
    .Y(_1748_));
 sky130_fd_sc_hd__and3_1 _5428_ (.A(_3381_[0]),
    .B(_3389_[0]),
    .C(_3396_[0]),
    .X(_1749_));
 sky130_fd_sc_hd__a21oi_1 _5429_ (.A1(_3388_[0]),
    .A2(_3381_[0]),
    .B1(_1749_),
    .Y(_1750_));
 sky130_fd_sc_hd__nor3_1 _5430_ (.A(_3372_[0]),
    .B(_3364_[0]),
    .C(_3380_[0]),
    .Y(_1751_));
 sky130_fd_sc_hd__o211ai_1 _5431_ (.A1(_1748_),
    .A2(_1747_),
    .B1(_1750_),
    .C1(_1751_),
    .Y(_1752_));
 sky130_fd_sc_hd__clkinv_1 _5432_ (.A(_3365_[0]),
    .Y(_1753_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_91 ();
 sky130_fd_sc_hd__nor2_2 _5434_ (.A(_3372_[0]),
    .B(_3373_[0]),
    .Y(_1755_));
 sky130_fd_sc_hd__o21bai_4 _5435_ (.A1(_1753_),
    .A2(_1755_),
    .B1_N(_3364_[0]),
    .Y(_1756_));
 sky130_fd_sc_hd__a211oi_1 _5436_ (.A1(_3308_[0]),
    .A2(_3301_[0]),
    .B1(_3300_[0]),
    .C1(_3316_[0]),
    .Y(_1757_));
 sky130_fd_sc_hd__nand2b_1 _5437_ (.A_N(_3356_[0]),
    .B(_1757_),
    .Y(_1758_));
 sky130_fd_sc_hd__inv_1 _5438_ (.A(_3333_[0]),
    .Y(_1759_));
 sky130_fd_sc_hd__a21oi_2 _5439_ (.A1(_3348_[0]),
    .A2(_3341_[0]),
    .B1(_3340_[0]),
    .Y(_1760_));
 sky130_fd_sc_hd__o21bai_1 _5440_ (.A1(_1760_),
    .A2(_1759_),
    .B1_N(_3332_[0]),
    .Y(_1761_));
 sky130_fd_sc_hd__a21o_1 _5441_ (.A1(_3325_[0]),
    .A2(_1761_),
    .B1(_3324_[0]),
    .X(_1762_));
 sky130_fd_sc_hd__a211o_4 _5442_ (.A1(net193),
    .A2(_1756_),
    .B1(_1758_),
    .C1(net269),
    .X(_1763_));
 sky130_fd_sc_hd__nand4_1 _5443_ (.A(_3325_[0]),
    .B(_3333_[0]),
    .C(net264),
    .D(_3349_[0]),
    .Y(_1764_));
 sky130_fd_sc_hd__nor2_1 _5444_ (.A(_3356_[0]),
    .B(_3357_[0]),
    .Y(_1765_));
 sky130_fd_sc_hd__a21oi_2 _5445_ (.A1(_3325_[0]),
    .A2(_1761_),
    .B1(_3324_[0]),
    .Y(_1766_));
 sky130_fd_sc_hd__o211ai_1 _5446_ (.A1(_1765_),
    .A2(_1764_),
    .B1(_1757_),
    .C1(_1766_),
    .Y(_1767_));
 sky130_fd_sc_hd__clkinv_2 _5447_ (.A(_3237_[0]),
    .Y(_1768_));
 sky130_fd_sc_hd__inv_4 _5448_ (.A(_3245_[0]),
    .Y(_1769_));
 sky130_fd_sc_hd__inv_4 _5449_ (.A(_3253_[0]),
    .Y(_1770_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_89 ();
 sky130_fd_sc_hd__nand2_1 _5452_ (.A(_3261_[0]),
    .B(_3269_[0]),
    .Y(_1773_));
 sky130_fd_sc_hd__nor4_4 _5453_ (.A(_1768_),
    .B(_1769_),
    .C(_1770_),
    .D(_1773_),
    .Y(_1774_));
 sky130_fd_sc_hd__and2_4 _5454_ (.A(_3277_[0]),
    .B(_3285_[0]),
    .X(_1775_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_88 ();
 sky130_fd_sc_hd__and3_1 _5456_ (.A(_3293_[0]),
    .B(_1774_),
    .C(_1775_),
    .X(_1777_));
 sky130_fd_sc_hd__nand4_1 _5457_ (.A(_1763_),
    .B(_1740_),
    .C(_1767_),
    .D(_1777_),
    .Y(_1778_));
 sky130_fd_sc_hd__a21o_1 _5458_ (.A1(_3292_[0]),
    .A2(_3285_[0]),
    .B1(_3284_[0]),
    .X(_1779_));
 sky130_fd_sc_hd__a21o_1 _5459_ (.A1(_3277_[0]),
    .A2(_1779_),
    .B1(_3276_[0]),
    .X(_1780_));
 sky130_fd_sc_hd__a21oi_2 _5460_ (.A1(_3269_[0]),
    .A2(_1780_),
    .B1(_3268_[0]),
    .Y(_1781_));
 sky130_fd_sc_hd__nand4_1 _5461_ (.A(net270),
    .B(_3261_[0]),
    .C(_3245_[0]),
    .D(_3253_[0]),
    .Y(_1782_));
 sky130_fd_sc_hd__a21oi_1 _5462_ (.A1(_3260_[0]),
    .A2(_3253_[0]),
    .B1(_3252_[0]),
    .Y(_1783_));
 sky130_fd_sc_hd__o21bai_1 _5463_ (.A1(_1769_),
    .A2(_1783_),
    .B1_N(_3244_[0]),
    .Y(_1784_));
 sky130_fd_sc_hd__a21oi_1 _5464_ (.A1(net252),
    .A2(_1784_),
    .B1(_3236_[0]),
    .Y(_1785_));
 sky130_fd_sc_hd__o21ai_2 _5465_ (.A1(_1781_),
    .A2(_1782_),
    .B1(_1785_),
    .Y(_1786_));
 sky130_fd_sc_hd__nor3_1 _5466_ (.A(_3220_[0]),
    .B(_3228_[0]),
    .C(_1786_),
    .Y(_1787_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_87 ();
 sky130_fd_sc_hd__nor3_1 _5468_ (.A(_3229_[0]),
    .B(_3220_[0]),
    .C(_3228_[0]),
    .Y(_1789_));
 sky130_fd_sc_hd__nor2_1 _5469_ (.A(_3221_[0]),
    .B(_3220_[0]),
    .Y(_1790_));
 sky130_fd_sc_hd__a211o_4 _5470_ (.A1(_1787_),
    .A2(_1778_),
    .B1(_1789_),
    .C1(_1790_),
    .X(_1791_));
 sky130_fd_sc_hd__nand2_1 _5471_ (.A(_3205_[0]),
    .B(_3213_[0]),
    .Y(_1792_));
 sky130_fd_sc_hd__a21oi_1 _5472_ (.A1(_3205_[0]),
    .A2(_3212_[0]),
    .B1(_3204_[0]),
    .Y(_1793_));
 sky130_fd_sc_hd__o21ai_4 _5473_ (.A1(_1792_),
    .A2(_1791_),
    .B1(_1793_),
    .Y(_1794_));
 sky130_fd_sc_hd__nand3b_1 _5474_ (.A_N(net814),
    .B(net815),
    .C(net5),
    .Y(_1795_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_86 ();
 sky130_fd_sc_hd__xnor2_1 _5476_ (.A(_0313_),
    .B(_0340_),
    .Y(_1796_));
 sky130_fd_sc_hd__o21ai_0 _5477_ (.A1(_1704_),
    .A2(_1795_),
    .B1(_1796_),
    .Y(_1797_));
 sky130_fd_sc_hd__xnor2_1 _5478_ (.A(_0151_),
    .B(_1797_),
    .Y(_1798_));
 sky130_fd_sc_hd__xnor2_2 _5479_ (.A(_1794_),
    .B(_1798_),
    .Y(_1799_));
 sky130_fd_sc_hd__nand2_2 _5480_ (.A(_1735_),
    .B(_1799_),
    .Y(_1800_));
 sky130_fd_sc_hd__mux2i_4 _5481_ (.A0(_3464_[0]),
    .A1(net159),
    .S(_0121_),
    .Y(_1801_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_85 ();
 sky130_fd_sc_hd__o21ai_4 _5483_ (.A1(_0121_),
    .A2(_3458_[0]),
    .B1(_1573_),
    .Y(_1803_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_84 ();
 sky130_fd_sc_hd__a31oi_4 _5485_ (.A1(net775),
    .A2(_0121_),
    .A3(_0351_),
    .B1(_1671_),
    .Y(_1805_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_82 ();
 sky130_fd_sc_hd__mux2i_1 _5488_ (.A0(_3342_[0]),
    .A1(net761),
    .S(net744),
    .Y(_1808_));
 sky130_fd_sc_hd__mux2i_2 _5489_ (.A0(net763),
    .A1(_1203_),
    .S(net744),
    .Y(_1809_));
 sky130_fd_sc_hd__a21o_4 _5490_ (.A1(net133),
    .A2(_0121_),
    .B1(_0149_),
    .X(_1810_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_80 ();
 sky130_fd_sc_hd__mux2i_2 _5493_ (.A0(_1808_),
    .A1(_1809_),
    .S(net742),
    .Y(_1813_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_78 ();
 sky130_fd_sc_hd__mux2i_1 _5496_ (.A0(net760),
    .A1(net758),
    .S(net744),
    .Y(_1816_));
 sky130_fd_sc_hd__mux2i_1 _5497_ (.A0(net759),
    .A1(net757),
    .S(net744),
    .Y(_1817_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_76 ();
 sky130_fd_sc_hd__mux2i_2 _5500_ (.A0(_1816_),
    .A1(_1817_),
    .S(net769),
    .Y(_1820_));
 sky130_fd_sc_hd__mux2i_4 _5501_ (.A0(_3454_[0]),
    .A1(net248),
    .S(_0121_),
    .Y(_1821_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_74 ();
 sky130_fd_sc_hd__mux2i_1 _5504_ (.A0(_1813_),
    .A1(_1820_),
    .S(net737),
    .Y(_1824_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_72 ();
 sky130_fd_sc_hd__clkinvlp_4 _5507_ (.A(_3398_[0]),
    .Y(_3394_[0]));
 sky130_fd_sc_hd__nand2_1 _5508_ (.A(net754),
    .B(net743),
    .Y(_1827_));
 sky130_fd_sc_hd__o21ai_0 _5509_ (.A1(_3394_[0]),
    .A2(net743),
    .B1(_1827_),
    .Y(_1828_));
 sky130_fd_sc_hd__inv_4 _5510_ (.A(net755),
    .Y(_3402_[0]));
 sky130_fd_sc_hd__nand2_1 _5511_ (.A(net753),
    .B(net743),
    .Y(_1829_));
 sky130_fd_sc_hd__o211ai_1 _5512_ (.A1(_3402_[0]),
    .A2(net743),
    .B1(_1829_),
    .C1(net768),
    .Y(_1830_));
 sky130_fd_sc_hd__o21ai_2 _5513_ (.A1(net768),
    .A2(_1828_),
    .B1(_1830_),
    .Y(_1831_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_70 ();
 sky130_fd_sc_hd__nor2_1 _5516_ (.A(net751),
    .B(_1699_),
    .Y(_1834_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_69 ();
 sky130_fd_sc_hd__a211oi_1 _5518_ (.A1(_3426_[0]),
    .A2(net751),
    .B1(_1834_),
    .C1(net768),
    .Y(_1836_));
 sky130_fd_sc_hd__nand2_1 _5519_ (.A(_3438_[0]),
    .B(net751),
    .Y(_1837_));
 sky130_fd_sc_hd__nand2_1 _5520_ (.A(_0237_),
    .B(net743),
    .Y(_1838_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_68 ();
 sky130_fd_sc_hd__a21oi_1 _5522_ (.A1(_1837_),
    .A2(_1838_),
    .B1(net742),
    .Y(_1840_));
 sky130_fd_sc_hd__nor3_1 _5523_ (.A(net740),
    .B(_1836_),
    .C(_1840_),
    .Y(_1841_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_67 ();
 sky130_fd_sc_hd__a211o_1 _5525_ (.A1(net740),
    .A2(_1831_),
    .B1(_1841_),
    .C1(net752),
    .X(_1843_));
 sky130_fd_sc_hd__o21ai_0 _5526_ (.A1(net747),
    .A2(_1824_),
    .B1(_1843_),
    .Y(_1844_));
 sky130_fd_sc_hd__mux2i_4 _5527_ (.A0(_3214_[0]),
    .A1(_3230_[0]),
    .S(net746),
    .Y(_1845_));
 sky130_fd_sc_hd__mux2i_4 _5528_ (.A0(_0314_),
    .A1(_3222_[0]),
    .S(net746),
    .Y(_1846_));
 sky130_fd_sc_hd__mux2_8 _5529_ (.A0(net343),
    .A1(_1846_),
    .S(net742),
    .X(_1847_));
 sky130_fd_sc_hd__mux2i_4 _5530_ (.A0(_3246_[0]),
    .A1(_3262_[0]),
    .S(net331),
    .Y(_1848_));
 sky130_fd_sc_hd__mux2i_4 _5531_ (.A0(net766),
    .A1(net285),
    .S(net746),
    .Y(_1849_));
 sky130_fd_sc_hd__mux2_8 _5532_ (.A0(_1848_),
    .A1(_1849_),
    .S(net742),
    .X(_1850_));
 sky130_fd_sc_hd__mux2i_1 _5533_ (.A0(_1847_),
    .A1(_1850_),
    .S(net738),
    .Y(_1851_));
 sky130_fd_sc_hd__mux2i_4 _5534_ (.A0(_3278_[0]),
    .A1(_3294_[0]),
    .S(net308),
    .Y(_1852_));
 sky130_fd_sc_hd__mux2i_2 _5535_ (.A0(net281),
    .A1(_3286_[0]),
    .S(net745),
    .Y(_1853_));
 sky130_fd_sc_hd__mux2_8 _5536_ (.A0(_1852_),
    .A1(_1853_),
    .S(net742),
    .X(_1854_));
 sky130_fd_sc_hd__mux2i_1 _5537_ (.A0(_3310_[0]),
    .A1(_3326_[0]),
    .S(net744),
    .Y(_1855_));
 sky130_fd_sc_hd__mux2i_2 _5538_ (.A0(net765),
    .A1(net764),
    .S(net744),
    .Y(_1856_));
 sky130_fd_sc_hd__mux2_8 _5539_ (.A0(_1855_),
    .A1(_1856_),
    .S(net742),
    .X(_1857_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_66 ();
 sky130_fd_sc_hd__mux2i_1 _5541_ (.A0(_1854_),
    .A1(_1857_),
    .S(net738),
    .Y(_1859_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_65 ();
 sky130_fd_sc_hd__mux2i_1 _5543_ (.A0(_1851_),
    .A1(_1859_),
    .S(net749),
    .Y(_1861_));
 sky130_fd_sc_hd__nor2_1 _5544_ (.A(net750),
    .B(_1861_),
    .Y(_1862_));
 sky130_fd_sc_hd__or3_4 _5545_ (.A(net5),
    .B(_1706_),
    .C(_1713_),
    .X(_1863_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_62 ();
 sky130_fd_sc_hd__a211oi_2 _5549_ (.A1(net750),
    .A2(_1844_),
    .B1(_1862_),
    .C1(_1863_),
    .Y(_1867_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_61 ();
 sky130_fd_sc_hd__nand3_4 _5551_ (.A(net768),
    .B(_3194_[0]),
    .C(net743),
    .Y(_1869_));
 sky130_fd_sc_hd__nand2_8 _5552_ (.A(_1801_),
    .B(_1863_),
    .Y(_1870_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_60 ();
 sky130_fd_sc_hd__nand2_4 _5554_ (.A(_1803_),
    .B(net739),
    .Y(_1872_));
 sky130_fd_sc_hd__nor3_2 _5555_ (.A(_1869_),
    .B(_1870_),
    .C(_1872_),
    .Y(_1873_));
 sky130_fd_sc_hd__nor3_4 _5556_ (.A(_1716_),
    .B(_1867_),
    .C(_1873_),
    .Y(_1874_));
 sky130_fd_sc_hd__a31oi_4 _5557_ (.A1(_1800_),
    .A2(_1734_),
    .A3(_1719_),
    .B1(_1874_),
    .Y(net66));
 sky130_fd_sc_hd__nand2_8 _5558_ (.A(_0044_),
    .B(_1713_),
    .Y(_1875_));
 sky130_fd_sc_hd__inv_16 _5559_ (.A(_1875_),
    .Y(net98));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_58 ();
 sky130_fd_sc_hd__mux2i_4 _5562_ (.A0(_3230_[0]),
    .A1(_3246_[0]),
    .S(net746),
    .Y(_1878_));
 sky130_fd_sc_hd__mux2i_4 _5563_ (.A0(_1849_),
    .A1(_1878_),
    .S(net742),
    .Y(_1879_));
 sky130_fd_sc_hd__nor2_2 _5564_ (.A(net337),
    .B(_3214_[0]),
    .Y(_1880_));
 sky130_fd_sc_hd__a22oi_2 _5565_ (.A1(_1846_),
    .A2(net771),
    .B1(_1880_),
    .B2(net746),
    .Y(_1881_));
 sky130_fd_sc_hd__mux2i_4 _5566_ (.A0(_1879_),
    .A1(_1881_),
    .S(net740),
    .Y(_1882_));
 sky130_fd_sc_hd__nor2_1 _5567_ (.A(net742),
    .B(_3222_[0]),
    .Y(_1883_));
 sky130_fd_sc_hd__nand2_1 _5568_ (.A(_0314_),
    .B(net751),
    .Y(_1884_));
 sky130_fd_sc_hd__o31ai_2 _5569_ (.A1(net751),
    .A2(_1883_),
    .A3(_1880_),
    .B1(_1884_),
    .Y(_1885_));
 sky130_fd_sc_hd__mux2i_4 _5570_ (.A0(_1879_),
    .A1(_1885_),
    .S(net740),
    .Y(_1886_));
 sky130_fd_sc_hd__mux2i_2 _5571_ (.A0(_1882_),
    .A1(_1886_),
    .S(net816),
    .Y(_1887_));
 sky130_fd_sc_hd__mux2i_4 _5572_ (.A0(_3262_[0]),
    .A1(_3278_[0]),
    .S(net745),
    .Y(_1888_));
 sky130_fd_sc_hd__mux2i_2 _5573_ (.A0(_1853_),
    .A1(_1888_),
    .S(net742),
    .Y(_1889_));
 sky130_fd_sc_hd__mux2i_1 _5574_ (.A0(_3294_[0]),
    .A1(_3310_[0]),
    .S(net744),
    .Y(_1890_));
 sky130_fd_sc_hd__mux2i_4 _5575_ (.A0(_1856_),
    .A1(_1890_),
    .S(net742),
    .Y(_1891_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_57 ();
 sky130_fd_sc_hd__mux2i_1 _5577_ (.A0(_1889_),
    .A1(_1891_),
    .S(net739),
    .Y(_1893_));
 sky130_fd_sc_hd__nand2_2 _5578_ (.A(net749),
    .B(_1893_),
    .Y(_1894_));
 sky130_fd_sc_hd__o21ai_4 _5579_ (.A1(_1887_),
    .A2(net749),
    .B1(_1894_),
    .Y(_1895_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_56 ();
 sky130_fd_sc_hd__mux2i_1 _5581_ (.A0(_3326_[0]),
    .A1(_3342_[0]),
    .S(net744),
    .Y(_1897_));
 sky130_fd_sc_hd__mux2i_4 _5582_ (.A0(_1809_),
    .A1(_1897_),
    .S(net742),
    .Y(_1898_));
 sky130_fd_sc_hd__mux2i_1 _5583_ (.A0(net761),
    .A1(net759),
    .S(net744),
    .Y(_1899_));
 sky130_fd_sc_hd__mux2i_2 _5584_ (.A0(_1816_),
    .A1(_1899_),
    .S(net742),
    .Y(_1900_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_55 ();
 sky130_fd_sc_hd__mux2i_2 _5586_ (.A0(_1898_),
    .A1(_1900_),
    .S(net737),
    .Y(_1902_));
 sky130_fd_sc_hd__nand2_1 _5587_ (.A(net752),
    .B(_1902_),
    .Y(_1903_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_54 ();
 sky130_fd_sc_hd__mux2i_1 _5589_ (.A0(net755),
    .A1(net754),
    .S(net768),
    .Y(_1905_));
 sky130_fd_sc_hd__mux2i_1 _5590_ (.A0(net757),
    .A1(net756),
    .S(net768),
    .Y(_1906_));
 sky130_fd_sc_hd__mux2_1 _5591_ (.A0(_1905_),
    .A1(_1906_),
    .S(net751),
    .X(_1907_));
 sky130_fd_sc_hd__nand2_1 _5592_ (.A(net742),
    .B(net753),
    .Y(_1908_));
 sky130_fd_sc_hd__o21ai_0 _5593_ (.A1(net742),
    .A2(_3426_[0]),
    .B1(_1908_),
    .Y(_1909_));
 sky130_fd_sc_hd__nand2_4 _5594_ (.A(net768),
    .B(_1699_),
    .Y(_1910_));
 sky130_fd_sc_hd__o211ai_1 _5595_ (.A1(net768),
    .A2(_3434_[0]),
    .B1(net743),
    .C1(_1910_),
    .Y(_1911_));
 sky130_fd_sc_hd__o211ai_1 _5596_ (.A1(net743),
    .A2(_1909_),
    .B1(_1911_),
    .C1(net737),
    .Y(_1912_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_53 ();
 sky130_fd_sc_hd__o211ai_1 _5598_ (.A1(net737),
    .A2(_1907_),
    .B1(_1912_),
    .C1(net747),
    .Y(_1914_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_52 ();
 sky130_fd_sc_hd__a21oi_1 _5600_ (.A1(_1903_),
    .A2(_1914_),
    .B1(net268),
    .Y(_1916_));
 sky130_fd_sc_hd__a21oi_2 _5601_ (.A1(net268),
    .A2(_1895_),
    .B1(_1916_),
    .Y(_1917_));
 sky130_fd_sc_hd__nor3_1 _5602_ (.A(net5),
    .B(_1706_),
    .C(_1713_),
    .Y(_1918_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_51 ();
 sky130_fd_sc_hd__nor2_4 _5604_ (.A(net268),
    .B(net778),
    .Y(_1920_));
 sky130_fd_sc_hd__nor2_4 _5605_ (.A(net752),
    .B(net740),
    .Y(_1921_));
 sky130_fd_sc_hd__nand2_2 _5606_ (.A(net742),
    .B(_0237_),
    .Y(_1922_));
 sky130_fd_sc_hd__and3_4 _5607_ (.A(net743),
    .B(_1910_),
    .C(_1922_),
    .X(_1923_));
 sky130_fd_sc_hd__a31oi_4 _5608_ (.A1(_1920_),
    .A2(_1921_),
    .A3(_1923_),
    .B1(_1716_),
    .Y(_1924_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_48 ();
 sky130_fd_sc_hd__nand2_1 _5612_ (.A(net5),
    .B(_3446_[0]),
    .Y(_1928_));
 sky130_fd_sc_hd__o21ai_0 _5613_ (.A1(net5),
    .A2(_3443_[0]),
    .B1(_1928_),
    .Y(_1929_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_47 ();
 sky130_fd_sc_hd__o21ai_0 _5615_ (.A1(_1721_),
    .A2(_1929_),
    .B1(_1716_),
    .Y(_1931_));
 sky130_fd_sc_hd__a221oi_2 _5616_ (.A1(_3442_[0]),
    .A2(net774),
    .B1(_1727_),
    .B2(_3188_[0]),
    .C1(_1931_),
    .Y(_1932_));
 sky130_fd_sc_hd__o22ai_4 _5617_ (.A1(_1863_),
    .A2(_1917_),
    .B1(_1924_),
    .B2(_1932_),
    .Y(net77));
 sky130_fd_sc_hd__mux2i_4 _5618_ (.A0(net285),
    .A1(net281),
    .S(net331),
    .Y(_1933_));
 sky130_fd_sc_hd__mux2_8 _5619_ (.A0(_1888_),
    .A1(_1933_),
    .S(net742),
    .X(_1934_));
 sky130_fd_sc_hd__mux2i_4 _5620_ (.A0(_3286_[0]),
    .A1(net765),
    .S(net308),
    .Y(_1935_));
 sky130_fd_sc_hd__mux2_4 _5621_ (.A0(_1890_),
    .A1(_1935_),
    .S(net742),
    .X(_1936_));
 sky130_fd_sc_hd__mux2i_2 _5622_ (.A0(_1934_),
    .A1(_1936_),
    .S(net738),
    .Y(_1937_));
 sky130_fd_sc_hd__nand2b_1 _5623_ (.A_N(_1937_),
    .B(net748),
    .Y(_1938_));
 sky130_fd_sc_hd__mux2i_4 _5624_ (.A0(_3222_[0]),
    .A1(net766),
    .S(net746),
    .Y(_1939_));
 sky130_fd_sc_hd__mux2_8 _5625_ (.A0(_1878_),
    .A1(_1939_),
    .S(net742),
    .X(_1940_));
 sky130_fd_sc_hd__nor2_1 _5626_ (.A(net771),
    .B(_0313_),
    .Y(_1941_));
 sky130_fd_sc_hd__a211oi_4 _5627_ (.A1(net771),
    .A2(_3214_[0]),
    .B1(net751),
    .C1(_1941_),
    .Y(_1942_));
 sky130_fd_sc_hd__mux2_8 _5628_ (.A0(_1940_),
    .A1(_1942_),
    .S(net740),
    .X(_1943_));
 sky130_fd_sc_hd__a21oi_1 _5629_ (.A1(net771),
    .A2(net746),
    .B1(_0313_),
    .Y(_1944_));
 sky130_fd_sc_hd__a311oi_1 _5630_ (.A1(net771),
    .A2(_3214_[0]),
    .A3(net746),
    .B1(_1944_),
    .C1(net739),
    .Y(_1945_));
 sky130_fd_sc_hd__a21oi_2 _5631_ (.A1(net739),
    .A2(_1940_),
    .B1(_1945_),
    .Y(_1946_));
 sky130_fd_sc_hd__nand2_1 _5632_ (.A(net816),
    .B(_1946_),
    .Y(_1947_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_46 ();
 sky130_fd_sc_hd__o211ai_1 _5634_ (.A1(net816),
    .A2(_1943_),
    .B1(_1947_),
    .C1(net752),
    .Y(_1949_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_45 ();
 sky130_fd_sc_hd__nand2_2 _5636_ (.A(net741),
    .B(net778),
    .Y(_1951_));
 sky130_fd_sc_hd__a21oi_2 _5637_ (.A1(_1938_),
    .A2(_1949_),
    .B1(_1951_),
    .Y(_1952_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_44 ();
 sky130_fd_sc_hd__nand2_1 _5639_ (.A(net758),
    .B(net751),
    .Y(_1954_));
 sky130_fd_sc_hd__nand2_1 _5640_ (.A(net756),
    .B(net744),
    .Y(_1955_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_43 ();
 sky130_fd_sc_hd__nand2_1 _5642_ (.A(net757),
    .B(net751),
    .Y(_1957_));
 sky130_fd_sc_hd__nand2_1 _5643_ (.A(net755),
    .B(net744),
    .Y(_1958_));
 sky130_fd_sc_hd__and3_1 _5644_ (.A(net768),
    .B(_1957_),
    .C(_1958_),
    .X(_1959_));
 sky130_fd_sc_hd__a31oi_1 _5645_ (.A1(net742),
    .A2(_1954_),
    .A3(_1955_),
    .B1(_1959_),
    .Y(_1960_));
 sky130_fd_sc_hd__nand2_1 _5646_ (.A(_3438_[0]),
    .B(net743),
    .Y(_1961_));
 sky130_fd_sc_hd__nand2_2 _5647_ (.A(_0237_),
    .B(net751),
    .Y(_1962_));
 sky130_fd_sc_hd__nor3_2 _5648_ (.A(net768),
    .B(net751),
    .C(_1699_),
    .Y(_1963_));
 sky130_fd_sc_hd__a31oi_4 _5649_ (.A1(net768),
    .A2(_1962_),
    .A3(_1961_),
    .B1(_1963_),
    .Y(_1964_));
 sky130_fd_sc_hd__nand2_1 _5650_ (.A(_1863_),
    .B(_1964_),
    .Y(_1965_));
 sky130_fd_sc_hd__a311oi_2 _5651_ (.A1(_0351_),
    .A2(_0121_),
    .A3(net775),
    .B1(_1671_),
    .C1(_3434_[0]),
    .Y(_1966_));
 sky130_fd_sc_hd__inv_4 _5652_ (.A(_3422_[0]),
    .Y(_3418_[0]));
 sky130_fd_sc_hd__nor2_1 _5653_ (.A(_3418_[0]),
    .B(net743),
    .Y(_1967_));
 sky130_fd_sc_hd__inv_1 _5654_ (.A(_3414_[0]),
    .Y(_3410_[0]));
 sky130_fd_sc_hd__nand3_4 _5655_ (.A(_1592_),
    .B(_1609_),
    .C(net379),
    .Y(_1968_));
 sky130_fd_sc_hd__o211ai_1 _5656_ (.A1(_3410_[0]),
    .A2(net743),
    .B1(_1968_),
    .C1(net742),
    .Y(_1969_));
 sky130_fd_sc_hd__o311ai_0 _5657_ (.A1(net742),
    .A2(_1966_),
    .A3(_1967_),
    .B1(net778),
    .C1(_1969_),
    .Y(_1970_));
 sky130_fd_sc_hd__nand3_1 _5658_ (.A(net737),
    .B(_1965_),
    .C(_1970_),
    .Y(_1971_));
 sky130_fd_sc_hd__o31ai_1 _5659_ (.A1(net737),
    .A2(_1863_),
    .A3(_1960_),
    .B1(_1971_),
    .Y(_1972_));
 sky130_fd_sc_hd__mux2i_1 _5660_ (.A0(net764),
    .A1(net763),
    .S(net744),
    .Y(_1973_));
 sky130_fd_sc_hd__mux2i_1 _5661_ (.A0(_1897_),
    .A1(_1973_),
    .S(net742),
    .Y(_1974_));
 sky130_fd_sc_hd__mux2i_2 _5662_ (.A0(_1203_),
    .A1(net760),
    .S(net744),
    .Y(_1975_));
 sky130_fd_sc_hd__mux2_1 _5663_ (.A0(_1899_),
    .A1(_1975_),
    .S(net742),
    .X(_1976_));
 sky130_fd_sc_hd__nor2_1 _5664_ (.A(net740),
    .B(_1976_),
    .Y(_1977_));
 sky130_fd_sc_hd__a21oi_1 _5665_ (.A1(net740),
    .A2(_1974_),
    .B1(_1977_),
    .Y(_1978_));
 sky130_fd_sc_hd__nor2_4 _5666_ (.A(net747),
    .B(_1863_),
    .Y(_1979_));
 sky130_fd_sc_hd__a22oi_1 _5667_ (.A1(net747),
    .A2(_1972_),
    .B1(_1978_),
    .B2(_1979_),
    .Y(_1980_));
 sky130_fd_sc_hd__nor2_1 _5668_ (.A(net741),
    .B(_1980_),
    .Y(_1981_));
 sky130_fd_sc_hd__xnor2_1 _5669_ (.A(_3187_[0]),
    .B(_3437_[0]),
    .Y(_1982_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_42 ();
 sky130_fd_sc_hd__inv_1 _5671_ (.A(_3437_[0]),
    .Y(_1984_));
 sky130_fd_sc_hd__mux2i_1 _5672_ (.A0(_1984_),
    .A1(_3440_[0]),
    .S(net5),
    .Y(_1985_));
 sky130_fd_sc_hd__a22oi_1 _5673_ (.A1(_3436_[0]),
    .A2(net774),
    .B1(net773),
    .B2(_1985_),
    .Y(_1986_));
 sky130_fd_sc_hd__o211ai_1 _5674_ (.A1(_1731_),
    .A2(_1982_),
    .B1(_1986_),
    .C1(_1716_),
    .Y(_1987_));
 sky130_fd_sc_hd__o31a_1 _5675_ (.A1(_1716_),
    .A2(_1981_),
    .A3(_1952_),
    .B1(_1987_),
    .X(net88));
 sky130_fd_sc_hd__a22oi_2 _5676_ (.A1(_0122_),
    .A2(_0150_),
    .B1(_0237_),
    .B2(_1810_),
    .Y(_3184_[0]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_41 ();
 sky130_fd_sc_hd__mux2i_1 _5678_ (.A0(_1742_),
    .A1(_3432_[0]),
    .S(net5),
    .Y(_1989_));
 sky130_fd_sc_hd__nand2_1 _5679_ (.A(_3443_[0]),
    .B(_3437_[0]),
    .Y(_1990_));
 sky130_fd_sc_hd__a221o_4 _5680_ (.A1(_0122_),
    .A2(_0150_),
    .B1(_0237_),
    .B2(net742),
    .C1(_1990_),
    .X(_1991_));
 sky130_fd_sc_hd__a21oi_2 _5681_ (.A1(net246),
    .A2(_3442_[0]),
    .B1(_3436_[0]),
    .Y(_1992_));
 sky130_fd_sc_hd__nand2_2 _5682_ (.A(_1992_),
    .B(_1991_),
    .Y(_1993_));
 sky130_fd_sc_hd__xnor2_1 _5683_ (.A(_1742_),
    .B(_1993_),
    .Y(_1994_));
 sky130_fd_sc_hd__a222oi_1 _5684_ (.A1(_3428_[0]),
    .A2(net774),
    .B1(net773),
    .B2(_1989_),
    .C1(_1994_),
    .C2(_1727_),
    .Y(_1995_));
 sky130_fd_sc_hd__nand2_2 _5685_ (.A(net751),
    .B(_1699_),
    .Y(_1996_));
 sky130_fd_sc_hd__a211oi_2 _5686_ (.A1(_0237_),
    .A2(net751),
    .B1(_1966_),
    .C1(net768),
    .Y(_1997_));
 sky130_fd_sc_hd__a31oi_4 _5687_ (.A1(net768),
    .A2(_1968_),
    .A3(_1996_),
    .B1(_1997_),
    .Y(_1998_));
 sky130_fd_sc_hd__inv_6 _5688_ (.A(_3374_[0]),
    .Y(_3370_[0]));
 sky130_fd_sc_hd__nand2_1 _5689_ (.A(net768),
    .B(net758),
    .Y(_1999_));
 sky130_fd_sc_hd__o21ai_2 _5690_ (.A1(net768),
    .A2(_3370_[0]),
    .B1(_1999_),
    .Y(_2000_));
 sky130_fd_sc_hd__nor2_1 _5691_ (.A(net751),
    .B(_1906_),
    .Y(_2001_));
 sky130_fd_sc_hd__a21oi_2 _5692_ (.A1(net751),
    .A2(_2000_),
    .B1(_2001_),
    .Y(_2002_));
 sky130_fd_sc_hd__nand2_1 _5693_ (.A(net751),
    .B(_1905_),
    .Y(_2003_));
 sky130_fd_sc_hd__o211ai_1 _5694_ (.A1(net751),
    .A2(_1909_),
    .B1(_2003_),
    .C1(net737),
    .Y(_2004_));
 sky130_fd_sc_hd__o211ai_1 _5695_ (.A1(net737),
    .A2(_2002_),
    .B1(_2004_),
    .C1(net778),
    .Y(_2005_));
 sky130_fd_sc_hd__o31ai_1 _5696_ (.A1(net740),
    .A2(net778),
    .A3(_1998_),
    .B1(_2005_),
    .Y(_2006_));
 sky130_fd_sc_hd__mux2i_2 _5697_ (.A0(_1855_),
    .A1(_1973_),
    .S(net769),
    .Y(_2007_));
 sky130_fd_sc_hd__mux2i_2 _5698_ (.A0(_1808_),
    .A1(_1975_),
    .S(net769),
    .Y(_2008_));
 sky130_fd_sc_hd__mux2i_2 _5699_ (.A0(_2007_),
    .A1(_2008_),
    .S(net737),
    .Y(_2009_));
 sky130_fd_sc_hd__a221o_1 _5700_ (.A1(net747),
    .A2(_2006_),
    .B1(_2009_),
    .B2(_1979_),
    .C1(net741),
    .X(_2010_));
 sky130_fd_sc_hd__nand2_8 _5701_ (.A(net816),
    .B(net778),
    .Y(_2011_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_39 ();
 sky130_fd_sc_hd__mux2i_2 _5704_ (.A0(_1848_),
    .A1(_1933_),
    .S(net770),
    .Y(_2014_));
 sky130_fd_sc_hd__mux2i_4 _5705_ (.A0(_1852_),
    .A1(_1935_),
    .S(net770),
    .Y(_2015_));
 sky130_fd_sc_hd__mux2i_2 _5706_ (.A0(_2014_),
    .A1(_2015_),
    .S(_1821_),
    .Y(_2016_));
 sky130_fd_sc_hd__mux2i_4 _5707_ (.A0(_1845_),
    .A1(_1939_),
    .S(net771),
    .Y(_2017_));
 sky130_fd_sc_hd__o21ai_2 _5708_ (.A1(_0313_),
    .A2(net739),
    .B1(net752),
    .Y(_2018_));
 sky130_fd_sc_hd__a21oi_1 _5709_ (.A1(net739),
    .A2(_2017_),
    .B1(_2018_),
    .Y(_2019_));
 sky130_fd_sc_hd__a21oi_2 _5710_ (.A1(_1803_),
    .A2(_2016_),
    .B1(_2019_),
    .Y(_2020_));
 sky130_fd_sc_hd__nor2_1 _5711_ (.A(net752),
    .B(_2016_),
    .Y(_2021_));
 sky130_fd_sc_hd__nor3_4 _5712_ (.A(net742),
    .B(_0314_),
    .C(net751),
    .Y(_2022_));
 sky130_fd_sc_hd__nor2_1 _5713_ (.A(_1821_),
    .B(_2022_),
    .Y(_2023_));
 sky130_fd_sc_hd__a21oi_2 _5714_ (.A1(_2017_),
    .A2(net739),
    .B1(_2023_),
    .Y(_2024_));
 sky130_fd_sc_hd__nor2_1 _5715_ (.A(_1803_),
    .B(_2024_),
    .Y(_2025_));
 sky130_fd_sc_hd__or4_4 _5716_ (.A(net816),
    .B(_1863_),
    .C(_2021_),
    .D(_2025_),
    .X(_2026_));
 sky130_fd_sc_hd__o211ai_1 _5717_ (.A1(_2011_),
    .A2(_2020_),
    .B1(net741),
    .C1(_2026_),
    .Y(_2027_));
 sky130_fd_sc_hd__a21oi_2 _5718_ (.A1(_2010_),
    .A2(_2027_),
    .B1(_1716_),
    .Y(_2028_));
 sky130_fd_sc_hd__a21oi_2 _5719_ (.A1(_1716_),
    .A2(_1995_),
    .B1(_2028_),
    .Y(net91));
 sky130_fd_sc_hd__nor4_1 _5720_ (.A(net799),
    .B(_1713_),
    .C(_1714_),
    .D(_1715_),
    .Y(_2029_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_36 ();
 sky130_fd_sc_hd__nand2_4 _5724_ (.A(net816),
    .B(_0313_),
    .Y(_2033_));
 sky130_fd_sc_hd__nand2_2 _5725_ (.A(net738),
    .B(_1847_),
    .Y(_2034_));
 sky130_fd_sc_hd__o21ai_2 _5726_ (.A1(net738),
    .A2(_2033_),
    .B1(_2034_),
    .Y(_2035_));
 sky130_fd_sc_hd__mux2i_1 _5727_ (.A0(_1850_),
    .A1(_1854_),
    .S(net738),
    .Y(_2036_));
 sky130_fd_sc_hd__nand2_1 _5728_ (.A(net749),
    .B(_2036_),
    .Y(_2037_));
 sky130_fd_sc_hd__o2111ai_4 _5729_ (.A1(net749),
    .A2(_2035_),
    .B1(_2037_),
    .C1(net778),
    .D1(net268),
    .Y(_2038_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_35 ();
 sky130_fd_sc_hd__nand2_1 _5731_ (.A(_1968_),
    .B(_1996_),
    .Y(_2040_));
 sky130_fd_sc_hd__mux2i_1 _5732_ (.A0(net753),
    .A1(_3438_[0]),
    .S(net751),
    .Y(_2041_));
 sky130_fd_sc_hd__nand2_1 _5733_ (.A(net768),
    .B(_2041_),
    .Y(_2042_));
 sky130_fd_sc_hd__o211a_1 _5734_ (.A1(net768),
    .A2(_2040_),
    .B1(_2042_),
    .C1(net737),
    .X(_2043_));
 sky130_fd_sc_hd__a21oi_2 _5735_ (.A1(net740),
    .A2(_1869_),
    .B1(_2043_),
    .Y(_2044_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_34 ();
 sky130_fd_sc_hd__nand2_1 _5737_ (.A(net740),
    .B(_1820_),
    .Y(_2046_));
 sky130_fd_sc_hd__o211a_1 _5738_ (.A1(net740),
    .A2(_1831_),
    .B1(_2046_),
    .C1(net778),
    .X(_2047_));
 sky130_fd_sc_hd__a21oi_1 _5739_ (.A1(_1863_),
    .A2(_2044_),
    .B1(_2047_),
    .Y(_2048_));
 sky130_fd_sc_hd__nor2_1 _5740_ (.A(net737),
    .B(_1857_),
    .Y(_2049_));
 sky130_fd_sc_hd__a21oi_1 _5741_ (.A1(net737),
    .A2(_1813_),
    .B1(_2049_),
    .Y(_2050_));
 sky130_fd_sc_hd__nand2_1 _5742_ (.A(_1979_),
    .B(_2050_),
    .Y(_2051_));
 sky130_fd_sc_hd__o21ai_0 _5743_ (.A1(net752),
    .A2(_2048_),
    .B1(_2051_),
    .Y(_2052_));
 sky130_fd_sc_hd__nand2_2 _5744_ (.A(net750),
    .B(_2052_),
    .Y(_2053_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_33 ();
 sky130_fd_sc_hd__o22ai_1 _5746_ (.A1(net5),
    .A2(_1721_),
    .B1(_1731_),
    .B2(net233),
    .Y(_2055_));
 sky130_fd_sc_hd__nand2_1 _5747_ (.A(_1727_),
    .B(net233),
    .Y(_2056_));
 sky130_fd_sc_hd__nand2_1 _5748_ (.A(_3420_[0]),
    .B(net774),
    .Y(_2057_));
 sky130_fd_sc_hd__o221ai_2 _5749_ (.A1(_3424_[0]),
    .A2(_1712_),
    .B1(_2056_),
    .B2(_3421_[0]),
    .C1(_2057_),
    .Y(_2058_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_32 ();
 sky130_fd_sc_hd__a211oi_2 _5751_ (.A1(_3421_[0]),
    .A2(_2055_),
    .B1(net777),
    .C1(_2058_),
    .Y(_2060_));
 sky130_fd_sc_hd__a31oi_4 _5752_ (.A1(net777),
    .A2(_2038_),
    .A3(_2053_),
    .B1(_2060_),
    .Y(net92));
 sky130_fd_sc_hd__a21o_1 _5753_ (.A1(_1993_),
    .A2(_3429_[0]),
    .B1(_3428_[0]),
    .X(_2061_));
 sky130_fd_sc_hd__a211oi_2 _5754_ (.A1(_2061_),
    .A2(_3421_[0]),
    .B1(_3420_[0]),
    .C1(_3413_[0]),
    .Y(_2062_));
 sky130_fd_sc_hd__nand3_1 _5755_ (.A(_3413_[0]),
    .B(_3421_[0]),
    .C(_3429_[0]),
    .Y(_2063_));
 sky130_fd_sc_hd__a21oi_4 _5756_ (.A1(_1991_),
    .A2(_1992_),
    .B1(_2063_),
    .Y(_2064_));
 sky130_fd_sc_hd__a21oi_1 _5757_ (.A1(_3428_[0]),
    .A2(_3421_[0]),
    .B1(_3420_[0]),
    .Y(_2065_));
 sky130_fd_sc_hd__nor2_1 _5758_ (.A(_1741_),
    .B(_2065_),
    .Y(_2066_));
 sky130_fd_sc_hd__nor3_1 _5759_ (.A(_2066_),
    .B(_2064_),
    .C(_2062_),
    .Y(_2067_));
 sky130_fd_sc_hd__mux2i_1 _5760_ (.A0(_1741_),
    .A1(_3416_[0]),
    .S(net5),
    .Y(_2068_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_31 ();
 sky130_fd_sc_hd__a222oi_1 _5762_ (.A1(_3412_[0]),
    .A2(net774),
    .B1(_1727_),
    .B2(_2067_),
    .C1(_2068_),
    .C2(net773),
    .Y(_2070_));
 sky130_fd_sc_hd__nand3_4 _5763_ (.A(net743),
    .B(_1910_),
    .C(_1922_),
    .Y(_2071_));
 sky130_fd_sc_hd__o21ai_2 _5764_ (.A1(_3426_[0]),
    .A2(net743),
    .B1(_1827_),
    .Y(_2072_));
 sky130_fd_sc_hd__nand2_1 _5765_ (.A(net742),
    .B(_2041_),
    .Y(_2073_));
 sky130_fd_sc_hd__o21a_4 _5766_ (.A1(net742),
    .A2(_2072_),
    .B1(_2073_),
    .X(_2074_));
 sky130_fd_sc_hd__mux2i_2 _5767_ (.A0(_2071_),
    .A1(_2074_),
    .S(net737),
    .Y(_2075_));
 sky130_fd_sc_hd__nand2_1 _5768_ (.A(net737),
    .B(_1907_),
    .Y(_2076_));
 sky130_fd_sc_hd__o211ai_1 _5769_ (.A1(net737),
    .A2(_1900_),
    .B1(_2076_),
    .C1(net778),
    .Y(_2077_));
 sky130_fd_sc_hd__o21ai_0 _5770_ (.A1(net778),
    .A2(_2075_),
    .B1(_2077_),
    .Y(_2078_));
 sky130_fd_sc_hd__mux2i_1 _5771_ (.A0(_1898_),
    .A1(_1891_),
    .S(net740),
    .Y(_2079_));
 sky130_fd_sc_hd__nand2_1 _5772_ (.A(_1979_),
    .B(_2079_),
    .Y(_2080_));
 sky130_fd_sc_hd__o21ai_2 _5773_ (.A1(net752),
    .A2(_2078_),
    .B1(_2080_),
    .Y(_2081_));
 sky130_fd_sc_hd__nand2_2 _5774_ (.A(net740),
    .B(_1879_),
    .Y(_2082_));
 sky130_fd_sc_hd__nand2_1 _5775_ (.A(net739),
    .B(_1889_),
    .Y(_2083_));
 sky130_fd_sc_hd__nand2_2 _5776_ (.A(_2082_),
    .B(_2083_),
    .Y(_2084_));
 sky130_fd_sc_hd__nor2_4 _5777_ (.A(net749),
    .B(net740),
    .Y(_2085_));
 sky130_fd_sc_hd__nand2b_2 _5778_ (.A_N(net307),
    .B(_2085_),
    .Y(_2086_));
 sky130_fd_sc_hd__a21oi_2 _5779_ (.A1(net739),
    .A2(_1885_),
    .B1(_2018_),
    .Y(_2087_));
 sky130_fd_sc_hd__nand2_1 _5780_ (.A(net816),
    .B(_2087_),
    .Y(_2088_));
 sky130_fd_sc_hd__o221ai_2 _5781_ (.A1(net752),
    .A2(_2084_),
    .B1(_2086_),
    .B2(net816),
    .C1(_2088_),
    .Y(_2089_));
 sky130_fd_sc_hd__nor2_2 _5782_ (.A(net750),
    .B(_1863_),
    .Y(_2090_));
 sky130_fd_sc_hd__a221oi_4 _5783_ (.A1(net750),
    .A2(_2081_),
    .B1(_2089_),
    .B2(_2090_),
    .C1(_1716_),
    .Y(_2091_));
 sky130_fd_sc_hd__a21oi_2 _5784_ (.A1(_1716_),
    .A2(_2070_),
    .B1(_2091_),
    .Y(net93));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_30 ();
 sky130_fd_sc_hd__nand2_1 _5786_ (.A(_3404_[0]),
    .B(net774),
    .Y(_2093_));
 sky130_fd_sc_hd__o21ai_0 _5787_ (.A1(_3408_[0]),
    .A2(_1712_),
    .B1(_2093_),
    .Y(_2094_));
 sky130_fd_sc_hd__o22a_1 _5788_ (.A1(net5),
    .A2(_1721_),
    .B1(_1731_),
    .B2(_1746_),
    .X(_2095_));
 sky130_fd_sc_hd__a21oi_1 _5789_ (.A1(_1727_),
    .A2(net238),
    .B1(_3405_[0]),
    .Y(_2096_));
 sky130_fd_sc_hd__a21oi_1 _5790_ (.A1(_3405_[0]),
    .A2(_2095_),
    .B1(_2096_),
    .Y(_2097_));
 sky130_fd_sc_hd__nand2_1 _5791_ (.A(net740),
    .B(_1976_),
    .Y(_2098_));
 sky130_fd_sc_hd__o21a_1 _5792_ (.A1(net740),
    .A2(_1960_),
    .B1(_2098_),
    .X(_2099_));
 sky130_fd_sc_hd__mux2i_1 _5793_ (.A0(net755),
    .A1(net753),
    .S(net751),
    .Y(_2100_));
 sky130_fd_sc_hd__nand2_1 _5794_ (.A(net768),
    .B(_2100_),
    .Y(_2101_));
 sky130_fd_sc_hd__o21ai_2 _5795_ (.A1(net768),
    .A2(_2072_),
    .B1(_2101_),
    .Y(_2102_));
 sky130_fd_sc_hd__nand2_1 _5796_ (.A(net740),
    .B(_1964_),
    .Y(_2103_));
 sky130_fd_sc_hd__o211ai_1 _5797_ (.A1(net740),
    .A2(_2102_),
    .B1(_2103_),
    .C1(_1863_),
    .Y(_2104_));
 sky130_fd_sc_hd__o21ai_0 _5798_ (.A1(_1863_),
    .A2(_2099_),
    .B1(_2104_),
    .Y(_2105_));
 sky130_fd_sc_hd__nor2_1 _5799_ (.A(net738),
    .B(_1936_),
    .Y(_2106_));
 sky130_fd_sc_hd__a21oi_1 _5800_ (.A1(net737),
    .A2(_1974_),
    .B1(_2106_),
    .Y(_2107_));
 sky130_fd_sc_hd__a22oi_1 _5801_ (.A1(_2105_),
    .A2(net747),
    .B1(_2107_),
    .B2(_1979_),
    .Y(_2108_));
 sky130_fd_sc_hd__nor2_1 _5802_ (.A(net739),
    .B(_1940_),
    .Y(_2109_));
 sky130_fd_sc_hd__nor2_1 _5803_ (.A(net740),
    .B(_1934_),
    .Y(_2110_));
 sky130_fd_sc_hd__nor2_2 _5804_ (.A(_2109_),
    .B(_2110_),
    .Y(_2111_));
 sky130_fd_sc_hd__nand2_2 _5805_ (.A(net739),
    .B(net746),
    .Y(_2112_));
 sky130_fd_sc_hd__a32oi_1 _5806_ (.A1(net816),
    .A2(_0313_),
    .A3(_2112_),
    .B1(_1942_),
    .B2(net739),
    .Y(_2113_));
 sky130_fd_sc_hd__nor2_1 _5807_ (.A(net748),
    .B(_2113_),
    .Y(_2114_));
 sky130_fd_sc_hd__a21oi_2 _5808_ (.A1(net748),
    .A2(_2111_),
    .B1(_2114_),
    .Y(_2115_));
 sky130_fd_sc_hd__o221ai_2 _5809_ (.A1(net741),
    .A2(_2108_),
    .B1(_2115_),
    .B2(_1951_),
    .C1(net777),
    .Y(_2116_));
 sky130_fd_sc_hd__o31a_1 _5810_ (.A1(net777),
    .A2(_2094_),
    .A3(_2097_),
    .B1(_2116_),
    .X(net94));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_29 ();
 sky130_fd_sc_hd__nor2_1 _5812_ (.A(_3412_[0]),
    .B(_2066_),
    .Y(_2118_));
 sky130_fd_sc_hd__nand2b_1 _5813_ (.A_N(_2064_),
    .B(_2118_),
    .Y(_2119_));
 sky130_fd_sc_hd__a21oi_1 _5814_ (.A1(_3405_[0]),
    .A2(_2119_),
    .B1(_3404_[0]),
    .Y(_2120_));
 sky130_fd_sc_hd__xnor2_1 _5815_ (.A(_3397_[0]),
    .B(_2120_),
    .Y(_2121_));
 sky130_fd_sc_hd__nand2_1 _5816_ (.A(_1727_),
    .B(_2121_),
    .Y(_2122_));
 sky130_fd_sc_hd__nand2_1 _5817_ (.A(_3396_[0]),
    .B(net774),
    .Y(_2123_));
 sky130_fd_sc_hd__inv_2 _5818_ (.A(_3397_[0]),
    .Y(_2124_));
 sky130_fd_sc_hd__mux2i_1 _5819_ (.A0(_2124_),
    .A1(_3400_[0]),
    .S(net5),
    .Y(_2125_));
 sky130_fd_sc_hd__a21oi_2 _5820_ (.A1(net773),
    .A2(_2125_),
    .B1(net777),
    .Y(_2126_));
 sky130_fd_sc_hd__mux2i_4 _5821_ (.A0(_2017_),
    .A1(_2014_),
    .S(_1821_),
    .Y(_2127_));
 sky130_fd_sc_hd__nor2_1 _5822_ (.A(net816),
    .B(net740),
    .Y(_2128_));
 sky130_fd_sc_hd__nand2_1 _5823_ (.A(_2022_),
    .B(_2128_),
    .Y(_2129_));
 sky130_fd_sc_hd__a31oi_1 _5824_ (.A1(net752),
    .A2(_2033_),
    .A3(_2129_),
    .B1(_1863_),
    .Y(_2130_));
 sky130_fd_sc_hd__o21ai_1 _5825_ (.A1(net752),
    .A2(_2127_),
    .B1(_2130_),
    .Y(_2131_));
 sky130_fd_sc_hd__nand2_1 _5826_ (.A(net740),
    .B(_1998_),
    .Y(_2132_));
 sky130_fd_sc_hd__mux2i_1 _5827_ (.A0(net756),
    .A1(net754),
    .S(net751),
    .Y(_2133_));
 sky130_fd_sc_hd__mux2i_2 _5828_ (.A0(_2100_),
    .A1(_2133_),
    .S(net339),
    .Y(_2134_));
 sky130_fd_sc_hd__nand2_1 _5829_ (.A(net737),
    .B(_2134_),
    .Y(_2135_));
 sky130_fd_sc_hd__nand2_4 _5830_ (.A(_2132_),
    .B(_2135_),
    .Y(_2136_));
 sky130_fd_sc_hd__nand2_1 _5831_ (.A(net740),
    .B(_2008_),
    .Y(_2137_));
 sky130_fd_sc_hd__o211ai_1 _5832_ (.A1(net740),
    .A2(_2002_),
    .B1(_2137_),
    .C1(net778),
    .Y(_2138_));
 sky130_fd_sc_hd__o21ai_0 _5833_ (.A1(net778),
    .A2(_2136_),
    .B1(_2138_),
    .Y(_2139_));
 sky130_fd_sc_hd__mux2i_1 _5834_ (.A0(_2007_),
    .A1(_2015_),
    .S(net740),
    .Y(_2140_));
 sky130_fd_sc_hd__a221oi_1 _5835_ (.A1(net747),
    .A2(_2139_),
    .B1(_2140_),
    .B2(_1979_),
    .C1(net268),
    .Y(_2141_));
 sky130_fd_sc_hd__a21o_4 _5836_ (.A1(net268),
    .A2(_2131_),
    .B1(_2141_),
    .X(_2142_));
 sky130_fd_sc_hd__a32oi_4 _5837_ (.A1(_2122_),
    .A2(_2123_),
    .A3(_2126_),
    .B1(_2142_),
    .B2(net777),
    .Y(net95));
 sky130_fd_sc_hd__inv_1 _5838_ (.A(net757),
    .Y(_3386_[0]));
 sky130_fd_sc_hd__nor2_1 _5839_ (.A(net749),
    .B(_2033_),
    .Y(_2143_));
 sky130_fd_sc_hd__nor2_1 _5840_ (.A(net752),
    .B(_1851_),
    .Y(_2144_));
 sky130_fd_sc_hd__o21a_4 _5841_ (.A1(_2143_),
    .A2(_2144_),
    .B1(net778),
    .X(_2145_));
 sky130_fd_sc_hd__o211ai_1 _5842_ (.A1(net768),
    .A2(_2040_),
    .B1(_2042_),
    .C1(net740),
    .Y(_2146_));
 sky130_fd_sc_hd__mux2i_1 _5843_ (.A0(net757),
    .A1(net755),
    .S(net751),
    .Y(_2147_));
 sky130_fd_sc_hd__mux2i_1 _5844_ (.A0(_2133_),
    .A1(_2147_),
    .S(net339),
    .Y(_2148_));
 sky130_fd_sc_hd__nand2_1 _5845_ (.A(net737),
    .B(_2148_),
    .Y(_2149_));
 sky130_fd_sc_hd__nand2_1 _5846_ (.A(net752),
    .B(net737),
    .Y(_2150_));
 sky130_fd_sc_hd__nor2_1 _5847_ (.A(_1869_),
    .B(_2150_),
    .Y(_2151_));
 sky130_fd_sc_hd__a31oi_1 _5848_ (.A1(net747),
    .A2(_2146_),
    .A3(_2149_),
    .B1(_2151_),
    .Y(_2152_));
 sky130_fd_sc_hd__nor2_1 _5849_ (.A(net749),
    .B(_1859_),
    .Y(_2153_));
 sky130_fd_sc_hd__a211oi_1 _5850_ (.A1(net747),
    .A2(_1824_),
    .B1(_2153_),
    .C1(_1863_),
    .Y(_2154_));
 sky130_fd_sc_hd__a211oi_2 _5851_ (.A1(_1863_),
    .A2(_2152_),
    .B1(_2154_),
    .C1(net268),
    .Y(_2155_));
 sky130_fd_sc_hd__a21oi_4 _5852_ (.A1(net268),
    .A2(_2145_),
    .B1(_2155_),
    .Y(_2156_));
 sky130_fd_sc_hd__nor2_1 _5853_ (.A(_1747_),
    .B(_2124_),
    .Y(_2157_));
 sky130_fd_sc_hd__nor2_1 _5854_ (.A(_3396_[0]),
    .B(_2157_),
    .Y(_2158_));
 sky130_fd_sc_hd__nand2_1 _5855_ (.A(_1727_),
    .B(_2158_),
    .Y(_2159_));
 sky130_fd_sc_hd__o21ai_2 _5856_ (.A1(net5),
    .A2(_1721_),
    .B1(_2159_),
    .Y(_2160_));
 sky130_fd_sc_hd__nor3_1 _5857_ (.A(_3389_[0]),
    .B(_1731_),
    .C(_2158_),
    .Y(_2161_));
 sky130_fd_sc_hd__nand2_1 _5858_ (.A(_3388_[0]),
    .B(net774),
    .Y(_2162_));
 sky130_fd_sc_hd__o21ai_0 _5859_ (.A1(_3392_[0]),
    .A2(_1712_),
    .B1(_2162_),
    .Y(_2163_));
 sky130_fd_sc_hd__a2111oi_4 _5860_ (.A1(_2160_),
    .A2(_3389_[0]),
    .B1(_2163_),
    .C1(net777),
    .D1(_2161_),
    .Y(_2164_));
 sky130_fd_sc_hd__a21oi_4 _5861_ (.A1(net777),
    .A2(_2156_),
    .B1(_2164_),
    .Y(net96));
 sky130_fd_sc_hd__inv_4 _5862_ (.A(_1364_),
    .Y(_3378_[0]));
 sky130_fd_sc_hd__inv_1 _5863_ (.A(_3381_[0]),
    .Y(_2165_));
 sky130_fd_sc_hd__nor4b_4 _5864_ (.A(_3404_[0]),
    .B(_3396_[0]),
    .C(_2064_),
    .D_N(_2118_),
    .Y(_2166_));
 sky130_fd_sc_hd__nor2_1 _5865_ (.A(_3404_[0]),
    .B(_3405_[0]),
    .Y(_2167_));
 sky130_fd_sc_hd__nor2_1 _5866_ (.A(_2124_),
    .B(_2167_),
    .Y(_2168_));
 sky130_fd_sc_hd__o21ai_2 _5867_ (.A1(_3396_[0]),
    .A2(_2168_),
    .B1(_3389_[0]),
    .Y(_2169_));
 sky130_fd_sc_hd__o21bai_2 _5868_ (.A1(_2169_),
    .A2(_2166_),
    .B1_N(_3388_[0]),
    .Y(_2170_));
 sky130_fd_sc_hd__xnor2_1 _5869_ (.A(_2165_),
    .B(net376),
    .Y(_2171_));
 sky130_fd_sc_hd__mux2i_1 _5870_ (.A0(_2165_),
    .A1(_3384_[0]),
    .S(net5),
    .Y(_2172_));
 sky130_fd_sc_hd__a222oi_1 _5871_ (.A1(_3380_[0]),
    .A2(net774),
    .B1(_2171_),
    .B2(_1727_),
    .C1(_2172_),
    .C2(net773),
    .Y(_2173_));
 sky130_fd_sc_hd__nand2_1 _5872_ (.A(net749),
    .B(_1902_),
    .Y(_2174_));
 sky130_fd_sc_hd__nand2_1 _5873_ (.A(net752),
    .B(_1893_),
    .Y(_2175_));
 sky130_fd_sc_hd__nand4_1 _5874_ (.A(net750),
    .B(net778),
    .C(_2174_),
    .D(_2175_),
    .Y(_2176_));
 sky130_fd_sc_hd__mux2i_2 _5875_ (.A0(net758),
    .A1(net756),
    .S(net751),
    .Y(_2177_));
 sky130_fd_sc_hd__mux2i_4 _5876_ (.A0(_2147_),
    .A1(_2177_),
    .S(net339),
    .Y(_2178_));
 sky130_fd_sc_hd__mux2i_2 _5877_ (.A0(_2074_),
    .A1(_2178_),
    .S(net737),
    .Y(_2179_));
 sky130_fd_sc_hd__a221o_1 _5878_ (.A1(_1923_),
    .A2(_2085_),
    .B1(_2179_),
    .B2(net749),
    .C1(_1870_),
    .X(_2180_));
 sky130_fd_sc_hd__nand2_1 _5879_ (.A(_0313_),
    .B(net752),
    .Y(_2181_));
 sky130_fd_sc_hd__a21boi_0 _5880_ (.A1(_1803_),
    .A2(_1886_),
    .B1_N(_2181_),
    .Y(_2182_));
 sky130_fd_sc_hd__nor3_4 _5881_ (.A(net816),
    .B(net752),
    .C(_1863_),
    .Y(_2183_));
 sky130_fd_sc_hd__a21oi_1 _5882_ (.A1(_1882_),
    .A2(_2183_),
    .B1(net750),
    .Y(_2184_));
 sky130_fd_sc_hd__o21ai_2 _5883_ (.A1(_2011_),
    .A2(_2182_),
    .B1(_2184_),
    .Y(_2185_));
 sky130_fd_sc_hd__nand4_1 _5884_ (.A(net777),
    .B(_2176_),
    .C(_2185_),
    .D(_2180_),
    .Y(_2186_));
 sky130_fd_sc_hd__o21ai_2 _5885_ (.A1(net777),
    .A2(_2173_),
    .B1(_2186_),
    .Y(net97));
 sky130_fd_sc_hd__mux2i_1 _5886_ (.A0(net759),
    .A1(net757),
    .S(net751),
    .Y(_2187_));
 sky130_fd_sc_hd__mux2i_1 _5887_ (.A0(_2177_),
    .A1(_2187_),
    .S(net339),
    .Y(_2188_));
 sky130_fd_sc_hd__nand2_1 _5888_ (.A(net737),
    .B(_2188_),
    .Y(_2189_));
 sky130_fd_sc_hd__o21ai_2 _5889_ (.A1(net737),
    .A2(_2102_),
    .B1(_2189_),
    .Y(_2190_));
 sky130_fd_sc_hd__o221ai_2 _5890_ (.A1(net313),
    .A2(_2150_),
    .B1(_2190_),
    .B2(net752),
    .C1(_1863_),
    .Y(_2191_));
 sky130_fd_sc_hd__nor2_1 _5891_ (.A(net747),
    .B(_1937_),
    .Y(_2192_));
 sky130_fd_sc_hd__a211o_1 _5892_ (.A1(net747),
    .A2(_1978_),
    .B1(_2192_),
    .C1(_1863_),
    .X(_2193_));
 sky130_fd_sc_hd__nand3_2 _5893_ (.A(net750),
    .B(_2191_),
    .C(_2193_),
    .Y(_2194_));
 sky130_fd_sc_hd__o21ai_1 _5894_ (.A1(net752),
    .A2(_1946_),
    .B1(_2181_),
    .Y(_2195_));
 sky130_fd_sc_hd__nor2_1 _5895_ (.A(net816),
    .B(net752),
    .Y(_2196_));
 sky130_fd_sc_hd__a22oi_2 _5896_ (.A1(net816),
    .A2(_2195_),
    .B1(_2196_),
    .B2(_1943_),
    .Y(_2197_));
 sky130_fd_sc_hd__or3_4 _5897_ (.A(_1801_),
    .B(_1863_),
    .C(_2197_),
    .X(_2198_));
 sky130_fd_sc_hd__o21ai_0 _5898_ (.A1(_1747_),
    .A2(_1748_),
    .B1(_1750_),
    .Y(_2199_));
 sky130_fd_sc_hd__nor2_1 _5899_ (.A(_2199_),
    .B(_3380_[0]),
    .Y(_2200_));
 sky130_fd_sc_hd__xnor2_1 _5900_ (.A(_2200_),
    .B(_3373_[0]),
    .Y(_2201_));
 sky130_fd_sc_hd__inv_1 _5901_ (.A(_3373_[0]),
    .Y(_2202_));
 sky130_fd_sc_hd__mux2i_1 _5902_ (.A0(_2202_),
    .A1(_3376_[0]),
    .S(net5),
    .Y(_2203_));
 sky130_fd_sc_hd__a221o_1 _5903_ (.A1(_3372_[0]),
    .A2(net774),
    .B1(net773),
    .B2(_2203_),
    .C1(net777),
    .X(_2204_));
 sky130_fd_sc_hd__a21oi_2 _5904_ (.A1(_2201_),
    .A2(_1727_),
    .B1(_2204_),
    .Y(_2205_));
 sky130_fd_sc_hd__a31oi_4 _5905_ (.A1(net777),
    .A2(_2198_),
    .A3(_2194_),
    .B1(_2205_),
    .Y(net67));
 sky130_fd_sc_hd__clkinv_1 _5906_ (.A(_3366_[0]),
    .Y(_3362_[0]));
 sky130_fd_sc_hd__a21o_1 _5907_ (.A1(_3373_[0]),
    .A2(_3380_[0]),
    .B1(_3372_[0]),
    .X(_2206_));
 sky130_fd_sc_hd__a31oi_2 _5908_ (.A1(_2170_),
    .A2(_3381_[0]),
    .A3(_3373_[0]),
    .B1(_2206_),
    .Y(_2207_));
 sky130_fd_sc_hd__xnor2_1 _5909_ (.A(_3365_[0]),
    .B(_2207_),
    .Y(_2208_));
 sky130_fd_sc_hd__mux2i_1 _5910_ (.A0(_1753_),
    .A1(_3368_[0]),
    .S(net5),
    .Y(_2209_));
 sky130_fd_sc_hd__a222oi_1 _5911_ (.A1(_3364_[0]),
    .A2(net774),
    .B1(_1727_),
    .B2(_2208_),
    .C1(_2209_),
    .C2(net773),
    .Y(_2210_));
 sky130_fd_sc_hd__nor2_1 _5912_ (.A(_1803_),
    .B(net298),
    .Y(_2211_));
 sky130_fd_sc_hd__nor2_1 _5913_ (.A(net752),
    .B(_2009_),
    .Y(_2212_));
 sky130_fd_sc_hd__mux2i_1 _5914_ (.A0(net760),
    .A1(net758),
    .S(net751),
    .Y(_2213_));
 sky130_fd_sc_hd__mux2i_2 _5915_ (.A0(_2187_),
    .A1(_2213_),
    .S(net339),
    .Y(_2214_));
 sky130_fd_sc_hd__mux2i_1 _5916_ (.A0(_2134_),
    .A1(_2214_),
    .S(_1821_),
    .Y(_2215_));
 sky130_fd_sc_hd__o21ai_0 _5917_ (.A1(net740),
    .A2(_1998_),
    .B1(net752),
    .Y(_2216_));
 sky130_fd_sc_hd__o211ai_1 _5918_ (.A1(net752),
    .A2(_2215_),
    .B1(_2216_),
    .C1(_1863_),
    .Y(_2217_));
 sky130_fd_sc_hd__o311ai_1 _5919_ (.A1(_1863_),
    .A2(_2211_),
    .A3(_2212_),
    .B1(_2217_),
    .C1(net750),
    .Y(_2218_));
 sky130_fd_sc_hd__a21oi_1 _5920_ (.A1(_1803_),
    .A2(net738),
    .B1(_0313_),
    .Y(_2219_));
 sky130_fd_sc_hd__a211oi_1 _5921_ (.A1(_1921_),
    .A2(_2017_),
    .B1(_2011_),
    .C1(_2219_),
    .Y(_2220_));
 sky130_fd_sc_hd__a21oi_1 _5922_ (.A1(net342),
    .A2(_2183_),
    .B1(_2220_),
    .Y(_2221_));
 sky130_fd_sc_hd__nand2_2 _5923_ (.A(net741),
    .B(_2221_),
    .Y(_2222_));
 sky130_fd_sc_hd__nand3_4 _5924_ (.A(net777),
    .B(_2218_),
    .C(_2222_),
    .Y(_2223_));
 sky130_fd_sc_hd__o21ai_2 _5925_ (.A1(net777),
    .A2(_2210_),
    .B1(_2223_),
    .Y(net68));
 sky130_fd_sc_hd__clkinv_1 _5926_ (.A(net761),
    .Y(_3354_[0]));
 sky130_fd_sc_hd__inv_1 _5927_ (.A(_3357_[0]),
    .Y(_2224_));
 sky130_fd_sc_hd__mux2i_1 _5928_ (.A0(_2224_),
    .A1(_3360_[0]),
    .S(net5),
    .Y(_2225_));
 sky130_fd_sc_hd__nand2_1 _5929_ (.A(net193),
    .B(_1756_),
    .Y(_2226_));
 sky130_fd_sc_hd__xnor2_1 _5930_ (.A(_3357_[0]),
    .B(_2226_),
    .Y(_2227_));
 sky130_fd_sc_hd__a222oi_1 _5931_ (.A1(_3356_[0]),
    .A2(net774),
    .B1(net773),
    .B2(_2225_),
    .C1(_2227_),
    .C2(_1727_),
    .Y(_2228_));
 sky130_fd_sc_hd__mux2i_2 _5932_ (.A0(net761),
    .A1(net759),
    .S(net751),
    .Y(_2229_));
 sky130_fd_sc_hd__mux2i_2 _5933_ (.A0(_2213_),
    .A1(_2229_),
    .S(net769),
    .Y(_2230_));
 sky130_fd_sc_hd__mux2i_1 _5934_ (.A0(_2148_),
    .A1(_2230_),
    .S(net737),
    .Y(_2231_));
 sky130_fd_sc_hd__mux2i_2 _5935_ (.A0(_2044_),
    .A1(_2231_),
    .S(net747),
    .Y(_2232_));
 sky130_fd_sc_hd__nand2_1 _5936_ (.A(net752),
    .B(_2036_),
    .Y(_2233_));
 sky130_fd_sc_hd__o21ai_0 _5937_ (.A1(net752),
    .A2(_2050_),
    .B1(_2233_),
    .Y(_2234_));
 sky130_fd_sc_hd__mux2i_1 _5938_ (.A0(_2232_),
    .A1(_2234_),
    .S(net778),
    .Y(_2235_));
 sky130_fd_sc_hd__nand2_1 _5939_ (.A(_1847_),
    .B(_1921_),
    .Y(_2236_));
 sky130_fd_sc_hd__o21ai_1 _5940_ (.A1(_1921_),
    .A2(_2033_),
    .B1(_2236_),
    .Y(_2237_));
 sky130_fd_sc_hd__a221oi_2 _5941_ (.A1(net750),
    .A2(_2235_),
    .B1(_2237_),
    .B2(_2090_),
    .C1(_1716_),
    .Y(_2238_));
 sky130_fd_sc_hd__a21oi_2 _5942_ (.A1(_2228_),
    .A2(_1716_),
    .B1(_2238_),
    .Y(net69));
 sky130_fd_sc_hd__inv_1 _5943_ (.A(_1203_),
    .Y(_3346_[0]));
 sky130_fd_sc_hd__a21oi_1 _5944_ (.A1(_1921_),
    .A2(_1885_),
    .B1(_2219_),
    .Y(_2239_));
 sky130_fd_sc_hd__nor2b_2 _5945_ (.A(_2011_),
    .B_N(_2239_),
    .Y(_2240_));
 sky130_fd_sc_hd__nand2_1 _5946_ (.A(net739),
    .B(_2183_),
    .Y(_2241_));
 sky130_fd_sc_hd__o21ai_2 _5947_ (.A1(net307),
    .A2(_2241_),
    .B1(net741),
    .Y(_2242_));
 sky130_fd_sc_hd__o21ai_4 _5948_ (.A1(_2240_),
    .A2(_2242_),
    .B1(net777),
    .Y(_2243_));
 sky130_fd_sc_hd__mux2i_2 _5949_ (.A0(_1203_),
    .A1(net760),
    .S(net751),
    .Y(_2244_));
 sky130_fd_sc_hd__mux2i_4 _5950_ (.A0(_2229_),
    .A1(_2244_),
    .S(net769),
    .Y(_2245_));
 sky130_fd_sc_hd__mux2i_4 _5951_ (.A0(_2178_),
    .A1(_2245_),
    .S(net737),
    .Y(_2246_));
 sky130_fd_sc_hd__mux2_4 _5952_ (.A0(_2075_),
    .A1(_2246_),
    .S(net749),
    .X(_2247_));
 sky130_fd_sc_hd__nand2_1 _5953_ (.A(net749),
    .B(_2079_),
    .Y(_2248_));
 sky130_fd_sc_hd__o2111ai_2 _5954_ (.A1(net749),
    .A2(_2084_),
    .B1(_2248_),
    .C1(net778),
    .D1(net750),
    .Y(_2249_));
 sky130_fd_sc_hd__o21ai_4 _5955_ (.A1(_1870_),
    .A2(_2247_),
    .B1(_2249_),
    .Y(_2250_));
 sky130_fd_sc_hd__inv_1 _5956_ (.A(_3349_[0]),
    .Y(_2251_));
 sky130_fd_sc_hd__mux2i_1 _5957_ (.A0(_2251_),
    .A1(_3352_[0]),
    .S(net5),
    .Y(_2252_));
 sky130_fd_sc_hd__nand4_1 _5958_ (.A(_3357_[0]),
    .B(_3365_[0]),
    .C(_3373_[0]),
    .D(_3381_[0]),
    .Y(_2253_));
 sky130_fd_sc_hd__nand2_1 _5959_ (.A(_3365_[0]),
    .B(_2206_),
    .Y(_2254_));
 sky130_fd_sc_hd__a41oi_1 _5960_ (.A1(_3388_[0]),
    .A2(_3365_[0]),
    .A3(_3373_[0]),
    .A4(_3381_[0]),
    .B1(_3364_[0]),
    .Y(_2255_));
 sky130_fd_sc_hd__nand2_1 _5961_ (.A(_2254_),
    .B(_2255_),
    .Y(_2256_));
 sky130_fd_sc_hd__a21oi_1 _5962_ (.A1(_3357_[0]),
    .A2(_2256_),
    .B1(_3356_[0]),
    .Y(_2257_));
 sky130_fd_sc_hd__o31a_1 _5963_ (.A1(_2253_),
    .A2(_2169_),
    .A3(_2166_),
    .B1(_2257_),
    .X(_2258_));
 sky130_fd_sc_hd__xnor2_1 _5964_ (.A(_3349_[0]),
    .B(net702),
    .Y(_2259_));
 sky130_fd_sc_hd__a222oi_1 _5965_ (.A1(_3348_[0]),
    .A2(net774),
    .B1(net773),
    .B2(_2252_),
    .C1(_2259_),
    .C2(_1727_),
    .Y(_2260_));
 sky130_fd_sc_hd__o22ai_4 _5966_ (.A1(_2243_),
    .A2(_2250_),
    .B1(net777),
    .B2(_2260_),
    .Y(net70));
 sky130_fd_sc_hd__inv_4 _5967_ (.A(_3342_[0]),
    .Y(_3338_[0]));
 sky130_fd_sc_hd__nand2_1 _5968_ (.A(net747),
    .B(_2107_),
    .Y(_2261_));
 sky130_fd_sc_hd__nand2_2 _5969_ (.A(net752),
    .B(_2111_),
    .Y(_2262_));
 sky130_fd_sc_hd__o211a_1 _5970_ (.A1(net740),
    .A2(_2102_),
    .B1(_2103_),
    .C1(net752),
    .X(_2263_));
 sky130_fd_sc_hd__mux2i_1 _5971_ (.A0(_3342_[0]),
    .A1(net761),
    .S(net751),
    .Y(_2264_));
 sky130_fd_sc_hd__mux2i_2 _5972_ (.A0(_2244_),
    .A1(_2264_),
    .S(net769),
    .Y(_2265_));
 sky130_fd_sc_hd__mux2i_2 _5973_ (.A0(_2188_),
    .A1(_2265_),
    .S(net737),
    .Y(_2266_));
 sky130_fd_sc_hd__and2_0 _5974_ (.A(net749),
    .B(_2266_),
    .X(_2267_));
 sky130_fd_sc_hd__nor3_1 _5975_ (.A(net778),
    .B(_2263_),
    .C(_2267_),
    .Y(_2268_));
 sky130_fd_sc_hd__a311oi_2 _5976_ (.A1(net778),
    .A2(_2261_),
    .A3(_2262_),
    .B1(_2268_),
    .C1(net741),
    .Y(_2269_));
 sky130_fd_sc_hd__a21oi_1 _5977_ (.A1(net745),
    .A2(_1921_),
    .B1(_0314_),
    .Y(_2270_));
 sky130_fd_sc_hd__a21oi_1 _5978_ (.A1(_1921_),
    .A2(_1942_),
    .B1(_2270_),
    .Y(_2271_));
 sky130_fd_sc_hd__nor2_2 _5979_ (.A(_2011_),
    .B(_2271_),
    .Y(_2272_));
 sky130_fd_sc_hd__a31oi_2 _5980_ (.A1(net739),
    .A2(_1942_),
    .A3(_2183_),
    .B1(_2272_),
    .Y(_2273_));
 sky130_fd_sc_hd__nor2_4 _5981_ (.A(_1801_),
    .B(_2273_),
    .Y(_2274_));
 sky130_fd_sc_hd__clkinv_1 _5982_ (.A(_3341_[0]),
    .Y(_2275_));
 sky130_fd_sc_hd__a31oi_1 _5983_ (.A1(_3357_[0]),
    .A2(net193),
    .A3(_1756_),
    .B1(_3356_[0]),
    .Y(_2276_));
 sky130_fd_sc_hd__o21ba_1 _5984_ (.A1(_2251_),
    .A2(_2276_),
    .B1_N(_3348_[0]),
    .X(_2277_));
 sky130_fd_sc_hd__xnor2_1 _5985_ (.A(_2275_),
    .B(_2277_),
    .Y(_2278_));
 sky130_fd_sc_hd__mux2i_1 _5986_ (.A0(_2275_),
    .A1(_3344_[0]),
    .S(net5),
    .Y(_2279_));
 sky130_fd_sc_hd__a22oi_1 _5987_ (.A1(_3340_[0]),
    .A2(net774),
    .B1(net773),
    .B2(_2279_),
    .Y(_2280_));
 sky130_fd_sc_hd__o211ai_1 _5988_ (.A1(_1731_),
    .A2(_2278_),
    .B1(_2280_),
    .C1(_1716_),
    .Y(_2281_));
 sky130_fd_sc_hd__o31a_1 _5989_ (.A1(_1716_),
    .A2(_2269_),
    .A3(_2274_),
    .B1(_2281_),
    .X(net71));
 sky130_fd_sc_hd__inv_1 _5990_ (.A(_3334_[0]),
    .Y(_3330_[0]));
 sky130_fd_sc_hd__nand2_1 _5991_ (.A(net264),
    .B(_3349_[0]),
    .Y(_2282_));
 sky130_fd_sc_hd__o21ai_0 _5992_ (.A1(_2282_),
    .A2(net702),
    .B1(_1760_),
    .Y(_2283_));
 sky130_fd_sc_hd__nor2_1 _5993_ (.A(_3333_[0]),
    .B(_1731_),
    .Y(_2284_));
 sky130_fd_sc_hd__o2111a_1 _5994_ (.A1(_2282_),
    .A2(net702),
    .B1(_3333_[0]),
    .C1(_1727_),
    .D1(_1760_),
    .X(_2285_));
 sky130_fd_sc_hd__mux2i_1 _5995_ (.A0(_1759_),
    .A1(_3336_[0]),
    .S(net5),
    .Y(_2286_));
 sky130_fd_sc_hd__a22o_1 _5996_ (.A1(_3332_[0]),
    .A2(net774),
    .B1(net773),
    .B2(_2286_),
    .X(_2287_));
 sky130_fd_sc_hd__a211oi_2 _5997_ (.A1(_2283_),
    .A2(_2284_),
    .B1(_2287_),
    .C1(_2285_),
    .Y(_2288_));
 sky130_fd_sc_hd__mux2i_1 _5998_ (.A0(net763),
    .A1(_1203_),
    .S(net751),
    .Y(_2289_));
 sky130_fd_sc_hd__mux2i_2 _5999_ (.A0(_2264_),
    .A1(_2289_),
    .S(net769),
    .Y(_2290_));
 sky130_fd_sc_hd__mux2i_1 _6000_ (.A0(_2214_),
    .A1(_2290_),
    .S(net738),
    .Y(_2291_));
 sky130_fd_sc_hd__nand2_1 _6001_ (.A(net748),
    .B(_2291_),
    .Y(_2292_));
 sky130_fd_sc_hd__o21ai_2 _6002_ (.A1(net748),
    .A2(_2136_),
    .B1(_2292_),
    .Y(_2293_));
 sky130_fd_sc_hd__nand2_1 _6003_ (.A(net749),
    .B(_2140_),
    .Y(_2294_));
 sky130_fd_sc_hd__nand2_1 _6004_ (.A(net752),
    .B(_2127_),
    .Y(_2295_));
 sky130_fd_sc_hd__or3_4 _6005_ (.A(net816),
    .B(net268),
    .C(_1863_),
    .X(_2296_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_28 ();
 sky130_fd_sc_hd__a21o_4 _6007_ (.A1(_0314_),
    .A2(net268),
    .B1(_2011_),
    .X(_2298_));
 sky130_fd_sc_hd__nand2_4 _6008_ (.A(_2296_),
    .B(_2298_),
    .Y(_2299_));
 sky130_fd_sc_hd__a31oi_2 _6009_ (.A1(net739),
    .A2(_2022_),
    .A3(_2183_),
    .B1(_2299_),
    .Y(_2300_));
 sky130_fd_sc_hd__a31oi_2 _6010_ (.A1(net750),
    .A2(_2294_),
    .A3(_2295_),
    .B1(_2300_),
    .Y(_2301_));
 sky130_fd_sc_hd__a211oi_4 _6011_ (.A1(_1920_),
    .A2(_2293_),
    .B1(_2301_),
    .C1(_1716_),
    .Y(_2302_));
 sky130_fd_sc_hd__a21oi_2 _6012_ (.A1(_2288_),
    .A2(_1716_),
    .B1(_2302_),
    .Y(net72));
 sky130_fd_sc_hd__inv_1 _6013_ (.A(_3326_[0]),
    .Y(_3322_[0]));
 sky130_fd_sc_hd__nor2_4 _6014_ (.A(_1801_),
    .B(net778),
    .Y(_2303_));
 sky130_fd_sc_hd__nand2_4 _6015_ (.A(_1921_),
    .B(_2303_),
    .Y(_2304_));
 sky130_fd_sc_hd__o21ai_0 _6016_ (.A1(net268),
    .A2(_1861_),
    .B1(_2299_),
    .Y(_2305_));
 sky130_fd_sc_hd__o211ai_1 _6017_ (.A1(_1869_),
    .A2(_2304_),
    .B1(_2305_),
    .C1(net777),
    .Y(_2306_));
 sky130_fd_sc_hd__nand3_2 _6018_ (.A(net752),
    .B(_2146_),
    .C(_2149_),
    .Y(_2307_));
 sky130_fd_sc_hd__mux2i_1 _6019_ (.A0(_3326_[0]),
    .A1(_3342_[0]),
    .S(net751),
    .Y(_2308_));
 sky130_fd_sc_hd__mux2i_1 _6020_ (.A0(_2289_),
    .A1(_2308_),
    .S(net769),
    .Y(_2309_));
 sky130_fd_sc_hd__mux2i_1 _6021_ (.A0(_2230_),
    .A1(_2309_),
    .S(net737),
    .Y(_2310_));
 sky130_fd_sc_hd__nand2_1 _6022_ (.A(net748),
    .B(_2310_),
    .Y(_2311_));
 sky130_fd_sc_hd__a21oi_1 _6023_ (.A1(_2307_),
    .A2(_2311_),
    .B1(_1870_),
    .Y(_2312_));
 sky130_fd_sc_hd__o21bai_1 _6024_ (.A1(_2275_),
    .A2(_2277_),
    .B1_N(_3340_[0]),
    .Y(_2313_));
 sky130_fd_sc_hd__a21oi_1 _6025_ (.A1(_3333_[0]),
    .A2(_2313_),
    .B1(_3332_[0]),
    .Y(_2314_));
 sky130_fd_sc_hd__xor2_1 _6026_ (.A(_3325_[0]),
    .B(_2314_),
    .X(_2315_));
 sky130_fd_sc_hd__nor2_1 _6027_ (.A(net5),
    .B(_3325_[0]),
    .Y(_2316_));
 sky130_fd_sc_hd__a21oi_1 _6028_ (.A1(net5),
    .A2(_3328_[0]),
    .B1(_2316_),
    .Y(_2317_));
 sky130_fd_sc_hd__a221oi_1 _6029_ (.A1(_3324_[0]),
    .A2(net774),
    .B1(net773),
    .B2(_2317_),
    .C1(net777),
    .Y(_2318_));
 sky130_fd_sc_hd__o21ai_0 _6030_ (.A1(_1731_),
    .A2(_2315_),
    .B1(_2318_),
    .Y(_2319_));
 sky130_fd_sc_hd__o21a_4 _6031_ (.A1(_2306_),
    .A2(_2312_),
    .B1(_2319_),
    .X(net73));
 sky130_fd_sc_hd__clkinv_1 _6032_ (.A(_3318_[0]),
    .Y(_3314_[0]));
 sky130_fd_sc_hd__inv_1 _6033_ (.A(_3317_[0]),
    .Y(_2320_));
 sky130_fd_sc_hd__o21ai_4 _6034_ (.A1(_1764_),
    .A2(net363),
    .B1(_1766_),
    .Y(_2321_));
 sky130_fd_sc_hd__xnor2_1 _6035_ (.A(_2321_),
    .B(_2320_),
    .Y(_2322_));
 sky130_fd_sc_hd__nand2_1 _6036_ (.A(_1727_),
    .B(_2322_),
    .Y(_2323_));
 sky130_fd_sc_hd__mux2i_1 _6037_ (.A0(_2320_),
    .A1(_3320_[0]),
    .S(net5),
    .Y(_2324_));
 sky130_fd_sc_hd__a221oi_2 _6038_ (.A1(_3316_[0]),
    .A2(net774),
    .B1(net773),
    .B2(_2324_),
    .C1(net777),
    .Y(_2325_));
 sky130_fd_sc_hd__nand2_1 _6039_ (.A(net752),
    .B(_2179_),
    .Y(_2326_));
 sky130_fd_sc_hd__mux2i_1 _6040_ (.A0(net764),
    .A1(net763),
    .S(net751),
    .Y(_2327_));
 sky130_fd_sc_hd__mux2i_1 _6041_ (.A0(_2308_),
    .A1(_2327_),
    .S(net769),
    .Y(_2328_));
 sky130_fd_sc_hd__mux2i_2 _6042_ (.A0(_2245_),
    .A1(_2328_),
    .S(net738),
    .Y(_2329_));
 sky130_fd_sc_hd__nand2_1 _6043_ (.A(net749),
    .B(_2329_),
    .Y(_2330_));
 sky130_fd_sc_hd__nand2_1 _6044_ (.A(_2326_),
    .B(_2330_),
    .Y(_2331_));
 sky130_fd_sc_hd__a21oi_1 _6045_ (.A1(net752),
    .A2(_1886_),
    .B1(net268),
    .Y(_2332_));
 sky130_fd_sc_hd__a21oi_1 _6046_ (.A1(_1894_),
    .A2(_2332_),
    .B1(_2298_),
    .Y(_2333_));
 sky130_fd_sc_hd__nand2_1 _6047_ (.A(net752),
    .B(_1882_),
    .Y(_2334_));
 sky130_fd_sc_hd__a21oi_1 _6048_ (.A1(_1894_),
    .A2(_2334_),
    .B1(_2296_),
    .Y(_2335_));
 sky130_fd_sc_hd__o21ai_1 _6049_ (.A1(_2071_),
    .A2(_2304_),
    .B1(net777),
    .Y(_2336_));
 sky130_fd_sc_hd__a2111oi_0 _6050_ (.A1(_1920_),
    .A2(_2331_),
    .B1(_2333_),
    .C1(_2335_),
    .D1(_2336_),
    .Y(_2337_));
 sky130_fd_sc_hd__a21oi_4 _6051_ (.A1(_2323_),
    .A2(_2325_),
    .B1(net703),
    .Y(net74));
 sky130_fd_sc_hd__clkinv_1 _6052_ (.A(_3310_[0]),
    .Y(_3306_[0]));
 sky130_fd_sc_hd__mux2i_1 _6053_ (.A0(_1937_),
    .A1(_1946_),
    .S(net752),
    .Y(_2338_));
 sky130_fd_sc_hd__a21oi_4 _6054_ (.A1(_0314_),
    .A2(net741),
    .B1(_2011_),
    .Y(_2339_));
 sky130_fd_sc_hd__o21ai_2 _6055_ (.A1(net741),
    .A2(_2338_),
    .B1(_2339_),
    .Y(_2340_));
 sky130_fd_sc_hd__or2_0 _6056_ (.A(net749),
    .B(_2190_),
    .X(_2341_));
 sky130_fd_sc_hd__mux2i_1 _6057_ (.A0(_3310_[0]),
    .A1(_3326_[0]),
    .S(net751),
    .Y(_2342_));
 sky130_fd_sc_hd__mux2_4 _6058_ (.A0(_2327_),
    .A1(_2342_),
    .S(net769),
    .X(_2343_));
 sky130_fd_sc_hd__nor2_1 _6059_ (.A(net740),
    .B(_2343_),
    .Y(_2344_));
 sky130_fd_sc_hd__a21oi_2 _6060_ (.A1(net740),
    .A2(_2265_),
    .B1(_2344_),
    .Y(_2345_));
 sky130_fd_sc_hd__nand2_1 _6061_ (.A(net748),
    .B(_2345_),
    .Y(_2346_));
 sky130_fd_sc_hd__a21oi_1 _6062_ (.A1(_2341_),
    .A2(_2346_),
    .B1(_1870_),
    .Y(_2347_));
 sky130_fd_sc_hd__o21ai_1 _6063_ (.A1(net314),
    .A2(_2304_),
    .B1(net777),
    .Y(_2348_));
 sky130_fd_sc_hd__nor3_2 _6064_ (.A(net816),
    .B(net268),
    .C(_1863_),
    .Y(_2349_));
 sky130_fd_sc_hd__o21ai_2 _6065_ (.A1(net748),
    .A2(_1943_),
    .B1(_2349_),
    .Y(_2350_));
 sky130_fd_sc_hd__a21oi_1 _6066_ (.A1(net748),
    .A2(_1937_),
    .B1(_2350_),
    .Y(_2351_));
 sky130_fd_sc_hd__nor3_2 _6067_ (.A(_2347_),
    .B(_2348_),
    .C(_2351_),
    .Y(_2352_));
 sky130_fd_sc_hd__o21ai_0 _6068_ (.A1(_1764_),
    .A2(_2276_),
    .B1(_1766_),
    .Y(_2353_));
 sky130_fd_sc_hd__a21oi_1 _6069_ (.A1(_3317_[0]),
    .A2(_2353_),
    .B1(_3316_[0]),
    .Y(_2354_));
 sky130_fd_sc_hd__xnor2_1 _6070_ (.A(_3309_[0]),
    .B(_2354_),
    .Y(_2355_));
 sky130_fd_sc_hd__nand2_1 _6071_ (.A(net5),
    .B(_3312_[0]),
    .Y(_2356_));
 sky130_fd_sc_hd__o21ai_0 _6072_ (.A1(net5),
    .A2(_3309_[0]),
    .B1(_2356_),
    .Y(_2357_));
 sky130_fd_sc_hd__o21ai_0 _6073_ (.A1(_1721_),
    .A2(_2357_),
    .B1(_1716_),
    .Y(_2358_));
 sky130_fd_sc_hd__a221oi_2 _6074_ (.A1(_3308_[0]),
    .A2(net774),
    .B1(_2355_),
    .B2(_1727_),
    .C1(_2358_),
    .Y(_2359_));
 sky130_fd_sc_hd__a21oi_4 _6075_ (.A1(_2340_),
    .A2(_2352_),
    .B1(_2359_),
    .Y(net75));
 sky130_fd_sc_hd__inv_4 _6076_ (.A(_3302_[0]),
    .Y(_3298_[0]));
 sky130_fd_sc_hd__nand2_1 _6077_ (.A(net750),
    .B(_2020_),
    .Y(_2360_));
 sky130_fd_sc_hd__mux2i_1 _6078_ (.A0(net765),
    .A1(net764),
    .S(net751),
    .Y(_2361_));
 sky130_fd_sc_hd__mux2i_2 _6079_ (.A0(_2342_),
    .A1(_2361_),
    .S(net769),
    .Y(_2362_));
 sky130_fd_sc_hd__mux2i_2 _6080_ (.A0(_2290_),
    .A1(_2362_),
    .S(net738),
    .Y(_2363_));
 sky130_fd_sc_hd__mux2i_1 _6081_ (.A0(_2215_),
    .A1(_2363_),
    .S(net749),
    .Y(_2364_));
 sky130_fd_sc_hd__o221ai_1 _6082_ (.A1(_1998_),
    .A2(_2304_),
    .B1(_2364_),
    .B2(_1870_),
    .C1(net777),
    .Y(_2365_));
 sky130_fd_sc_hd__a21oi_1 _6083_ (.A1(_2339_),
    .A2(_2360_),
    .B1(_2365_),
    .Y(_2366_));
 sky130_fd_sc_hd__o21ai_2 _6084_ (.A1(net741),
    .A2(_2026_),
    .B1(_2366_),
    .Y(_2367_));
 sky130_fd_sc_hd__inv_1 _6085_ (.A(_3301_[0]),
    .Y(_2368_));
 sky130_fd_sc_hd__mux2i_1 _6086_ (.A0(_2368_),
    .A1(_3304_[0]),
    .S(net5),
    .Y(_2369_));
 sky130_fd_sc_hd__a221o_1 _6087_ (.A1(_3300_[0]),
    .A2(net774),
    .B1(net773),
    .B2(_2369_),
    .C1(net777),
    .X(_2370_));
 sky130_fd_sc_hd__nand3_1 _6088_ (.A(_3309_[0]),
    .B(_3301_[0]),
    .C(_3317_[0]),
    .Y(_2371_));
 sky130_fd_sc_hd__nor3_2 _6089_ (.A(_1764_),
    .B(net702),
    .C(_2371_),
    .Y(_2372_));
 sky130_fd_sc_hd__a21oi_2 _6090_ (.A1(_1762_),
    .A2(_3317_[0]),
    .B1(_3316_[0]),
    .Y(_2373_));
 sky130_fd_sc_hd__nor2_1 _6091_ (.A(_1736_),
    .B(_2373_),
    .Y(_2374_));
 sky130_fd_sc_hd__nor2_1 _6092_ (.A(_3308_[0]),
    .B(_2374_),
    .Y(_2375_));
 sky130_fd_sc_hd__nor2_1 _6093_ (.A(_2368_),
    .B(_2375_),
    .Y(_2376_));
 sky130_fd_sc_hd__nor3_1 _6094_ (.A(_1731_),
    .B(_2372_),
    .C(_2376_),
    .Y(_2377_));
 sky130_fd_sc_hd__or2_4 _6095_ (.A(_2370_),
    .B(_2377_),
    .X(_2378_));
 sky130_fd_sc_hd__a21oi_1 _6096_ (.A1(_3317_[0]),
    .A2(_2321_),
    .B1(_3316_[0]),
    .Y(_2379_));
 sky130_fd_sc_hd__nor3_1 _6097_ (.A(_3308_[0]),
    .B(_3301_[0]),
    .C(_2370_),
    .Y(_2380_));
 sky130_fd_sc_hd__o21ai_1 _6098_ (.A1(_1736_),
    .A2(_2379_),
    .B1(_2380_),
    .Y(_2381_));
 sky130_fd_sc_hd__and3_1 _6099_ (.A(_2367_),
    .B(_2378_),
    .C(_2381_),
    .X(net76));
 sky130_fd_sc_hd__clkinv_1 _6100_ (.A(_3294_[0]),
    .Y(_3290_[0]));
 sky130_fd_sc_hd__nor2_1 _6101_ (.A(net740),
    .B(_1847_),
    .Y(_2382_));
 sky130_fd_sc_hd__o21ai_2 _6102_ (.A1(_2018_),
    .A2(_2382_),
    .B1(net750),
    .Y(_2383_));
 sky130_fd_sc_hd__nand2_1 _6103_ (.A(net749),
    .B(_2299_),
    .Y(_2384_));
 sky130_fd_sc_hd__o32ai_1 _6104_ (.A1(net749),
    .A2(_2034_),
    .A3(_2296_),
    .B1(_2384_),
    .B2(_2036_),
    .Y(_2385_));
 sky130_fd_sc_hd__a211oi_4 _6105_ (.A1(_2339_),
    .A2(_2383_),
    .B1(_2385_),
    .C1(_1716_),
    .Y(_2386_));
 sky130_fd_sc_hd__and2_0 _6106_ (.A(net752),
    .B(_2231_),
    .X(_2387_));
 sky130_fd_sc_hd__mux2_1 _6107_ (.A0(_2289_),
    .A1(_2308_),
    .S(net769),
    .X(_2388_));
 sky130_fd_sc_hd__mux2i_1 _6108_ (.A0(_3294_[0]),
    .A1(_3310_[0]),
    .S(net751),
    .Y(_2389_));
 sky130_fd_sc_hd__mux2_1 _6109_ (.A0(_2361_),
    .A1(_2389_),
    .S(net769),
    .X(_2390_));
 sky130_fd_sc_hd__mux2i_2 _6110_ (.A0(_2388_),
    .A1(_2390_),
    .S(net738),
    .Y(_2391_));
 sky130_fd_sc_hd__nor2_1 _6111_ (.A(net752),
    .B(_2391_),
    .Y(_2392_));
 sky130_fd_sc_hd__o21ai_0 _6112_ (.A1(_2387_),
    .A2(_2392_),
    .B1(net750),
    .Y(_2393_));
 sky130_fd_sc_hd__nand3_1 _6113_ (.A(net741),
    .B(net747),
    .C(_2044_),
    .Y(_2394_));
 sky130_fd_sc_hd__a21o_4 _6114_ (.A1(_2393_),
    .A2(_2394_),
    .B1(net778),
    .X(_2395_));
 sky130_fd_sc_hd__nand3_1 _6115_ (.A(_1740_),
    .B(_1763_),
    .C(net262),
    .Y(_2396_));
 sky130_fd_sc_hd__xnor2_1 _6116_ (.A(_3293_[0]),
    .B(_2396_),
    .Y(_2397_));
 sky130_fd_sc_hd__nand2_1 _6117_ (.A(net5),
    .B(_3296_[0]),
    .Y(_2398_));
 sky130_fd_sc_hd__o21ai_0 _6118_ (.A1(net5),
    .A2(_3293_[0]),
    .B1(_2398_),
    .Y(_2399_));
 sky130_fd_sc_hd__o21ai_0 _6119_ (.A1(_1721_),
    .A2(_2399_),
    .B1(_1716_),
    .Y(_2400_));
 sky130_fd_sc_hd__a221oi_2 _6120_ (.A1(_3292_[0]),
    .A2(net774),
    .B1(_2397_),
    .B2(_1727_),
    .C1(_2400_),
    .Y(_2401_));
 sky130_fd_sc_hd__a21oi_2 _6121_ (.A1(_2386_),
    .A2(_2395_),
    .B1(_2401_),
    .Y(net78));
 sky130_fd_sc_hd__clkinv_1 _6122_ (.A(_3286_[0]),
    .Y(_3282_[0]));
 sky130_fd_sc_hd__inv_1 _6123_ (.A(_3285_[0]),
    .Y(_2402_));
 sky130_fd_sc_hd__mux2i_1 _6124_ (.A0(_2402_),
    .A1(_3288_[0]),
    .S(net5),
    .Y(_2403_));
 sky130_fd_sc_hd__a221oi_1 _6125_ (.A1(_3284_[0]),
    .A2(net774),
    .B1(net773),
    .B2(_2403_),
    .C1(net777),
    .Y(_2404_));
 sky130_fd_sc_hd__nor2_1 _6126_ (.A(_1764_),
    .B(_2371_),
    .Y(_2405_));
 sky130_fd_sc_hd__nand2_1 _6127_ (.A(_3293_[0]),
    .B(_2405_),
    .Y(_2406_));
 sky130_fd_sc_hd__o21ai_2 _6128_ (.A1(_3300_[0]),
    .A2(_2376_),
    .B1(_3293_[0]),
    .Y(_2407_));
 sky130_fd_sc_hd__inv_1 _6129_ (.A(_3292_[0]),
    .Y(_2408_));
 sky130_fd_sc_hd__o211ai_1 _6130_ (.A1(_2406_),
    .A2(_2258_),
    .B1(_2407_),
    .C1(_2408_),
    .Y(_2409_));
 sky130_fd_sc_hd__xnor2_1 _6131_ (.A(_2402_),
    .B(net220),
    .Y(_2410_));
 sky130_fd_sc_hd__nand2_1 _6132_ (.A(_1727_),
    .B(_2410_),
    .Y(_2411_));
 sky130_fd_sc_hd__o21ai_0 _6133_ (.A1(net741),
    .A2(_2087_),
    .B1(_2339_),
    .Y(_2412_));
 sky130_fd_sc_hd__o211ai_1 _6134_ (.A1(_2086_),
    .A2(_2296_),
    .B1(_2412_),
    .C1(net777),
    .Y(_2413_));
 sky130_fd_sc_hd__mux2i_1 _6135_ (.A0(_3286_[0]),
    .A1(net765),
    .S(net751),
    .Y(_2414_));
 sky130_fd_sc_hd__mux2i_1 _6136_ (.A0(_2389_),
    .A1(_2414_),
    .S(net770),
    .Y(_2415_));
 sky130_fd_sc_hd__mux2i_1 _6137_ (.A0(_2328_),
    .A1(_2415_),
    .S(net738),
    .Y(_2416_));
 sky130_fd_sc_hd__a22oi_2 _6138_ (.A1(_2075_),
    .A2(_2303_),
    .B1(_2416_),
    .B2(_1920_),
    .Y(_2417_));
 sky130_fd_sc_hd__nand3_1 _6139_ (.A(_2082_),
    .B(_2083_),
    .C(_2299_),
    .Y(_2418_));
 sky130_fd_sc_hd__a21oi_1 _6140_ (.A1(_2417_),
    .A2(_2418_),
    .B1(net752),
    .Y(_2419_));
 sky130_fd_sc_hd__a311oi_4 _6141_ (.A1(net752),
    .A2(_1920_),
    .A3(_2246_),
    .B1(_2413_),
    .C1(_2419_),
    .Y(_2420_));
 sky130_fd_sc_hd__a21oi_4 _6142_ (.A1(_2411_),
    .A2(_2404_),
    .B1(_2420_),
    .Y(net79));
 sky130_fd_sc_hd__inv_1 _6143_ (.A(_3278_[0]),
    .Y(_3274_[0]));
 sky130_fd_sc_hd__a41o_1 _6144_ (.A1(_1763_),
    .A2(_1740_),
    .A3(_3293_[0]),
    .A4(net258),
    .B1(_3292_[0]),
    .X(_2421_));
 sky130_fd_sc_hd__a21oi_2 _6145_ (.A1(net260),
    .A2(_3285_[0]),
    .B1(_3284_[0]),
    .Y(_2422_));
 sky130_fd_sc_hd__xnor2_1 _6146_ (.A(_3277_[0]),
    .B(_2422_),
    .Y(_2423_));
 sky130_fd_sc_hd__nand2_1 _6147_ (.A(net5),
    .B(_3280_[0]),
    .Y(_2424_));
 sky130_fd_sc_hd__o21ai_0 _6148_ (.A1(net5),
    .A2(_3277_[0]),
    .B1(_2424_),
    .Y(_2425_));
 sky130_fd_sc_hd__o21ai_0 _6149_ (.A1(_1721_),
    .A2(_2425_),
    .B1(_1716_),
    .Y(_2426_));
 sky130_fd_sc_hd__a221oi_2 _6150_ (.A1(_3276_[0]),
    .A2(net774),
    .B1(_2423_),
    .B2(_1727_),
    .C1(_2426_),
    .Y(_2427_));
 sky130_fd_sc_hd__nor2_4 _6151_ (.A(_0314_),
    .B(_2011_),
    .Y(_2428_));
 sky130_fd_sc_hd__nor2_1 _6152_ (.A(_1801_),
    .B(_2428_),
    .Y(_2429_));
 sky130_fd_sc_hd__mux2i_1 _6153_ (.A0(_3278_[0]),
    .A1(_3294_[0]),
    .S(net751),
    .Y(_2430_));
 sky130_fd_sc_hd__mux2_1 _6154_ (.A0(_2414_),
    .A1(_2430_),
    .S(net770),
    .X(_2431_));
 sky130_fd_sc_hd__mux2i_1 _6155_ (.A0(_2343_),
    .A1(_2431_),
    .S(net738),
    .Y(_2432_));
 sky130_fd_sc_hd__nand2_1 _6156_ (.A(_1920_),
    .B(_2432_),
    .Y(_2433_));
 sky130_fd_sc_hd__o21ai_0 _6157_ (.A1(_1863_),
    .A2(_2111_),
    .B1(_2433_),
    .Y(_2434_));
 sky130_fd_sc_hd__a21oi_2 _6158_ (.A1(net374),
    .A2(_2429_),
    .B1(_2434_),
    .Y(_2435_));
 sky130_fd_sc_hd__a22oi_1 _6159_ (.A1(_1920_),
    .A2(_2266_),
    .B1(_2428_),
    .B2(_2112_),
    .Y(_2436_));
 sky130_fd_sc_hd__a31oi_1 _6160_ (.A1(_2111_),
    .A2(_2112_),
    .A3(_2428_),
    .B1(net752),
    .Y(_2437_));
 sky130_fd_sc_hd__a32oi_1 _6161_ (.A1(_1942_),
    .A2(_2085_),
    .A3(_2299_),
    .B1(_2339_),
    .B2(net741),
    .Y(_2438_));
 sky130_fd_sc_hd__o211ai_1 _6162_ (.A1(_2436_),
    .A2(_2437_),
    .B1(_2438_),
    .C1(net777),
    .Y(_2439_));
 sky130_fd_sc_hd__a21oi_4 _6163_ (.A1(net748),
    .A2(_2435_),
    .B1(_2439_),
    .Y(_2440_));
 sky130_fd_sc_hd__nor2_2 _6164_ (.A(_2440_),
    .B(_2427_),
    .Y(net80));
 sky130_fd_sc_hd__clkinvlp_4 _6165_ (.A(_3270_[0]),
    .Y(_3266_[0]));
 sky130_fd_sc_hd__nand2_1 _6166_ (.A(net752),
    .B(_2291_),
    .Y(_2441_));
 sky130_fd_sc_hd__mux2i_1 _6167_ (.A0(net281),
    .A1(_3286_[0]),
    .S(net751),
    .Y(_2442_));
 sky130_fd_sc_hd__mux2i_1 _6168_ (.A0(_2430_),
    .A1(_2442_),
    .S(net770),
    .Y(_2443_));
 sky130_fd_sc_hd__mux2i_1 _6169_ (.A0(_2362_),
    .A1(_2443_),
    .S(net738),
    .Y(_2444_));
 sky130_fd_sc_hd__nand2_1 _6170_ (.A(net748),
    .B(_2444_),
    .Y(_2445_));
 sky130_fd_sc_hd__a21oi_1 _6171_ (.A1(_2441_),
    .A2(_2445_),
    .B1(_1870_),
    .Y(_2446_));
 sky130_fd_sc_hd__a22oi_1 _6172_ (.A1(_2022_),
    .A2(_2085_),
    .B1(_2127_),
    .B2(net749),
    .Y(_2447_));
 sky130_fd_sc_hd__a21oi_1 _6173_ (.A1(net750),
    .A2(net749),
    .B1(_0314_),
    .Y(_2448_));
 sky130_fd_sc_hd__a31oi_1 _6174_ (.A1(net750),
    .A2(net749),
    .A3(_2127_),
    .B1(_2448_),
    .Y(_2449_));
 sky130_fd_sc_hd__o22ai_2 _6175_ (.A1(_2296_),
    .A2(_2447_),
    .B1(_2449_),
    .B2(_2011_),
    .Y(_2450_));
 sky130_fd_sc_hd__nand2_1 _6176_ (.A(net741),
    .B(_1863_),
    .Y(_2451_));
 sky130_fd_sc_hd__o31ai_1 _6177_ (.A1(net752),
    .A2(_2136_),
    .A3(_2451_),
    .B1(net777),
    .Y(_2452_));
 sky130_fd_sc_hd__nor3_2 _6178_ (.A(_2446_),
    .B(_2450_),
    .C(_2452_),
    .Y(_2453_));
 sky130_fd_sc_hd__inv_1 _6179_ (.A(_3269_[0]),
    .Y(_2454_));
 sky130_fd_sc_hd__mux2i_1 _6180_ (.A0(_2454_),
    .A1(_3272_[0]),
    .S(net5),
    .Y(_2455_));
 sky130_fd_sc_hd__a221o_1 _6181_ (.A1(_3268_[0]),
    .A2(net774),
    .B1(net773),
    .B2(_2455_),
    .C1(net777),
    .X(_2456_));
 sky130_fd_sc_hd__a21o_4 _6182_ (.A1(_3277_[0]),
    .A2(_3284_[0]),
    .B1(_3276_[0]),
    .X(_2457_));
 sky130_fd_sc_hd__a21oi_1 _6183_ (.A1(_1775_),
    .A2(net219),
    .B1(_2457_),
    .Y(_2458_));
 sky130_fd_sc_hd__nor3_1 _6184_ (.A(_2454_),
    .B(_2456_),
    .C(_2458_),
    .Y(_2459_));
 sky130_fd_sc_hd__nor3b_1 _6185_ (.A(_3269_[0]),
    .B(_2456_),
    .C_N(_2458_),
    .Y(_2460_));
 sky130_fd_sc_hd__nor2_1 _6186_ (.A(_1727_),
    .B(_2456_),
    .Y(_2461_));
 sky130_fd_sc_hd__nor4_2 _6187_ (.A(_2453_),
    .B(_2461_),
    .C(_2460_),
    .D(_2459_),
    .Y(net81));
 sky130_fd_sc_hd__clkinv_1 _6188_ (.A(_3262_[0]),
    .Y(_3258_[0]));
 sky130_fd_sc_hd__nand2_1 _6189_ (.A(_3260_[0]),
    .B(net774),
    .Y(_2462_));
 sky130_fd_sc_hd__nand2_1 _6190_ (.A(net5),
    .B(_3264_[0]),
    .Y(_2463_));
 sky130_fd_sc_hd__o211ai_1 _6191_ (.A1(net5),
    .A2(_3261_[0]),
    .B1(net773),
    .C1(_2463_),
    .Y(_2464_));
 sky130_fd_sc_hd__nand4_1 _6192_ (.A(_1763_),
    .B(_1740_),
    .C(_3293_[0]),
    .D(net258),
    .Y(_2465_));
 sky130_fd_sc_hd__nand2_1 _6193_ (.A(_3269_[0]),
    .B(_1775_),
    .Y(_2466_));
 sky130_fd_sc_hd__o21ai_2 _6194_ (.A1(_2466_),
    .A2(_2465_),
    .B1(_1781_),
    .Y(_2467_));
 sky130_fd_sc_hd__xnor2_1 _6195_ (.A(_3261_[0]),
    .B(_2467_),
    .Y(_2468_));
 sky130_fd_sc_hd__or2_0 _6196_ (.A(_1731_),
    .B(_2468_),
    .X(_2469_));
 sky130_fd_sc_hd__mux2i_1 _6197_ (.A0(_3262_[0]),
    .A1(_3278_[0]),
    .S(net751),
    .Y(_2470_));
 sky130_fd_sc_hd__mux2i_1 _6198_ (.A0(_2442_),
    .A1(_2470_),
    .S(net770),
    .Y(_2471_));
 sky130_fd_sc_hd__nor2_1 _6199_ (.A(net740),
    .B(_2471_),
    .Y(_2472_));
 sky130_fd_sc_hd__a21oi_1 _6200_ (.A1(net740),
    .A2(_2390_),
    .B1(_2472_),
    .Y(_2473_));
 sky130_fd_sc_hd__nand2_1 _6201_ (.A(net752),
    .B(_2310_),
    .Y(_2474_));
 sky130_fd_sc_hd__o21ai_0 _6202_ (.A1(net752),
    .A2(_2473_),
    .B1(_2474_),
    .Y(_2475_));
 sky130_fd_sc_hd__a211oi_2 _6203_ (.A1(_1863_),
    .A2(_2475_),
    .B1(_2145_),
    .C1(net741),
    .Y(_2476_));
 sky130_fd_sc_hd__nor2_2 _6204_ (.A(net778),
    .B(_2152_),
    .Y(_2477_));
 sky130_fd_sc_hd__nor3_1 _6205_ (.A(_1801_),
    .B(_2428_),
    .C(_2477_),
    .Y(_2478_));
 sky130_fd_sc_hd__o21a_4 _6206_ (.A1(_2476_),
    .A2(_2478_),
    .B1(net777),
    .X(_2479_));
 sky130_fd_sc_hd__a41oi_2 _6207_ (.A1(_1716_),
    .A2(_2462_),
    .A3(_2464_),
    .A4(_2469_),
    .B1(_2479_),
    .Y(net82));
 sky130_fd_sc_hd__clkinv_1 _6208_ (.A(_3254_[0]),
    .Y(_3250_[0]));
 sky130_fd_sc_hd__mux2i_1 _6209_ (.A0(_1770_),
    .A1(_3256_[0]),
    .S(net5),
    .Y(_2480_));
 sky130_fd_sc_hd__a22oi_2 _6210_ (.A1(_3252_[0]),
    .A2(net774),
    .B1(net773),
    .B2(_2480_),
    .Y(_2481_));
 sky130_fd_sc_hd__nand3_1 _6211_ (.A(_3253_[0]),
    .B(_1716_),
    .C(_2481_),
    .Y(_2482_));
 sky130_fd_sc_hd__nand3_1 _6212_ (.A(_1770_),
    .B(_1716_),
    .C(_2481_),
    .Y(_2483_));
 sky130_fd_sc_hd__a21o_1 _6213_ (.A1(_3269_[0]),
    .A2(_2457_),
    .B1(_3268_[0]),
    .X(_2484_));
 sky130_fd_sc_hd__a21o_4 _6214_ (.A1(_3261_[0]),
    .A2(_2484_),
    .B1(_3260_[0]),
    .X(_2485_));
 sky130_fd_sc_hd__a41oi_2 _6215_ (.A1(net219),
    .A2(_3269_[0]),
    .A3(_1775_),
    .A4(_3261_[0]),
    .B1(_2485_),
    .Y(_2486_));
 sky130_fd_sc_hd__mux2i_1 _6216_ (.A0(_2482_),
    .A1(_2483_),
    .S(_2486_),
    .Y(_2487_));
 sky130_fd_sc_hd__a31oi_1 _6217_ (.A1(net750),
    .A2(net749),
    .A3(_1886_),
    .B1(_2448_),
    .Y(_2488_));
 sky130_fd_sc_hd__nor2_2 _6218_ (.A(_2011_),
    .B(_2488_),
    .Y(_2489_));
 sky130_fd_sc_hd__nand2_1 _6219_ (.A(net740),
    .B(_2415_),
    .Y(_2490_));
 sky130_fd_sc_hd__mux2i_1 _6220_ (.A0(net285),
    .A1(net281),
    .S(net751),
    .Y(_2491_));
 sky130_fd_sc_hd__mux2i_1 _6221_ (.A0(_2470_),
    .A1(_2491_),
    .S(net770),
    .Y(_2492_));
 sky130_fd_sc_hd__nand2_1 _6222_ (.A(net738),
    .B(_2492_),
    .Y(_2493_));
 sky130_fd_sc_hd__and3_4 _6223_ (.A(_1801_),
    .B(_2490_),
    .C(_2493_),
    .X(_2494_));
 sky130_fd_sc_hd__a21oi_1 _6224_ (.A1(net268),
    .A2(_2179_),
    .B1(_2494_),
    .Y(_2495_));
 sky130_fd_sc_hd__nor3_2 _6225_ (.A(net752),
    .B(net778),
    .C(_2495_),
    .Y(_2496_));
 sky130_fd_sc_hd__nand3_1 _6226_ (.A(net752),
    .B(_1920_),
    .C(_2329_),
    .Y(_2497_));
 sky130_fd_sc_hd__nand3_1 _6227_ (.A(net749),
    .B(_1882_),
    .C(_2349_),
    .Y(_2498_));
 sky130_fd_sc_hd__a31oi_2 _6228_ (.A1(_1923_),
    .A2(_2085_),
    .A3(_2303_),
    .B1(_1716_),
    .Y(_2499_));
 sky130_fd_sc_hd__nand3_2 _6229_ (.A(_2497_),
    .B(_2498_),
    .C(_2499_),
    .Y(_2500_));
 sky130_fd_sc_hd__nor3_4 _6230_ (.A(_2489_),
    .B(_2496_),
    .C(_2500_),
    .Y(_2501_));
 sky130_fd_sc_hd__a211oi_2 _6231_ (.A1(_1731_),
    .A2(_2481_),
    .B1(_2501_),
    .C1(_2487_),
    .Y(net83));
 sky130_fd_sc_hd__clkinv_1 _6232_ (.A(_3246_[0]),
    .Y(_3242_[0]));
 sky130_fd_sc_hd__mux2i_1 _6233_ (.A0(_3246_[0]),
    .A1(_3262_[0]),
    .S(net751),
    .Y(_2502_));
 sky130_fd_sc_hd__mux2i_1 _6234_ (.A0(_2491_),
    .A1(_2502_),
    .S(net770),
    .Y(_2503_));
 sky130_fd_sc_hd__nor2_1 _6235_ (.A(net738),
    .B(_2431_),
    .Y(_2504_));
 sky130_fd_sc_hd__a211oi_1 _6236_ (.A1(net738),
    .A2(_2503_),
    .B1(_2504_),
    .C1(net752),
    .Y(_2505_));
 sky130_fd_sc_hd__a21oi_1 _6237_ (.A1(net752),
    .A2(_2345_),
    .B1(_2505_),
    .Y(_2506_));
 sky130_fd_sc_hd__mux2i_1 _6238_ (.A0(_2197_),
    .A1(_2506_),
    .S(_1863_),
    .Y(_2507_));
 sky130_fd_sc_hd__nand2_1 _6239_ (.A(net778),
    .B(_2033_),
    .Y(_2508_));
 sky130_fd_sc_hd__and3_4 _6240_ (.A(net741),
    .B(_2191_),
    .C(_2508_),
    .X(_2509_));
 sky130_fd_sc_hd__a21oi_2 _6241_ (.A1(_1801_),
    .A2(_2507_),
    .B1(_2509_),
    .Y(_2510_));
 sky130_fd_sc_hd__a41o_1 _6242_ (.A1(_2421_),
    .A2(_3269_[0]),
    .A3(_1775_),
    .A4(_3261_[0]),
    .B1(_2485_),
    .X(_2511_));
 sky130_fd_sc_hd__a21oi_2 _6243_ (.A1(_2511_),
    .A2(_3253_[0]),
    .B1(_3252_[0]),
    .Y(_2512_));
 sky130_fd_sc_hd__xnor2_1 _6244_ (.A(_2512_),
    .B(_1769_),
    .Y(_2513_));
 sky130_fd_sc_hd__nor2_1 _6245_ (.A(_1731_),
    .B(_2513_),
    .Y(_2514_));
 sky130_fd_sc_hd__mux2i_1 _6246_ (.A0(_1769_),
    .A1(_3248_[0]),
    .S(net5),
    .Y(_2515_));
 sky130_fd_sc_hd__a221o_4 _6247_ (.A1(_3244_[0]),
    .A2(net774),
    .B1(net773),
    .B2(_2515_),
    .C1(net777),
    .X(_2516_));
 sky130_fd_sc_hd__o2bb2ai_2 _6248_ (.A1_N(net777),
    .A2_N(_2510_),
    .B1(_2516_),
    .B2(_2514_),
    .Y(_2517_));
 sky130_fd_sc_hd__inv_1 _6249_ (.A(_2517_),
    .Y(net84));
 sky130_fd_sc_hd__inv_1 _6250_ (.A(_3238_[0]),
    .Y(_3234_[0]));
 sky130_fd_sc_hd__a21oi_1 _6251_ (.A1(_3261_[0]),
    .A2(_3268_[0]),
    .B1(_3260_[0]),
    .Y(_2518_));
 sky130_fd_sc_hd__o21bai_1 _6252_ (.A1(_1770_),
    .A2(_2518_),
    .B1_N(_3252_[0]),
    .Y(_2519_));
 sky130_fd_sc_hd__a21oi_2 _6253_ (.A1(_3245_[0]),
    .A2(_2519_),
    .B1(_3244_[0]),
    .Y(_2520_));
 sky130_fd_sc_hd__nor2_1 _6254_ (.A(_3292_[0]),
    .B(_2457_),
    .Y(_2521_));
 sky130_fd_sc_hd__o2111ai_4 _6255_ (.A1(net362),
    .A2(_2406_),
    .B1(net286),
    .C1(_2520_),
    .D1(_2521_),
    .Y(_2522_));
 sky130_fd_sc_hd__nor2_1 _6256_ (.A(_1775_),
    .B(_2457_),
    .Y(_2523_));
 sky130_fd_sc_hd__o41ai_1 _6257_ (.A1(_1769_),
    .A2(_1770_),
    .A3(_1773_),
    .A4(_2523_),
    .B1(_2520_),
    .Y(_2524_));
 sky130_fd_sc_hd__nand2_1 _6258_ (.A(net5),
    .B(_3240_[0]),
    .Y(_2525_));
 sky130_fd_sc_hd__o21ai_0 _6259_ (.A1(net5),
    .A2(net270),
    .B1(_2525_),
    .Y(_2526_));
 sky130_fd_sc_hd__nand2_1 _6260_ (.A(_3236_[0]),
    .B(net774),
    .Y(_2527_));
 sky130_fd_sc_hd__o21ai_2 _6261_ (.A1(_1721_),
    .A2(_2526_),
    .B1(_2527_),
    .Y(_2528_));
 sky130_fd_sc_hd__nor3_1 _6262_ (.A(_1768_),
    .B(net777),
    .C(_2528_),
    .Y(_2529_));
 sky130_fd_sc_hd__and3_1 _6263_ (.A(_2522_),
    .B(_2524_),
    .C(_2529_),
    .X(_2530_));
 sky130_fd_sc_hd__or3_1 _6264_ (.A(net253),
    .B(net777),
    .C(_2528_),
    .X(_2531_));
 sky130_fd_sc_hd__a21oi_1 _6265_ (.A1(_2522_),
    .A2(_2524_),
    .B1(_2531_),
    .Y(_2532_));
 sky130_fd_sc_hd__nand2_1 _6266_ (.A(net752),
    .B(_2363_),
    .Y(_2533_));
 sky130_fd_sc_hd__mux2_1 _6267_ (.A0(net766),
    .A1(net285),
    .S(net751),
    .X(_2534_));
 sky130_fd_sc_hd__nor2_1 _6268_ (.A(net742),
    .B(_2534_),
    .Y(_2535_));
 sky130_fd_sc_hd__and2_4 _6269_ (.A(net742),
    .B(_2502_),
    .X(_2536_));
 sky130_fd_sc_hd__nand2_1 _6270_ (.A(net740),
    .B(_2443_),
    .Y(_2537_));
 sky130_fd_sc_hd__o311ai_0 _6271_ (.A1(net740),
    .A2(_2535_),
    .A3(_2536_),
    .B1(_2537_),
    .C1(net748),
    .Y(_2538_));
 sky130_fd_sc_hd__a21oi_1 _6272_ (.A1(_2533_),
    .A2(_2538_),
    .B1(_1870_),
    .Y(_2539_));
 sky130_fd_sc_hd__nand3_1 _6273_ (.A(_1803_),
    .B(net341),
    .C(_2349_),
    .Y(_2540_));
 sky130_fd_sc_hd__nand2_1 _6274_ (.A(net777),
    .B(_2540_),
    .Y(_2541_));
 sky130_fd_sc_hd__nor2_1 _6275_ (.A(net741),
    .B(_2220_),
    .Y(_2542_));
 sky130_fd_sc_hd__a21oi_1 _6276_ (.A1(_2217_),
    .A2(_2298_),
    .B1(_2542_),
    .Y(_2543_));
 sky130_fd_sc_hd__o32ai_1 _6277_ (.A1(_2539_),
    .A2(_2541_),
    .A3(_2543_),
    .B1(_2528_),
    .B2(_1727_),
    .Y(_2544_));
 sky130_fd_sc_hd__nor3_4 _6278_ (.A(_2532_),
    .B(_2530_),
    .C(_2544_),
    .Y(net85));
 sky130_fd_sc_hd__nand2b_1 _6279_ (.A_N(_1786_),
    .B(net326),
    .Y(_2545_));
 sky130_fd_sc_hd__xor2_1 _6280_ (.A(_2545_),
    .B(_3229_[0]),
    .X(_2546_));
 sky130_fd_sc_hd__nand2_1 _6281_ (.A(net5),
    .B(_3232_[0]),
    .Y(_2547_));
 sky130_fd_sc_hd__o21ai_0 _6282_ (.A1(net5),
    .A2(_3229_[0]),
    .B1(_2547_),
    .Y(_2548_));
 sky130_fd_sc_hd__o21ai_0 _6283_ (.A1(_1721_),
    .A2(_2548_),
    .B1(_1716_),
    .Y(_2549_));
 sky130_fd_sc_hd__a221oi_2 _6284_ (.A1(_3228_[0]),
    .A2(net774),
    .B1(_2546_),
    .B2(_1727_),
    .C1(_2549_),
    .Y(_2550_));
 sky130_fd_sc_hd__nor2_1 _6285_ (.A(_3226_[0]),
    .B(net751),
    .Y(_2551_));
 sky130_fd_sc_hd__a21oi_1 _6286_ (.A1(_3246_[0]),
    .A2(net751),
    .B1(_2551_),
    .Y(_2552_));
 sky130_fd_sc_hd__nand2_1 _6287_ (.A(net770),
    .B(_2552_),
    .Y(_2553_));
 sky130_fd_sc_hd__o21ai_1 _6288_ (.A1(net770),
    .A2(_2534_),
    .B1(_2553_),
    .Y(_2554_));
 sky130_fd_sc_hd__nor2_1 _6289_ (.A(net738),
    .B(_2471_),
    .Y(_2555_));
 sky130_fd_sc_hd__a21oi_1 _6290_ (.A1(net738),
    .A2(_2554_),
    .B1(_2555_),
    .Y(_2556_));
 sky130_fd_sc_hd__o22ai_1 _6291_ (.A1(_2034_),
    .A2(_2296_),
    .B1(_2556_),
    .B2(_1870_),
    .Y(_2557_));
 sky130_fd_sc_hd__nor3_1 _6292_ (.A(net748),
    .B(_1870_),
    .C(_2391_),
    .Y(_2558_));
 sky130_fd_sc_hd__o21ai_0 _6293_ (.A1(net741),
    .A2(_1872_),
    .B1(_0314_),
    .Y(_2559_));
 sky130_fd_sc_hd__o31ai_1 _6294_ (.A1(net741),
    .A2(_1847_),
    .A3(_1872_),
    .B1(_2559_),
    .Y(_2560_));
 sky130_fd_sc_hd__o221ai_1 _6295_ (.A1(_2232_),
    .A2(_2451_),
    .B1(_2560_),
    .B2(_2011_),
    .C1(net777),
    .Y(_2561_));
 sky130_fd_sc_hd__a211oi_2 _6296_ (.A1(net748),
    .A2(_2557_),
    .B1(_2558_),
    .C1(_2561_),
    .Y(_2562_));
 sky130_fd_sc_hd__nor2_2 _6297_ (.A(_2562_),
    .B(_2550_),
    .Y(net86));
 sky130_fd_sc_hd__a21oi_1 _6298_ (.A1(_3253_[0]),
    .A2(_2485_),
    .B1(_3252_[0]),
    .Y(_2563_));
 sky130_fd_sc_hd__nor2_1 _6299_ (.A(_1769_),
    .B(_2563_),
    .Y(_2564_));
 sky130_fd_sc_hd__o21ai_0 _6300_ (.A1(_3244_[0]),
    .A2(_2564_),
    .B1(net252),
    .Y(_2565_));
 sky130_fd_sc_hd__nand2b_1 _6301_ (.A_N(_3236_[0]),
    .B(_2565_),
    .Y(_2566_));
 sky130_fd_sc_hd__a21o_1 _6302_ (.A1(_3229_[0]),
    .A2(_2566_),
    .B1(_3228_[0]),
    .X(_2567_));
 sky130_fd_sc_hd__a41oi_2 _6303_ (.A1(_3229_[0]),
    .A2(_1774_),
    .A3(_1775_),
    .A4(net219),
    .B1(_2567_),
    .Y(_2568_));
 sky130_fd_sc_hd__xnor2_1 _6304_ (.A(_3221_[0]),
    .B(_2568_),
    .Y(_2569_));
 sky130_fd_sc_hd__o21ai_1 _6305_ (.A1(net777),
    .A2(_2569_),
    .B1(_1727_),
    .Y(_2570_));
 sky130_fd_sc_hd__nor2_1 _6306_ (.A(net5),
    .B(_3221_[0]),
    .Y(_2571_));
 sky130_fd_sc_hd__a21oi_1 _6307_ (.A1(net5),
    .A2(_3224_[0]),
    .B1(_2571_),
    .Y(_2572_));
 sky130_fd_sc_hd__a22oi_1 _6308_ (.A1(_3220_[0]),
    .A2(net774),
    .B1(net773),
    .B2(_2572_),
    .Y(_2573_));
 sky130_fd_sc_hd__o21ai_0 _6309_ (.A1(net741),
    .A2(_2239_),
    .B1(_2339_),
    .Y(_2574_));
 sky130_fd_sc_hd__o311a_1 _6310_ (.A1(_1872_),
    .A2(net307),
    .A3(_2296_),
    .B1(_2574_),
    .C1(net777),
    .X(_2575_));
 sky130_fd_sc_hd__nor2_1 _6311_ (.A(_0490_),
    .B(net751),
    .Y(_2576_));
 sky130_fd_sc_hd__a21oi_1 _6312_ (.A1(net766),
    .A2(net751),
    .B1(_2576_),
    .Y(_2577_));
 sky130_fd_sc_hd__mux2_1 _6313_ (.A0(_2552_),
    .A1(_2577_),
    .S(net770),
    .X(_2578_));
 sky130_fd_sc_hd__nor2_1 _6314_ (.A(net738),
    .B(_2492_),
    .Y(_2579_));
 sky130_fd_sc_hd__a21oi_1 _6315_ (.A1(net738),
    .A2(_2578_),
    .B1(_2579_),
    .Y(_2580_));
 sky130_fd_sc_hd__nand2_1 _6316_ (.A(net741),
    .B(_2246_),
    .Y(_2581_));
 sky130_fd_sc_hd__o21ai_0 _6317_ (.A1(net741),
    .A2(_2580_),
    .B1(_2581_),
    .Y(_2582_));
 sky130_fd_sc_hd__nand3_1 _6318_ (.A(_1803_),
    .B(_1863_),
    .C(_2582_),
    .Y(_2583_));
 sky130_fd_sc_hd__o211ai_1 _6319_ (.A1(_1803_),
    .A2(_2417_),
    .B1(_2575_),
    .C1(_2583_),
    .Y(_2584_));
 sky130_fd_sc_hd__a21boi_1 _6320_ (.A1(_2573_),
    .A2(_2570_),
    .B1_N(_2584_),
    .Y(net87));
 sky130_fd_sc_hd__inv_2 _6321_ (.A(net767),
    .Y(_3210_[0]));
 sky130_fd_sc_hd__o21a_1 _6322_ (.A1(_2263_),
    .A2(_2267_),
    .B1(_1863_),
    .X(_2585_));
 sky130_fd_sc_hd__o22ai_2 _6323_ (.A1(net741),
    .A2(_2272_),
    .B1(_2339_),
    .B2(_2585_),
    .Y(_2586_));
 sky130_fd_sc_hd__nor2_2 _6324_ (.A(_1872_),
    .B(_2296_),
    .Y(_2587_));
 sky130_fd_sc_hd__nor2_1 _6325_ (.A(_3226_[0]),
    .B(net745),
    .Y(_2588_));
 sky130_fd_sc_hd__a21oi_1 _6326_ (.A1(net767),
    .A2(net745),
    .B1(_2588_),
    .Y(_2589_));
 sky130_fd_sc_hd__mux2_1 _6327_ (.A0(_2577_),
    .A1(_2589_),
    .S(net770),
    .X(_2590_));
 sky130_fd_sc_hd__nand2_1 _6328_ (.A(net740),
    .B(_2503_),
    .Y(_2591_));
 sky130_fd_sc_hd__o211ai_1 _6329_ (.A1(net740),
    .A2(_2590_),
    .B1(_2591_),
    .C1(net748),
    .Y(_2592_));
 sky130_fd_sc_hd__o21ai_0 _6330_ (.A1(net748),
    .A2(_2432_),
    .B1(_2592_),
    .Y(_2593_));
 sky130_fd_sc_hd__a221oi_2 _6331_ (.A1(_1942_),
    .A2(_2587_),
    .B1(_2593_),
    .B2(_1920_),
    .C1(_1716_),
    .Y(_2594_));
 sky130_fd_sc_hd__xnor2_2 _6332_ (.A(_3213_[0]),
    .B(_1791_),
    .Y(_2595_));
 sky130_fd_sc_hd__inv_1 _6333_ (.A(_3216_[0]),
    .Y(_2596_));
 sky130_fd_sc_hd__mux2i_1 _6334_ (.A0(_3213_[0]),
    .A1(_2596_),
    .S(net5),
    .Y(_2597_));
 sky130_fd_sc_hd__o21ai_0 _6335_ (.A1(_1721_),
    .A2(_2597_),
    .B1(_1716_),
    .Y(_2598_));
 sky130_fd_sc_hd__a221oi_2 _6336_ (.A1(_3212_[0]),
    .A2(net774),
    .B1(_2595_),
    .B2(_1727_),
    .C1(_2598_),
    .Y(_2599_));
 sky130_fd_sc_hd__a21oi_1 _6337_ (.A1(_2586_),
    .A2(_2594_),
    .B1(_2599_),
    .Y(net89));
 sky130_fd_sc_hd__nor2_1 _6338_ (.A(net777),
    .B(_1792_),
    .Y(_2600_));
 sky130_fd_sc_hd__nor3_1 _6339_ (.A(_3205_[0]),
    .B(_3212_[0]),
    .C(net777),
    .Y(_2601_));
 sky130_fd_sc_hd__o21bai_1 _6340_ (.A1(_1768_),
    .A2(_2520_),
    .B1_N(_3236_[0]),
    .Y(_2602_));
 sky130_fd_sc_hd__a21o_1 _6341_ (.A1(_3229_[0]),
    .A2(_2602_),
    .B1(_3228_[0]),
    .X(_2603_));
 sky130_fd_sc_hd__a21oi_1 _6342_ (.A1(_3221_[0]),
    .A2(_2603_),
    .B1(_3220_[0]),
    .Y(_2604_));
 sky130_fd_sc_hd__o2111ai_1 _6343_ (.A1(net702),
    .A2(_2406_),
    .B1(net267),
    .C1(_2521_),
    .D1(_2604_),
    .Y(_2605_));
 sky130_fd_sc_hd__nand3_1 _6344_ (.A(_3221_[0]),
    .B(_3229_[0]),
    .C(_1774_),
    .Y(_2606_));
 sky130_fd_sc_hd__o21ai_0 _6345_ (.A1(_2523_),
    .A2(_2606_),
    .B1(_2604_),
    .Y(_2607_));
 sky130_fd_sc_hd__nand2_1 _6346_ (.A(_2607_),
    .B(_2605_),
    .Y(_2608_));
 sky130_fd_sc_hd__mux2i_1 _6347_ (.A0(_2600_),
    .A1(_2601_),
    .S(_2608_),
    .Y(_2609_));
 sky130_fd_sc_hd__nor4_1 _6348_ (.A(_3205_[0]),
    .B(_3213_[0]),
    .C(_3212_[0]),
    .D(net777),
    .Y(_2610_));
 sky130_fd_sc_hd__a31oi_1 _6349_ (.A1(_3205_[0]),
    .A2(_3212_[0]),
    .A3(_1716_),
    .B1(_2610_),
    .Y(_2611_));
 sky130_fd_sc_hd__nand3_1 _6350_ (.A(_1727_),
    .B(_2609_),
    .C(_2611_),
    .Y(_2612_));
 sky130_fd_sc_hd__nor2_1 _6351_ (.A(net5),
    .B(_3205_[0]),
    .Y(_2613_));
 sky130_fd_sc_hd__a21oi_1 _6352_ (.A1(net5),
    .A2(_3208_[0]),
    .B1(_2613_),
    .Y(_2614_));
 sky130_fd_sc_hd__a22oi_1 _6353_ (.A1(_3204_[0]),
    .A2(net774),
    .B1(net773),
    .B2(_2614_),
    .Y(_2615_));
 sky130_fd_sc_hd__nor2_1 _6354_ (.A(_2535_),
    .B(_2536_),
    .Y(_2616_));
 sky130_fd_sc_hd__nor2_1 _6355_ (.A(_0490_),
    .B(net745),
    .Y(_2617_));
 sky130_fd_sc_hd__a211oi_1 _6356_ (.A1(_0314_),
    .A2(net745),
    .B1(_2617_),
    .C1(net742),
    .Y(_2618_));
 sky130_fd_sc_hd__a211oi_1 _6357_ (.A1(net742),
    .A2(_2589_),
    .B1(_2618_),
    .C1(net740),
    .Y(_2619_));
 sky130_fd_sc_hd__a211oi_1 _6358_ (.A1(net740),
    .A2(_2616_),
    .B1(_2619_),
    .C1(net752),
    .Y(_2620_));
 sky130_fd_sc_hd__a21oi_1 _6359_ (.A1(net752),
    .A2(_2444_),
    .B1(_2620_),
    .Y(_2621_));
 sky130_fd_sc_hd__a211oi_1 _6360_ (.A1(_2022_),
    .A2(_2587_),
    .B1(_2428_),
    .C1(_1716_),
    .Y(_2622_));
 sky130_fd_sc_hd__o21ai_2 _6361_ (.A1(_1870_),
    .A2(_2621_),
    .B1(_2622_),
    .Y(_2623_));
 sky130_fd_sc_hd__a21oi_2 _6362_ (.A1(_2293_),
    .A2(_2303_),
    .B1(_2623_),
    .Y(_2624_));
 sky130_fd_sc_hd__a21oi_2 _6363_ (.A1(_2615_),
    .A2(_2612_),
    .B1(_2624_),
    .Y(net90));
 sky130_fd_sc_hd__nand2b_4 _6364_ (.A_N(net30),
    .B(net31),
    .Y(_2625_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_27 ();
 sky130_fd_sc_hd__or2_4 _6366_ (.A(net31),
    .B(net30),
    .X(_2627_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_26 ();
 sky130_fd_sc_hd__nor2_2 _6368_ (.A(_0036_),
    .B(_0130_),
    .Y(_2629_));
 sky130_fd_sc_hd__nor3_4 _6369_ (.A(_0137_),
    .B(_0896_),
    .C(_2629_),
    .Y(_2630_));
 sky130_fd_sc_hd__nor2_4 _6370_ (.A(net32),
    .B(_2630_),
    .Y(_2631_));
 sky130_fd_sc_hd__nor2_4 _6371_ (.A(net3),
    .B(net2),
    .Y(_2632_));
 sky130_fd_sc_hd__nand3_4 _6372_ (.A(_2627_),
    .B(_2631_),
    .C(_2632_),
    .Y(_2633_));
 sky130_fd_sc_hd__nor2_4 _6373_ (.A(_2625_),
    .B(_2633_),
    .Y(_0021_));
 sky130_fd_sc_hd__nand2_8 _6374_ (.A(net31),
    .B(net30),
    .Y(_2634_));
 sky130_fd_sc_hd__nand3b_1 _6375_ (.A_N(net3),
    .B(net2),
    .C(_2631_),
    .Y(_2635_));
 sky130_fd_sc_hd__nor2_4 _6376_ (.A(_2634_),
    .B(_2635_),
    .Y(_0001_));
 sky130_fd_sc_hd__nor2b_4 _6377_ (.A(_2630_),
    .B_N(net32),
    .Y(_2636_));
 sky130_fd_sc_hd__nand3b_1 _6378_ (.A_N(net2),
    .B(_2636_),
    .C(net3),
    .Y(_2637_));
 sky130_fd_sc_hd__nor2_4 _6379_ (.A(_2627_),
    .B(_2637_),
    .Y(_0011_));
 sky130_fd_sc_hd__nor2_4 _6380_ (.A(_2625_),
    .B(_2635_),
    .Y(_0000_));
 sky130_fd_sc_hd__nand2b_4 _6381_ (.A_N(net31),
    .B(net30),
    .Y(_2638_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__nor2_4 _6383_ (.A(_2635_),
    .B(_2638_),
    .Y(_0030_));
 sky130_fd_sc_hd__nand3b_1 _6384_ (.A_N(net2),
    .B(_2631_),
    .C(net3),
    .Y(_2640_));
 sky130_fd_sc_hd__nor2_4 _6385_ (.A(_2634_),
    .B(_2640_),
    .Y(_0009_));
 sky130_fd_sc_hd__nor2_4 _6386_ (.A(_2627_),
    .B(_2635_),
    .Y(_0029_));
 sky130_fd_sc_hd__nor2_4 _6387_ (.A(_2625_),
    .B(_2640_),
    .Y(_0008_));
 sky130_fd_sc_hd__nor2_4 _6388_ (.A(_2638_),
    .B(_2640_),
    .Y(_0007_));
 sky130_fd_sc_hd__nand2_8 _6389_ (.A(_2632_),
    .B(_2636_),
    .Y(_2641_));
 sky130_fd_sc_hd__nor2_4 _6390_ (.A(_2634_),
    .B(_2641_),
    .Y(_0028_));
 sky130_fd_sc_hd__nor2_4 _6391_ (.A(_2627_),
    .B(_2640_),
    .Y(_0006_));
 sky130_fd_sc_hd__nor2_4 _6392_ (.A(_2625_),
    .B(_2641_),
    .Y(_0027_));
 sky130_fd_sc_hd__nor2_4 _6393_ (.A(_2638_),
    .B(_2641_),
    .Y(_0026_));
 sky130_fd_sc_hd__nand3b_1 _6394_ (.A_N(net3),
    .B(net2),
    .C(_2636_),
    .Y(_2642_));
 sky130_fd_sc_hd__nor2_4 _6395_ (.A(_2634_),
    .B(_2642_),
    .Y(_0005_));
 sky130_fd_sc_hd__nor2_4 _6396_ (.A(_2627_),
    .B(_2641_),
    .Y(_0025_));
 sky130_fd_sc_hd__nor2_4 _6397_ (.A(_2625_),
    .B(_2642_),
    .Y(_0004_));
 sky130_fd_sc_hd__nor2_4 _6398_ (.A(_2638_),
    .B(_2642_),
    .Y(_0003_));
 sky130_fd_sc_hd__nand2_1 _6399_ (.A(_2631_),
    .B(_2632_),
    .Y(_2643_));
 sky130_fd_sc_hd__nor2_4 _6400_ (.A(_2643_),
    .B(_2634_),
    .Y(_0024_));
 sky130_fd_sc_hd__nor2_4 _6401_ (.A(_2627_),
    .B(_2642_),
    .Y(_0002_));
 sky130_fd_sc_hd__nor2_4 _6402_ (.A(_2633_),
    .B(_2638_),
    .Y(_0010_));
 sky130_fd_sc_hd__nand3_4 _6403_ (.A(net3),
    .B(net2),
    .C(_2636_),
    .Y(_2644_));
 sky130_fd_sc_hd__nor2_4 _6404_ (.A(_2634_),
    .B(_2644_),
    .Y(_0023_));
 sky130_fd_sc_hd__nor2_4 _6405_ (.A(_2625_),
    .B(_2644_),
    .Y(_0022_));
 sky130_fd_sc_hd__nor2_4 _6406_ (.A(_2638_),
    .B(_2644_),
    .Y(_0020_));
 sky130_fd_sc_hd__nand3_4 _6407_ (.A(net3),
    .B(net2),
    .C(_2631_),
    .Y(_2645_));
 sky130_fd_sc_hd__nor2_4 _6408_ (.A(_2638_),
    .B(_2645_),
    .Y(_0016_));
 sky130_fd_sc_hd__nor2_4 _6409_ (.A(_2627_),
    .B(_2644_),
    .Y(_0019_));
 sky130_fd_sc_hd__nor2_4 _6410_ (.A(_2625_),
    .B(_2645_),
    .Y(_0017_));
 sky130_fd_sc_hd__nor2_4 _6411_ (.A(_2634_),
    .B(_2645_),
    .Y(_0018_));
 sky130_fd_sc_hd__nor2_4 _6412_ (.A(_2627_),
    .B(_2645_),
    .Y(_0015_));
 sky130_fd_sc_hd__nor2_4 _6413_ (.A(_2634_),
    .B(_2637_),
    .Y(_0014_));
 sky130_fd_sc_hd__nor2_4 _6414_ (.A(_2637_),
    .B(_2638_),
    .Y(_0012_));
 sky130_fd_sc_hd__nor2_4 _6415_ (.A(_2625_),
    .B(_2637_),
    .Y(_0013_));
 sky130_fd_sc_hd__clkinv_16 _6416_ (.A(net65),
    .Y(_0031_));
 sky130_fd_sc_hd__or3_4 _6417_ (.A(net28),
    .B(_0134_),
    .C(_0135_),
    .X(_2646_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__nand3_4 _6419_ (.A(_0901_),
    .B(_0897_),
    .C(_2646_),
    .Y(_2648_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_22 ();
 sky130_fd_sc_hd__nand2_1 _6422_ (.A(net100),
    .B(_2648_),
    .Y(_2651_));
 sky130_fd_sc_hd__o21ai_0 _6423_ (.A1(_0237_),
    .A2(_2648_),
    .B1(_2651_),
    .Y(_3448_[0]));
 sky130_fd_sc_hd__nand2_1 _6424_ (.A(net111),
    .B(_2648_),
    .Y(_2652_));
 sky130_fd_sc_hd__o21ai_2 _6425_ (.A1(_1699_),
    .A2(_2648_),
    .B1(_2652_),
    .Y(_3190_[0]));
 sky130_fd_sc_hd__nand2_1 _6426_ (.A(net122),
    .B(_2648_),
    .Y(_2653_));
 sky130_fd_sc_hd__o21ai_0 _6427_ (.A1(_3438_[0]),
    .A2(_2648_),
    .B1(_2653_),
    .Y(_3453_[0]));
 sky130_fd_sc_hd__nand2_1 _6428_ (.A(net125),
    .B(_2648_),
    .Y(_2654_));
 sky130_fd_sc_hd__o21ai_0 _6429_ (.A1(_3430_[0]),
    .A2(_2648_),
    .B1(_2654_),
    .Y(_3457_[0]));
 sky130_fd_sc_hd__nand2_1 _6430_ (.A(net126),
    .B(_2648_),
    .Y(_2655_));
 sky130_fd_sc_hd__o21ai_2 _6431_ (.A1(_3422_[0]),
    .A2(_2648_),
    .B1(_2655_),
    .Y(_3463_[0]));
 sky130_fd_sc_hd__nand2_1 _6432_ (.A(net127),
    .B(_2648_),
    .Y(_2656_));
 sky130_fd_sc_hd__o21ai_2 _6433_ (.A1(_3414_[0]),
    .A2(_2648_),
    .B1(_2656_),
    .Y(_3467_[0]));
 sky130_fd_sc_hd__nand2_1 _6434_ (.A(net128),
    .B(_2648_),
    .Y(_2657_));
 sky130_fd_sc_hd__o21ai_2 _6435_ (.A1(_3406_[0]),
    .A2(_2648_),
    .B1(_2657_),
    .Y(_3471_[0]));
 sky130_fd_sc_hd__nand2_1 _6436_ (.A(net129),
    .B(_2648_),
    .Y(_2658_));
 sky130_fd_sc_hd__o21ai_2 _6437_ (.A1(_3398_[0]),
    .A2(_2648_),
    .B1(_2658_),
    .Y(_3475_[0]));
 sky130_fd_sc_hd__nand2_1 _6438_ (.A(net130),
    .B(_2648_),
    .Y(_2659_));
 sky130_fd_sc_hd__o21ai_0 _6439_ (.A1(_1405_),
    .A2(_2648_),
    .B1(_2659_),
    .Y(_3479_[0]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_21 ();
 sky130_fd_sc_hd__nand2_1 _6441_ (.A(net131),
    .B(_2648_),
    .Y(_2661_));
 sky130_fd_sc_hd__o21ai_0 _6442_ (.A1(_1364_),
    .A2(_2648_),
    .B1(_2661_),
    .Y(_3483_[0]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_20 ();
 sky130_fd_sc_hd__nand2_1 _6444_ (.A(net101),
    .B(_2648_),
    .Y(_2663_));
 sky130_fd_sc_hd__o21ai_0 _6445_ (.A1(_3374_[0]),
    .A2(_2648_),
    .B1(_2663_),
    .Y(_3487_[0]));
 sky130_fd_sc_hd__nand2_1 _6446_ (.A(net102),
    .B(_2648_),
    .Y(_2664_));
 sky130_fd_sc_hd__o21ai_0 _6447_ (.A1(_3366_[0]),
    .A2(_2648_),
    .B1(_2664_),
    .Y(_3491_[0]));
 sky130_fd_sc_hd__nand2_1 _6448_ (.A(net103),
    .B(_2648_),
    .Y(_2665_));
 sky130_fd_sc_hd__o21ai_0 _6449_ (.A1(_3358_[0]),
    .A2(_2648_),
    .B1(_2665_),
    .Y(_3495_[0]));
 sky130_fd_sc_hd__nand2_1 _6450_ (.A(net104),
    .B(_2648_),
    .Y(_2666_));
 sky130_fd_sc_hd__o21ai_0 _6451_ (.A1(_1203_),
    .A2(_2648_),
    .B1(_2666_),
    .Y(_3499_[0]));
 sky130_fd_sc_hd__nand2_1 _6452_ (.A(net105),
    .B(_2648_),
    .Y(_2667_));
 sky130_fd_sc_hd__o21ai_0 _6453_ (.A1(_3342_[0]),
    .A2(_2648_),
    .B1(_2667_),
    .Y(_3503_[0]));
 sky130_fd_sc_hd__nand2_1 _6454_ (.A(net106),
    .B(_2648_),
    .Y(_2668_));
 sky130_fd_sc_hd__o21ai_0 _6455_ (.A1(_3334_[0]),
    .A2(_2648_),
    .B1(_2668_),
    .Y(_3507_[0]));
 sky130_fd_sc_hd__nand2_1 _6456_ (.A(net107),
    .B(_2648_),
    .Y(_2669_));
 sky130_fd_sc_hd__o21ai_2 _6457_ (.A1(_3326_[0]),
    .A2(_2648_),
    .B1(_2669_),
    .Y(_3511_[0]));
 sky130_fd_sc_hd__nand2_1 _6458_ (.A(net108),
    .B(_2648_),
    .Y(_2670_));
 sky130_fd_sc_hd__o21ai_0 _6459_ (.A1(_3318_[0]),
    .A2(_2648_),
    .B1(_2670_),
    .Y(_3515_[0]));
 sky130_fd_sc_hd__nand2_1 _6460_ (.A(net109),
    .B(_2648_),
    .Y(_2671_));
 sky130_fd_sc_hd__o21ai_2 _6461_ (.A1(_3310_[0]),
    .A2(_2648_),
    .B1(_2671_),
    .Y(_3519_[0]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_19 ();
 sky130_fd_sc_hd__nand2_1 _6463_ (.A(net110),
    .B(_2648_),
    .Y(_2673_));
 sky130_fd_sc_hd__o21ai_0 _6464_ (.A1(_3302_[0]),
    .A2(_2648_),
    .B1(_2673_),
    .Y(_3523_[0]));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_18 ();
 sky130_fd_sc_hd__nand2_1 _6466_ (.A(net112),
    .B(_2648_),
    .Y(_2675_));
 sky130_fd_sc_hd__o21ai_0 _6467_ (.A1(_3294_[0]),
    .A2(_2648_),
    .B1(_2675_),
    .Y(_3527_[0]));
 sky130_fd_sc_hd__nand2_1 _6468_ (.A(net113),
    .B(_2648_),
    .Y(_2676_));
 sky130_fd_sc_hd__o21ai_0 _6469_ (.A1(_3286_[0]),
    .A2(_2648_),
    .B1(_2676_),
    .Y(_3531_[0]));
 sky130_fd_sc_hd__nand2_1 _6470_ (.A(net114),
    .B(_2648_),
    .Y(_2677_));
 sky130_fd_sc_hd__o21ai_0 _6471_ (.A1(_3278_[0]),
    .A2(_2648_),
    .B1(_2677_),
    .Y(_3535_[0]));
 sky130_fd_sc_hd__nand2_1 _6472_ (.A(net115),
    .B(net776),
    .Y(_2678_));
 sky130_fd_sc_hd__o21ai_0 _6473_ (.A1(_3270_[0]),
    .A2(net776),
    .B1(_2678_),
    .Y(_3539_[0]));
 sky130_fd_sc_hd__nand2_1 _6474_ (.A(net116),
    .B(net776),
    .Y(_2679_));
 sky130_fd_sc_hd__o21ai_0 _6475_ (.A1(_3262_[0]),
    .A2(net776),
    .B1(_2679_),
    .Y(_3543_[0]));
 sky130_fd_sc_hd__nand2_1 _6476_ (.A(net117),
    .B(net776),
    .Y(_2680_));
 sky130_fd_sc_hd__o21ai_0 _6477_ (.A1(_3254_[0]),
    .A2(net776),
    .B1(_2680_),
    .Y(_3547_[0]));
 sky130_fd_sc_hd__nand2_1 _6478_ (.A(net118),
    .B(net776),
    .Y(_2681_));
 sky130_fd_sc_hd__o21ai_2 _6479_ (.A1(_3246_[0]),
    .A2(net776),
    .B1(_2681_),
    .Y(_3551_[0]));
 sky130_fd_sc_hd__nand2_1 _6480_ (.A(net119),
    .B(net776),
    .Y(_2682_));
 sky130_fd_sc_hd__o21ai_2 _6481_ (.A1(net766),
    .A2(net776),
    .B1(_2682_),
    .Y(_3555_[0]));
 sky130_fd_sc_hd__nand2_1 _6482_ (.A(net120),
    .B(net776),
    .Y(_2683_));
 sky130_fd_sc_hd__o21ai_2 _6483_ (.A1(_3230_[0]),
    .A2(net776),
    .B1(_2683_),
    .Y(_3559_[0]));
 sky130_fd_sc_hd__nand2_1 _6484_ (.A(net121),
    .B(net776),
    .Y(_2684_));
 sky130_fd_sc_hd__o21ai_2 _6485_ (.A1(_3222_[0]),
    .A2(net776),
    .B1(_2684_),
    .Y(_3563_[0]));
 sky130_fd_sc_hd__nand2_1 _6486_ (.A(net123),
    .B(net776),
    .Y(_2685_));
 sky130_fd_sc_hd__o21ai_0 _6487_ (.A1(net767),
    .A2(net776),
    .B1(_2685_),
    .Y(_3567_[0]));
 sky130_fd_sc_hd__nand2_1 _6488_ (.A(_1216_),
    .B(_1217_),
    .Y(_3496_[0]));
 sky130_fd_sc_hd__nand2_8 _6489_ (.A(_0143_),
    .B(_0118_),
    .Y(_2686_));
 sky130_fd_sc_hd__nand2_2 _6490_ (.A(net159),
    .B(net753),
    .Y(_2687_));
 sky130_fd_sc_hd__nand2_1 _6491_ (.A(net247),
    .B(_3438_[0]),
    .Y(_2688_));
 sky130_fd_sc_hd__nand2_1 _6492_ (.A(net144),
    .B(_1699_),
    .Y(_2689_));
 sky130_fd_sc_hd__o22ai_1 _6493_ (.A1(net133),
    .A2(_0237_),
    .B1(net144),
    .B2(_1699_),
    .Y(_2690_));
 sky130_fd_sc_hd__nand3_1 _6494_ (.A(_2688_),
    .B(_2689_),
    .C(_2690_),
    .Y(_2691_));
 sky130_fd_sc_hd__o221ai_1 _6495_ (.A1(net222),
    .A2(_3430_[0]),
    .B1(net240),
    .B2(_3438_[0]),
    .C1(_2691_),
    .Y(_2692_));
 sky130_fd_sc_hd__nand2_1 _6496_ (.A(net223),
    .B(_3430_[0]),
    .Y(_2693_));
 sky130_fd_sc_hd__o22ai_2 _6497_ (.A1(net160),
    .A2(net754),
    .B1(net330),
    .B2(net753),
    .Y(_2694_));
 sky130_fd_sc_hd__a31oi_2 _6498_ (.A1(_2687_),
    .A2(_2692_),
    .A3(_2693_),
    .B1(_2694_),
    .Y(_2695_));
 sky130_fd_sc_hd__nor2_2 _6499_ (.A(_1253_),
    .B(_3366_[0]),
    .Y(_2696_));
 sky130_fd_sc_hd__o21ai_2 _6500_ (.A1(_0492_),
    .A2(_1329_),
    .B1(_1335_),
    .Y(_2697_));
 sky130_fd_sc_hd__clkinv_1 _6501_ (.A(_1377_),
    .Y(_2698_));
 sky130_fd_sc_hd__a221oi_1 _6502_ (.A1(_2697_),
    .A2(_1364_),
    .B1(_2698_),
    .B2(net757),
    .C1(_3374_[0]),
    .Y(_2699_));
 sky130_fd_sc_hd__nor3_1 _6503_ (.A(_3374_[0]),
    .B(_2697_),
    .C(_1364_),
    .Y(_2700_));
 sky130_fd_sc_hd__nor4_2 _6504_ (.A(_1295_),
    .B(_2696_),
    .C(_2699_),
    .D(_2700_),
    .Y(_2701_));
 sky130_fd_sc_hd__a21oi_1 _6505_ (.A1(_2698_),
    .A2(net757),
    .B1(_1364_),
    .Y(_2702_));
 sky130_fd_sc_hd__a31oi_1 _6506_ (.A1(_1364_),
    .A2(_2698_),
    .A3(net757),
    .B1(_2697_),
    .Y(_2703_));
 sky130_fd_sc_hd__nand2_2 _6507_ (.A(_1253_),
    .B(_3366_[0]),
    .Y(_2704_));
 sky130_fd_sc_hd__o41ai_2 _6508_ (.A1(_3370_[0]),
    .A2(_2696_),
    .A3(_2702_),
    .A4(_2703_),
    .B1(_2704_),
    .Y(_2705_));
 sky130_fd_sc_hd__nor2_2 _6509_ (.A(_2701_),
    .B(_2705_),
    .Y(_2706_));
 sky130_fd_sc_hd__nand2_4 _6510_ (.A(net160),
    .B(net754),
    .Y(_2707_));
 sky130_fd_sc_hd__nand2_2 _6511_ (.A(net162),
    .B(net756),
    .Y(_2708_));
 sky130_fd_sc_hd__nand2_1 _6512_ (.A(net161),
    .B(net755),
    .Y(_2709_));
 sky130_fd_sc_hd__nand4_1 _6513_ (.A(_2706_),
    .B(_2707_),
    .C(_2708_),
    .D(_2709_),
    .Y(_2710_));
 sky130_fd_sc_hd__nor2_4 _6514_ (.A(net162),
    .B(net756),
    .Y(_2711_));
 sky130_fd_sc_hd__nor2_1 _6515_ (.A(net160),
    .B(net754),
    .Y(_2712_));
 sky130_fd_sc_hd__o21a_1 _6516_ (.A1(_2712_),
    .A2(_2687_),
    .B1(_2707_),
    .X(_2713_));
 sky130_fd_sc_hd__nor3_1 _6517_ (.A(_3402_[0]),
    .B(_2711_),
    .C(_2713_),
    .Y(_2714_));
 sky130_fd_sc_hd__nand2_1 _6518_ (.A(_3418_[0]),
    .B(_2707_),
    .Y(_2715_));
 sky130_fd_sc_hd__nand2_1 _6519_ (.A(net209),
    .B(_3426_[0]),
    .Y(_2716_));
 sky130_fd_sc_hd__o211ai_1 _6520_ (.A1(net240),
    .A2(_3438_[0]),
    .B1(net144),
    .C1(_1699_),
    .Y(_2717_));
 sky130_fd_sc_hd__o2111ai_1 _6521_ (.A1(net775),
    .A2(_1699_),
    .B1(net133),
    .C1(_0237_),
    .D1(_3438_[0]),
    .Y(_2718_));
 sky130_fd_sc_hd__o2111ai_1 _6522_ (.A1(net775),
    .A2(_1699_),
    .B1(net133),
    .C1(_0237_),
    .D1(net240),
    .Y(_2719_));
 sky130_fd_sc_hd__a32oi_2 _6523_ (.A1(_1592_),
    .A2(net158),
    .A3(_1609_),
    .B1(net240),
    .B2(_3438_[0]),
    .Y(_2720_));
 sky130_fd_sc_hd__nand4_1 _6524_ (.A(_2717_),
    .B(_2718_),
    .C(_2719_),
    .D(_2720_),
    .Y(_2721_));
 sky130_fd_sc_hd__nor3_1 _6525_ (.A(_3402_[0]),
    .B(_2712_),
    .C(_2711_),
    .Y(_2722_));
 sky130_fd_sc_hd__o2111a_4 _6526_ (.A1(net159),
    .A2(_2715_),
    .B1(_2716_),
    .C1(_2721_),
    .D1(_2722_),
    .X(_2723_));
 sky130_fd_sc_hd__nand4_1 _6527_ (.A(_3402_[0]),
    .B(_2687_),
    .C(_2707_),
    .D(_2708_),
    .Y(_2724_));
 sky130_fd_sc_hd__a21oi_1 _6528_ (.A1(_1592_),
    .A2(_1609_),
    .B1(net222),
    .Y(_2725_));
 sky130_fd_sc_hd__a41oi_2 _6529_ (.A1(_2720_),
    .A2(_2718_),
    .A3(_2719_),
    .A4(_2717_),
    .B1(_2725_),
    .Y(_2726_));
 sky130_fd_sc_hd__o21ai_0 _6530_ (.A1(net162),
    .A2(net756),
    .B1(net161),
    .Y(_2727_));
 sky130_fd_sc_hd__a31o_1 _6531_ (.A1(_3402_[0]),
    .A2(_2694_),
    .A3(_2707_),
    .B1(_2727_),
    .X(_2728_));
 sky130_fd_sc_hd__a2bb2oi_2 _6532_ (.A1_N(_2726_),
    .A2_N(_2724_),
    .B1(_2708_),
    .B2(_2728_),
    .Y(_2729_));
 sky130_fd_sc_hd__nor3_4 _6533_ (.A(_2714_),
    .B(_2729_),
    .C(_2723_),
    .Y(_2730_));
 sky130_fd_sc_hd__nor2_1 _6534_ (.A(_2698_),
    .B(net757),
    .Y(_2731_));
 sky130_fd_sc_hd__maj3_1 _6535_ (.A(_1336_),
    .B(_3378_[0]),
    .C(_2731_),
    .X(_2732_));
 sky130_fd_sc_hd__a211o_1 _6536_ (.A1(_1295_),
    .A2(_3370_[0]),
    .B1(_2696_),
    .C1(_2732_),
    .X(_2733_));
 sky130_fd_sc_hd__or3_1 _6537_ (.A(_1295_),
    .B(_3370_[0]),
    .C(_2696_),
    .X(_2734_));
 sky130_fd_sc_hd__o21ai_0 _6538_ (.A1(_1215_),
    .A2(net761),
    .B1(_1203_),
    .Y(_2735_));
 sky130_fd_sc_hd__o31ai_1 _6539_ (.A1(_1203_),
    .A2(_1215_),
    .A3(net761),
    .B1(_1173_),
    .Y(_2736_));
 sky130_fd_sc_hd__nor2_1 _6540_ (.A(_1088_),
    .B(_3334_[0]),
    .Y(_2737_));
 sky130_fd_sc_hd__a311oi_1 _6541_ (.A1(_3338_[0]),
    .A2(_2735_),
    .A3(_2736_),
    .B1(_2737_),
    .C1(_1125_),
    .Y(_2738_));
 sky130_fd_sc_hd__a211oi_1 _6542_ (.A1(_2735_),
    .A2(_2736_),
    .B1(_3338_[0]),
    .C1(_2737_),
    .Y(_2739_));
 sky130_fd_sc_hd__a211oi_2 _6543_ (.A1(_1088_),
    .A2(net763),
    .B1(_2738_),
    .C1(_2739_),
    .Y(_2740_));
 sky130_fd_sc_hd__a31oi_2 _6544_ (.A1(_2704_),
    .A2(_2733_),
    .A3(_2734_),
    .B1(_2740_),
    .Y(_2741_));
 sky130_fd_sc_hd__nor2_2 _6545_ (.A(_0732_),
    .B(_3266_[0]),
    .Y(_2742_));
 sky130_fd_sc_hd__a21oi_4 _6546_ (.A1(_0774_),
    .A2(_0780_),
    .B1(_0111_),
    .Y(_2743_));
 sky130_fd_sc_hd__o21ai_0 _6547_ (.A1(_0886_),
    .A2(_0895_),
    .B1(_0866_),
    .Y(_2744_));
 sky130_fd_sc_hd__maj3_1 _6548_ (.A(_0821_),
    .B(_3286_[0]),
    .C(_2744_),
    .X(_2745_));
 sky130_fd_sc_hd__maj3_1 _6549_ (.A(_2743_),
    .B(_3278_[0]),
    .C(_2745_),
    .X(_2746_));
 sky130_fd_sc_hd__nand2_2 _6550_ (.A(_0732_),
    .B(_3266_[0]),
    .Y(_2747_));
 sky130_fd_sc_hd__o21ai_2 _6551_ (.A1(_2742_),
    .A2(_2746_),
    .B1(_2747_),
    .Y(_2748_));
 sky130_fd_sc_hd__clkinvlp_2 _6552_ (.A(_0917_),
    .Y(_2749_));
 sky130_fd_sc_hd__nor2b_1 _6553_ (.A(_0952_),
    .B_N(_3310_[0]),
    .Y(_2750_));
 sky130_fd_sc_hd__a21oi_4 _6554_ (.A1(_0986_),
    .A2(_0992_),
    .B1(_0111_),
    .Y(_2751_));
 sky130_fd_sc_hd__nor3_1 _6555_ (.A(_1039_),
    .B(_1063_),
    .C(_1072_),
    .Y(_2752_));
 sky130_fd_sc_hd__maj3_1 _6556_ (.A(_2751_),
    .B(net764),
    .C(_2752_),
    .X(_2753_));
 sky130_fd_sc_hd__nand2b_1 _6557_ (.A_N(_3310_[0]),
    .B(_0952_),
    .Y(_2754_));
 sky130_fd_sc_hd__o21ai_0 _6558_ (.A1(_2750_),
    .A2(_2753_),
    .B1(_2754_),
    .Y(_2755_));
 sky130_fd_sc_hd__maj3_1 _6559_ (.A(_2749_),
    .B(_3298_[0]),
    .C(_2755_),
    .X(_2756_));
 sky130_fd_sc_hd__inv_1 _6560_ (.A(_1125_),
    .Y(_2757_));
 sky130_fd_sc_hd__a22o_1 _6561_ (.A1(_1173_),
    .A2(_1203_),
    .B1(_1215_),
    .B2(net761),
    .X(_2758_));
 sky130_fd_sc_hd__o22a_1 _6562_ (.A1(_2757_),
    .A2(_3342_[0]),
    .B1(_1173_),
    .B2(_1203_),
    .X(_2759_));
 sky130_fd_sc_hd__a222oi_1 _6563_ (.A1(_1088_),
    .A2(net763),
    .B1(_2757_),
    .B2(_3342_[0]),
    .C1(_2758_),
    .C2(_2759_),
    .Y(_2760_));
 sky130_fd_sc_hd__or2_4 _6564_ (.A(_2737_),
    .B(_2760_),
    .X(_2761_));
 sky130_fd_sc_hd__nor2_2 _6565_ (.A(net161),
    .B(net755),
    .Y(_2762_));
 sky130_fd_sc_hd__nor4_2 _6566_ (.A(_2701_),
    .B(_2705_),
    .C(_2711_),
    .D(_2762_),
    .Y(_2763_));
 sky130_fd_sc_hd__nor3_1 _6567_ (.A(_0866_),
    .B(_0886_),
    .C(_0895_),
    .Y(_2764_));
 sky130_fd_sc_hd__maj3_1 _6568_ (.A(_0821_),
    .B(_3286_[0]),
    .C(_2764_),
    .X(_2765_));
 sky130_fd_sc_hd__maj3_2 _6569_ (.A(_2743_),
    .B(_3278_[0]),
    .C(_2765_),
    .X(_2766_));
 sky130_fd_sc_hd__a21oi_2 _6570_ (.A1(_2747_),
    .A2(_2766_),
    .B1(_2742_),
    .Y(_2767_));
 sky130_fd_sc_hd__o2111a_4 _6571_ (.A1(_2748_),
    .A2(_2756_),
    .B1(_2761_),
    .C1(_2763_),
    .D1(_2767_),
    .X(_2768_));
 sky130_fd_sc_hd__o2111ai_4 _6572_ (.A1(_2695_),
    .A2(_2710_),
    .B1(_2768_),
    .C1(_2741_),
    .D1(_2730_),
    .Y(_2769_));
 sky130_fd_sc_hd__xnor2_1 _6573_ (.A(_0314_),
    .B(_0338_),
    .Y(_2770_));
 sky130_fd_sc_hd__nor2_1 _6574_ (.A(_0369_),
    .B(_3210_[0]),
    .Y(_2771_));
 sky130_fd_sc_hd__nand2_1 _6575_ (.A(net5),
    .B(_0139_),
    .Y(_2772_));
 sky130_fd_sc_hd__nor2_1 _6576_ (.A(_0338_),
    .B(_2772_),
    .Y(_2773_));
 sky130_fd_sc_hd__and3_1 _6577_ (.A(_0313_),
    .B(_0338_),
    .C(_2772_),
    .X(_2774_));
 sky130_fd_sc_hd__a221oi_1 _6578_ (.A1(_2770_),
    .A2(_2771_),
    .B1(_2773_),
    .B2(_0314_),
    .C1(_2774_),
    .Y(_2775_));
 sky130_fd_sc_hd__inv_1 _6579_ (.A(_0369_),
    .Y(_2776_));
 sky130_fd_sc_hd__o21ai_0 _6580_ (.A1(_0610_),
    .A2(_0622_),
    .B1(_0598_),
    .Y(_2777_));
 sky130_fd_sc_hd__maj3_1 _6581_ (.A(_0543_),
    .B(net766),
    .C(_2777_),
    .X(_2778_));
 sky130_fd_sc_hd__nor3_1 _6582_ (.A(_0690_),
    .B(_0706_),
    .C(_0719_),
    .Y(_2779_));
 sky130_fd_sc_hd__maj3_1 _6583_ (.A(_0637_),
    .B(_3254_[0]),
    .C(_2779_),
    .X(_2780_));
 sky130_fd_sc_hd__o21ai_0 _6584_ (.A1(_0447_),
    .A2(_0490_),
    .B1(_3226_[0]),
    .Y(_2781_));
 sky130_fd_sc_hd__o21a_4 _6585_ (.A1(_0492_),
    .A2(_0501_),
    .B1(_0507_),
    .X(_2782_));
 sky130_fd_sc_hd__o21ai_0 _6586_ (.A1(_0447_),
    .A2(_0490_),
    .B1(_2782_),
    .Y(_2783_));
 sky130_fd_sc_hd__nor3_1 _6587_ (.A(_0598_),
    .B(_0610_),
    .C(_0622_),
    .Y(_2784_));
 sky130_fd_sc_hd__maj3_2 _6588_ (.A(_0543_),
    .B(net766),
    .C(_2784_),
    .X(_2785_));
 sky130_fd_sc_hd__a221oi_2 _6589_ (.A1(_2778_),
    .A2(_2780_),
    .B1(_2781_),
    .B2(_2783_),
    .C1(_2785_),
    .Y(_2786_));
 sky130_fd_sc_hd__nor2_1 _6590_ (.A(_0447_),
    .B(_0490_),
    .Y(_2787_));
 sky130_fd_sc_hd__nand2_1 _6591_ (.A(_0447_),
    .B(_0490_),
    .Y(_2788_));
 sky130_fd_sc_hd__o31ai_1 _6592_ (.A1(_0508_),
    .A2(_3230_[0]),
    .A3(_2787_),
    .B1(_2788_),
    .Y(_2789_));
 sky130_fd_sc_hd__nor2_2 _6593_ (.A(_2786_),
    .B(_2789_),
    .Y(_2790_));
 sky130_fd_sc_hd__o211ai_1 _6594_ (.A1(_2776_),
    .A2(net767),
    .B1(_2770_),
    .C1(_2790_),
    .Y(_2791_));
 sky130_fd_sc_hd__nand2_1 _6595_ (.A(_2775_),
    .B(_2791_),
    .Y(_2792_));
 sky130_fd_sc_hd__o21ai_0 _6596_ (.A1(_0706_),
    .A2(_0719_),
    .B1(_0690_),
    .Y(_2793_));
 sky130_fd_sc_hd__maj3_1 _6597_ (.A(_0637_),
    .B(_3254_[0]),
    .C(_2793_),
    .X(_2794_));
 sky130_fd_sc_hd__a21oi_1 _6598_ (.A1(_0447_),
    .A2(_0490_),
    .B1(_3226_[0]),
    .Y(_2795_));
 sky130_fd_sc_hd__a21oi_1 _6599_ (.A1(_0447_),
    .A2(_0490_),
    .B1(_2782_),
    .Y(_2796_));
 sky130_fd_sc_hd__o221a_4 _6600_ (.A1(_2785_),
    .A2(_2794_),
    .B1(_2795_),
    .B2(_2796_),
    .C1(_2778_),
    .X(_2797_));
 sky130_fd_sc_hd__a311oi_2 _6601_ (.A1(_0508_),
    .A2(_3230_[0]),
    .A3(_2788_),
    .B1(_2787_),
    .C1(_2797_),
    .Y(_2798_));
 sky130_fd_sc_hd__o21ai_0 _6602_ (.A1(_2776_),
    .A2(net767),
    .B1(_2770_),
    .Y(_2799_));
 sky130_fd_sc_hd__o21ai_0 _6603_ (.A1(_2798_),
    .A2(_2799_),
    .B1(_2775_),
    .Y(_2800_));
 sky130_fd_sc_hd__o21ai_0 _6604_ (.A1(_1063_),
    .A2(_1072_),
    .B1(_1039_),
    .Y(_2801_));
 sky130_fd_sc_hd__maj3_1 _6605_ (.A(_2751_),
    .B(net764),
    .C(_2801_),
    .X(_2802_));
 sky130_fd_sc_hd__a211oi_1 _6606_ (.A1(_0917_),
    .A2(net765),
    .B1(_2750_),
    .C1(_2802_),
    .Y(_2803_));
 sky130_fd_sc_hd__a21oi_1 _6607_ (.A1(_0917_),
    .A2(net765),
    .B1(_2754_),
    .Y(_2804_));
 sky130_fd_sc_hd__a211o_1 _6608_ (.A1(_2749_),
    .A2(_3298_[0]),
    .B1(_2803_),
    .C1(_2804_),
    .X(_2805_));
 sky130_fd_sc_hd__a21oi_1 _6609_ (.A1(_2767_),
    .A2(_2805_),
    .B1(_2748_),
    .Y(_2806_));
 sky130_fd_sc_hd__nand2_1 _6610_ (.A(_2800_),
    .B(_2806_),
    .Y(_2807_));
 sky130_fd_sc_hd__o31ai_1 _6611_ (.A1(_2769_),
    .A2(_2792_),
    .A3(_2807_),
    .B1(net815),
    .Y(_2808_));
 sky130_fd_sc_hd__or4_1 _6612_ (.A(net815),
    .B(_2792_),
    .C(_2769_),
    .D(_2807_),
    .X(_2809_));
 sky130_fd_sc_hd__a2111o_1 _6613_ (.A1(_2809_),
    .A2(_2808_),
    .B1(net814),
    .C1(net5),
    .D1(_0901_),
    .X(_2810_));
 sky130_fd_sc_hd__nor2_1 _6614_ (.A(_0901_),
    .B(_1706_),
    .Y(_2811_));
 sky130_fd_sc_hd__nor3b_1 _6615_ (.A(net815),
    .B(_0901_),
    .C_N(net814),
    .Y(_2812_));
 sky130_fd_sc_hd__or3_4 _6616_ (.A(_2714_),
    .B(_2723_),
    .C(_2729_),
    .X(_2813_));
 sky130_fd_sc_hd__o21ai_0 _6617_ (.A1(_2706_),
    .A2(_2740_),
    .B1(_2761_),
    .Y(_2814_));
 sky130_fd_sc_hd__a21oi_2 _6618_ (.A1(_2813_),
    .A2(_2741_),
    .B1(_2814_),
    .Y(_2815_));
 sky130_fd_sc_hd__o21ai_0 _6619_ (.A1(_2748_),
    .A2(_2756_),
    .B1(_2767_),
    .Y(_2816_));
 sky130_fd_sc_hd__nand2_1 _6620_ (.A(_2816_),
    .B(_2800_),
    .Y(_2817_));
 sky130_fd_sc_hd__and2_0 _6621_ (.A(_2775_),
    .B(_2791_),
    .X(_2818_));
 sky130_fd_sc_hd__o211ai_1 _6622_ (.A1(_2807_),
    .A2(_2815_),
    .B1(_2817_),
    .C1(_2818_),
    .Y(_2819_));
 sky130_fd_sc_hd__mux2i_1 _6623_ (.A0(_2811_),
    .A1(_2812_),
    .S(_2819_),
    .Y(_2820_));
 sky130_fd_sc_hd__nand3_4 _6624_ (.A(_2686_),
    .B(_2810_),
    .C(_2820_),
    .Y(_2821_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_17 ();
 sky130_fd_sc_hd__mux2_1 _6626_ (.A0(net100),
    .A1(_3450_[0]),
    .S(net241),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _6627_ (.A0(net111),
    .A1(_3193_[0]),
    .S(net241),
    .X(_0033_));
 sky130_fd_sc_hd__nand3_4 _6628_ (.A(net126),
    .B(_3461_[0]),
    .C(net127),
    .Y(_2823_));
 sky130_fd_sc_hd__nand2_2 _6629_ (.A(net128),
    .B(net129),
    .Y(_2824_));
 sky130_fd_sc_hd__nor2_2 _6630_ (.A(_2823_),
    .B(_2824_),
    .Y(_2825_));
 sky130_fd_sc_hd__nand3_1 _6631_ (.A(net130),
    .B(net131),
    .C(_2825_),
    .Y(_2826_));
 sky130_fd_sc_hd__xor2_1 _6632_ (.A(net101),
    .B(_2826_),
    .X(_2827_));
 sky130_fd_sc_hd__a21o_1 _6633_ (.A1(_3482_[0]),
    .A2(_3477_[0]),
    .B1(_3481_[0]),
    .X(_2828_));
 sky130_fd_sc_hd__a21oi_2 _6634_ (.A1(_3486_[0]),
    .A2(_2828_),
    .B1(_3485_[0]),
    .Y(_2829_));
 sky130_fd_sc_hd__o21a_4 _6635_ (.A1(_3470_[0]),
    .A2(_3469_[0]),
    .B1(_3474_[0]),
    .X(_2830_));
 sky130_fd_sc_hd__o21ai_2 _6636_ (.A1(_3473_[0]),
    .A2(_2830_),
    .B1(_3478_[0]),
    .Y(_2831_));
 sky130_fd_sc_hd__nand2_1 _6637_ (.A(_3482_[0]),
    .B(_3486_[0]),
    .Y(_2832_));
 sky130_fd_sc_hd__nor2_1 _6638_ (.A(_2831_),
    .B(_2832_),
    .Y(_2833_));
 sky130_fd_sc_hd__inv_2 _6639_ (.A(_3466_[0]),
    .Y(_2834_));
 sky130_fd_sc_hd__a21o_1 _6640_ (.A1(_3192_[0]),
    .A2(_3456_[0]),
    .B1(_3455_[0]),
    .X(_2835_));
 sky130_fd_sc_hd__a21oi_4 _6641_ (.A1(_3460_[0]),
    .A2(_2835_),
    .B1(_3459_[0]),
    .Y(_2836_));
 sky130_fd_sc_hd__nor3_4 _6642_ (.A(_3465_[0]),
    .B(_3469_[0]),
    .C(_3473_[0]),
    .Y(_2837_));
 sky130_fd_sc_hd__o21ai_4 _6643_ (.A1(_2834_),
    .A2(_2836_),
    .B1(_2837_),
    .Y(_2838_));
 sky130_fd_sc_hd__nand2_1 _6644_ (.A(_2833_),
    .B(_2838_),
    .Y(_2839_));
 sky130_fd_sc_hd__nand2_1 _6645_ (.A(_2829_),
    .B(_2839_),
    .Y(_2840_));
 sky130_fd_sc_hd__xnor2_1 _6646_ (.A(_3490_[0]),
    .B(_2840_),
    .Y(_2841_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_16 ();
 sky130_fd_sc_hd__mux2i_1 _6648_ (.A0(_2827_),
    .A1(_2841_),
    .S(net701),
    .Y(\dp.ISRmux.d0[10] ));
 sky130_fd_sc_hd__nand3_2 _6649_ (.A(net126),
    .B(net127),
    .C(net128),
    .Y(_2843_));
 sky130_fd_sc_hd__nand2_2 _6650_ (.A(net122),
    .B(net125),
    .Y(_2844_));
 sky130_fd_sc_hd__nor2_4 _6651_ (.A(_2843_),
    .B(_2844_),
    .Y(_2845_));
 sky130_fd_sc_hd__nand2_2 _6652_ (.A(net129),
    .B(_2845_),
    .Y(_2846_));
 sky130_fd_sc_hd__nand3_1 _6653_ (.A(net130),
    .B(net131),
    .C(net101),
    .Y(_2847_));
 sky130_fd_sc_hd__nor2_1 _6654_ (.A(_2846_),
    .B(_2847_),
    .Y(_2848_));
 sky130_fd_sc_hd__xnor2_1 _6655_ (.A(net102),
    .B(_2848_),
    .Y(_2849_));
 sky130_fd_sc_hd__o2111ai_2 _6656_ (.A1(_3473_[0]),
    .A2(_2830_),
    .B1(_3478_[0]),
    .C1(_3482_[0]),
    .D1(_3486_[0]),
    .Y(_2850_));
 sky130_fd_sc_hd__a21oi_1 _6657_ (.A1(_3189_[0]),
    .A2(_3452_[0]),
    .B1(_3451_[0]),
    .Y(_2851_));
 sky130_fd_sc_hd__nand4b_1 _6658_ (.A_N(_2851_),
    .B(_3466_[0]),
    .C(_3460_[0]),
    .D(_3456_[0]),
    .Y(_2852_));
 sky130_fd_sc_hd__a21o_4 _6659_ (.A1(_3460_[0]),
    .A2(_3455_[0]),
    .B1(_3459_[0]),
    .X(_2853_));
 sky130_fd_sc_hd__nand2_4 _6660_ (.A(_3466_[0]),
    .B(_2853_),
    .Y(_2854_));
 sky130_fd_sc_hd__and3_4 _6661_ (.A(_2837_),
    .B(_2852_),
    .C(_2854_),
    .X(_2855_));
 sky130_fd_sc_hd__o21ai_1 _6662_ (.A1(_2850_),
    .A2(_2855_),
    .B1(_2829_),
    .Y(_2856_));
 sky130_fd_sc_hd__a21oi_1 _6663_ (.A1(_3490_[0]),
    .A2(_2856_),
    .B1(_3489_[0]),
    .Y(_2857_));
 sky130_fd_sc_hd__xor2_1 _6664_ (.A(_3494_[0]),
    .B(_2857_),
    .X(_2858_));
 sky130_fd_sc_hd__mux2i_1 _6665_ (.A0(_2849_),
    .A1(_2858_),
    .S(net237),
    .Y(\dp.ISRmux.d0[11] ));
 sky130_fd_sc_hd__nand4_1 _6666_ (.A(net130),
    .B(net131),
    .C(net101),
    .D(net102),
    .Y(_2859_));
 sky130_fd_sc_hd__nor3_4 _6667_ (.A(_2823_),
    .B(_2824_),
    .C(_2859_),
    .Y(_2860_));
 sky130_fd_sc_hd__xnor2_1 _6668_ (.A(net103),
    .B(_2860_),
    .Y(_2861_));
 sky130_fd_sc_hd__nor2_1 _6669_ (.A(_3489_[0]),
    .B(_3493_[0]),
    .Y(_2862_));
 sky130_fd_sc_hd__nand2_4 _6670_ (.A(_2829_),
    .B(_2862_),
    .Y(_2863_));
 sky130_fd_sc_hd__a21oi_4 _6671_ (.A1(_2833_),
    .A2(_2838_),
    .B1(_2863_),
    .Y(_2864_));
 sky130_fd_sc_hd__o21a_4 _6672_ (.A1(_3490_[0]),
    .A2(_3489_[0]),
    .B1(_3494_[0]),
    .X(_2865_));
 sky130_fd_sc_hd__nor2_1 _6673_ (.A(_3493_[0]),
    .B(_2865_),
    .Y(_2866_));
 sky130_fd_sc_hd__nor2_1 _6674_ (.A(_2864_),
    .B(_2866_),
    .Y(_2867_));
 sky130_fd_sc_hd__xnor2_1 _6675_ (.A(_3498_[0]),
    .B(_2867_),
    .Y(_2868_));
 sky130_fd_sc_hd__mux2i_1 _6676_ (.A0(_2861_),
    .A1(_2868_),
    .S(net701),
    .Y(\dp.ISRmux.d0[12] ));
 sky130_fd_sc_hd__nor2_2 _6677_ (.A(_2846_),
    .B(_2859_),
    .Y(_2869_));
 sky130_fd_sc_hd__nand2_1 _6678_ (.A(net103),
    .B(_2869_),
    .Y(_2870_));
 sky130_fd_sc_hd__xor2_1 _6679_ (.A(net104),
    .B(_2870_),
    .X(_2871_));
 sky130_fd_sc_hd__o21ai_0 _6680_ (.A1(_3493_[0]),
    .A2(_2865_),
    .B1(_3498_[0]),
    .Y(_2872_));
 sky130_fd_sc_hd__a31oi_4 _6681_ (.A1(_2837_),
    .A2(_2852_),
    .A3(_2854_),
    .B1(_2850_),
    .Y(_2873_));
 sky130_fd_sc_hd__nor2_1 _6682_ (.A(_2873_),
    .B(_2863_),
    .Y(_2874_));
 sky130_fd_sc_hd__nor2_1 _6683_ (.A(_2872_),
    .B(_2874_),
    .Y(_2875_));
 sky130_fd_sc_hd__nor2_1 _6684_ (.A(_3497_[0]),
    .B(_2875_),
    .Y(_2876_));
 sky130_fd_sc_hd__xor2_1 _6685_ (.A(_3502_[0]),
    .B(_2876_),
    .X(_2877_));
 sky130_fd_sc_hd__mux2i_1 _6686_ (.A0(_2871_),
    .A1(_2877_),
    .S(net701),
    .Y(\dp.ISRmux.d0[13] ));
 sky130_fd_sc_hd__nand3_1 _6687_ (.A(net103),
    .B(net104),
    .C(_2860_),
    .Y(_2878_));
 sky130_fd_sc_hd__xor2_1 _6688_ (.A(net105),
    .B(_2878_),
    .X(_2879_));
 sky130_fd_sc_hd__inv_1 _6689_ (.A(_3506_[0]),
    .Y(_2880_));
 sky130_fd_sc_hd__o21bai_1 _6690_ (.A1(_2864_),
    .A2(_2872_),
    .B1_N(_3497_[0]),
    .Y(_2881_));
 sky130_fd_sc_hd__a21oi_1 _6691_ (.A1(_3502_[0]),
    .A2(_2881_),
    .B1(_3501_[0]),
    .Y(_2882_));
 sky130_fd_sc_hd__xnor2_1 _6692_ (.A(_2880_),
    .B(_2882_),
    .Y(_2883_));
 sky130_fd_sc_hd__mux2i_1 _6693_ (.A0(_2879_),
    .A1(_2883_),
    .S(net225),
    .Y(\dp.ISRmux.d0[14] ));
 sky130_fd_sc_hd__nand4_1 _6694_ (.A(net103),
    .B(net104),
    .C(net105),
    .D(_2869_),
    .Y(_2884_));
 sky130_fd_sc_hd__xor2_1 _6695_ (.A(net106),
    .B(_2884_),
    .X(_2885_));
 sky130_fd_sc_hd__o211ai_1 _6696_ (.A1(_3493_[0]),
    .A2(_2865_),
    .B1(_3498_[0]),
    .C1(_3502_[0]),
    .Y(_2886_));
 sky130_fd_sc_hd__nor2_1 _6697_ (.A(_3506_[0]),
    .B(_3505_[0]),
    .Y(_2887_));
 sky130_fd_sc_hd__a21o_1 _6698_ (.A1(_3502_[0]),
    .A2(_3497_[0]),
    .B1(_3501_[0]),
    .X(_2888_));
 sky130_fd_sc_hd__a21oi_1 _6699_ (.A1(_3506_[0]),
    .A2(_2888_),
    .B1(_3505_[0]),
    .Y(_2889_));
 sky130_fd_sc_hd__o31ai_1 _6700_ (.A1(_2874_),
    .A2(_2886_),
    .A3(_2887_),
    .B1(_2889_),
    .Y(_2890_));
 sky130_fd_sc_hd__xnor2_1 _6701_ (.A(_3510_[0]),
    .B(_2890_),
    .Y(_2891_));
 sky130_fd_sc_hd__mux2i_1 _6702_ (.A0(_2885_),
    .A1(_2891_),
    .S(net225),
    .Y(\dp.ISRmux.d0[15] ));
 sky130_fd_sc_hd__and4_4 _6703_ (.A(net103),
    .B(net104),
    .C(net105),
    .D(_2860_),
    .X(_2892_));
 sky130_fd_sc_hd__nand2_1 _6704_ (.A(net106),
    .B(_2892_),
    .Y(_2893_));
 sky130_fd_sc_hd__xor2_1 _6705_ (.A(net107),
    .B(_2893_),
    .X(_2894_));
 sky130_fd_sc_hd__inv_1 _6706_ (.A(_3514_[0]),
    .Y(_2895_));
 sky130_fd_sc_hd__o31ai_1 _6707_ (.A1(_2880_),
    .A2(_2864_),
    .A3(_2886_),
    .B1(_2889_),
    .Y(_2896_));
 sky130_fd_sc_hd__a21oi_2 _6708_ (.A1(_2896_),
    .A2(_3510_[0]),
    .B1(_3509_[0]),
    .Y(_2897_));
 sky130_fd_sc_hd__xnor2_1 _6709_ (.A(_2895_),
    .B(_2897_),
    .Y(_2898_));
 sky130_fd_sc_hd__mux2i_1 _6710_ (.A0(_2894_),
    .A1(_2898_),
    .S(net701),
    .Y(\dp.ISRmux.d0[16] ));
 sky130_fd_sc_hd__nand2_1 _6711_ (.A(net106),
    .B(net107),
    .Y(_2899_));
 sky130_fd_sc_hd__nor2_1 _6712_ (.A(_2884_),
    .B(_2899_),
    .Y(_2900_));
 sky130_fd_sc_hd__xnor2_1 _6713_ (.A(net108),
    .B(_2900_),
    .Y(_2901_));
 sky130_fd_sc_hd__nand2_1 _6714_ (.A(_3510_[0]),
    .B(_3514_[0]),
    .Y(_2902_));
 sky130_fd_sc_hd__nor3_1 _6715_ (.A(_2886_),
    .B(_2887_),
    .C(_2902_),
    .Y(_2903_));
 sky130_fd_sc_hd__o21ai_2 _6716_ (.A1(_2873_),
    .A2(_2863_),
    .B1(_2903_),
    .Y(_2904_));
 sky130_fd_sc_hd__nor2_1 _6717_ (.A(_2889_),
    .B(_2902_),
    .Y(_2905_));
 sky130_fd_sc_hd__a21oi_2 _6718_ (.A1(_3514_[0]),
    .A2(_3509_[0]),
    .B1(_2905_),
    .Y(_2906_));
 sky130_fd_sc_hd__nand3b_1 _6719_ (.A_N(_3513_[0]),
    .B(_2904_),
    .C(_2906_),
    .Y(_2907_));
 sky130_fd_sc_hd__xnor2_1 _6720_ (.A(_3518_[0]),
    .B(_2907_),
    .Y(_2908_));
 sky130_fd_sc_hd__mux2i_1 _6721_ (.A0(_2901_),
    .A1(_2908_),
    .S(net224),
    .Y(\dp.ISRmux.d0[17] ));
 sky130_fd_sc_hd__nand4_1 _6722_ (.A(net106),
    .B(net107),
    .C(net108),
    .D(_2892_),
    .Y(_2909_));
 sky130_fd_sc_hd__xor2_1 _6723_ (.A(net109),
    .B(_2909_),
    .X(_2910_));
 sky130_fd_sc_hd__nand3_1 _6724_ (.A(_3514_[0]),
    .B(_3518_[0]),
    .C(_3522_[0]),
    .Y(_2911_));
 sky130_fd_sc_hd__nand2_1 _6725_ (.A(_3522_[0]),
    .B(_3517_[0]),
    .Y(_2912_));
 sky130_fd_sc_hd__nand3_1 _6726_ (.A(_3518_[0]),
    .B(_3522_[0]),
    .C(_3513_[0]),
    .Y(_2913_));
 sky130_fd_sc_hd__o211a_4 _6727_ (.A1(_2897_),
    .A2(_2911_),
    .B1(_2912_),
    .C1(_2913_),
    .X(_2914_));
 sky130_fd_sc_hd__o21bai_1 _6728_ (.A1(_2895_),
    .A2(_2897_),
    .B1_N(_3513_[0]),
    .Y(_2915_));
 sky130_fd_sc_hd__a211o_1 _6729_ (.A1(_3518_[0]),
    .A2(_2915_),
    .B1(_3517_[0]),
    .C1(_3522_[0]),
    .X(_2916_));
 sky130_fd_sc_hd__nand2_1 _6730_ (.A(_2914_),
    .B(_2916_),
    .Y(_2917_));
 sky130_fd_sc_hd__mux2i_1 _6731_ (.A0(_2910_),
    .A1(_2917_),
    .S(net701),
    .Y(\dp.ISRmux.d0[18] ));
 sky130_fd_sc_hd__nand4_1 _6732_ (.A(net106),
    .B(net107),
    .C(net108),
    .D(net109),
    .Y(_2918_));
 sky130_fd_sc_hd__nor2_1 _6733_ (.A(_2884_),
    .B(_2918_),
    .Y(_2919_));
 sky130_fd_sc_hd__xnor2_1 _6734_ (.A(net110),
    .B(_2919_),
    .Y(_2920_));
 sky130_fd_sc_hd__nor3_1 _6735_ (.A(_3513_[0]),
    .B(_3517_[0]),
    .C(_3521_[0]),
    .Y(_2921_));
 sky130_fd_sc_hd__or2_0 _6736_ (.A(_3518_[0]),
    .B(_3517_[0]),
    .X(_2922_));
 sky130_fd_sc_hd__a21oi_1 _6737_ (.A1(_3522_[0]),
    .A2(_2922_),
    .B1(_3521_[0]),
    .Y(_2923_));
 sky130_fd_sc_hd__a31oi_1 _6738_ (.A1(_2904_),
    .A2(_2906_),
    .A3(_2921_),
    .B1(_2923_),
    .Y(_2924_));
 sky130_fd_sc_hd__xnor2_1 _6739_ (.A(_3526_[0]),
    .B(_2924_),
    .Y(_2925_));
 sky130_fd_sc_hd__mux2i_1 _6740_ (.A0(_2920_),
    .A1(_2925_),
    .S(net225),
    .Y(\dp.ISRmux.d0[19] ));
 sky130_fd_sc_hd__inv_1 _6741_ (.A(net110),
    .Y(_2926_));
 sky130_fd_sc_hd__nand4_1 _6742_ (.A(net103),
    .B(net104),
    .C(net105),
    .D(_2860_),
    .Y(_2927_));
 sky130_fd_sc_hd__nor3_1 _6743_ (.A(_2926_),
    .B(_2927_),
    .C(_2918_),
    .Y(_2928_));
 sky130_fd_sc_hd__xnor2_1 _6744_ (.A(net112),
    .B(_2928_),
    .Y(_2929_));
 sky130_fd_sc_hd__nand2b_1 _6745_ (.A_N(_3521_[0]),
    .B(_2914_),
    .Y(_2930_));
 sky130_fd_sc_hd__a21oi_1 _6746_ (.A1(_3526_[0]),
    .A2(_2930_),
    .B1(_3525_[0]),
    .Y(_2931_));
 sky130_fd_sc_hd__xor2_1 _6747_ (.A(_3530_[0]),
    .B(_2931_),
    .X(_2932_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_15 ();
 sky130_fd_sc_hd__mux2i_1 _6749_ (.A0(_2929_),
    .A1(_2932_),
    .S(net225),
    .Y(\dp.ISRmux.d0[20] ));
 sky130_fd_sc_hd__nor2_2 _6750_ (.A(_2926_),
    .B(_2918_),
    .Y(_2934_));
 sky130_fd_sc_hd__nand2_1 _6751_ (.A(net112),
    .B(_2934_),
    .Y(_2935_));
 sky130_fd_sc_hd__nor2_1 _6752_ (.A(_2884_),
    .B(_2935_),
    .Y(_2936_));
 sky130_fd_sc_hd__xnor2_1 _6753_ (.A(net113),
    .B(_2936_),
    .Y(_2937_));
 sky130_fd_sc_hd__nand2_1 _6754_ (.A(_3526_[0]),
    .B(_3530_[0]),
    .Y(_2938_));
 sky130_fd_sc_hd__a311oi_2 _6755_ (.A1(_2904_),
    .A2(_2906_),
    .A3(_2921_),
    .B1(_2923_),
    .C1(_2938_),
    .Y(_2939_));
 sky130_fd_sc_hd__a21o_1 _6756_ (.A1(_3530_[0]),
    .A2(_3525_[0]),
    .B1(_3529_[0]),
    .X(_2940_));
 sky130_fd_sc_hd__nor2_1 _6757_ (.A(_2939_),
    .B(_2940_),
    .Y(_2941_));
 sky130_fd_sc_hd__xor2_1 _6758_ (.A(_3534_[0]),
    .B(_2941_),
    .X(_2942_));
 sky130_fd_sc_hd__mux2i_1 _6759_ (.A0(_2937_),
    .A1(_2942_),
    .S(net225),
    .Y(\dp.ISRmux.d0[21] ));
 sky130_fd_sc_hd__nand4_1 _6760_ (.A(net112),
    .B(net113),
    .C(_2892_),
    .D(_2934_),
    .Y(_2943_));
 sky130_fd_sc_hd__xor2_1 _6761_ (.A(net114),
    .B(_2943_),
    .X(_2944_));
 sky130_fd_sc_hd__nor3_1 _6762_ (.A(_3521_[0]),
    .B(_3525_[0]),
    .C(_3529_[0]),
    .Y(_2945_));
 sky130_fd_sc_hd__or2_0 _6763_ (.A(_3526_[0]),
    .B(_3525_[0]),
    .X(_2946_));
 sky130_fd_sc_hd__a21oi_1 _6764_ (.A1(_3530_[0]),
    .A2(_2946_),
    .B1(_3529_[0]),
    .Y(_2947_));
 sky130_fd_sc_hd__a21oi_1 _6765_ (.A1(_2914_),
    .A2(_2945_),
    .B1(_2947_),
    .Y(_2948_));
 sky130_fd_sc_hd__a21oi_1 _6766_ (.A1(_3534_[0]),
    .A2(_2948_),
    .B1(_3533_[0]),
    .Y(_2949_));
 sky130_fd_sc_hd__xor2_1 _6767_ (.A(_3538_[0]),
    .B(_2949_),
    .X(_2950_));
 sky130_fd_sc_hd__mux2i_2 _6768_ (.A0(_2944_),
    .A1(_2950_),
    .S(net701),
    .Y(\dp.ISRmux.d0[22] ));
 sky130_fd_sc_hd__nand4_1 _6769_ (.A(net112),
    .B(net113),
    .C(net114),
    .D(_2934_),
    .Y(_2951_));
 sky130_fd_sc_hd__nor2_4 _6770_ (.A(_2884_),
    .B(_2951_),
    .Y(_2952_));
 sky130_fd_sc_hd__xnor2_1 _6771_ (.A(net115),
    .B(_2952_),
    .Y(_2953_));
 sky130_fd_sc_hd__o21ai_2 _6772_ (.A1(_2939_),
    .A2(_2940_),
    .B1(_3534_[0]),
    .Y(_2954_));
 sky130_fd_sc_hd__nand2b_1 _6773_ (.A_N(_3533_[0]),
    .B(_2954_),
    .Y(_2955_));
 sky130_fd_sc_hd__a21oi_1 _6774_ (.A1(_3538_[0]),
    .A2(_2955_),
    .B1(_3537_[0]),
    .Y(_2956_));
 sky130_fd_sc_hd__xor2_1 _6775_ (.A(_3542_[0]),
    .B(_2956_),
    .X(_2957_));
 sky130_fd_sc_hd__mux2i_1 _6776_ (.A0(_2953_),
    .A1(_2957_),
    .S(net225),
    .Y(\dp.ISRmux.d0[23] ));
 sky130_fd_sc_hd__nor2_4 _6777_ (.A(_2927_),
    .B(_2951_),
    .Y(_2958_));
 sky130_fd_sc_hd__nand2_1 _6778_ (.A(net115),
    .B(_2958_),
    .Y(_2959_));
 sky130_fd_sc_hd__xor2_1 _6779_ (.A(net116),
    .B(_2959_),
    .X(_2960_));
 sky130_fd_sc_hd__nand3_1 _6780_ (.A(_3534_[0]),
    .B(_3538_[0]),
    .C(_3542_[0]),
    .Y(_2961_));
 sky130_fd_sc_hd__a211o_4 _6781_ (.A1(_2914_),
    .A2(_2945_),
    .B1(_2947_),
    .C1(_2961_),
    .X(_2962_));
 sky130_fd_sc_hd__and3_1 _6782_ (.A(_3538_[0]),
    .B(_3542_[0]),
    .C(_3533_[0]),
    .X(_2963_));
 sky130_fd_sc_hd__a21oi_1 _6783_ (.A1(_3542_[0]),
    .A2(_3537_[0]),
    .B1(_2963_),
    .Y(_2964_));
 sky130_fd_sc_hd__nand3b_1 _6784_ (.A_N(_3541_[0]),
    .B(_2962_),
    .C(_2964_),
    .Y(_2965_));
 sky130_fd_sc_hd__xnor2_1 _6785_ (.A(_3546_[0]),
    .B(_2965_),
    .Y(_2966_));
 sky130_fd_sc_hd__mux2i_1 _6786_ (.A0(_2960_),
    .A1(_2966_),
    .S(net237),
    .Y(\dp.ISRmux.d0[24] ));
 sky130_fd_sc_hd__nand3_1 _6787_ (.A(net115),
    .B(net116),
    .C(_2952_),
    .Y(_2967_));
 sky130_fd_sc_hd__xor2_1 _6788_ (.A(net117),
    .B(_2967_),
    .X(_2968_));
 sky130_fd_sc_hd__nor3_1 _6789_ (.A(_3533_[0]),
    .B(_3537_[0]),
    .C(_3541_[0]),
    .Y(_2969_));
 sky130_fd_sc_hd__or2_0 _6790_ (.A(_3538_[0]),
    .B(_3537_[0]),
    .X(_2970_));
 sky130_fd_sc_hd__a21oi_1 _6791_ (.A1(_3542_[0]),
    .A2(_2970_),
    .B1(_3541_[0]),
    .Y(_2971_));
 sky130_fd_sc_hd__a21oi_1 _6792_ (.A1(_2954_),
    .A2(_2969_),
    .B1(_2971_),
    .Y(_2972_));
 sky130_fd_sc_hd__a21oi_1 _6793_ (.A1(_3546_[0]),
    .A2(_2972_),
    .B1(_3545_[0]),
    .Y(_2973_));
 sky130_fd_sc_hd__xor2_1 _6794_ (.A(_3550_[0]),
    .B(_2973_),
    .X(_2974_));
 sky130_fd_sc_hd__mux2i_1 _6795_ (.A0(_2968_),
    .A1(_2974_),
    .S(net237),
    .Y(\dp.ISRmux.d0[25] ));
 sky130_fd_sc_hd__and3_4 _6796_ (.A(net115),
    .B(net116),
    .C(net117),
    .X(_2975_));
 sky130_fd_sc_hd__nand2_1 _6797_ (.A(_2958_),
    .B(_2975_),
    .Y(_2976_));
 sky130_fd_sc_hd__xor2_1 _6798_ (.A(net118),
    .B(_2976_),
    .X(_2977_));
 sky130_fd_sc_hd__nor3_1 _6799_ (.A(_3541_[0]),
    .B(_3545_[0]),
    .C(_3549_[0]),
    .Y(_2978_));
 sky130_fd_sc_hd__or2_0 _6800_ (.A(_3546_[0]),
    .B(_3545_[0]),
    .X(_2979_));
 sky130_fd_sc_hd__a21oi_1 _6801_ (.A1(_3550_[0]),
    .A2(_2979_),
    .B1(_3549_[0]),
    .Y(_2980_));
 sky130_fd_sc_hd__a31oi_2 _6802_ (.A1(_2962_),
    .A2(_2964_),
    .A3(_2978_),
    .B1(_2980_),
    .Y(_2981_));
 sky130_fd_sc_hd__xnor2_1 _6803_ (.A(_3554_[0]),
    .B(_2981_),
    .Y(_2982_));
 sky130_fd_sc_hd__mux2i_1 _6804_ (.A0(_2977_),
    .A1(_2982_),
    .S(net237),
    .Y(\dp.ISRmux.d0[26] ));
 sky130_fd_sc_hd__and3_4 _6805_ (.A(net118),
    .B(_2952_),
    .C(_2975_),
    .X(_2983_));
 sky130_fd_sc_hd__xnor2_1 _6806_ (.A(net119),
    .B(_2983_),
    .Y(_2984_));
 sky130_fd_sc_hd__nand3_1 _6807_ (.A(_3546_[0]),
    .B(_3550_[0]),
    .C(_3554_[0]),
    .Y(_2985_));
 sky130_fd_sc_hd__a211oi_2 _6808_ (.A1(_2954_),
    .A2(_2969_),
    .B1(_2971_),
    .C1(_2985_),
    .Y(_2986_));
 sky130_fd_sc_hd__nand2_1 _6809_ (.A(_3554_[0]),
    .B(_3549_[0]),
    .Y(_2987_));
 sky130_fd_sc_hd__nand3_1 _6810_ (.A(_3550_[0]),
    .B(_3554_[0]),
    .C(_3545_[0]),
    .Y(_2988_));
 sky130_fd_sc_hd__nand2_2 _6811_ (.A(_2987_),
    .B(_2988_),
    .Y(_2989_));
 sky130_fd_sc_hd__nor3_1 _6812_ (.A(_3553_[0]),
    .B(_2986_),
    .C(_2989_),
    .Y(_2990_));
 sky130_fd_sc_hd__xor2_1 _6813_ (.A(_3558_[0]),
    .B(_2990_),
    .X(_2991_));
 sky130_fd_sc_hd__mux2i_1 _6814_ (.A0(_2984_),
    .A1(_2991_),
    .S(net237),
    .Y(\dp.ISRmux.d0[27] ));
 sky130_fd_sc_hd__nand4_1 _6815_ (.A(net118),
    .B(net119),
    .C(_2958_),
    .D(_2975_),
    .Y(_2992_));
 sky130_fd_sc_hd__xor2_1 _6816_ (.A(net120),
    .B(_2992_),
    .X(_2993_));
 sky130_fd_sc_hd__a21o_1 _6817_ (.A1(_3554_[0]),
    .A2(_2981_),
    .B1(_3553_[0]),
    .X(_2994_));
 sky130_fd_sc_hd__a21oi_1 _6818_ (.A1(_3558_[0]),
    .A2(_2994_),
    .B1(_3557_[0]),
    .Y(_2995_));
 sky130_fd_sc_hd__xor2_1 _6819_ (.A(_3562_[0]),
    .B(_2995_),
    .X(_2996_));
 sky130_fd_sc_hd__mux2i_1 _6820_ (.A0(_2993_),
    .A1(_2996_),
    .S(net237),
    .Y(\dp.ISRmux.d0[28] ));
 sky130_fd_sc_hd__nand3_1 _6821_ (.A(net119),
    .B(net120),
    .C(_2983_),
    .Y(_2997_));
 sky130_fd_sc_hd__xor2_1 _6822_ (.A(net121),
    .B(_2997_),
    .X(_2998_));
 sky130_fd_sc_hd__or3_4 _6823_ (.A(_3553_[0]),
    .B(_3557_[0]),
    .C(_3561_[0]),
    .X(_2999_));
 sky130_fd_sc_hd__nor3_1 _6824_ (.A(_3558_[0]),
    .B(_3557_[0]),
    .C(_3561_[0]),
    .Y(_3000_));
 sky130_fd_sc_hd__nor2_1 _6825_ (.A(_3562_[0]),
    .B(_3561_[0]),
    .Y(_3001_));
 sky130_fd_sc_hd__nor2_2 _6826_ (.A(_3000_),
    .B(_3001_),
    .Y(_3002_));
 sky130_fd_sc_hd__o31ai_4 _6827_ (.A1(_2986_),
    .A2(_2989_),
    .A3(_2999_),
    .B1(_3002_),
    .Y(_3003_));
 sky130_fd_sc_hd__xor2_1 _6828_ (.A(_3566_[0]),
    .B(_3003_),
    .X(_3004_));
 sky130_fd_sc_hd__mux2i_1 _6829_ (.A0(_2998_),
    .A1(_3004_),
    .S(net237),
    .Y(\dp.ISRmux.d0[29] ));
 sky130_fd_sc_hd__xnor2_1 _6830_ (.A(_3192_[0]),
    .B(_3456_[0]),
    .Y(_3005_));
 sky130_fd_sc_hd__mux2i_1 _6831_ (.A0(net122),
    .A1(_3005_),
    .S(net241),
    .Y(\dp.ISRmux.d0[2] ));
 sky130_fd_sc_hd__and3_4 _6832_ (.A(net119),
    .B(net120),
    .C(net121),
    .X(_3006_));
 sky130_fd_sc_hd__nand4_1 _6833_ (.A(net118),
    .B(_2958_),
    .C(_2975_),
    .D(_3006_),
    .Y(_3007_));
 sky130_fd_sc_hd__xor2_2 _6834_ (.A(net123),
    .B(_3007_),
    .X(_3008_));
 sky130_fd_sc_hd__nand4_1 _6835_ (.A(_3554_[0]),
    .B(_3558_[0]),
    .C(_3562_[0]),
    .D(_2981_),
    .Y(_3009_));
 sky130_fd_sc_hd__nand2_1 _6836_ (.A(_3562_[0]),
    .B(_3557_[0]),
    .Y(_3010_));
 sky130_fd_sc_hd__nand3_1 _6837_ (.A(_3558_[0]),
    .B(_3562_[0]),
    .C(_3553_[0]),
    .Y(_3011_));
 sky130_fd_sc_hd__nand4b_1 _6838_ (.A_N(_3561_[0]),
    .B(_3009_),
    .C(_3010_),
    .D(_3011_),
    .Y(_3012_));
 sky130_fd_sc_hd__a21oi_2 _6839_ (.A1(_3566_[0]),
    .A2(_3012_),
    .B1(_3565_[0]),
    .Y(_3013_));
 sky130_fd_sc_hd__xor2_2 _6840_ (.A(_3013_),
    .B(_3570_[0]),
    .X(_3014_));
 sky130_fd_sc_hd__mux2i_1 _6841_ (.A0(_3008_),
    .A1(_3014_),
    .S(net237),
    .Y(\dp.ISRmux.d0[30] ));
 sky130_fd_sc_hd__nand3_1 _6842_ (.A(net123),
    .B(_2983_),
    .C(_3006_),
    .Y(_3015_));
 sky130_fd_sc_hd__xor2_1 _6843_ (.A(net124),
    .B(_3015_),
    .X(_3016_));
 sky130_fd_sc_hd__nand2_1 _6844_ (.A(net124),
    .B(net776),
    .Y(_3017_));
 sky130_fd_sc_hd__o21ai_0 _6845_ (.A1(_0314_),
    .A2(net776),
    .B1(_3017_),
    .Y(_3018_));
 sky130_fd_sc_hd__xor2_1 _6846_ (.A(net25),
    .B(_3018_),
    .X(_3019_));
 sky130_fd_sc_hd__and3_1 _6847_ (.A(_3566_[0]),
    .B(_3570_[0]),
    .C(_3019_),
    .X(_3020_));
 sky130_fd_sc_hd__nor3_1 _6848_ (.A(_3565_[0]),
    .B(_3569_[0]),
    .C(_3019_),
    .Y(_3021_));
 sky130_fd_sc_hd__mux2i_1 _6849_ (.A0(_3020_),
    .A1(_3021_),
    .S(_3003_),
    .Y(_3022_));
 sky130_fd_sc_hd__nand2_1 _6850_ (.A(_3569_[0]),
    .B(_3019_),
    .Y(_3023_));
 sky130_fd_sc_hd__nand3_1 _6851_ (.A(_3570_[0]),
    .B(_3565_[0]),
    .C(_3019_),
    .Y(_3024_));
 sky130_fd_sc_hd__nor4_1 _6852_ (.A(_3566_[0]),
    .B(_3565_[0]),
    .C(_3569_[0]),
    .D(_3019_),
    .Y(_3025_));
 sky130_fd_sc_hd__nor3_1 _6853_ (.A(_3570_[0]),
    .B(_3569_[0]),
    .C(_3019_),
    .Y(_3026_));
 sky130_fd_sc_hd__nor2_1 _6854_ (.A(_3025_),
    .B(_3026_),
    .Y(_3027_));
 sky130_fd_sc_hd__nand4_1 _6855_ (.A(_3022_),
    .B(_3023_),
    .C(_3024_),
    .D(_3027_),
    .Y(_3028_));
 sky130_fd_sc_hd__mux2i_1 _6856_ (.A0(_3016_),
    .A1(_3028_),
    .S(net237),
    .Y(\dp.ISRmux.d0[31] ));
 sky130_fd_sc_hd__nor2b_1 _6857_ (.A(_2851_),
    .B_N(_3456_[0]),
    .Y(_3029_));
 sky130_fd_sc_hd__nor2_1 _6858_ (.A(_3455_[0]),
    .B(_3029_),
    .Y(_3030_));
 sky130_fd_sc_hd__xnor2_1 _6859_ (.A(_3460_[0]),
    .B(_3030_),
    .Y(_3031_));
 sky130_fd_sc_hd__mux2_1 _6860_ (.A0(_3462_[0]),
    .A1(_3031_),
    .S(net241),
    .X(\dp.ISRmux.d0[3] ));
 sky130_fd_sc_hd__xnor2_1 _6861_ (.A(net126),
    .B(_3461_[0]),
    .Y(_3032_));
 sky130_fd_sc_hd__xnor2_1 _6862_ (.A(_2834_),
    .B(_2836_),
    .Y(_3033_));
 sky130_fd_sc_hd__mux2i_1 _6863_ (.A0(_3032_),
    .A1(_3033_),
    .S(net243),
    .Y(\dp.ISRmux.d0[4] ));
 sky130_fd_sc_hd__nand3_1 _6864_ (.A(net122),
    .B(net125),
    .C(net126),
    .Y(_3034_));
 sky130_fd_sc_hd__xor2_1 _6865_ (.A(net127),
    .B(_3034_),
    .X(_3035_));
 sky130_fd_sc_hd__nand2_1 _6866_ (.A(_2852_),
    .B(_2854_),
    .Y(_3036_));
 sky130_fd_sc_hd__nor2_1 _6867_ (.A(_3465_[0]),
    .B(_3036_),
    .Y(_3037_));
 sky130_fd_sc_hd__xor2_1 _6868_ (.A(_3470_[0]),
    .B(_3037_),
    .X(_3038_));
 sky130_fd_sc_hd__mux2i_1 _6869_ (.A0(_3035_),
    .A1(_3038_),
    .S(net241),
    .Y(\dp.ISRmux.d0[5] ));
 sky130_fd_sc_hd__xor2_1 _6870_ (.A(net128),
    .B(_2823_),
    .X(_3039_));
 sky130_fd_sc_hd__o21bai_1 _6871_ (.A1(_2834_),
    .A2(_2836_),
    .B1_N(_3465_[0]),
    .Y(_3040_));
 sky130_fd_sc_hd__a21oi_1 _6872_ (.A1(_3470_[0]),
    .A2(_3040_),
    .B1(_3469_[0]),
    .Y(_3041_));
 sky130_fd_sc_hd__xor2_1 _6873_ (.A(_3474_[0]),
    .B(_3041_),
    .X(_3042_));
 sky130_fd_sc_hd__mux2i_1 _6874_ (.A0(_3039_),
    .A1(_3042_),
    .S(net242),
    .Y(\dp.ISRmux.d0[6] ));
 sky130_fd_sc_hd__xnor2_1 _6875_ (.A(net129),
    .B(_2845_),
    .Y(_3043_));
 sky130_fd_sc_hd__nor2_1 _6876_ (.A(_3473_[0]),
    .B(_2830_),
    .Y(_3044_));
 sky130_fd_sc_hd__nor2_1 _6877_ (.A(_3044_),
    .B(_2855_),
    .Y(_3045_));
 sky130_fd_sc_hd__xnor2_1 _6878_ (.A(_3478_[0]),
    .B(_3045_),
    .Y(_3046_));
 sky130_fd_sc_hd__mux2i_1 _6879_ (.A0(_3043_),
    .A1(_3046_),
    .S(net237),
    .Y(\dp.ISRmux.d0[7] ));
 sky130_fd_sc_hd__xnor2_1 _6880_ (.A(net130),
    .B(_2825_),
    .Y(_3047_));
 sky130_fd_sc_hd__inv_1 _6881_ (.A(_2831_),
    .Y(_3048_));
 sky130_fd_sc_hd__a21oi_1 _6882_ (.A1(_3048_),
    .A2(_2838_),
    .B1(_3477_[0]),
    .Y(_3049_));
 sky130_fd_sc_hd__xor2_1 _6883_ (.A(_3482_[0]),
    .B(_3049_),
    .X(_3050_));
 sky130_fd_sc_hd__mux2i_1 _6884_ (.A0(_3047_),
    .A1(_3050_),
    .S(net237),
    .Y(\dp.ISRmux.d0[8] ));
 sky130_fd_sc_hd__nand3_1 _6885_ (.A(net129),
    .B(net130),
    .C(_2845_),
    .Y(_3051_));
 sky130_fd_sc_hd__xor2_1 _6886_ (.A(net131),
    .B(_3051_),
    .X(_3052_));
 sky130_fd_sc_hd__o21bai_1 _6887_ (.A1(_2831_),
    .A2(_2855_),
    .B1_N(_3477_[0]),
    .Y(_3053_));
 sky130_fd_sc_hd__a21oi_1 _6888_ (.A1(_3482_[0]),
    .A2(_3053_),
    .B1(_3481_[0]),
    .Y(_3054_));
 sky130_fd_sc_hd__xor2_1 _6889_ (.A(_3486_[0]),
    .B(_3054_),
    .X(_3055_));
 sky130_fd_sc_hd__mux2i_1 _6890_ (.A0(_3052_),
    .A1(_3055_),
    .S(net237),
    .Y(\dp.ISRmux.d0[9] ));
 sky130_fd_sc_hd__nor2_4 _6891_ (.A(net28),
    .B(_0347_),
    .Y(_3056_));
 sky130_fd_sc_hd__nor2_4 _6892_ (.A(_0896_),
    .B(_3056_),
    .Y(_3057_));
 sky130_fd_sc_hd__nand2_8 _6893_ (.A(_1875_),
    .B(_3057_),
    .Y(_3058_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__o22a_1 _6896_ (.A1(net100),
    .A2(_2686_),
    .B1(_2646_),
    .B2(_3450_[0]),
    .X(_3061_));
 sky130_fd_sc_hd__o221a_4 _6897_ (.A1(net33),
    .A2(_1875_),
    .B1(_3058_),
    .B2(net244),
    .C1(_3061_),
    .X(\dp.result2[0] ));
 sky130_fd_sc_hd__nor4_1 _6898_ (.A(net815),
    .B(net5),
    .C(net99),
    .D(_1700_),
    .Y(_3062_));
 sky130_fd_sc_hd__nand3b_1 _6899_ (.A_N(net6),
    .B(net62),
    .C(_3062_),
    .Y(_3063_));
 sky130_fd_sc_hd__and2_4 _6900_ (.A(net98),
    .B(_3063_),
    .X(_3064_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__nor2_2 _6902_ (.A(net815),
    .B(net5),
    .Y(_3066_));
 sky130_fd_sc_hd__nand3_4 _6903_ (.A(_0044_),
    .B(_3066_),
    .C(_1713_),
    .Y(_3067_));
 sky130_fd_sc_hd__nand2_1 _6904_ (.A(net34),
    .B(_3067_),
    .Y(_3068_));
 sky130_fd_sc_hd__nand2_4 _6905_ (.A(_2686_),
    .B(_2646_),
    .Y(_3069_));
 sky130_fd_sc_hd__a21oi_1 _6906_ (.A1(_3064_),
    .A2(_3068_),
    .B1(_3069_),
    .Y(_3070_));
 sky130_fd_sc_hd__o21ai_4 _6907_ (.A1(net98),
    .A2(net373),
    .B1(_3070_),
    .Y(_3071_));
 sky130_fd_sc_hd__o221ai_4 _6908_ (.A1(_2686_),
    .A2(_2827_),
    .B1(_2841_),
    .B2(_2646_),
    .C1(_3071_),
    .Y(\dp.result2[10] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__nand2_1 _6911_ (.A(net35),
    .B(_3067_),
    .Y(_3074_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__a222oi_1 _6913_ (.A1(_0896_),
    .A2(_2849_),
    .B1(_3064_),
    .B2(_3074_),
    .C1(_2858_),
    .C2(_3056_),
    .Y(_3076_));
 sky130_fd_sc_hd__o21a_4 _6914_ (.A1(net375),
    .A2(_3058_),
    .B1(_3076_),
    .X(\dp.result2[11] ));
 sky130_fd_sc_hd__nand2_1 _6915_ (.A(net36),
    .B(_3067_),
    .Y(_3077_));
 sky130_fd_sc_hd__a222oi_1 _6916_ (.A1(_0896_),
    .A2(_2861_),
    .B1(_3064_),
    .B2(_3077_),
    .C1(_2868_),
    .C2(_3056_),
    .Y(_3078_));
 sky130_fd_sc_hd__o21a_4 _6917_ (.A1(net367),
    .A2(_3058_),
    .B1(_3078_),
    .X(\dp.result2[12] ));
 sky130_fd_sc_hd__nor2_1 _6918_ (.A(net98),
    .B(net361),
    .Y(_3079_));
 sky130_fd_sc_hd__nand2_2 _6919_ (.A(net98),
    .B(_3063_),
    .Y(_3080_));
 sky130_fd_sc_hd__and2_0 _6920_ (.A(net37),
    .B(_3067_),
    .X(_3081_));
 sky130_fd_sc_hd__o21ai_2 _6921_ (.A1(_3080_),
    .A2(_3081_),
    .B1(_3057_),
    .Y(_3082_));
 sky130_fd_sc_hd__o22ai_1 _6922_ (.A1(_2686_),
    .A2(_2871_),
    .B1(_2877_),
    .B2(_2646_),
    .Y(_3083_));
 sky130_fd_sc_hd__o21bai_4 _6923_ (.A1(_3079_),
    .A2(_3082_),
    .B1_N(_3083_),
    .Y(\dp.result2[13] ));
 sky130_fd_sc_hd__a21oi_1 _6924_ (.A1(net38),
    .A2(_3067_),
    .B1(_3080_),
    .Y(_3084_));
 sky130_fd_sc_hd__a221oi_1 _6925_ (.A1(_0896_),
    .A2(_2879_),
    .B1(_2883_),
    .B2(_3056_),
    .C1(_3084_),
    .Y(_3085_));
 sky130_fd_sc_hd__o21a_4 _6926_ (.A1(net332),
    .A2(_3058_),
    .B1(_3085_),
    .X(\dp.result2[14] ));
 sky130_fd_sc_hd__nand2_1 _6927_ (.A(net39),
    .B(_3067_),
    .Y(_3086_));
 sky130_fd_sc_hd__a21oi_1 _6928_ (.A1(_3064_),
    .A2(_3086_),
    .B1(_3069_),
    .Y(_3087_));
 sky130_fd_sc_hd__o21ai_2 _6929_ (.A1(net98),
    .A2(net368),
    .B1(_3087_),
    .Y(_3088_));
 sky130_fd_sc_hd__o221ai_4 _6930_ (.A1(_2686_),
    .A2(_2885_),
    .B1(_2891_),
    .B2(_2646_),
    .C1(_3088_),
    .Y(\dp.result2[15] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__or3_4 _6932_ (.A(net28),
    .B(_1700_),
    .C(_1715_),
    .X(_3090_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__nor3b_4 _6935_ (.A(_3090_),
    .B(net814),
    .C_N(net39),
    .Y(_3093_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__a21oi_1 _6937_ (.A1(net40),
    .A2(_3090_),
    .B1(_3093_),
    .Y(_3095_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__o21ai_0 _6939_ (.A1(net772),
    .A2(_3095_),
    .B1(_3064_),
    .Y(_3097_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__a22oi_1 _6942_ (.A1(_0896_),
    .A2(_2894_),
    .B1(_2898_),
    .B2(_3056_),
    .Y(_3100_));
 sky130_fd_sc_hd__o211a_4 _6943_ (.A1(net73),
    .A2(_3058_),
    .B1(_3097_),
    .C1(_3100_),
    .X(\dp.result2[16] ));
 sky130_fd_sc_hd__o22ai_1 _6944_ (.A1(_2686_),
    .A2(_2901_),
    .B1(_2908_),
    .B2(_2646_),
    .Y(_3101_));
 sky130_fd_sc_hd__a21oi_1 _6945_ (.A1(net41),
    .A2(_3090_),
    .B1(_3093_),
    .Y(_3102_));
 sky130_fd_sc_hd__o21ai_0 _6946_ (.A1(net772),
    .A2(_3102_),
    .B1(_3064_),
    .Y(_3103_));
 sky130_fd_sc_hd__a21o_1 _6947_ (.A1(_3057_),
    .A2(_3103_),
    .B1(_3101_),
    .X(_3104_));
 sky130_fd_sc_hd__o31a_1 _6948_ (.A1(net98),
    .A2(net358),
    .A3(_3101_),
    .B1(_3104_),
    .X(\dp.result2[17] ));
 sky130_fd_sc_hd__nand2_1 _6949_ (.A(_3056_),
    .B(_2917_),
    .Y(_3105_));
 sky130_fd_sc_hd__a21oi_1 _6950_ (.A1(net42),
    .A2(_3090_),
    .B1(_3093_),
    .Y(_3106_));
 sky130_fd_sc_hd__o21ai_0 _6951_ (.A1(net772),
    .A2(_3106_),
    .B1(_3064_),
    .Y(_3107_));
 sky130_fd_sc_hd__nand2_1 _6952_ (.A(_0896_),
    .B(_2910_),
    .Y(_3108_));
 sky130_fd_sc_hd__o2111a_4 _6953_ (.A1(net75),
    .A2(_3058_),
    .B1(_3105_),
    .C1(_3107_),
    .D1(_3108_),
    .X(\dp.result2[18] ));
 sky130_fd_sc_hd__a21oi_1 _6954_ (.A1(net43),
    .A2(_3090_),
    .B1(_3093_),
    .Y(_3109_));
 sky130_fd_sc_hd__o21ai_0 _6955_ (.A1(net772),
    .A2(_3109_),
    .B1(_3064_),
    .Y(_3110_));
 sky130_fd_sc_hd__nand2_1 _6956_ (.A(_3057_),
    .B(_3110_),
    .Y(_3111_));
 sky130_fd_sc_hd__a31oi_2 _6957_ (.A1(_2367_),
    .A2(_2378_),
    .A3(net364),
    .B1(net98),
    .Y(_3112_));
 sky130_fd_sc_hd__o22ai_1 _6958_ (.A1(_2686_),
    .A2(_2920_),
    .B1(_2925_),
    .B2(_2646_),
    .Y(_3113_));
 sky130_fd_sc_hd__o21bai_2 _6959_ (.A1(_3111_),
    .A2(_3112_),
    .B1_N(_3113_),
    .Y(\dp.result2[19] ));
 sky130_fd_sc_hd__o22a_1 _6960_ (.A1(net111),
    .A2(_2686_),
    .B1(_2646_),
    .B2(_3193_[0]),
    .X(_3114_));
 sky130_fd_sc_hd__o221a_4 _6961_ (.A1(net44),
    .A2(_1875_),
    .B1(net380),
    .B2(_3058_),
    .C1(_3114_),
    .X(\dp.result2[1] ));
 sky130_fd_sc_hd__a21oi_1 _6962_ (.A1(net45),
    .A2(_3090_),
    .B1(_3093_),
    .Y(_3115_));
 sky130_fd_sc_hd__o21ai_0 _6963_ (.A1(net772),
    .A2(_3115_),
    .B1(_3064_),
    .Y(_3116_));
 sky130_fd_sc_hd__o211ai_1 _6964_ (.A1(net98),
    .A2(net335),
    .B1(_3057_),
    .C1(_3116_),
    .Y(_3117_));
 sky130_fd_sc_hd__o221ai_4 _6965_ (.A1(_2686_),
    .A2(_2929_),
    .B1(_2932_),
    .B2(_2646_),
    .C1(_3117_),
    .Y(\dp.result2[20] ));
 sky130_fd_sc_hd__a21oi_1 _6966_ (.A1(net46),
    .A2(_3090_),
    .B1(_3093_),
    .Y(_3118_));
 sky130_fd_sc_hd__o21ai_0 _6967_ (.A1(net772),
    .A2(_3118_),
    .B1(_3064_),
    .Y(_3119_));
 sky130_fd_sc_hd__a22oi_1 _6968_ (.A1(_0896_),
    .A2(_2937_),
    .B1(_2942_),
    .B2(_3056_),
    .Y(_3120_));
 sky130_fd_sc_hd__o211a_4 _6969_ (.A1(net334),
    .A2(_3058_),
    .B1(_3119_),
    .C1(_3120_),
    .X(\dp.result2[21] ));
 sky130_fd_sc_hd__nand2_1 _6970_ (.A(_3056_),
    .B(_2950_),
    .Y(_3121_));
 sky130_fd_sc_hd__a21oi_1 _6971_ (.A1(net47),
    .A2(_3090_),
    .B1(_3093_),
    .Y(_3122_));
 sky130_fd_sc_hd__o21ai_0 _6972_ (.A1(net772),
    .A2(_3122_),
    .B1(_3064_),
    .Y(_3123_));
 sky130_fd_sc_hd__nand2_1 _6973_ (.A(_0896_),
    .B(_2944_),
    .Y(_3124_));
 sky130_fd_sc_hd__o2111a_4 _6974_ (.A1(net259),
    .A2(_3058_),
    .B1(_3121_),
    .C1(_3123_),
    .D1(_3124_),
    .X(\dp.result2[22] ));
 sky130_fd_sc_hd__a21oi_1 _6975_ (.A1(net48),
    .A2(_3090_),
    .B1(_3093_),
    .Y(_3125_));
 sky130_fd_sc_hd__o21ai_0 _6976_ (.A1(net772),
    .A2(_3125_),
    .B1(_3064_),
    .Y(_3126_));
 sky130_fd_sc_hd__nand2_1 _6977_ (.A(_0896_),
    .B(_2953_),
    .Y(_3127_));
 sky130_fd_sc_hd__nand2_1 _6978_ (.A(_3056_),
    .B(_2957_),
    .Y(_3128_));
 sky130_fd_sc_hd__o2111a_4 _6979_ (.A1(net254),
    .A2(_3058_),
    .B1(_3126_),
    .C1(_3127_),
    .D1(_3128_),
    .X(\dp.result2[23] ));
 sky130_fd_sc_hd__nand2_1 _6980_ (.A(_3056_),
    .B(_2966_),
    .Y(_3129_));
 sky130_fd_sc_hd__a21oi_1 _6981_ (.A1(net49),
    .A2(_3090_),
    .B1(_3093_),
    .Y(_3130_));
 sky130_fd_sc_hd__o21ai_0 _6982_ (.A1(net772),
    .A2(_3130_),
    .B1(_3064_),
    .Y(_3131_));
 sky130_fd_sc_hd__nand2_1 _6983_ (.A(_0896_),
    .B(_2960_),
    .Y(_3132_));
 sky130_fd_sc_hd__o2111a_4 _6984_ (.A1(net257),
    .A2(_3058_),
    .B1(_3129_),
    .C1(_3131_),
    .D1(_3132_),
    .X(\dp.result2[24] ));
 sky130_fd_sc_hd__a21oi_1 _6985_ (.A1(net50),
    .A2(_3090_),
    .B1(_3093_),
    .Y(_3133_));
 sky130_fd_sc_hd__o21ai_0 _6986_ (.A1(net772),
    .A2(_3133_),
    .B1(_3064_),
    .Y(_3134_));
 sky130_fd_sc_hd__a22oi_1 _6987_ (.A1(_0896_),
    .A2(_2968_),
    .B1(_2974_),
    .B2(_3056_),
    .Y(_3135_));
 sky130_fd_sc_hd__o211a_4 _6988_ (.A1(net255),
    .A2(_3058_),
    .B1(_3134_),
    .C1(_3135_),
    .X(\dp.result2[25] ));
 sky130_fd_sc_hd__nor2_4 _6989_ (.A(net98),
    .B(_3069_),
    .Y(_3136_));
 sky130_fd_sc_hd__a21oi_1 _6990_ (.A1(net51),
    .A2(_3090_),
    .B1(_3093_),
    .Y(_3137_));
 sky130_fd_sc_hd__o21ai_0 _6991_ (.A1(net772),
    .A2(_3137_),
    .B1(_3064_),
    .Y(_3138_));
 sky130_fd_sc_hd__nand2_1 _6992_ (.A(_0896_),
    .B(_2977_),
    .Y(_3139_));
 sky130_fd_sc_hd__nand2_1 _6993_ (.A(_3138_),
    .B(_3139_),
    .Y(_3140_));
 sky130_fd_sc_hd__a221oi_2 _6994_ (.A1(_3056_),
    .A2(_2982_),
    .B1(_3136_),
    .B2(net221),
    .C1(_3140_),
    .Y(\dp.result2[26] ));
 sky130_fd_sc_hd__a21oi_1 _6995_ (.A1(net52),
    .A2(_3090_),
    .B1(_3093_),
    .Y(_3141_));
 sky130_fd_sc_hd__o21ai_0 _6996_ (.A1(net772),
    .A2(_3141_),
    .B1(_3064_),
    .Y(_3142_));
 sky130_fd_sc_hd__o211ai_1 _6997_ (.A1(net98),
    .A2(net85),
    .B1(_3057_),
    .C1(_3142_),
    .Y(_3143_));
 sky130_fd_sc_hd__o221ai_2 _6998_ (.A1(_2686_),
    .A2(_2984_),
    .B1(_2991_),
    .B2(_2646_),
    .C1(_3143_),
    .Y(\dp.result2[27] ));
 sky130_fd_sc_hd__a21oi_1 _6999_ (.A1(net53),
    .A2(_3090_),
    .B1(_3093_),
    .Y(_3144_));
 sky130_fd_sc_hd__o21ai_0 _7000_ (.A1(net772),
    .A2(_3144_),
    .B1(_3064_),
    .Y(_3145_));
 sky130_fd_sc_hd__nand2_2 _7001_ (.A(_0896_),
    .B(_2993_),
    .Y(_3146_));
 sky130_fd_sc_hd__nand2_1 _7002_ (.A(_3056_),
    .B(_2996_),
    .Y(_3147_));
 sky130_fd_sc_hd__o2111a_4 _7003_ (.A1(net327),
    .A2(_3058_),
    .B1(_3145_),
    .C1(_3146_),
    .D1(_3147_),
    .X(\dp.result2[28] ));
 sky130_fd_sc_hd__o22ai_2 _7004_ (.A1(_2686_),
    .A2(_2998_),
    .B1(_3004_),
    .B2(_2646_),
    .Y(_3148_));
 sky130_fd_sc_hd__nor3b_1 _7005_ (.A(_3148_),
    .B(net98),
    .C_N(_2573_),
    .Y(_3149_));
 sky130_fd_sc_hd__a21oi_1 _7006_ (.A1(net54),
    .A2(_3090_),
    .B1(_3093_),
    .Y(_3150_));
 sky130_fd_sc_hd__o21ai_0 _7007_ (.A1(net772),
    .A2(_3150_),
    .B1(_3064_),
    .Y(_3151_));
 sky130_fd_sc_hd__a31oi_1 _7008_ (.A1(_2584_),
    .A2(_3057_),
    .A3(_3151_),
    .B1(_3148_),
    .Y(_3152_));
 sky130_fd_sc_hd__a21oi_2 _7009_ (.A1(_2570_),
    .A2(_3149_),
    .B1(_3152_),
    .Y(\dp.result2[29] ));
 sky130_fd_sc_hd__a22oi_1 _7010_ (.A1(net122),
    .A2(_0896_),
    .B1(_3056_),
    .B2(_3005_),
    .Y(_3153_));
 sky130_fd_sc_hd__o221a_4 _7011_ (.A1(net55),
    .A2(_1875_),
    .B1(net378),
    .B2(_3058_),
    .C1(_3153_),
    .X(\dp.result2[2] ));
 sky130_fd_sc_hd__a21oi_1 _7012_ (.A1(net56),
    .A2(_3090_),
    .B1(_3093_),
    .Y(_3154_));
 sky130_fd_sc_hd__o21ai_0 _7013_ (.A1(net772),
    .A2(_3154_),
    .B1(_3064_),
    .Y(_3155_));
 sky130_fd_sc_hd__o211ai_1 _7014_ (.A1(net98),
    .A2(net261),
    .B1(_3057_),
    .C1(_3155_),
    .Y(_3156_));
 sky130_fd_sc_hd__o221ai_4 _7015_ (.A1(_2686_),
    .A2(_3008_),
    .B1(_3014_),
    .B2(_2646_),
    .C1(_3156_),
    .Y(\dp.result2[30] ));
 sky130_fd_sc_hd__o22a_4 _7016_ (.A1(_2686_),
    .A2(_3016_),
    .B1(_3028_),
    .B2(_2646_),
    .X(_3157_));
 sky130_fd_sc_hd__nand3_1 _7017_ (.A(_1875_),
    .B(_2615_),
    .C(_3157_),
    .Y(_3158_));
 sky130_fd_sc_hd__a31oi_1 _7018_ (.A1(_1727_),
    .A2(_2609_),
    .A3(_2611_),
    .B1(_3158_),
    .Y(_3159_));
 sky130_fd_sc_hd__a21oi_1 _7019_ (.A1(net57),
    .A2(_3090_),
    .B1(_3093_),
    .Y(_3160_));
 sky130_fd_sc_hd__o21ai_0 _7020_ (.A1(net772),
    .A2(_3160_),
    .B1(_3064_),
    .Y(_3161_));
 sky130_fd_sc_hd__nand2_1 _7021_ (.A(_3057_),
    .B(_3161_),
    .Y(_3162_));
 sky130_fd_sc_hd__o21a_1 _7022_ (.A1(_2624_),
    .A2(_3162_),
    .B1(_3157_),
    .X(_3163_));
 sky130_fd_sc_hd__nor2_2 _7023_ (.A(_3159_),
    .B(_3163_),
    .Y(\dp.result2[31] ));
 sky130_fd_sc_hd__a22o_1 _7024_ (.A1(net58),
    .A2(net98),
    .B1(_3056_),
    .B2(_3031_),
    .X(_3164_));
 sky130_fd_sc_hd__a221o_4 _7025_ (.A1(_3462_[0]),
    .A2(_0896_),
    .B1(net340),
    .B2(_3136_),
    .C1(_3164_),
    .X(\dp.result2[3] ));
 sky130_fd_sc_hd__nand2_1 _7026_ (.A(_0896_),
    .B(_3032_),
    .Y(_3165_));
 sky130_fd_sc_hd__nor2_1 _7027_ (.A(net59),
    .B(_1875_),
    .Y(_3166_));
 sky130_fd_sc_hd__a21oi_1 _7028_ (.A1(_3056_),
    .A2(_3033_),
    .B1(_3166_),
    .Y(_3167_));
 sky130_fd_sc_hd__o211a_4 _7029_ (.A1(net381),
    .A2(_3058_),
    .B1(_3165_),
    .C1(_3167_),
    .X(\dp.result2[4] ));
 sky130_fd_sc_hd__a22oi_1 _7030_ (.A1(_0896_),
    .A2(_3035_),
    .B1(_3038_),
    .B2(_3056_),
    .Y(_3168_));
 sky130_fd_sc_hd__o221a_4 _7031_ (.A1(net60),
    .A2(_1875_),
    .B1(net377),
    .B2(_3058_),
    .C1(_3168_),
    .X(\dp.result2[5] ));
 sky130_fd_sc_hd__a22oi_2 _7032_ (.A1(_0896_),
    .A2(_3039_),
    .B1(_3042_),
    .B2(_3056_),
    .Y(_3169_));
 sky130_fd_sc_hd__o221a_4 _7033_ (.A1(net61),
    .A2(_1875_),
    .B1(net312),
    .B2(_3058_),
    .C1(_3169_),
    .X(\dp.result2[6] ));
 sky130_fd_sc_hd__nor2_1 _7034_ (.A(net62),
    .B(_1875_),
    .Y(_3170_));
 sky130_fd_sc_hd__a221oi_1 _7035_ (.A1(_0896_),
    .A2(_3043_),
    .B1(_3046_),
    .B2(_3056_),
    .C1(_3170_),
    .Y(_3171_));
 sky130_fd_sc_hd__o21a_4 _7036_ (.A1(net382),
    .A2(_3058_),
    .B1(_3171_),
    .X(\dp.result2[7] ));
 sky130_fd_sc_hd__nand2_1 _7037_ (.A(net63),
    .B(_3067_),
    .Y(_3172_));
 sky130_fd_sc_hd__a222oi_1 _7038_ (.A1(_0896_),
    .A2(_3047_),
    .B1(_3064_),
    .B2(_3172_),
    .C1(_3050_),
    .C2(_3056_),
    .Y(_3173_));
 sky130_fd_sc_hd__o21a_4 _7039_ (.A1(net360),
    .A2(_3058_),
    .B1(_3173_),
    .X(\dp.result2[8] ));
 sky130_fd_sc_hd__nand2_1 _7040_ (.A(net64),
    .B(_3067_),
    .Y(_3174_));
 sky130_fd_sc_hd__a21oi_1 _7041_ (.A1(_3064_),
    .A2(_3174_),
    .B1(_3069_),
    .Y(_3175_));
 sky130_fd_sc_hd__o21ai_2 _7042_ (.A1(net98),
    .A2(net371),
    .B1(_3175_),
    .Y(_3176_));
 sky130_fd_sc_hd__o221ai_4 _7043_ (.A1(_2686_),
    .A2(_3052_),
    .B1(_3055_),
    .B2(_2646_),
    .C1(_3176_),
    .Y(\dp.result2[9] ));
 sky130_fd_sc_hd__and4_1 _7044_ (.A(net27),
    .B(net28),
    .C(net29),
    .D(net803),
    .X(net132));
 sky130_fd_sc_hd__and3_4 _7045_ (.A(net99),
    .B(_3066_),
    .C(_1713_),
    .X(_3177_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__nor2_1 _7047_ (.A(_1295_),
    .B(_3177_),
    .Y(net134));
 sky130_fd_sc_hd__inv_1 _7048_ (.A(_3177_),
    .Y(_3179_));
 sky130_fd_sc_hd__and2_0 _7049_ (.A(_1253_),
    .B(_3179_),
    .X(net135));
 sky130_fd_sc_hd__nor3_1 _7050_ (.A(_0111_),
    .B(_1214_),
    .C(_3177_),
    .Y(net136));
 sky130_fd_sc_hd__nor2b_1 _7051_ (.A(_3177_),
    .B_N(_1173_),
    .Y(net137));
 sky130_fd_sc_hd__nor2_1 _7052_ (.A(_1125_),
    .B(_3177_),
    .Y(net138));
 sky130_fd_sc_hd__nor2b_1 _7053_ (.A(_3177_),
    .B_N(_1088_),
    .Y(net139));
 sky130_fd_sc_hd__nor2_4 _7054_ (.A(net5),
    .B(_0044_),
    .Y(_3180_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__nor2_1 _7056_ (.A(_1039_),
    .B(_3180_),
    .Y(net140));
 sky130_fd_sc_hd__nor2_1 _7057_ (.A(_0994_),
    .B(_3180_),
    .Y(net141));
 sky130_fd_sc_hd__nor2_1 _7058_ (.A(_0952_),
    .B(_3180_),
    .Y(net142));
 sky130_fd_sc_hd__nor2_1 _7059_ (.A(_2749_),
    .B(_3180_),
    .Y(net143));
 sky130_fd_sc_hd__nor2_1 _7060_ (.A(_0866_),
    .B(_3180_),
    .Y(net145));
 sky130_fd_sc_hd__o21a_1 _7061_ (.A1(net5),
    .A2(_0044_),
    .B1(_0821_),
    .X(net146));
 sky130_fd_sc_hd__nor2_1 _7062_ (.A(_0782_),
    .B(_3180_),
    .Y(net147));
 sky130_fd_sc_hd__nor2_1 _7063_ (.A(_0732_),
    .B(_3180_),
    .Y(net148));
 sky130_fd_sc_hd__nor2_1 _7064_ (.A(_0690_),
    .B(_3180_),
    .Y(net149));
 sky130_fd_sc_hd__inv_1 _7065_ (.A(_0637_),
    .Y(_3182_));
 sky130_fd_sc_hd__nor2_1 _7066_ (.A(_3182_),
    .B(_3180_),
    .Y(net150));
 sky130_fd_sc_hd__nor2_1 _7067_ (.A(_0598_),
    .B(_3180_),
    .Y(net151));
 sky130_fd_sc_hd__inv_1 _7068_ (.A(_0543_),
    .Y(_3183_));
 sky130_fd_sc_hd__nor2_1 _7069_ (.A(_3183_),
    .B(_3180_),
    .Y(net152));
 sky130_fd_sc_hd__nor2_1 _7070_ (.A(_2782_),
    .B(_3180_),
    .Y(net153));
 sky130_fd_sc_hd__nor2_1 _7071_ (.A(_0447_),
    .B(_3180_),
    .Y(net154));
 sky130_fd_sc_hd__nor2_1 _7072_ (.A(_0369_),
    .B(_3180_),
    .Y(net156));
 sky130_fd_sc_hd__nor2_1 _7073_ (.A(_0338_),
    .B(_3180_),
    .Y(net157));
 sky130_fd_sc_hd__nor2_1 _7074_ (.A(_1377_),
    .B(_3177_),
    .Y(net163));
 sky130_fd_sc_hd__nor2_1 _7075_ (.A(_1336_),
    .B(_3177_),
    .Y(net164));
 sky130_fd_sc_hd__fa_2 _7076_ (.A(_3184_[0]),
    .B(_3185_[0]),
    .CIN(_3186_[0]),
    .COUT(_3187_[0]),
    .SUM(_3188_[0]));
 sky130_fd_sc_hd__fa_1 _7077_ (.A(_3189_[0]),
    .B(_3190_[0]),
    .CIN(_3191_[0]),
    .COUT(_3192_[0]),
    .SUM(_3193_[0]));
 sky130_fd_sc_hd__ha_1 _7078_ (.A(_3194_[0]),
    .B(_3195_[0]),
    .COUT(_3196_[0]),
    .SUM(_3197_[0]));
 sky130_fd_sc_hd__ha_1 _7079_ (.A(_0237_),
    .B(_3199_[0]),
    .COUT(_3200_[0]),
    .SUM(_3201_[0]));
 sky130_fd_sc_hd__ha_1 _7080_ (.A(_3202_[0]),
    .B(_0313_),
    .COUT(_3204_[0]),
    .SUM(_3205_[0]));
 sky130_fd_sc_hd__ha_1 _7081_ (.A(_3206_[0]),
    .B(_0314_),
    .COUT(_3208_[0]),
    .SUM(_3209_[0]));
 sky130_fd_sc_hd__ha_4 _7082_ (.A(_3210_[0]),
    .B(_3211_[0]),
    .COUT(_3212_[0]),
    .SUM(_3213_[0]));
 sky130_fd_sc_hd__ha_1 _7083_ (.A(net767),
    .B(_3215_[0]),
    .COUT(_3216_[0]),
    .SUM(_3217_[0]));
 sky130_fd_sc_hd__ha_4 _7084_ (.A(_0490_),
    .B(_3219_[0]),
    .COUT(_3220_[0]),
    .SUM(_3221_[0]));
 sky130_fd_sc_hd__ha_1 _7085_ (.A(_3222_[0]),
    .B(_3223_[0]),
    .COUT(_3224_[0]),
    .SUM(_3225_[0]));
 sky130_fd_sc_hd__ha_4 _7086_ (.A(_3226_[0]),
    .B(_3227_[0]),
    .COUT(_3228_[0]),
    .SUM(_3229_[0]));
 sky130_fd_sc_hd__ha_1 _7087_ (.A(_3230_[0]),
    .B(_3231_[0]),
    .COUT(_3232_[0]),
    .SUM(_3233_[0]));
 sky130_fd_sc_hd__ha_1 _7088_ (.A(_3234_[0]),
    .B(_3235_[0]),
    .COUT(_3236_[0]),
    .SUM(_3237_[0]));
 sky130_fd_sc_hd__ha_1 _7089_ (.A(net766),
    .B(_3239_[0]),
    .COUT(_3240_[0]),
    .SUM(_3241_[0]));
 sky130_fd_sc_hd__ha_4 _7090_ (.A(_3242_[0]),
    .B(_3243_[0]),
    .COUT(_3244_[0]),
    .SUM(_3245_[0]));
 sky130_fd_sc_hd__ha_1 _7091_ (.A(_3246_[0]),
    .B(_3247_[0]),
    .COUT(_3248_[0]),
    .SUM(_3249_[0]));
 sky130_fd_sc_hd__ha_4 _7092_ (.A(_3250_[0]),
    .B(_3251_[0]),
    .COUT(_3252_[0]),
    .SUM(_3253_[0]));
 sky130_fd_sc_hd__ha_1 _7093_ (.A(_3254_[0]),
    .B(_3255_[0]),
    .COUT(_3256_[0]),
    .SUM(_3257_[0]));
 sky130_fd_sc_hd__ha_4 _7094_ (.A(_3258_[0]),
    .B(_3259_[0]),
    .COUT(_3260_[0]),
    .SUM(_3261_[0]));
 sky130_fd_sc_hd__ha_1 _7095_ (.A(_3262_[0]),
    .B(_3263_[0]),
    .COUT(_3264_[0]),
    .SUM(_3265_[0]));
 sky130_fd_sc_hd__ha_4 _7096_ (.A(_3266_[0]),
    .B(_3267_[0]),
    .COUT(_3268_[0]),
    .SUM(_3269_[0]));
 sky130_fd_sc_hd__ha_1 _7097_ (.A(net281),
    .B(_3271_[0]),
    .COUT(_3272_[0]),
    .SUM(_3273_[0]));
 sky130_fd_sc_hd__ha_2 _7098_ (.A(_3274_[0]),
    .B(_3275_[0]),
    .COUT(_3276_[0]),
    .SUM(_3277_[0]));
 sky130_fd_sc_hd__ha_1 _7099_ (.A(_3278_[0]),
    .B(_3279_[0]),
    .COUT(_3280_[0]),
    .SUM(_3281_[0]));
 sky130_fd_sc_hd__ha_4 _7100_ (.A(_3282_[0]),
    .B(_3283_[0]),
    .COUT(_3284_[0]),
    .SUM(_3285_[0]));
 sky130_fd_sc_hd__ha_1 _7101_ (.A(_3286_[0]),
    .B(_3287_[0]),
    .COUT(_3288_[0]),
    .SUM(_3289_[0]));
 sky130_fd_sc_hd__ha_4 _7102_ (.A(_3290_[0]),
    .B(_3291_[0]),
    .COUT(_3292_[0]),
    .SUM(_3293_[0]));
 sky130_fd_sc_hd__ha_1 _7103_ (.A(_3294_[0]),
    .B(_3295_[0]),
    .COUT(_3296_[0]),
    .SUM(_3297_[0]));
 sky130_fd_sc_hd__ha_4 _7104_ (.A(_3298_[0]),
    .B(_3299_[0]),
    .COUT(_3300_[0]),
    .SUM(_3301_[0]));
 sky130_fd_sc_hd__ha_1 _7105_ (.A(net765),
    .B(_3303_[0]),
    .COUT(_3304_[0]),
    .SUM(_3305_[0]));
 sky130_fd_sc_hd__ha_4 _7106_ (.A(_3306_[0]),
    .B(_3307_[0]),
    .COUT(_3308_[0]),
    .SUM(_3309_[0]));
 sky130_fd_sc_hd__ha_1 _7107_ (.A(_3310_[0]),
    .B(_3311_[0]),
    .COUT(_3312_[0]),
    .SUM(_3313_[0]));
 sky130_fd_sc_hd__ha_4 _7108_ (.A(_3314_[0]),
    .B(_3315_[0]),
    .COUT(_3316_[0]),
    .SUM(_3317_[0]));
 sky130_fd_sc_hd__ha_1 _7109_ (.A(net764),
    .B(_3319_[0]),
    .COUT(_3320_[0]),
    .SUM(_3321_[0]));
 sky130_fd_sc_hd__ha_1 _7110_ (.A(_3322_[0]),
    .B(_3323_[0]),
    .COUT(_3324_[0]),
    .SUM(_3325_[0]));
 sky130_fd_sc_hd__ha_1 _7111_ (.A(_3326_[0]),
    .B(_3327_[0]),
    .COUT(_3328_[0]),
    .SUM(_3329_[0]));
 sky130_fd_sc_hd__ha_1 _7112_ (.A(_3330_[0]),
    .B(_3331_[0]),
    .COUT(_3332_[0]),
    .SUM(_3333_[0]));
 sky130_fd_sc_hd__ha_1 _7113_ (.A(net763),
    .B(_3335_[0]),
    .COUT(_3336_[0]),
    .SUM(_3337_[0]));
 sky130_fd_sc_hd__ha_1 _7114_ (.A(_3339_[0]),
    .B(_3338_[0]),
    .COUT(_3340_[0]),
    .SUM(_3341_[0]));
 sky130_fd_sc_hd__ha_1 _7115_ (.A(_3342_[0]),
    .B(_3343_[0]),
    .COUT(_3344_[0]),
    .SUM(_3345_[0]));
 sky130_fd_sc_hd__ha_1 _7116_ (.A(_3346_[0]),
    .B(_3347_[0]),
    .COUT(_3348_[0]),
    .SUM(_3349_[0]));
 sky130_fd_sc_hd__ha_1 _7117_ (.A(_1203_),
    .B(_3351_[0]),
    .COUT(_3352_[0]),
    .SUM(_3353_[0]));
 sky130_fd_sc_hd__ha_4 _7118_ (.A(_3354_[0]),
    .B(_3355_[0]),
    .COUT(_3356_[0]),
    .SUM(_3357_[0]));
 sky130_fd_sc_hd__ha_1 _7119_ (.A(net761),
    .B(_3359_[0]),
    .COUT(_3360_[0]),
    .SUM(_3361_[0]));
 sky130_fd_sc_hd__ha_4 _7120_ (.A(_3362_[0]),
    .B(_3363_[0]),
    .COUT(_3364_[0]),
    .SUM(_3365_[0]));
 sky130_fd_sc_hd__ha_1 _7121_ (.A(net760),
    .B(_3367_[0]),
    .COUT(_3368_[0]),
    .SUM(_3369_[0]));
 sky130_fd_sc_hd__ha_4 _7122_ (.A(_3370_[0]),
    .B(_3371_[0]),
    .COUT(_3372_[0]),
    .SUM(_3373_[0]));
 sky130_fd_sc_hd__ha_1 _7123_ (.A(net759),
    .B(_3375_[0]),
    .COUT(_3376_[0]),
    .SUM(_3377_[0]));
 sky130_fd_sc_hd__ha_2 _7124_ (.A(_3378_[0]),
    .B(_3379_[0]),
    .COUT(_3380_[0]),
    .SUM(_3381_[0]));
 sky130_fd_sc_hd__ha_1 _7125_ (.A(net758),
    .B(_3383_[0]),
    .COUT(_3384_[0]),
    .SUM(_3385_[0]));
 sky130_fd_sc_hd__ha_2 _7126_ (.A(_3386_[0]),
    .B(_3387_[0]),
    .COUT(_3388_[0]),
    .SUM(_3389_[0]));
 sky130_fd_sc_hd__ha_1 _7127_ (.A(net757),
    .B(_3391_[0]),
    .COUT(_3392_[0]),
    .SUM(_3393_[0]));
 sky130_fd_sc_hd__ha_4 _7128_ (.A(_3394_[0]),
    .B(_3395_[0]),
    .COUT(_3396_[0]),
    .SUM(_3397_[0]));
 sky130_fd_sc_hd__ha_1 _7129_ (.A(net756),
    .B(_3399_[0]),
    .COUT(_3400_[0]),
    .SUM(_3401_[0]));
 sky130_fd_sc_hd__ha_4 _7130_ (.A(_3402_[0]),
    .B(_3403_[0]),
    .COUT(_3404_[0]),
    .SUM(_3405_[0]));
 sky130_fd_sc_hd__ha_1 _7131_ (.A(net755),
    .B(_3407_[0]),
    .COUT(_3408_[0]),
    .SUM(_3409_[0]));
 sky130_fd_sc_hd__ha_1 _7132_ (.A(_3410_[0]),
    .B(_3411_[0]),
    .COUT(_3412_[0]),
    .SUM(_3413_[0]));
 sky130_fd_sc_hd__ha_1 _7133_ (.A(net754),
    .B(_3415_[0]),
    .COUT(_3416_[0]),
    .SUM(_3417_[0]));
 sky130_fd_sc_hd__ha_4 _7134_ (.A(_3418_[0]),
    .B(_3419_[0]),
    .COUT(_3420_[0]),
    .SUM(_3421_[0]));
 sky130_fd_sc_hd__ha_1 _7135_ (.A(net753),
    .B(_3423_[0]),
    .COUT(_3424_[0]),
    .SUM(_3425_[0]));
 sky130_fd_sc_hd__ha_4 _7136_ (.A(_3427_[0]),
    .B(_3426_[0]),
    .COUT(_3428_[0]),
    .SUM(_3429_[0]));
 sky130_fd_sc_hd__ha_1 _7137_ (.A(_3430_[0]),
    .B(_3431_[0]),
    .COUT(_3432_[0]),
    .SUM(_3433_[0]));
 sky130_fd_sc_hd__ha_4 _7138_ (.A(_3434_[0]),
    .B(_3435_[0]),
    .COUT(_3436_[0]),
    .SUM(_3437_[0]));
 sky130_fd_sc_hd__ha_1 _7139_ (.A(_3438_[0]),
    .B(_3439_[0]),
    .COUT(_3440_[0]),
    .SUM(_3441_[0]));
 sky130_fd_sc_hd__ha_4 _7140_ (.A(_3185_[0]),
    .B(_3186_[0]),
    .COUT(_3442_[0]),
    .SUM(_3443_[0]));
 sky130_fd_sc_hd__ha_1 _7141_ (.A(_1699_),
    .B(_3445_[0]),
    .COUT(_3446_[0]),
    .SUM(_3447_[0]));
 sky130_fd_sc_hd__ha_1 _7142_ (.A(_3448_[0]),
    .B(_3449_[0]),
    .COUT(_3189_[0]),
    .SUM(_3450_[0]));
 sky130_fd_sc_hd__ha_1 _7143_ (.A(_3190_[0]),
    .B(_3191_[0]),
    .COUT(_3451_[0]),
    .SUM(_3452_[0]));
 sky130_fd_sc_hd__ha_2 _7144_ (.A(_3453_[0]),
    .B(_3454_[0]),
    .COUT(_3455_[0]),
    .SUM(_3456_[0]));
 sky130_fd_sc_hd__ha_1 _7145_ (.A(_3457_[0]),
    .B(_3458_[0]),
    .COUT(_3459_[0]),
    .SUM(_3460_[0]));
 sky130_fd_sc_hd__ha_4 _7146_ (.A(net122),
    .B(net125),
    .COUT(_3461_[0]),
    .SUM(_3462_[0]));
 sky130_fd_sc_hd__ha_4 _7147_ (.A(_3463_[0]),
    .B(_3464_[0]),
    .COUT(_3465_[0]),
    .SUM(_3466_[0]));
 sky130_fd_sc_hd__ha_4 _7148_ (.A(_3467_[0]),
    .B(_3468_[0]),
    .COUT(_3469_[0]),
    .SUM(_3470_[0]));
 sky130_fd_sc_hd__ha_4 _7149_ (.A(_3471_[0]),
    .B(_3472_[0]),
    .COUT(_3473_[0]),
    .SUM(_3474_[0]));
 sky130_fd_sc_hd__ha_4 _7150_ (.A(_3475_[0]),
    .B(_3476_[0]),
    .COUT(_3477_[0]),
    .SUM(_3478_[0]));
 sky130_fd_sc_hd__ha_1 _7151_ (.A(_3479_[0]),
    .B(_3480_[0]),
    .COUT(_3481_[0]),
    .SUM(_3482_[0]));
 sky130_fd_sc_hd__ha_1 _7152_ (.A(_3483_[0]),
    .B(_3484_[0]),
    .COUT(_3485_[0]),
    .SUM(_3486_[0]));
 sky130_fd_sc_hd__ha_1 _7153_ (.A(_3487_[0]),
    .B(_3488_[0]),
    .COUT(_3489_[0]),
    .SUM(_3490_[0]));
 sky130_fd_sc_hd__ha_2 _7154_ (.A(_3491_[0]),
    .B(_3492_[0]),
    .COUT(_3493_[0]),
    .SUM(_3494_[0]));
 sky130_fd_sc_hd__ha_1 _7155_ (.A(_3495_[0]),
    .B(_3496_[0]),
    .COUT(_3497_[0]),
    .SUM(_3498_[0]));
 sky130_fd_sc_hd__ha_1 _7156_ (.A(_3499_[0]),
    .B(_3500_[0]),
    .COUT(_3501_[0]),
    .SUM(_3502_[0]));
 sky130_fd_sc_hd__ha_1 _7157_ (.A(_3503_[0]),
    .B(_3504_[0]),
    .COUT(_3505_[0]),
    .SUM(_3506_[0]));
 sky130_fd_sc_hd__ha_1 _7158_ (.A(_3507_[0]),
    .B(_3508_[0]),
    .COUT(_3509_[0]),
    .SUM(_3510_[0]));
 sky130_fd_sc_hd__ha_4 _7159_ (.A(_3511_[0]),
    .B(_3512_[0]),
    .COUT(_3513_[0]),
    .SUM(_3514_[0]));
 sky130_fd_sc_hd__ha_2 _7160_ (.A(_3515_[0]),
    .B(_3516_[0]),
    .COUT(_3517_[0]),
    .SUM(_3518_[0]));
 sky130_fd_sc_hd__ha_4 _7161_ (.A(_3519_[0]),
    .B(_3520_[0]),
    .COUT(_3521_[0]),
    .SUM(_3522_[0]));
 sky130_fd_sc_hd__ha_2 _7162_ (.A(_3523_[0]),
    .B(_3524_[0]),
    .COUT(_3525_[0]),
    .SUM(_3526_[0]));
 sky130_fd_sc_hd__ha_1 _7163_ (.A(_3527_[0]),
    .B(_3528_[0]),
    .COUT(_3529_[0]),
    .SUM(_3530_[0]));
 sky130_fd_sc_hd__ha_2 _7164_ (.A(_3531_[0]),
    .B(_3532_[0]),
    .COUT(_3533_[0]),
    .SUM(_3534_[0]));
 sky130_fd_sc_hd__ha_2 _7165_ (.A(_3535_[0]),
    .B(_3536_[0]),
    .COUT(_3537_[0]),
    .SUM(_3538_[0]));
 sky130_fd_sc_hd__ha_2 _7166_ (.A(_3539_[0]),
    .B(_3540_[0]),
    .COUT(_3541_[0]),
    .SUM(_3542_[0]));
 sky130_fd_sc_hd__ha_2 _7167_ (.A(_3543_[0]),
    .B(_3544_[0]),
    .COUT(_3545_[0]),
    .SUM(_3546_[0]));
 sky130_fd_sc_hd__ha_1 _7168_ (.A(_3547_[0]),
    .B(_3548_[0]),
    .COUT(_3549_[0]),
    .SUM(_3550_[0]));
 sky130_fd_sc_hd__ha_4 _7169_ (.A(_3551_[0]),
    .B(_3552_[0]),
    .COUT(_3553_[0]),
    .SUM(_3554_[0]));
 sky130_fd_sc_hd__ha_4 _7170_ (.A(_3555_[0]),
    .B(_3556_[0]),
    .COUT(_3557_[0]),
    .SUM(_3558_[0]));
 sky130_fd_sc_hd__ha_4 _7171_ (.A(_3559_[0]),
    .B(_3560_[0]),
    .COUT(_3561_[0]),
    .SUM(_3562_[0]));
 sky130_fd_sc_hd__ha_4 _7172_ (.A(_3563_[0]),
    .B(_3564_[0]),
    .COUT(_3565_[0]),
    .SUM(_3566_[0]));
 sky130_fd_sc_hd__ha_2 _7173_ (.A(_3567_[0]),
    .B(_3568_[0]),
    .COUT(_3569_[0]),
    .SUM(_3570_[0]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[0]$_DFFE_PP0P_  (.D(_0032_),
    .Q(net100),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[10]$_DFF_PP0_  (.D(\dp.ISRmux.d0[10] ),
    .Q(net101),
    .RESET_B(_0031_),
    .CLK(clknet_5_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[11]$_DFF_PP0_  (.D(\dp.ISRmux.d0[11] ),
    .Q(net102),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[12]$_DFF_PP0_  (.D(\dp.ISRmux.d0[12] ),
    .Q(net103),
    .RESET_B(_0031_),
    .CLK(clknet_5_7__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[13]$_DFF_PP0_  (.D(\dp.ISRmux.d0[13] ),
    .Q(net104),
    .RESET_B(_0031_),
    .CLK(clknet_5_26__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[14]$_DFF_PP0_  (.D(\dp.ISRmux.d0[14] ),
    .Q(net105),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[15]$_DFF_PP0_  (.D(\dp.ISRmux.d0[15] ),
    .Q(net106),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[16]$_DFF_PP0_  (.D(\dp.ISRmux.d0[16] ),
    .Q(net107),
    .RESET_B(_0031_),
    .CLK(clknet_5_27__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[17]$_DFF_PP0_  (.D(\dp.ISRmux.d0[17] ),
    .Q(net108),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[18]$_DFF_PP0_  (.D(\dp.ISRmux.d0[18] ),
    .Q(net109),
    .RESET_B(_0031_),
    .CLK(clknet_5_27__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[19]$_DFF_PP0_  (.D(\dp.ISRmux.d0[19] ),
    .Q(net110),
    .RESET_B(_0031_),
    .CLK(clknet_5_27__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[1]$_DFFE_PP0P_  (.D(_0033_),
    .Q(net111),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[20]$_DFF_PP0_  (.D(\dp.ISRmux.d0[20] ),
    .Q(net112),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[21]$_DFF_PP0_  (.D(\dp.ISRmux.d0[21] ),
    .Q(net113),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[22]$_DFF_PP0_  (.D(\dp.ISRmux.d0[22] ),
    .Q(net114),
    .RESET_B(_0031_),
    .CLK(clknet_5_30__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[23]$_DFF_PP0_  (.D(\dp.ISRmux.d0[23] ),
    .Q(net115),
    .RESET_B(_0031_),
    .CLK(clknet_5_30__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[24]$_DFF_PP0_  (.D(\dp.ISRmux.d0[24] ),
    .Q(net116),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[25]$_DFF_PP0_  (.D(\dp.ISRmux.d0[25] ),
    .Q(net117),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[26]$_DFF_PP0_  (.D(\dp.ISRmux.d0[26] ),
    .Q(net118),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[27]$_DFF_PP0_  (.D(\dp.ISRmux.d0[27] ),
    .Q(net119),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[28]$_DFF_PP0_  (.D(\dp.ISRmux.d0[28] ),
    .Q(net120),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[29]$_DFF_PP0_  (.D(\dp.ISRmux.d0[29] ),
    .Q(net121),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[2]$_DFF_PP0_  (.D(\dp.ISRmux.d0[2] ),
    .Q(net122),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[30]$_DFF_PP0_  (.D(\dp.ISRmux.d0[30] ),
    .Q(net123),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[31]$_DFF_PP0_  (.D(\dp.ISRmux.d0[31] ),
    .Q(net124),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[3]$_DFF_PP0_  (.D(\dp.ISRmux.d0[3] ),
    .Q(net125),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[4]$_DFF_PP0_  (.D(\dp.ISRmux.d0[4] ),
    .Q(net126),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[5]$_DFF_PP0_  (.D(\dp.ISRmux.d0[5] ),
    .Q(net127),
    .RESET_B(_0031_),
    .CLK(clknet_5_13__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[6]$_DFF_PP0_  (.D(\dp.ISRmux.d0[6] ),
    .Q(net128),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[7]$_DFF_PP0_  (.D(\dp.ISRmux.d0[7] ),
    .Q(net129),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[8]$_DFF_PP0_  (.D(\dp.ISRmux.d0[8] ),
    .Q(net130),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__dfrtp_4 \dp.pcreg.q[9]$_DFF_PP0_  (.D(\dp.ISRmux.d0[9] ),
    .Q(net131),
    .RESET_B(_0031_),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(net165),
    .Q(\dp.rf.rf[0][0] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net166),
    .Q(\dp.rf.rf[0][10] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(net167),
    .Q(\dp.rf.rf[0][11] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(net168),
    .Q(\dp.rf.rf[0][12] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net169),
    .Q(\dp.rf.rf[0][13] ),
    .CLK(clknet_leaf_300_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(net170),
    .Q(\dp.rf.rf[0][14] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net171),
    .Q(\dp.rf.rf[0][15] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][17]$_DFFE_PP_  (.D(net700),
    .DE(net172),
    .Q(\dp.rf.rf[0][17] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net173),
    .Q(\dp.rf.rf[0][18] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][19]$_DFFE_PP_  (.D(net699),
    .DE(net174),
    .Q(\dp.rf.rf[0][19] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(net175),
    .Q(\dp.rf.rf[0][1] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net176),
    .Q(\dp.rf.rf[0][21] ),
    .CLK(clknet_5_17__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net177),
    .Q(\dp.rf.rf[0][22] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net178),
    .Q(\dp.rf.rf[0][23] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net179),
    .Q(\dp.rf.rf[0][24] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net180),
    .Q(\dp.rf.rf[0][25] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][27]$_DFFE_PP_  (.D(net697),
    .DE(net181),
    .Q(\dp.rf.rf[0][27] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net182),
    .Q(\dp.rf.rf[0][28] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][29]$_DFFE_PP_  (.D(net696),
    .DE(net183),
    .Q(\dp.rf.rf[0][29] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][30]$_DFFE_PP_  (.D(net695),
    .DE(net184),
    .Q(\dp.rf.rf[0][30] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][31]$_DFFE_PP_  (.D(net694),
    .DE(net185),
    .Q(\dp.rf.rf[0][31] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net186),
    .Q(\dp.rf.rf[0][3] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(net187),
    .Q(\dp.rf.rf[0][4] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(net188),
    .Q(\dp.rf.rf[0][5] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(net189),
    .Q(\dp.rf.rf[0][6] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(net190),
    .Q(\dp.rf.rf[0][7] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net191),
    .Q(\dp.rf.rf[0][8] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[0][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net192),
    .Q(\dp.rf.rf[0][9] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][0] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net733),
    .Q(\dp.rf.rf[10][10] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][11] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][12] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net733),
    .Q(\dp.rf.rf[10][13] ),
    .CLK(clknet_leaf_299_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(net733),
    .Q(\dp.rf.rf[10][14] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net733),
    .Q(\dp.rf.rf[10][15] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net733),
    .Q(\dp.rf.rf[10][16] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][17]$_DFFE_PP_  (.D(net700),
    .DE(net733),
    .Q(\dp.rf.rf[10][17] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net733),
    .Q(\dp.rf.rf[10][18] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][19]$_DFFE_PP_  (.D(net699),
    .DE(net733),
    .Q(\dp.rf.rf[10][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][1] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net733),
    .Q(\dp.rf.rf[10][20] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net733),
    .Q(\dp.rf.rf[10][21] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net733),
    .Q(\dp.rf.rf[10][22] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net733),
    .Q(\dp.rf.rf[10][23] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net733),
    .Q(\dp.rf.rf[10][24] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net733),
    .Q(\dp.rf.rf[10][25] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][26]$_DFFE_PP_  (.D(net698),
    .DE(net733),
    .Q(\dp.rf.rf[10][26] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][27]$_DFFE_PP_  (.D(net697),
    .DE(net733),
    .Q(\dp.rf.rf[10][27] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net733),
    .Q(\dp.rf.rf[10][28] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][29]$_DFFE_PP_  (.D(net696),
    .DE(net733),
    .Q(\dp.rf.rf[10][29] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][2] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][30]$_DFFE_PP_  (.D(net695),
    .DE(net733),
    .Q(\dp.rf.rf[10][30] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][31]$_DFFE_PP_  (.D(net694),
    .DE(net733),
    .Q(\dp.rf.rf[10][31] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net733),
    .Q(\dp.rf.rf[10][3] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(net733),
    .Q(\dp.rf.rf[10][4] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][5] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0000_),
    .Q(\dp.rf.rf[10][6] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(net733),
    .Q(\dp.rf.rf[10][7] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net733),
    .Q(\dp.rf.rf[10][8] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[10][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net733),
    .Q(\dp.rf.rf[10][9] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][0] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net735),
    .Q(\dp.rf.rf[11][10] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][11] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][12] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net735),
    .Q(\dp.rf.rf[11][13] ),
    .CLK(clknet_leaf_299_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(net735),
    .Q(\dp.rf.rf[11][14] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net735),
    .Q(\dp.rf.rf[11][15] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net735),
    .Q(\dp.rf.rf[11][16] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][17]$_DFFE_PP_  (.D(net700),
    .DE(net735),
    .Q(\dp.rf.rf[11][17] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net735),
    .Q(\dp.rf.rf[11][18] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][19]$_DFFE_PP_  (.D(net699),
    .DE(net735),
    .Q(\dp.rf.rf[11][19] ),
    .CLK(clknet_leaf_302_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][1] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net735),
    .Q(\dp.rf.rf[11][20] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net735),
    .Q(\dp.rf.rf[11][21] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net735),
    .Q(\dp.rf.rf[11][22] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net735),
    .Q(\dp.rf.rf[11][23] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net735),
    .Q(\dp.rf.rf[11][24] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net735),
    .Q(\dp.rf.rf[11][25] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][26]$_DFFE_PP_  (.D(net698),
    .DE(net735),
    .Q(\dp.rf.rf[11][26] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][27]$_DFFE_PP_  (.D(net697),
    .DE(net735),
    .Q(\dp.rf.rf[11][27] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net735),
    .Q(\dp.rf.rf[11][28] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][29]$_DFFE_PP_  (.D(net696),
    .DE(net735),
    .Q(\dp.rf.rf[11][29] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][2] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][30]$_DFFE_PP_  (.D(net695),
    .DE(net735),
    .Q(\dp.rf.rf[11][30] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][31]$_DFFE_PP_  (.D(net694),
    .DE(net735),
    .Q(\dp.rf.rf[11][31] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net735),
    .Q(\dp.rf.rf[11][3] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(net735),
    .Q(\dp.rf.rf[11][4] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][5] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0001_),
    .Q(\dp.rf.rf[11][6] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(net735),
    .Q(\dp.rf.rf[11][7] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net735),
    .Q(\dp.rf.rf[11][8] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[11][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net735),
    .Q(\dp.rf.rf[11][9] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][0] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net718),
    .Q(\dp.rf.rf[12][10] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][11] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][12] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net718),
    .Q(\dp.rf.rf[12][13] ),
    .CLK(clknet_leaf_299_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(net718),
    .Q(\dp.rf.rf[12][14] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net718),
    .Q(\dp.rf.rf[12][15] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net718),
    .Q(\dp.rf.rf[12][16] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][17]$_DFFE_PP_  (.D(net700),
    .DE(net718),
    .Q(\dp.rf.rf[12][17] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net718),
    .Q(\dp.rf.rf[12][18] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][19]$_DFFE_PP_  (.D(net699),
    .DE(net718),
    .Q(\dp.rf.rf[12][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][1] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net718),
    .Q(\dp.rf.rf[12][20] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net718),
    .Q(\dp.rf.rf[12][21] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net718),
    .Q(\dp.rf.rf[12][22] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net718),
    .Q(\dp.rf.rf[12][23] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net718),
    .Q(\dp.rf.rf[12][24] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net718),
    .Q(\dp.rf.rf[12][25] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][26]$_DFFE_PP_  (.D(net698),
    .DE(net718),
    .Q(\dp.rf.rf[12][26] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][27]$_DFFE_PP_  (.D(net697),
    .DE(net718),
    .Q(\dp.rf.rf[12][27] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net718),
    .Q(\dp.rf.rf[12][28] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][29]$_DFFE_PP_  (.D(net696),
    .DE(net718),
    .Q(\dp.rf.rf[12][29] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][2] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][30]$_DFFE_PP_  (.D(net695),
    .DE(net718),
    .Q(\dp.rf.rf[12][30] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][31]$_DFFE_PP_  (.D(net694),
    .DE(net718),
    .Q(\dp.rf.rf[12][31] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net718),
    .Q(\dp.rf.rf[12][3] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(net718),
    .Q(\dp.rf.rf[12][4] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][5] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0002_),
    .Q(\dp.rf.rf[12][6] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(net718),
    .Q(\dp.rf.rf[12][7] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net718),
    .Q(\dp.rf.rf[12][8] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[12][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net718),
    .Q(\dp.rf.rf[12][9] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][0] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net720),
    .Q(\dp.rf.rf[13][10] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][11] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][12] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net720),
    .Q(\dp.rf.rf[13][13] ),
    .CLK(clknet_leaf_299_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(net720),
    .Q(\dp.rf.rf[13][14] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net720),
    .Q(\dp.rf.rf[13][15] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net720),
    .Q(\dp.rf.rf[13][16] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][17]$_DFFE_PP_  (.D(net700),
    .DE(net720),
    .Q(\dp.rf.rf[13][17] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net720),
    .Q(\dp.rf.rf[13][18] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][19]$_DFFE_PP_  (.D(net699),
    .DE(net720),
    .Q(\dp.rf.rf[13][19] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][1] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net720),
    .Q(\dp.rf.rf[13][20] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net720),
    .Q(\dp.rf.rf[13][21] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net720),
    .Q(\dp.rf.rf[13][22] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net720),
    .Q(\dp.rf.rf[13][23] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net720),
    .Q(\dp.rf.rf[13][24] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net720),
    .Q(\dp.rf.rf[13][25] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][26]$_DFFE_PP_  (.D(net698),
    .DE(net720),
    .Q(\dp.rf.rf[13][26] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][27]$_DFFE_PP_  (.D(net697),
    .DE(net720),
    .Q(\dp.rf.rf[13][27] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net720),
    .Q(\dp.rf.rf[13][28] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][29]$_DFFE_PP_  (.D(net696),
    .DE(net720),
    .Q(\dp.rf.rf[13][29] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][2] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][30]$_DFFE_PP_  (.D(net695),
    .DE(net720),
    .Q(\dp.rf.rf[13][30] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][31]$_DFFE_PP_  (.D(net694),
    .DE(net720),
    .Q(\dp.rf.rf[13][31] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net720),
    .Q(\dp.rf.rf[13][3] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(net720),
    .Q(\dp.rf.rf[13][4] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][5] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0003_),
    .Q(\dp.rf.rf[13][6] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(net720),
    .Q(\dp.rf.rf[13][7] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net720),
    .Q(\dp.rf.rf[13][8] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[13][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net720),
    .Q(\dp.rf.rf[13][9] ),
    .CLK(clknet_5_18__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][0] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net721),
    .Q(\dp.rf.rf[14][10] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][11] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][12] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net721),
    .Q(\dp.rf.rf[14][13] ),
    .CLK(clknet_leaf_299_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(net721),
    .Q(\dp.rf.rf[14][14] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net721),
    .Q(\dp.rf.rf[14][15] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net721),
    .Q(\dp.rf.rf[14][16] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][17]$_DFFE_PP_  (.D(net700),
    .DE(net721),
    .Q(\dp.rf.rf[14][17] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net721),
    .Q(\dp.rf.rf[14][18] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][19]$_DFFE_PP_  (.D(net699),
    .DE(net721),
    .Q(\dp.rf.rf[14][19] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][1] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net721),
    .Q(\dp.rf.rf[14][20] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net721),
    .Q(\dp.rf.rf[14][21] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net721),
    .Q(\dp.rf.rf[14][22] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net721),
    .Q(\dp.rf.rf[14][23] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net721),
    .Q(\dp.rf.rf[14][24] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net721),
    .Q(\dp.rf.rf[14][25] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][26]$_DFFE_PP_  (.D(net698),
    .DE(net721),
    .Q(\dp.rf.rf[14][26] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][27]$_DFFE_PP_  (.D(net697),
    .DE(net721),
    .Q(\dp.rf.rf[14][27] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net721),
    .Q(\dp.rf.rf[14][28] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][29]$_DFFE_PP_  (.D(net696),
    .DE(net721),
    .Q(\dp.rf.rf[14][29] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][2] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][30]$_DFFE_PP_  (.D(net695),
    .DE(net721),
    .Q(\dp.rf.rf[14][30] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][31]$_DFFE_PP_  (.D(net694),
    .DE(net721),
    .Q(\dp.rf.rf[14][31] ),
    .CLK(clknet_5_19__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net721),
    .Q(\dp.rf.rf[14][3] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(net721),
    .Q(\dp.rf.rf[14][4] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][5] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0004_),
    .Q(\dp.rf.rf[14][6] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(net721),
    .Q(\dp.rf.rf[14][7] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net721),
    .Q(\dp.rf.rf[14][8] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[14][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net721),
    .Q(\dp.rf.rf[14][9] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][0] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net723),
    .Q(\dp.rf.rf[15][10] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][11] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][12] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net723),
    .Q(\dp.rf.rf[15][13] ),
    .CLK(clknet_leaf_299_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(net723),
    .Q(\dp.rf.rf[15][14] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net723),
    .Q(\dp.rf.rf[15][15] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net723),
    .Q(\dp.rf.rf[15][16] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][17]$_DFFE_PP_  (.D(net700),
    .DE(net723),
    .Q(\dp.rf.rf[15][17] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net723),
    .Q(\dp.rf.rf[15][18] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][19]$_DFFE_PP_  (.D(net699),
    .DE(net723),
    .Q(\dp.rf.rf[15][19] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][1] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net723),
    .Q(\dp.rf.rf[15][20] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net723),
    .Q(\dp.rf.rf[15][21] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net723),
    .Q(\dp.rf.rf[15][22] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net723),
    .Q(\dp.rf.rf[15][23] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net723),
    .Q(\dp.rf.rf[15][24] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net723),
    .Q(\dp.rf.rf[15][25] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][26]$_DFFE_PP_  (.D(net698),
    .DE(net723),
    .Q(\dp.rf.rf[15][26] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][27]$_DFFE_PP_  (.D(net697),
    .DE(net723),
    .Q(\dp.rf.rf[15][27] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net723),
    .Q(\dp.rf.rf[15][28] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][29]$_DFFE_PP_  (.D(net696),
    .DE(net723),
    .Q(\dp.rf.rf[15][29] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][2] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][30]$_DFFE_PP_  (.D(net695),
    .DE(net723),
    .Q(\dp.rf.rf[15][30] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][31]$_DFFE_PP_  (.D(net694),
    .DE(net723),
    .Q(\dp.rf.rf[15][31] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net723),
    .Q(\dp.rf.rf[15][3] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(net723),
    .Q(\dp.rf.rf[15][4] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][5] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0005_),
    .Q(\dp.rf.rf[15][6] ),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(net723),
    .Q(\dp.rf.rf[15][7] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net723),
    .Q(\dp.rf.rf[15][8] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[15][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net723),
    .Q(\dp.rf.rf[15][9] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][0] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net726),
    .Q(\dp.rf.rf[16][10] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][11] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][12] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net726),
    .Q(\dp.rf.rf[16][13] ),
    .CLK(clknet_leaf_295_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(net726),
    .Q(\dp.rf.rf[16][14] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net726),
    .Q(\dp.rf.rf[16][15] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net726),
    .Q(\dp.rf.rf[16][16] ),
    .CLK(clknet_5_25__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][17]$_DFFE_PP_  (.D(net700),
    .DE(net726),
    .Q(\dp.rf.rf[16][17] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net726),
    .Q(\dp.rf.rf[16][18] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][19]$_DFFE_PP_  (.D(net699),
    .DE(net726),
    .Q(\dp.rf.rf[16][19] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][1] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net726),
    .Q(\dp.rf.rf[16][20] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net726),
    .Q(\dp.rf.rf[16][21] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net726),
    .Q(\dp.rf.rf[16][22] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net726),
    .Q(\dp.rf.rf[16][23] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net726),
    .Q(\dp.rf.rf[16][24] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net726),
    .Q(\dp.rf.rf[16][25] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][26]$_DFFE_PP_  (.D(net698),
    .DE(net726),
    .Q(\dp.rf.rf[16][26] ),
    .CLK(clknet_5_29__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][27]$_DFFE_PP_  (.D(net697),
    .DE(net726),
    .Q(\dp.rf.rf[16][27] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net726),
    .Q(\dp.rf.rf[16][28] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][29]$_DFFE_PP_  (.D(net696),
    .DE(net726),
    .Q(\dp.rf.rf[16][29] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][2] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][30]$_DFFE_PP_  (.D(net695),
    .DE(net726),
    .Q(\dp.rf.rf[16][30] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][31]$_DFFE_PP_  (.D(net694),
    .DE(net726),
    .Q(\dp.rf.rf[16][31] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net726),
    .Q(\dp.rf.rf[16][3] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][4] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][5] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0006_),
    .Q(\dp.rf.rf[16][6] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(net726),
    .Q(\dp.rf.rf[16][7] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net726),
    .Q(\dp.rf.rf[16][8] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[16][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net726),
    .Q(\dp.rf.rf[16][9] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][0] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][10] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][11] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][12] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][13] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][14] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][15] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net728),
    .Q(\dp.rf.rf[17][16] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][17]$_DFFE_PP_  (.D(net700),
    .DE(net728),
    .Q(\dp.rf.rf[17][17] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net728),
    .Q(\dp.rf.rf[17][18] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][19]$_DFFE_PP_  (.D(net699),
    .DE(net728),
    .Q(\dp.rf.rf[17][19] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][1] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net728),
    .Q(\dp.rf.rf[17][20] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net728),
    .Q(\dp.rf.rf[17][21] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net728),
    .Q(\dp.rf.rf[17][22] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net728),
    .Q(\dp.rf.rf[17][23] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net728),
    .Q(\dp.rf.rf[17][24] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net728),
    .Q(\dp.rf.rf[17][25] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][26]$_DFFE_PP_  (.D(net698),
    .DE(net728),
    .Q(\dp.rf.rf[17][26] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][27]$_DFFE_PP_  (.D(net697),
    .DE(net728),
    .Q(\dp.rf.rf[17][27] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net728),
    .Q(\dp.rf.rf[17][28] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][29]$_DFFE_PP_  (.D(net696),
    .DE(net728),
    .Q(\dp.rf.rf[17][29] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][2] ),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][30]$_DFFE_PP_  (.D(net695),
    .DE(net728),
    .Q(\dp.rf.rf[17][30] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][31]$_DFFE_PP_  (.D(net694),
    .DE(net728),
    .Q(\dp.rf.rf[17][31] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][3] ),
    .CLK(clknet_5_13__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][4] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][5] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][6] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][7] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net728),
    .Q(\dp.rf.rf[17][8] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[17][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0007_),
    .Q(\dp.rf.rf[17][9] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][0] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net729),
    .Q(\dp.rf.rf[18][10] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][12] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net729),
    .Q(\dp.rf.rf[18][13] ),
    .CLK(clknet_leaf_295_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(net729),
    .Q(\dp.rf.rf[18][14] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net729),
    .Q(\dp.rf.rf[18][15] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net729),
    .Q(\dp.rf.rf[18][16] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][17]$_DFFE_PP_  (.D(net700),
    .DE(net729),
    .Q(\dp.rf.rf[18][17] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net729),
    .Q(\dp.rf.rf[18][18] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][19]$_DFFE_PP_  (.D(net699),
    .DE(net729),
    .Q(\dp.rf.rf[18][19] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][1] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net729),
    .Q(\dp.rf.rf[18][20] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net729),
    .Q(\dp.rf.rf[18][21] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net729),
    .Q(\dp.rf.rf[18][22] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net729),
    .Q(\dp.rf.rf[18][23] ),
    .CLK(clknet_5_23__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net729),
    .Q(\dp.rf.rf[18][24] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net729),
    .Q(\dp.rf.rf[18][25] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][26]$_DFFE_PP_  (.D(net698),
    .DE(net729),
    .Q(\dp.rf.rf[18][26] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][27]$_DFFE_PP_  (.D(net697),
    .DE(net729),
    .Q(\dp.rf.rf[18][27] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net729),
    .Q(\dp.rf.rf[18][28] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][29]$_DFFE_PP_  (.D(net696),
    .DE(net729),
    .Q(\dp.rf.rf[18][29] ),
    .CLK(clknet_5_16__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][2] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][30]$_DFFE_PP_  (.D(net695),
    .DE(net729),
    .Q(\dp.rf.rf[18][30] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][31]$_DFFE_PP_  (.D(net694),
    .DE(net729),
    .Q(\dp.rf.rf[18][31] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net729),
    .Q(\dp.rf.rf[18][3] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][4] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][5] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0008_),
    .Q(\dp.rf.rf[18][6] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(net729),
    .Q(\dp.rf.rf[18][7] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net729),
    .Q(\dp.rf.rf[18][8] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[18][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net729),
    .Q(\dp.rf.rf[18][9] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][0] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net731),
    .Q(\dp.rf.rf[19][10] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][11] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][12] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net731),
    .Q(\dp.rf.rf[19][13] ),
    .CLK(clknet_leaf_295_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(net731),
    .Q(\dp.rf.rf[19][14] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net731),
    .Q(\dp.rf.rf[19][15] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net731),
    .Q(\dp.rf.rf[19][16] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][17]$_DFFE_PP_  (.D(net700),
    .DE(net731),
    .Q(\dp.rf.rf[19][17] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net731),
    .Q(\dp.rf.rf[19][18] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][19]$_DFFE_PP_  (.D(net699),
    .DE(net731),
    .Q(\dp.rf.rf[19][19] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][1] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net731),
    .Q(\dp.rf.rf[19][20] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net731),
    .Q(\dp.rf.rf[19][21] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net731),
    .Q(\dp.rf.rf[19][22] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net731),
    .Q(\dp.rf.rf[19][23] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net731),
    .Q(\dp.rf.rf[19][24] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net731),
    .Q(\dp.rf.rf[19][25] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][26]$_DFFE_PP_  (.D(net698),
    .DE(net731),
    .Q(\dp.rf.rf[19][26] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][27]$_DFFE_PP_  (.D(net697),
    .DE(net731),
    .Q(\dp.rf.rf[19][27] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net731),
    .Q(\dp.rf.rf[19][28] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][29]$_DFFE_PP_  (.D(net696),
    .DE(net731),
    .Q(\dp.rf.rf[19][29] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][2] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][30]$_DFFE_PP_  (.D(net695),
    .DE(net731),
    .Q(\dp.rf.rf[19][30] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][31]$_DFFE_PP_  (.D(net694),
    .DE(net731),
    .Q(\dp.rf.rf[19][31] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net731),
    .Q(\dp.rf.rf[19][3] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][4] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][5] ),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0009_),
    .Q(\dp.rf.rf[19][6] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(net731),
    .Q(\dp.rf.rf[19][7] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net731),
    .Q(\dp.rf.rf[19][8] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[19][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net731),
    .Q(\dp.rf.rf[19][9] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][0] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net717),
    .Q(\dp.rf.rf[1][10] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][11] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][12] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net717),
    .Q(\dp.rf.rf[1][13] ),
    .CLK(clknet_leaf_301_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(net717),
    .Q(\dp.rf.rf[1][14] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net717),
    .Q(\dp.rf.rf[1][15] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net717),
    .Q(\dp.rf.rf[1][16] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][17]$_DFFE_PP_  (.D(net700),
    .DE(net717),
    .Q(\dp.rf.rf[1][17] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net717),
    .Q(\dp.rf.rf[1][18] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][19]$_DFFE_PP_  (.D(net699),
    .DE(net717),
    .Q(\dp.rf.rf[1][19] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][1] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net717),
    .Q(\dp.rf.rf[1][20] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net717),
    .Q(\dp.rf.rf[1][21] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net717),
    .Q(\dp.rf.rf[1][22] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net717),
    .Q(\dp.rf.rf[1][23] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net717),
    .Q(\dp.rf.rf[1][24] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net717),
    .Q(\dp.rf.rf[1][25] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][26]$_DFFE_PP_  (.D(net698),
    .DE(net717),
    .Q(\dp.rf.rf[1][26] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][27]$_DFFE_PP_  (.D(net697),
    .DE(net717),
    .Q(\dp.rf.rf[1][27] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net717),
    .Q(\dp.rf.rf[1][28] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][29]$_DFFE_PP_  (.D(net696),
    .DE(net717),
    .Q(\dp.rf.rf[1][29] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][2] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][30]$_DFFE_PP_  (.D(net695),
    .DE(net717),
    .Q(\dp.rf.rf[1][30] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][31]$_DFFE_PP_  (.D(net694),
    .DE(net717),
    .Q(\dp.rf.rf[1][31] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net717),
    .Q(\dp.rf.rf[1][3] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][4] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][5] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0010_),
    .Q(\dp.rf.rf[1][6] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(net717),
    .Q(\dp.rf.rf[1][7] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net717),
    .Q(\dp.rf.rf[1][8] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[1][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net717),
    .Q(\dp.rf.rf[1][9] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][0] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net734),
    .Q(\dp.rf.rf[20][10] ),
    .CLK(clknet_leaf_291_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][11] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][12] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net734),
    .Q(\dp.rf.rf[20][13] ),
    .CLK(clknet_leaf_295_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(net734),
    .Q(\dp.rf.rf[20][14] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net734),
    .Q(\dp.rf.rf[20][15] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net734),
    .Q(\dp.rf.rf[20][16] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][17]$_DFFE_PP_  (.D(net700),
    .DE(net734),
    .Q(\dp.rf.rf[20][17] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net734),
    .Q(\dp.rf.rf[20][18] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][19]$_DFFE_PP_  (.D(net699),
    .DE(net734),
    .Q(\dp.rf.rf[20][19] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][1] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net734),
    .Q(\dp.rf.rf[20][20] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net734),
    .Q(\dp.rf.rf[20][21] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net734),
    .Q(\dp.rf.rf[20][22] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net734),
    .Q(\dp.rf.rf[20][23] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net734),
    .Q(\dp.rf.rf[20][24] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net734),
    .Q(\dp.rf.rf[20][25] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][26]$_DFFE_PP_  (.D(net698),
    .DE(net734),
    .Q(\dp.rf.rf[20][26] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][27]$_DFFE_PP_  (.D(net697),
    .DE(net734),
    .Q(\dp.rf.rf[20][27] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net734),
    .Q(\dp.rf.rf[20][28] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][29]$_DFFE_PP_  (.D(net696),
    .DE(net734),
    .Q(\dp.rf.rf[20][29] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][2] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][30]$_DFFE_PP_  (.D(net695),
    .DE(net734),
    .Q(\dp.rf.rf[20][30] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][31]$_DFFE_PP_  (.D(net694),
    .DE(net734),
    .Q(\dp.rf.rf[20][31] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net734),
    .Q(\dp.rf.rf[20][3] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(net734),
    .Q(\dp.rf.rf[20][4] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][5] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0011_),
    .Q(\dp.rf.rf[20][6] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(net734),
    .Q(\dp.rf.rf[20][7] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net734),
    .Q(\dp.rf.rf[20][8] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[20][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net734),
    .Q(\dp.rf.rf[20][9] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][0] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net706),
    .Q(\dp.rf.rf[21][10] ),
    .CLK(clknet_leaf_291_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][11] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][12] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net706),
    .Q(\dp.rf.rf[21][13] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(net706),
    .Q(\dp.rf.rf[21][14] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net706),
    .Q(\dp.rf.rf[21][15] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net706),
    .Q(\dp.rf.rf[21][16] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][17]$_DFFE_PP_  (.D(net700),
    .DE(net706),
    .Q(\dp.rf.rf[21][17] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net706),
    .Q(\dp.rf.rf[21][18] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][19]$_DFFE_PP_  (.D(net699),
    .DE(net706),
    .Q(\dp.rf.rf[21][19] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][1] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net706),
    .Q(\dp.rf.rf[21][20] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net706),
    .Q(\dp.rf.rf[21][21] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net706),
    .Q(\dp.rf.rf[21][22] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net706),
    .Q(\dp.rf.rf[21][23] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net706),
    .Q(\dp.rf.rf[21][24] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net706),
    .Q(\dp.rf.rf[21][25] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][26]$_DFFE_PP_  (.D(net698),
    .DE(net706),
    .Q(\dp.rf.rf[21][26] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][27]$_DFFE_PP_  (.D(net697),
    .DE(net706),
    .Q(\dp.rf.rf[21][27] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net706),
    .Q(\dp.rf.rf[21][28] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][29]$_DFFE_PP_  (.D(net696),
    .DE(net706),
    .Q(\dp.rf.rf[21][29] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][2] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][30]$_DFFE_PP_  (.D(net695),
    .DE(net706),
    .Q(\dp.rf.rf[21][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][31]$_DFFE_PP_  (.D(net694),
    .DE(net706),
    .Q(\dp.rf.rf[21][31] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net706),
    .Q(\dp.rf.rf[21][3] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(net706),
    .Q(\dp.rf.rf[21][4] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][5] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0012_),
    .Q(\dp.rf.rf[21][6] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(net706),
    .Q(\dp.rf.rf[21][7] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net706),
    .Q(\dp.rf.rf[21][8] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[21][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net706),
    .Q(\dp.rf.rf[21][9] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][0] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][10] ),
    .CLK(clknet_leaf_292_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][12] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][13] ),
    .CLK(clknet_leaf_295_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][14] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net705),
    .Q(\dp.rf.rf[22][15] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net705),
    .Q(\dp.rf.rf[22][16] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][17]$_DFFE_PP_  (.D(net700),
    .DE(net705),
    .Q(\dp.rf.rf[22][17] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net705),
    .Q(\dp.rf.rf[22][18] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][19]$_DFFE_PP_  (.D(net699),
    .DE(net705),
    .Q(\dp.rf.rf[22][19] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][1] ),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net705),
    .Q(\dp.rf.rf[22][20] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net705),
    .Q(\dp.rf.rf[22][21] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net705),
    .Q(\dp.rf.rf[22][22] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net705),
    .Q(\dp.rf.rf[22][23] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net705),
    .Q(\dp.rf.rf[22][24] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net705),
    .Q(\dp.rf.rf[22][25] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][26]$_DFFE_PP_  (.D(net698),
    .DE(net705),
    .Q(\dp.rf.rf[22][26] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][27]$_DFFE_PP_  (.D(net697),
    .DE(net705),
    .Q(\dp.rf.rf[22][27] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net705),
    .Q(\dp.rf.rf[22][28] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][29]$_DFFE_PP_  (.D(net696),
    .DE(net705),
    .Q(\dp.rf.rf[22][29] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][2] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][30]$_DFFE_PP_  (.D(net695),
    .DE(net705),
    .Q(\dp.rf.rf[22][30] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][31]$_DFFE_PP_  (.D(net694),
    .DE(net705),
    .Q(\dp.rf.rf[22][31] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net705),
    .Q(\dp.rf.rf[22][3] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][4] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][5] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][6] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(_0013_),
    .Q(\dp.rf.rf[22][7] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net705),
    .Q(\dp.rf.rf[22][8] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[22][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net705),
    .Q(\dp.rf.rf[22][9] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][0] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][10] ),
    .CLK(clknet_leaf_291_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][12] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][13] ),
    .CLK(clknet_leaf_294_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][14] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net707),
    .Q(\dp.rf.rf[23][15] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net707),
    .Q(\dp.rf.rf[23][16] ),
    .CLK(clknet_5_25__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][17]$_DFFE_PP_  (.D(net700),
    .DE(net707),
    .Q(\dp.rf.rf[23][17] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net707),
    .Q(\dp.rf.rf[23][18] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][19]$_DFFE_PP_  (.D(net699),
    .DE(net707),
    .Q(\dp.rf.rf[23][19] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][1] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net707),
    .Q(\dp.rf.rf[23][20] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net707),
    .Q(\dp.rf.rf[23][21] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net707),
    .Q(\dp.rf.rf[23][22] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net707),
    .Q(\dp.rf.rf[23][23] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net707),
    .Q(\dp.rf.rf[23][24] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net707),
    .Q(\dp.rf.rf[23][25] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][26]$_DFFE_PP_  (.D(net698),
    .DE(net707),
    .Q(\dp.rf.rf[23][26] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][27]$_DFFE_PP_  (.D(net697),
    .DE(net707),
    .Q(\dp.rf.rf[23][27] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net707),
    .Q(\dp.rf.rf[23][28] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][29]$_DFFE_PP_  (.D(net696),
    .DE(net707),
    .Q(\dp.rf.rf[23][29] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][2] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][30]$_DFFE_PP_  (.D(net695),
    .DE(net707),
    .Q(\dp.rf.rf[23][30] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][31]$_DFFE_PP_  (.D(net694),
    .DE(net707),
    .Q(\dp.rf.rf[23][31] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net707),
    .Q(\dp.rf.rf[23][3] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][4] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][5] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][6] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(_0014_),
    .Q(\dp.rf.rf[23][7] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net707),
    .Q(\dp.rf.rf[23][8] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[23][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net707),
    .Q(\dp.rf.rf[23][9] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][0] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][10] ),
    .CLK(clknet_leaf_294_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(net708),
    .Q(\dp.rf.rf[24][11] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(net708),
    .Q(\dp.rf.rf[24][12] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][13] ),
    .CLK(clknet_leaf_297_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][14] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][15] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net709),
    .Q(\dp.rf.rf[24][16] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][17]$_DFFE_PP_  (.D(net700),
    .DE(net709),
    .Q(\dp.rf.rf[24][17] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net709),
    .Q(\dp.rf.rf[24][18] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][19]$_DFFE_PP_  (.D(net699),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][19] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(net708),
    .Q(\dp.rf.rf[24][1] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net709),
    .Q(\dp.rf.rf[24][20] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net709),
    .Q(\dp.rf.rf[24][21] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net709),
    .Q(\dp.rf.rf[24][22] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net709),
    .Q(\dp.rf.rf[24][23] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net709),
    .Q(\dp.rf.rf[24][24] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net709),
    .Q(\dp.rf.rf[24][25] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][26]$_DFFE_PP_  (.D(net698),
    .DE(net709),
    .Q(\dp.rf.rf[24][26] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][27]$_DFFE_PP_  (.D(net697),
    .DE(net709),
    .Q(\dp.rf.rf[24][27] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net709),
    .Q(\dp.rf.rf[24][28] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][29]$_DFFE_PP_  (.D(net696),
    .DE(net709),
    .Q(\dp.rf.rf[24][29] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(net708),
    .Q(\dp.rf.rf[24][2] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][30]$_DFFE_PP_  (.D(net695),
    .DE(net709),
    .Q(\dp.rf.rf[24][30] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][31]$_DFFE_PP_  (.D(net694),
    .DE(net709),
    .Q(\dp.rf.rf[24][31] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][3] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][4] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(net708),
    .Q(\dp.rf.rf[24][5] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(net708),
    .Q(\dp.rf.rf[24][6] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][7] ),
    .CLK(clknet_leaf_290_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0015_),
    .Q(\dp.rf.rf[24][8] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[24][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net709),
    .Q(\dp.rf.rf[24][9] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][0] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net713),
    .Q(\dp.rf.rf[25][10] ),
    .CLK(clknet_leaf_291_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(net713),
    .Q(\dp.rf.rf[25][11] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(net713),
    .Q(\dp.rf.rf[25][12] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net713),
    .Q(\dp.rf.rf[25][13] ),
    .CLK(clknet_leaf_297_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(net713),
    .Q(\dp.rf.rf[25][14] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net713),
    .Q(\dp.rf.rf[25][15] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][16] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][17]$_DFFE_PP_  (.D(net700),
    .DE(net713),
    .Q(\dp.rf.rf[25][17] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net713),
    .Q(\dp.rf.rf[25][18] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][19]$_DFFE_PP_  (.D(net699),
    .DE(net713),
    .Q(\dp.rf.rf[25][19] ),
    .CLK(clknet_leaf_302_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(net713),
    .Q(\dp.rf.rf[25][1] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][20] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][21] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net713),
    .Q(\dp.rf.rf[25][22] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net713),
    .Q(\dp.rf.rf[25][23] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][24] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][25] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][26]$_DFFE_PP_  (.D(net698),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][26] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][27]$_DFFE_PP_  (.D(net697),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][27] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net713),
    .Q(\dp.rf.rf[25][28] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][29]$_DFFE_PP_  (.D(net696),
    .DE(net713),
    .Q(\dp.rf.rf[25][29] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(net713),
    .Q(\dp.rf.rf[25][2] ),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][30]$_DFFE_PP_  (.D(net695),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][30] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][31]$_DFFE_PP_  (.D(net694),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][31] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][3] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(net713),
    .Q(\dp.rf.rf[25][4] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(net713),
    .Q(\dp.rf.rf[25][5] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(net713),
    .Q(\dp.rf.rf[25][6] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(net713),
    .Q(\dp.rf.rf[25][7] ),
    .CLK(clknet_leaf_290_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net713),
    .Q(\dp.rf.rf[25][8] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[25][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(_0016_),
    .Q(\dp.rf.rf[25][9] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(net711),
    .Q(\dp.rf.rf[26][0] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][10] ),
    .CLK(clknet_leaf_293_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][11] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][12] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][13] ),
    .CLK(clknet_leaf_297_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][14] ),
    .CLK(clknet_leaf_289_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][15] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net711),
    .Q(\dp.rf.rf[26][16] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][17]$_DFFE_PP_  (.D(net700),
    .DE(net711),
    .Q(\dp.rf.rf[26][17] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net711),
    .Q(\dp.rf.rf[26][18] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][19]$_DFFE_PP_  (.D(net699),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][19] ),
    .CLK(clknet_leaf_301_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(net711),
    .Q(\dp.rf.rf[26][1] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net711),
    .Q(\dp.rf.rf[26][20] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net711),
    .Q(\dp.rf.rf[26][21] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net711),
    .Q(\dp.rf.rf[26][22] ),
    .CLK(clknet_5_17__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net711),
    .Q(\dp.rf.rf[26][23] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net711),
    .Q(\dp.rf.rf[26][24] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net711),
    .Q(\dp.rf.rf[26][25] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][26]$_DFFE_PP_  (.D(net698),
    .DE(net711),
    .Q(\dp.rf.rf[26][26] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][27]$_DFFE_PP_  (.D(net697),
    .DE(net711),
    .Q(\dp.rf.rf[26][27] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net711),
    .Q(\dp.rf.rf[26][28] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][29]$_DFFE_PP_  (.D(net696),
    .DE(net711),
    .Q(\dp.rf.rf[26][29] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(net711),
    .Q(\dp.rf.rf[26][2] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][30]$_DFFE_PP_  (.D(net695),
    .DE(net711),
    .Q(\dp.rf.rf[26][30] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][31]$_DFFE_PP_  (.D(net694),
    .DE(net711),
    .Q(\dp.rf.rf[26][31] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net711),
    .Q(\dp.rf.rf[26][3] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][4] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(net711),
    .Q(\dp.rf.rf[26][5] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][6] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][7] ),
    .CLK(clknet_leaf_290_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(_0017_),
    .Q(\dp.rf.rf[26][8] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[26][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net711),
    .Q(\dp.rf.rf[26][9] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(net710),
    .Q(\dp.rf.rf[27][0] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][10] ),
    .CLK(clknet_leaf_293_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][12] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][13] ),
    .CLK(clknet_leaf_297_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][14] ),
    .CLK(clknet_leaf_289_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][15] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net710),
    .Q(\dp.rf.rf[27][16] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][17]$_DFFE_PP_  (.D(net700),
    .DE(net710),
    .Q(\dp.rf.rf[27][17] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net710),
    .Q(\dp.rf.rf[27][18] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][19]$_DFFE_PP_  (.D(net699),
    .DE(net710),
    .Q(\dp.rf.rf[27][19] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(net710),
    .Q(\dp.rf.rf[27][1] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net710),
    .Q(\dp.rf.rf[27][20] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net710),
    .Q(\dp.rf.rf[27][21] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net710),
    .Q(\dp.rf.rf[27][22] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net710),
    .Q(\dp.rf.rf[27][23] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net710),
    .Q(\dp.rf.rf[27][24] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net710),
    .Q(\dp.rf.rf[27][25] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][26]$_DFFE_PP_  (.D(net698),
    .DE(net710),
    .Q(\dp.rf.rf[27][26] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][27]$_DFFE_PP_  (.D(net697),
    .DE(net710),
    .Q(\dp.rf.rf[27][27] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net710),
    .Q(\dp.rf.rf[27][28] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][29]$_DFFE_PP_  (.D(net696),
    .DE(net710),
    .Q(\dp.rf.rf[27][29] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(net710),
    .Q(\dp.rf.rf[27][2] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][30]$_DFFE_PP_  (.D(net695),
    .DE(net710),
    .Q(\dp.rf.rf[27][30] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][31]$_DFFE_PP_  (.D(net694),
    .DE(net710),
    .Q(\dp.rf.rf[27][31] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net710),
    .Q(\dp.rf.rf[27][3] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][4] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(net710),
    .Q(\dp.rf.rf[27][5] ),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][6] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(_0018_),
    .Q(\dp.rf.rf[27][7] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net710),
    .Q(\dp.rf.rf[27][8] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[27][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net710),
    .Q(\dp.rf.rf[27][9] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][0] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][10] ),
    .CLK(clknet_leaf_292_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][11] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][12] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][13] ),
    .CLK(clknet_leaf_296_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][14] ),
    .CLK(clknet_leaf_289_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][15] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net712),
    .Q(\dp.rf.rf[28][16] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][17]$_DFFE_PP_  (.D(net700),
    .DE(net712),
    .Q(\dp.rf.rf[28][17] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net712),
    .Q(\dp.rf.rf[28][18] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][19]$_DFFE_PP_  (.D(net699),
    .DE(net712),
    .Q(\dp.rf.rf[28][19] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][1] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net712),
    .Q(\dp.rf.rf[28][20] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net712),
    .Q(\dp.rf.rf[28][21] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net712),
    .Q(\dp.rf.rf[28][22] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net712),
    .Q(\dp.rf.rf[28][23] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net712),
    .Q(\dp.rf.rf[28][24] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net712),
    .Q(\dp.rf.rf[28][25] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][26]$_DFFE_PP_  (.D(net698),
    .DE(net712),
    .Q(\dp.rf.rf[28][26] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][27]$_DFFE_PP_  (.D(net697),
    .DE(net712),
    .Q(\dp.rf.rf[28][27] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net712),
    .Q(\dp.rf.rf[28][28] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][29]$_DFFE_PP_  (.D(net696),
    .DE(net712),
    .Q(\dp.rf.rf[28][29] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][2] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][30]$_DFFE_PP_  (.D(net695),
    .DE(net712),
    .Q(\dp.rf.rf[28][30] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][31]$_DFFE_PP_  (.D(net694),
    .DE(net712),
    .Q(\dp.rf.rf[28][31] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net712),
    .Q(\dp.rf.rf[28][3] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][4] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][5] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][6] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(_0019_),
    .Q(\dp.rf.rf[28][7] ),
    .CLK(clknet_leaf_290_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net712),
    .Q(\dp.rf.rf[28][8] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[28][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net712),
    .Q(\dp.rf.rf[28][9] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(net714),
    .Q(\dp.rf.rf[29][0] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net714),
    .Q(\dp.rf.rf[29][10] ),
    .CLK(clknet_leaf_294_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][11] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][12] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net714),
    .Q(\dp.rf.rf[29][13] ),
    .CLK(clknet_leaf_298_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][14] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][15] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net714),
    .Q(\dp.rf.rf[29][16] ),
    .CLK(clknet_5_27__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][17]$_DFFE_PP_  (.D(net700),
    .DE(net714),
    .Q(\dp.rf.rf[29][17] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net714),
    .Q(\dp.rf.rf[29][18] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][19]$_DFFE_PP_  (.D(net699),
    .DE(net714),
    .Q(\dp.rf.rf[29][19] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(net714),
    .Q(\dp.rf.rf[29][1] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net714),
    .Q(\dp.rf.rf[29][20] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net714),
    .Q(\dp.rf.rf[29][21] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net714),
    .Q(\dp.rf.rf[29][22] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net714),
    .Q(\dp.rf.rf[29][23] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net714),
    .Q(\dp.rf.rf[29][24] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net714),
    .Q(\dp.rf.rf[29][25] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][26]$_DFFE_PP_  (.D(net698),
    .DE(net714),
    .Q(\dp.rf.rf[29][26] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][27]$_DFFE_PP_  (.D(net697),
    .DE(net714),
    .Q(\dp.rf.rf[29][27] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net714),
    .Q(\dp.rf.rf[29][28] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][29]$_DFFE_PP_  (.D(net696),
    .DE(net714),
    .Q(\dp.rf.rf[29][29] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][2] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][30]$_DFFE_PP_  (.D(net695),
    .DE(net714),
    .Q(\dp.rf.rf[29][30] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][31]$_DFFE_PP_  (.D(net694),
    .DE(net714),
    .Q(\dp.rf.rf[29][31] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net714),
    .Q(\dp.rf.rf[29][3] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][4] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][5] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][6] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(_0020_),
    .Q(\dp.rf.rf[29][7] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net714),
    .Q(\dp.rf.rf[29][8] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[29][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net714),
    .Q(\dp.rf.rf[29][9] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(net736),
    .Q(\dp.rf.rf[2][0] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net736),
    .Q(\dp.rf.rf[2][10] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][11] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][12] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net736),
    .Q(\dp.rf.rf[2][13] ),
    .CLK(clknet_leaf_301_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][14] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net736),
    .Q(\dp.rf.rf[2][15] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net736),
    .Q(\dp.rf.rf[2][16] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][17]$_DFFE_PP_  (.D(net700),
    .DE(net736),
    .Q(\dp.rf.rf[2][17] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net736),
    .Q(\dp.rf.rf[2][18] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][19]$_DFFE_PP_  (.D(net699),
    .DE(net736),
    .Q(\dp.rf.rf[2][19] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(net736),
    .Q(\dp.rf.rf[2][1] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net736),
    .Q(\dp.rf.rf[2][20] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net736),
    .Q(\dp.rf.rf[2][21] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net736),
    .Q(\dp.rf.rf[2][22] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net736),
    .Q(\dp.rf.rf[2][23] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net736),
    .Q(\dp.rf.rf[2][24] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net736),
    .Q(\dp.rf.rf[2][25] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][26]$_DFFE_PP_  (.D(net698),
    .DE(net736),
    .Q(\dp.rf.rf[2][26] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][27]$_DFFE_PP_  (.D(net697),
    .DE(net736),
    .Q(\dp.rf.rf[2][27] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net736),
    .Q(\dp.rf.rf[2][28] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][29]$_DFFE_PP_  (.D(net696),
    .DE(net736),
    .Q(\dp.rf.rf[2][29] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(net736),
    .Q(\dp.rf.rf[2][2] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][30]$_DFFE_PP_  (.D(net695),
    .DE(net736),
    .Q(\dp.rf.rf[2][30] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][31]$_DFFE_PP_  (.D(net694),
    .DE(net736),
    .Q(\dp.rf.rf[2][31] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net736),
    .Q(\dp.rf.rf[2][3] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][4] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][5] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][6] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(_0021_),
    .Q(\dp.rf.rf[2][7] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net736),
    .Q(\dp.rf.rf[2][8] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[2][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net736),
    .Q(\dp.rf.rf[2][9] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][0] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][10] ),
    .CLK(clknet_leaf_293_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][11] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][12] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][13] ),
    .CLK(clknet_leaf_296_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][14] ),
    .CLK(clknet_leaf_289_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][15] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net715),
    .Q(\dp.rf.rf[30][16] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][17]$_DFFE_PP_  (.D(net700),
    .DE(net715),
    .Q(\dp.rf.rf[30][17] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net715),
    .Q(\dp.rf.rf[30][18] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][19]$_DFFE_PP_  (.D(net699),
    .DE(net715),
    .Q(\dp.rf.rf[30][19] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][1] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net715),
    .Q(\dp.rf.rf[30][20] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net715),
    .Q(\dp.rf.rf[30][21] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net715),
    .Q(\dp.rf.rf[30][22] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net715),
    .Q(\dp.rf.rf[30][23] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net715),
    .Q(\dp.rf.rf[30][24] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net715),
    .Q(\dp.rf.rf[30][25] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][26]$_DFFE_PP_  (.D(net698),
    .DE(net715),
    .Q(\dp.rf.rf[30][26] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][27]$_DFFE_PP_  (.D(net697),
    .DE(net715),
    .Q(\dp.rf.rf[30][27] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net715),
    .Q(\dp.rf.rf[30][28] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][29]$_DFFE_PP_  (.D(net696),
    .DE(net715),
    .Q(\dp.rf.rf[30][29] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][2] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][30]$_DFFE_PP_  (.D(net695),
    .DE(net715),
    .Q(\dp.rf.rf[30][30] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][31]$_DFFE_PP_  (.D(net694),
    .DE(net715),
    .Q(\dp.rf.rf[30][31] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net715),
    .Q(\dp.rf.rf[30][3] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][4] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][5] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][6] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(_0022_),
    .Q(\dp.rf.rf[30][7] ),
    .CLK(clknet_leaf_290_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net715),
    .Q(\dp.rf.rf[30][8] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[30][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net715),
    .Q(\dp.rf.rf[30][9] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][0] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][10] ),
    .CLK(clknet_leaf_295_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][11] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][12] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][13] ),
    .CLK(clknet_leaf_295_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][14] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][15] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net716),
    .Q(\dp.rf.rf[31][16] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][17]$_DFFE_PP_  (.D(net700),
    .DE(net716),
    .Q(\dp.rf.rf[31][17] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net716),
    .Q(\dp.rf.rf[31][18] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][19]$_DFFE_PP_  (.D(net699),
    .DE(net716),
    .Q(\dp.rf.rf[31][19] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][1] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net716),
    .Q(\dp.rf.rf[31][20] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net716),
    .Q(\dp.rf.rf[31][21] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net716),
    .Q(\dp.rf.rf[31][22] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net716),
    .Q(\dp.rf.rf[31][23] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net716),
    .Q(\dp.rf.rf[31][24] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net716),
    .Q(\dp.rf.rf[31][25] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][26]$_DFFE_PP_  (.D(net698),
    .DE(net716),
    .Q(\dp.rf.rf[31][26] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][27]$_DFFE_PP_  (.D(net697),
    .DE(net716),
    .Q(\dp.rf.rf[31][27] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net716),
    .Q(\dp.rf.rf[31][28] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][29]$_DFFE_PP_  (.D(net696),
    .DE(net716),
    .Q(\dp.rf.rf[31][29] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][2] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][30]$_DFFE_PP_  (.D(net695),
    .DE(net716),
    .Q(\dp.rf.rf[31][30] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][31]$_DFFE_PP_  (.D(net694),
    .DE(net716),
    .Q(\dp.rf.rf[31][31] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net716),
    .Q(\dp.rf.rf[31][3] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][4] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][5] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][6] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(_0023_),
    .Q(\dp.rf.rf[31][7] ),
    .CLK(clknet_leaf_291_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net716),
    .Q(\dp.rf.rf[31][8] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[31][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net716),
    .Q(\dp.rf.rf[31][9] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][0] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][10] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][11] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][12] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][13] ),
    .CLK(clknet_leaf_301_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][14] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][15] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][16] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][17]$_DFFE_PP_  (.D(net700),
    .DE(net719),
    .Q(\dp.rf.rf[3][17] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][18] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][19]$_DFFE_PP_  (.D(net699),
    .DE(net719),
    .Q(\dp.rf.rf[3][19] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][1] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][20] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][21] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][22] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][23] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][24] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][25] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][26]$_DFFE_PP_  (.D(net698),
    .DE(net719),
    .Q(\dp.rf.rf[3][26] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][27]$_DFFE_PP_  (.D(net697),
    .DE(net719),
    .Q(\dp.rf.rf[3][27] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][28] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][29]$_DFFE_PP_  (.D(net696),
    .DE(net719),
    .Q(\dp.rf.rf[3][29] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][2] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][30]$_DFFE_PP_  (.D(net695),
    .DE(net719),
    .Q(\dp.rf.rf[3][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][31]$_DFFE_PP_  (.D(net694),
    .DE(net719),
    .Q(\dp.rf.rf[3][31] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][3] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][4] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0024_),
    .Q(\dp.rf.rf[3][5] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][6] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][7] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][8] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[3][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net719),
    .Q(\dp.rf.rf[3][9] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][0] ),
    .CLK(clknet_5_13__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net722),
    .Q(\dp.rf.rf[4][10] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][11] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][12] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net722),
    .Q(\dp.rf.rf[4][13] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(net722),
    .Q(\dp.rf.rf[4][14] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net722),
    .Q(\dp.rf.rf[4][15] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net722),
    .Q(\dp.rf.rf[4][16] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][17]$_DFFE_PP_  (.D(net700),
    .DE(net722),
    .Q(\dp.rf.rf[4][17] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net722),
    .Q(\dp.rf.rf[4][18] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][19]$_DFFE_PP_  (.D(net699),
    .DE(net722),
    .Q(\dp.rf.rf[4][19] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][1] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net722),
    .Q(\dp.rf.rf[4][20] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net722),
    .Q(\dp.rf.rf[4][21] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net722),
    .Q(\dp.rf.rf[4][22] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net722),
    .Q(\dp.rf.rf[4][23] ),
    .CLK(clknet_5_21__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net722),
    .Q(\dp.rf.rf[4][24] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net722),
    .Q(\dp.rf.rf[4][25] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][26]$_DFFE_PP_  (.D(net698),
    .DE(net722),
    .Q(\dp.rf.rf[4][26] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][27]$_DFFE_PP_  (.D(net697),
    .DE(net722),
    .Q(\dp.rf.rf[4][27] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net722),
    .Q(\dp.rf.rf[4][28] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][29]$_DFFE_PP_  (.D(net696),
    .DE(net722),
    .Q(\dp.rf.rf[4][29] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][2] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][30]$_DFFE_PP_  (.D(net695),
    .DE(net722),
    .Q(\dp.rf.rf[4][30] ),
    .CLK(clknet_5_26__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][31]$_DFFE_PP_  (.D(net694),
    .DE(net722),
    .Q(\dp.rf.rf[4][31] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net722),
    .Q(\dp.rf.rf[4][3] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(net722),
    .Q(\dp.rf.rf[4][4] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][5] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0025_),
    .Q(\dp.rf.rf[4][6] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(net722),
    .Q(\dp.rf.rf[4][7] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net722),
    .Q(\dp.rf.rf[4][8] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[4][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net722),
    .Q(\dp.rf.rf[4][9] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][0] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net724),
    .Q(\dp.rf.rf[5][10] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][11] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][12] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net724),
    .Q(\dp.rf.rf[5][13] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][14] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net724),
    .Q(\dp.rf.rf[5][15] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net724),
    .Q(\dp.rf.rf[5][16] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][17]$_DFFE_PP_  (.D(net700),
    .DE(net724),
    .Q(\dp.rf.rf[5][17] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net724),
    .Q(\dp.rf.rf[5][18] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][19]$_DFFE_PP_  (.D(net699),
    .DE(net724),
    .Q(\dp.rf.rf[5][19] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][1] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net724),
    .Q(\dp.rf.rf[5][20] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net724),
    .Q(\dp.rf.rf[5][21] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net724),
    .Q(\dp.rf.rf[5][22] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net724),
    .Q(\dp.rf.rf[5][23] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net724),
    .Q(\dp.rf.rf[5][24] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net724),
    .Q(\dp.rf.rf[5][25] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][26]$_DFFE_PP_  (.D(net698),
    .DE(net724),
    .Q(\dp.rf.rf[5][26] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][27]$_DFFE_PP_  (.D(net697),
    .DE(net724),
    .Q(\dp.rf.rf[5][27] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net724),
    .Q(\dp.rf.rf[5][28] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][29]$_DFFE_PP_  (.D(net696),
    .DE(net724),
    .Q(\dp.rf.rf[5][29] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][2] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][30]$_DFFE_PP_  (.D(net695),
    .DE(net724),
    .Q(\dp.rf.rf[5][30] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][31]$_DFFE_PP_  (.D(net694),
    .DE(net724),
    .Q(\dp.rf.rf[5][31] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net724),
    .Q(\dp.rf.rf[5][3] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][4] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][5] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][6] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(_0026_),
    .Q(\dp.rf.rf[5][7] ),
    .CLK(clknet_5_12__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net724),
    .Q(\dp.rf.rf[5][8] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[5][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net724),
    .Q(\dp.rf.rf[5][9] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][0] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net725),
    .Q(\dp.rf.rf[6][10] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][11] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][12] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net725),
    .Q(\dp.rf.rf[6][13] ),
    .CLK(clknet_leaf_300_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(net725),
    .Q(\dp.rf.rf[6][14] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net725),
    .Q(\dp.rf.rf[6][15] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net725),
    .Q(\dp.rf.rf[6][16] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][17]$_DFFE_PP_  (.D(net700),
    .DE(net725),
    .Q(\dp.rf.rf[6][17] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net725),
    .Q(\dp.rf.rf[6][18] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][19]$_DFFE_PP_  (.D(net699),
    .DE(net725),
    .Q(\dp.rf.rf[6][19] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][1] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net725),
    .Q(\dp.rf.rf[6][20] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net725),
    .Q(\dp.rf.rf[6][21] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net725),
    .Q(\dp.rf.rf[6][22] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net725),
    .Q(\dp.rf.rf[6][23] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net725),
    .Q(\dp.rf.rf[6][24] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net725),
    .Q(\dp.rf.rf[6][25] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][26]$_DFFE_PP_  (.D(net698),
    .DE(net725),
    .Q(\dp.rf.rf[6][26] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][27]$_DFFE_PP_  (.D(net697),
    .DE(net725),
    .Q(\dp.rf.rf[6][27] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net725),
    .Q(\dp.rf.rf[6][28] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][29]$_DFFE_PP_  (.D(net696),
    .DE(net725),
    .Q(\dp.rf.rf[6][29] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][2] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][30]$_DFFE_PP_  (.D(net695),
    .DE(net725),
    .Q(\dp.rf.rf[6][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][31]$_DFFE_PP_  (.D(net694),
    .DE(net725),
    .Q(\dp.rf.rf[6][31] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net725),
    .Q(\dp.rf.rf[6][3] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(net725),
    .Q(\dp.rf.rf[6][4] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][5] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0027_),
    .Q(\dp.rf.rf[6][6] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(net725),
    .Q(\dp.rf.rf[6][7] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net725),
    .Q(\dp.rf.rf[6][8] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[6][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net725),
    .Q(\dp.rf.rf[6][9] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][0] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net727),
    .Q(\dp.rf.rf[7][10] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][11] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][12] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net727),
    .Q(\dp.rf.rf[7][13] ),
    .CLK(clknet_leaf_300_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(net727),
    .Q(\dp.rf.rf[7][14] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net727),
    .Q(\dp.rf.rf[7][15] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net727),
    .Q(\dp.rf.rf[7][16] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][17]$_DFFE_PP_  (.D(net700),
    .DE(net727),
    .Q(\dp.rf.rf[7][17] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net727),
    .Q(\dp.rf.rf[7][18] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][19]$_DFFE_PP_  (.D(net699),
    .DE(net727),
    .Q(\dp.rf.rf[7][19] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][1] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net727),
    .Q(\dp.rf.rf[7][20] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net727),
    .Q(\dp.rf.rf[7][21] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net727),
    .Q(\dp.rf.rf[7][22] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net727),
    .Q(\dp.rf.rf[7][23] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net727),
    .Q(\dp.rf.rf[7][24] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net727),
    .Q(\dp.rf.rf[7][25] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][26]$_DFFE_PP_  (.D(net698),
    .DE(net727),
    .Q(\dp.rf.rf[7][26] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][27]$_DFFE_PP_  (.D(net697),
    .DE(net727),
    .Q(\dp.rf.rf[7][27] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net727),
    .Q(\dp.rf.rf[7][28] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][29]$_DFFE_PP_  (.D(net696),
    .DE(net727),
    .Q(\dp.rf.rf[7][29] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][2] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][30]$_DFFE_PP_  (.D(net695),
    .DE(net727),
    .Q(\dp.rf.rf[7][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][31]$_DFFE_PP_  (.D(net694),
    .DE(net727),
    .Q(\dp.rf.rf[7][31] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net727),
    .Q(\dp.rf.rf[7][3] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(net727),
    .Q(\dp.rf.rf[7][4] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][5] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0028_),
    .Q(\dp.rf.rf[7][6] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(net727),
    .Q(\dp.rf.rf[7][7] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net727),
    .Q(\dp.rf.rf[7][8] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[7][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net727),
    .Q(\dp.rf.rf[7][9] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][0] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net730),
    .Q(\dp.rf.rf[8][10] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][11] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][12] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net730),
    .Q(\dp.rf.rf[8][13] ),
    .CLK(clknet_leaf_300_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][14] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net730),
    .Q(\dp.rf.rf[8][15] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net730),
    .Q(\dp.rf.rf[8][16] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][17]$_DFFE_PP_  (.D(net700),
    .DE(net730),
    .Q(\dp.rf.rf[8][17] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net730),
    .Q(\dp.rf.rf[8][18] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][19]$_DFFE_PP_  (.D(net699),
    .DE(net730),
    .Q(\dp.rf.rf[8][19] ),
    .CLK(clknet_leaf_302_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][1] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net730),
    .Q(\dp.rf.rf[8][20] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net730),
    .Q(\dp.rf.rf[8][21] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net730),
    .Q(\dp.rf.rf[8][22] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net730),
    .Q(\dp.rf.rf[8][23] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net730),
    .Q(\dp.rf.rf[8][24] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net730),
    .Q(\dp.rf.rf[8][25] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][26]$_DFFE_PP_  (.D(net698),
    .DE(net730),
    .Q(\dp.rf.rf[8][26] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][27]$_DFFE_PP_  (.D(net697),
    .DE(net730),
    .Q(\dp.rf.rf[8][27] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net730),
    .Q(\dp.rf.rf[8][28] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][29]$_DFFE_PP_  (.D(net696),
    .DE(net730),
    .Q(\dp.rf.rf[8][29] ),
    .CLK(clknet_5_16__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][2] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][30]$_DFFE_PP_  (.D(net695),
    .DE(net730),
    .Q(\dp.rf.rf[8][30] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][31]$_DFFE_PP_  (.D(net694),
    .DE(net730),
    .Q(\dp.rf.rf[8][31] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net730),
    .Q(\dp.rf.rf[8][3] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][4] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][5] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][6] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(_0029_),
    .Q(\dp.rf.rf[8][7] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net730),
    .Q(\dp.rf.rf[8][8] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[8][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net730),
    .Q(\dp.rf.rf[8][9] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][0]$_DFFE_PP_  (.D(\dp.result2[0] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][0] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][10]$_DFFE_PP_  (.D(\dp.result2[10] ),
    .DE(net732),
    .Q(\dp.rf.rf[9][10] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][11]$_DFFE_PP_  (.D(\dp.result2[11] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][11] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][12]$_DFFE_PP_  (.D(\dp.result2[12] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][12] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][13]$_DFFE_PP_  (.D(\dp.result2[13] ),
    .DE(net732),
    .Q(\dp.rf.rf[9][13] ),
    .CLK(clknet_leaf_298_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][14]$_DFFE_PP_  (.D(\dp.result2[14] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][14] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][15]$_DFFE_PP_  (.D(\dp.result2[15] ),
    .DE(net732),
    .Q(\dp.rf.rf[9][15] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][16]$_DFFE_PP_  (.D(\dp.result2[16] ),
    .DE(net732),
    .Q(\dp.rf.rf[9][16] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][17]$_DFFE_PP_  (.D(net700),
    .DE(net732),
    .Q(\dp.rf.rf[9][17] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][18]$_DFFE_PP_  (.D(\dp.result2[18] ),
    .DE(net732),
    .Q(\dp.rf.rf[9][18] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][19]$_DFFE_PP_  (.D(net699),
    .DE(net732),
    .Q(\dp.rf.rf[9][19] ),
    .CLK(clknet_leaf_302_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][1]$_DFFE_PP_  (.D(\dp.result2[1] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][1] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][20]$_DFFE_PP_  (.D(\dp.result2[20] ),
    .DE(net732),
    .Q(\dp.rf.rf[9][20] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][21]$_DFFE_PP_  (.D(\dp.result2[21] ),
    .DE(net732),
    .Q(\dp.rf.rf[9][21] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][22]$_DFFE_PP_  (.D(\dp.result2[22] ),
    .DE(net732),
    .Q(\dp.rf.rf[9][22] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][23]$_DFFE_PP_  (.D(\dp.result2[23] ),
    .DE(net732),
    .Q(\dp.rf.rf[9][23] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][24]$_DFFE_PP_  (.D(\dp.result2[24] ),
    .DE(net732),
    .Q(\dp.rf.rf[9][24] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][25]$_DFFE_PP_  (.D(\dp.result2[25] ),
    .DE(net732),
    .Q(\dp.rf.rf[9][25] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][26]$_DFFE_PP_  (.D(net698),
    .DE(net732),
    .Q(\dp.rf.rf[9][26] ),
    .CLK(clknet_5_29__leaf_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][27]$_DFFE_PP_  (.D(net697),
    .DE(net732),
    .Q(\dp.rf.rf[9][27] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][28]$_DFFE_PP_  (.D(\dp.result2[28] ),
    .DE(net732),
    .Q(\dp.rf.rf[9][28] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][29]$_DFFE_PP_  (.D(net696),
    .DE(net732),
    .Q(\dp.rf.rf[9][29] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][2]$_DFFE_PP_  (.D(\dp.result2[2] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][2] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][30]$_DFFE_PP_  (.D(net695),
    .DE(net732),
    .Q(\dp.rf.rf[9][30] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][31]$_DFFE_PP_  (.D(net694),
    .DE(net732),
    .Q(\dp.rf.rf[9][31] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][3]$_DFFE_PP_  (.D(\dp.result2[3] ),
    .DE(net732),
    .Q(\dp.rf.rf[9][3] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][4]$_DFFE_PP_  (.D(\dp.result2[4] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][4] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][5]$_DFFE_PP_  (.D(\dp.result2[5] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][5] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][6]$_DFFE_PP_  (.D(\dp.result2[6] ),
    .DE(_0030_),
    .Q(\dp.rf.rf[9][6] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][7]$_DFFE_PP_  (.D(\dp.result2[7] ),
    .DE(net732),
    .Q(\dp.rf.rf[9][7] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][8]$_DFFE_PP_  (.D(\dp.result2[8] ),
    .DE(net732),
    .Q(\dp.rf.rf[9][8] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \dp.rf.rf[9][9]$_DFFE_PP_  (.D(\dp.result2[9] ),
    .DE(net732),
    .Q(\dp.rf.rf[9][9] ),
    .CLK(clknet_5_18__leaf_clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_1780 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(instr[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(instr[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(instr[11]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(instr[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_12 input5 (.A(instr[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(instr[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_12 input7 (.A(instr[15]),
    .X(net7));
 sky130_fd_sc_hd__buf_12 input8 (.A(instr[16]),
    .X(net8));
 sky130_fd_sc_hd__buf_12 input9 (.A(instr[17]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 input10 (.A(instr[18]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(instr[19]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(instr[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_12 input13 (.A(instr[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_12 input14 (.A(instr[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_12 input15 (.A(instr[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_12 input16 (.A(instr[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_12 input17 (.A(instr[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(instr[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(instr[26]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(instr[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(instr[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(instr[29]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(instr[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(instr[30]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(instr[31]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(instr[3]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(instr[4]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(instr[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(instr[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(instr[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(instr[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(instr[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(readdata[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(readdata[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(readdata[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(readdata[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(readdata[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(readdata[14]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(readdata[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input40 (.A(readdata[16]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(readdata[17]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(readdata[18]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(readdata[19]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(readdata[1]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(readdata[20]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(readdata[21]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(readdata[22]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(readdata[23]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(readdata[24]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input50 (.A(readdata[25]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(readdata[26]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(readdata[27]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(readdata[28]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(readdata[29]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(readdata[2]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(readdata[30]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(readdata[31]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(readdata[3]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(readdata[4]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input60 (.A(readdata[5]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(readdata[6]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(readdata[7]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(readdata[8]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(readdata[9]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input65 (.A(reset),
    .X(net65));
 sky130_fd_sc_hd__buf_6 output66 (.A(net66),
    .X(aluout[0]));
 sky130_fd_sc_hd__buf_6 output67 (.A(net67),
    .X(aluout[10]));
 sky130_fd_sc_hd__clkbuf_2 output68 (.A(net68),
    .X(aluout[11]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(aluout[12]));
 sky130_fd_sc_hd__buf_6 output70 (.A(net70),
    .X(aluout[13]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(aluout[14]));
 sky130_fd_sc_hd__buf_6 output72 (.A(net72),
    .X(aluout[15]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(aluout[16]));
 sky130_fd_sc_hd__buf_6 output74 (.A(net74),
    .X(aluout[17]));
 sky130_fd_sc_hd__buf_4 output75 (.A(net75),
    .X(aluout[18]));
 sky130_fd_sc_hd__buf_6 output76 (.A(net76),
    .X(aluout[19]));
 sky130_fd_sc_hd__clkbuf_2 output77 (.A(net77),
    .X(aluout[1]));
 sky130_fd_sc_hd__buf_6 output78 (.A(net78),
    .X(aluout[20]));
 sky130_fd_sc_hd__buf_6 output79 (.A(net79),
    .X(aluout[21]));
 sky130_fd_sc_hd__buf_6 output80 (.A(net80),
    .X(aluout[22]));
 sky130_fd_sc_hd__buf_4 output81 (.A(net81),
    .X(aluout[23]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(aluout[24]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(aluout[25]));
 sky130_fd_sc_hd__buf_1 output84 (.A(net84),
    .X(aluout[26]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(aluout[27]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(aluout[28]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(aluout[29]));
 sky130_fd_sc_hd__buf_1 output88 (.A(net88),
    .X(aluout[2]));
 sky130_fd_sc_hd__buf_4 output89 (.A(net89),
    .X(aluout[30]));
 sky130_fd_sc_hd__buf_6 output90 (.A(net90),
    .X(aluout[31]));
 sky130_fd_sc_hd__buf_6 output91 (.A(net91),
    .X(aluout[3]));
 sky130_fd_sc_hd__buf_6 output92 (.A(net92),
    .X(aluout[4]));
 sky130_fd_sc_hd__buf_6 output93 (.A(net93),
    .X(aluout[5]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(aluout[6]));
 sky130_fd_sc_hd__buf_6 output95 (.A(net95),
    .X(aluout[7]));
 sky130_fd_sc_hd__buf_6 output96 (.A(net96),
    .X(aluout[8]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(aluout[9]));
 sky130_fd_sc_hd__buf_1 output98 (.A(net98),
    .X(memread));
 sky130_fd_sc_hd__buf_1 output99 (.A(net99),
    .X(memwrite));
 sky130_fd_sc_hd__buf_1 output100 (.A(net100),
    .X(pc[0]));
 sky130_fd_sc_hd__buf_1 output101 (.A(net101),
    .X(pc[10]));
 sky130_fd_sc_hd__buf_1 output102 (.A(net102),
    .X(pc[11]));
 sky130_fd_sc_hd__buf_1 output103 (.A(net103),
    .X(pc[12]));
 sky130_fd_sc_hd__buf_1 output104 (.A(net104),
    .X(pc[13]));
 sky130_fd_sc_hd__buf_1 output105 (.A(net105),
    .X(pc[14]));
 sky130_fd_sc_hd__buf_1 output106 (.A(net106),
    .X(pc[15]));
 sky130_fd_sc_hd__buf_1 output107 (.A(net107),
    .X(pc[16]));
 sky130_fd_sc_hd__buf_1 output108 (.A(net108),
    .X(pc[17]));
 sky130_fd_sc_hd__buf_1 output109 (.A(net109),
    .X(pc[18]));
 sky130_fd_sc_hd__buf_1 output110 (.A(net110),
    .X(pc[19]));
 sky130_fd_sc_hd__buf_1 output111 (.A(net111),
    .X(pc[1]));
 sky130_fd_sc_hd__buf_1 output112 (.A(net112),
    .X(pc[20]));
 sky130_fd_sc_hd__buf_1 output113 (.A(net113),
    .X(pc[21]));
 sky130_fd_sc_hd__buf_1 output114 (.A(net114),
    .X(pc[22]));
 sky130_fd_sc_hd__buf_1 output115 (.A(net115),
    .X(pc[23]));
 sky130_fd_sc_hd__buf_1 output116 (.A(net116),
    .X(pc[24]));
 sky130_fd_sc_hd__buf_1 output117 (.A(net117),
    .X(pc[25]));
 sky130_fd_sc_hd__buf_1 output118 (.A(net118),
    .X(pc[26]));
 sky130_fd_sc_hd__buf_1 output119 (.A(net119),
    .X(pc[27]));
 sky130_fd_sc_hd__buf_1 output120 (.A(net120),
    .X(pc[28]));
 sky130_fd_sc_hd__buf_1 output121 (.A(net121),
    .X(pc[29]));
 sky130_fd_sc_hd__buf_1 output122 (.A(net122),
    .X(pc[2]));
 sky130_fd_sc_hd__buf_1 output123 (.A(net123),
    .X(pc[30]));
 sky130_fd_sc_hd__buf_1 output124 (.A(net124),
    .X(pc[31]));
 sky130_fd_sc_hd__buf_1 output125 (.A(net125),
    .X(pc[3]));
 sky130_fd_sc_hd__buf_1 output126 (.A(net126),
    .X(pc[4]));
 sky130_fd_sc_hd__buf_1 output127 (.A(net127),
    .X(pc[5]));
 sky130_fd_sc_hd__buf_1 output128 (.A(net128),
    .X(pc[6]));
 sky130_fd_sc_hd__buf_1 output129 (.A(net129),
    .X(pc[7]));
 sky130_fd_sc_hd__buf_1 output130 (.A(net130),
    .X(pc[8]));
 sky130_fd_sc_hd__buf_1 output131 (.A(net131),
    .X(pc[9]));
 sky130_fd_sc_hd__buf_1 output132 (.A(net132),
    .X(suspend));
 sky130_fd_sc_hd__buf_1 output133 (.A(net133),
    .X(writedata[0]));
 sky130_fd_sc_hd__buf_1 output134 (.A(net134),
    .X(writedata[10]));
 sky130_fd_sc_hd__buf_1 output135 (.A(net135),
    .X(writedata[11]));
 sky130_fd_sc_hd__buf_1 output136 (.A(net136),
    .X(writedata[12]));
 sky130_fd_sc_hd__buf_1 output137 (.A(net137),
    .X(writedata[13]));
 sky130_fd_sc_hd__buf_1 output138 (.A(net138),
    .X(writedata[14]));
 sky130_fd_sc_hd__buf_1 output139 (.A(net139),
    .X(writedata[15]));
 sky130_fd_sc_hd__buf_1 output140 (.A(net140),
    .X(writedata[16]));
 sky130_fd_sc_hd__buf_1 output141 (.A(net141),
    .X(writedata[17]));
 sky130_fd_sc_hd__buf_1 output142 (.A(net142),
    .X(writedata[18]));
 sky130_fd_sc_hd__buf_1 output143 (.A(net143),
    .X(writedata[19]));
 sky130_fd_sc_hd__buf_1 output144 (.A(net144),
    .X(writedata[1]));
 sky130_fd_sc_hd__buf_1 output145 (.A(net145),
    .X(writedata[20]));
 sky130_fd_sc_hd__buf_1 output146 (.A(net146),
    .X(writedata[21]));
 sky130_fd_sc_hd__buf_1 output147 (.A(net147),
    .X(writedata[22]));
 sky130_fd_sc_hd__buf_1 output148 (.A(net148),
    .X(writedata[23]));
 sky130_fd_sc_hd__buf_1 output149 (.A(net149),
    .X(writedata[24]));
 sky130_fd_sc_hd__buf_1 output150 (.A(net150),
    .X(writedata[25]));
 sky130_fd_sc_hd__buf_1 output151 (.A(net151),
    .X(writedata[26]));
 sky130_fd_sc_hd__buf_1 output152 (.A(net152),
    .X(writedata[27]));
 sky130_fd_sc_hd__buf_1 output153 (.A(net153),
    .X(writedata[28]));
 sky130_fd_sc_hd__buf_1 output154 (.A(net154),
    .X(writedata[29]));
 sky130_fd_sc_hd__buf_1 output155 (.A(net239),
    .X(writedata[2]));
 sky130_fd_sc_hd__buf_1 output156 (.A(net156),
    .X(writedata[30]));
 sky130_fd_sc_hd__buf_1 output157 (.A(net157),
    .X(writedata[31]));
 sky130_fd_sc_hd__buf_1 output158 (.A(net158),
    .X(writedata[3]));
 sky130_fd_sc_hd__buf_1 output159 (.A(net159),
    .X(writedata[4]));
 sky130_fd_sc_hd__buf_1 output160 (.A(net160),
    .X(writedata[5]));
 sky130_fd_sc_hd__buf_1 output161 (.A(net161),
    .X(writedata[6]));
 sky130_fd_sc_hd__buf_1 output162 (.A(net162),
    .X(writedata[7]));
 sky130_fd_sc_hd__buf_1 output163 (.A(net163),
    .X(writedata[8]));
 sky130_fd_sc_hd__buf_1 output164 (.A(net164),
    .X(writedata[9]));
 sky130_fd_sc_hd__buf_2 place766 (.A(_3238_[0]),
    .X(net766));
 sky130_fd_sc_hd__buf_1 place776 (.A(_2648_),
    .X(net776));
 sky130_fd_sc_hd__buf_12 place778 (.A(_1918_),
    .X(net778));
 sky130_fd_sc_hd__buf_1 place792 (.A(_0259_),
    .X(net792));
 sky130_fd_sc_hd__buf_1 place787 (.A(_0298_),
    .X(net787));
 sky130_fd_sc_hd__buf_12 place784 (.A(_0412_),
    .X(net784));
 sky130_fd_sc_hd__buf_1 place790 (.A(_0265_),
    .X(net790));
 sky130_fd_sc_hd__buf_1 place795 (.A(_0224_),
    .X(net795));
 sky130_fd_sc_hd__clkbuf_2 place759 (.A(_3374_[0]),
    .X(net759));
 sky130_fd_sc_hd__buf_12 place796 (.A(_0193_),
    .X(net796));
 sky130_fd_sc_hd__buf_12 place805 (.A(net804),
    .X(net805));
 sky130_fd_sc_hd__buf_12 place800 (.A(_0231_),
    .X(net800));
 sky130_fd_sc_hd__buf_12 place802 (.A(_0116_),
    .X(net802));
 sky130_fd_sc_hd__buf_12 place826 (.A(net13),
    .X(net826));
 sky130_fd_sc_hd__buf_12 place811 (.A(net810),
    .X(net811));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][15]$_DFFE_PP__7  (.LO(net171));
 sky130_fd_sc_hd__buf_1 place757 (.A(_1405_),
    .X(net757));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][21]$_DFFE_PP__12  (.LO(net176));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][12]$_DFFE_PP__4  (.LO(net168));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][11]$_DFFE_PP__3  (.LO(net167));
 sky130_fd_sc_hd__buf_12 place824 (.A(net823),
    .X(net824));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][14]$_DFFE_PP__6  (.LO(net170));
 sky130_fd_sc_hd__buf_12 place747 (.A(_1803_),
    .X(net747));
 sky130_fd_sc_hd__buf_12 place807 (.A(net806),
    .X(net807));
 sky130_fd_sc_hd__buf_12 place812 (.A(net7),
    .X(net812));
 sky130_fd_sc_hd__buf_12 place707 (.A(_0014_),
    .X(net707));
 sky130_fd_sc_hd__buf_12 place818 (.A(net15),
    .X(net818));
 sky130_fd_sc_hd__buf_12 place706 (.A(_0012_),
    .X(net706));
 sky130_fd_sc_hd__buf_12 place696 (.A(\dp.result2[29] ),
    .X(net696));
 sky130_fd_sc_hd__buf_12 place738 (.A(_1821_),
    .X(net738));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][0]$_DFFE_PP__1  (.LO(net165));
 sky130_fd_sc_hd__buf_12 place699 (.A(\dp.result2[19] ),
    .X(net699));
 sky130_fd_sc_hd__buf_12 place819 (.A(net14),
    .X(net819));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][13]$_DFFE_PP__5  (.LO(net169));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][19]$_DFFE_PP__10  (.LO(net174));
 sky130_fd_sc_hd__buf_12 place694 (.A(\dp.result2[31] ),
    .X(net694));
 sky130_fd_sc_hd__buf_12 place695 (.A(\dp.result2[30] ),
    .X(net695));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][22]$_DFFE_PP__13  (.LO(net177));
 sky130_fd_sc_hd__buf_1 place755 (.A(_3406_[0]),
    .X(net755));
 sky130_fd_sc_hd__buf_12 place769 (.A(net337),
    .X(net769));
 sky130_fd_sc_hd__buf_1 rebuffer132 (.A(net78),
    .X(net325));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][1]$_DFFE_PP__11  (.LO(net175));
 sky130_fd_sc_hd__buf_12 place797 (.A(_0193_),
    .X(net797));
 sky130_fd_sc_hd__buf_12 place705 (.A(_0013_),
    .X(net705));
 sky130_fd_sc_hd__buf_1 place708 (.A(_0015_),
    .X(net708));
 sky130_fd_sc_hd__clkbuf_2 place771 (.A(net337),
    .X(net771));
 sky130_fd_sc_hd__buf_12 place698 (.A(\dp.result2[26] ),
    .X(net698));
 sky130_fd_sc_hd__buf_12 place700 (.A(\dp.result2[17] ),
    .X(net700));
 sky130_fd_sc_hd__buf_1 place703 (.A(_2337_),
    .X(net703));
 sky130_fd_sc_hd__buf_12 place701 (.A(_2821_),
    .X(net701));
 sky130_fd_sc_hd__buf_12 place709 (.A(_0015_),
    .X(net709));
 sky130_fd_sc_hd__buf_12 place746 (.A(net331),
    .X(net746));
 sky130_fd_sc_hd__buf_12 place710 (.A(_0018_),
    .X(net710));
 sky130_fd_sc_hd__buf_12 place711 (.A(_0017_),
    .X(net711));
 sky130_fd_sc_hd__buf_12 place712 (.A(_0019_),
    .X(net712));
 sky130_fd_sc_hd__buf_12 place713 (.A(_0016_),
    .X(net713));
 sky130_fd_sc_hd__buf_12 place714 (.A(_0020_),
    .X(net714));
 sky130_fd_sc_hd__buf_12 place715 (.A(_0022_),
    .X(net715));
 sky130_fd_sc_hd__buf_2 place745 (.A(net331),
    .X(net745));
 sky130_fd_sc_hd__buf_12 place744 (.A(net331),
    .X(net744));
 sky130_fd_sc_hd__buf_12 place718 (.A(_0002_),
    .X(net718));
 sky130_fd_sc_hd__buf_12 place719 (.A(_0024_),
    .X(net719));
 sky130_fd_sc_hd__buf_12 place720 (.A(_0003_),
    .X(net720));
 sky130_fd_sc_hd__buf_12 place721 (.A(_0004_),
    .X(net721));
 sky130_fd_sc_hd__buf_12 place722 (.A(_0025_),
    .X(net722));
 sky130_fd_sc_hd__buf_12 place723 (.A(_0005_),
    .X(net723));
 sky130_fd_sc_hd__buf_12 place724 (.A(_0026_),
    .X(net724));
 sky130_fd_sc_hd__buf_12 place725 (.A(_0027_),
    .X(net725));
 sky130_fd_sc_hd__buf_12 place726 (.A(_0006_),
    .X(net726));
 sky130_fd_sc_hd__buf_12 place727 (.A(_0028_),
    .X(net727));
 sky130_fd_sc_hd__buf_12 place728 (.A(_0007_),
    .X(net728));
 sky130_fd_sc_hd__buf_12 place729 (.A(_0008_),
    .X(net729));
 sky130_fd_sc_hd__buf_12 place730 (.A(_0029_),
    .X(net730));
 sky130_fd_sc_hd__buf_12 place731 (.A(_0009_),
    .X(net731));
 sky130_fd_sc_hd__buf_12 place732 (.A(_0030_),
    .X(net732));
 sky130_fd_sc_hd__buf_12 place733 (.A(_0000_),
    .X(net733));
 sky130_fd_sc_hd__buf_12 place734 (.A(_0011_),
    .X(net734));
 sky130_fd_sc_hd__buf_12 place735 (.A(_0001_),
    .X(net735));
 sky130_fd_sc_hd__buf_12 place736 (.A(_0021_),
    .X(net736));
 sky130_fd_sc_hd__buf_12 place737 (.A(_1821_),
    .X(net737));
 sky130_fd_sc_hd__buf_12 place740 (.A(net271),
    .X(net740));
 sky130_fd_sc_hd__buf_12 place748 (.A(_1803_),
    .X(net748));
 sky130_fd_sc_hd__buf_1 place781 (.A(_0185_),
    .X(net781));
 sky130_fd_sc_hd__buf_12 place788 (.A(_0298_),
    .X(net788));
 sky130_fd_sc_hd__buf_1 rebuffer32 (.A(net701),
    .X(net224));
 sky130_fd_sc_hd__buf_12 place751 (.A(net249),
    .X(net751));
 sky130_fd_sc_hd__buf_12 place743 (.A(net308),
    .X(net743));
 sky130_fd_sc_hd__buf_12 place750 (.A(_1801_),
    .X(net750));
 sky130_fd_sc_hd__buf_1 place753 (.A(_3422_[0]),
    .X(net753));
 sky130_fd_sc_hd__buf_12 place752 (.A(net245),
    .X(net752));
 sky130_fd_sc_hd__buf_2 rebuffer60 (.A(net270),
    .X(net252));
 sky130_fd_sc_hd__buf_1 place756 (.A(_3398_[0]),
    .X(net756));
 sky130_fd_sc_hd__buf_12 place820 (.A(net14),
    .X(net820));
 sky130_fd_sc_hd__buf_1 place767 (.A(_3214_[0]),
    .X(net767));
 sky130_fd_sc_hd__buf_1 place763 (.A(_3334_[0]),
    .X(net763));
 sky130_fd_sc_hd__clkbuf_2 place761 (.A(_3358_[0]),
    .X(net761));
 sky130_fd_sc_hd__buf_4 place775 (.A(_1670_),
    .X(net775));
 sky130_fd_sc_hd__buf_1 place793 (.A(_0255_),
    .X(net793));
 sky130_fd_sc_hd__buf_12 place780 (.A(_0185_),
    .X(net780));
 sky130_fd_sc_hd__buf_1 place782 (.A(_0148_),
    .X(net782));
 sky130_fd_sc_hd__buf_1 place760 (.A(_3366_[0]),
    .X(net760));
 sky130_fd_sc_hd__buf_12 place810 (.A(net7),
    .X(net810));
 sky130_fd_sc_hd__buf_12 place808 (.A(net8),
    .X(net808));
 sky130_fd_sc_hd__buf_1 place758 (.A(_1364_),
    .X(net758));
 sky130_fd_sc_hd__buf_12 place804 (.A(net9),
    .X(net804));
 sky130_fd_sc_hd__buf_2 place754 (.A(_3414_[0]),
    .X(net754));
 sky130_fd_sc_hd__buf_12 place823 (.A(net822),
    .X(net823));
 sky130_fd_sc_hd__buf_12 place717 (.A(_0010_),
    .X(net717));
 sky130_fd_sc_hd__buf_12 place716 (.A(_0023_),
    .X(net716));
 sky130_fd_sc_hd__buf_12 place817 (.A(net16),
    .X(net817));
 sky130_fd_sc_hd__buf_12 place770 (.A(net337),
    .X(net770));
 sky130_fd_sc_hd__buf_12 place749 (.A(_1803_),
    .X(net749));
 sky130_fd_sc_hd__buf_12 place741 (.A(net268),
    .X(net741));
 sky130_fd_sc_hd__buf_12 place697 (.A(\dp.result2[27] ),
    .X(net697));
 sky130_fd_sc_hd__buf_12 place742 (.A(_1810_),
    .X(net742));
 sky130_fd_sc_hd__buf_12 place777 (.A(_2029_),
    .X(net777));
 sky130_fd_sc_hd__clkbuf_2 place764 (.A(_3318_[0]),
    .X(net764));
 sky130_fd_sc_hd__buf_2 place765 (.A(_3302_[0]),
    .X(net765));
 sky130_fd_sc_hd__buf_12 place768 (.A(net338),
    .X(net768));
 sky130_fd_sc_hd__buf_1 place772 (.A(_3062_),
    .X(net772));
 sky130_fd_sc_hd__buf_1 place814 (.A(net6),
    .X(net814));
 sky130_fd_sc_hd__buf_12 place825 (.A(net13),
    .X(net825));
 sky130_fd_sc_hd__buf_12 place816 (.A(net24),
    .X(net816));
 sky130_fd_sc_hd__buf_12 place774 (.A(_1708_),
    .X(net774));
 sky130_fd_sc_hd__buf_12 place773 (.A(_1711_),
    .X(net773));
 sky130_fd_sc_hd__buf_12 place789 (.A(_0265_),
    .X(net789));
 sky130_fd_sc_hd__buf_1 place783 (.A(_0620_),
    .X(net783));
 sky130_fd_sc_hd__buf_1 place785 (.A(_0389_),
    .X(net785));
 sky130_fd_sc_hd__buf_12 place786 (.A(_0304_),
    .X(net786));
 sky130_fd_sc_hd__buf_12 place791 (.A(_0259_),
    .X(net791));
 sky130_fd_sc_hd__buf_12 place794 (.A(_0224_),
    .X(net794));
 sky130_fd_sc_hd__buf_12 place806 (.A(net804),
    .X(net806));
 sky130_fd_sc_hd__buf_1 place798 (.A(_0166_),
    .X(net798));
 sky130_fd_sc_hd__buf_12 place799 (.A(_0137_),
    .X(net799));
 sky130_fd_sc_hd__buf_12 place801 (.A(_0173_),
    .X(net801));
 sky130_fd_sc_hd__buf_1 place803 (.A(_0040_),
    .X(net803));
 sky130_fd_sc_hd__buf_12 place821 (.A(net14),
    .X(net821));
 sky130_fd_sc_hd__buf_12 place809 (.A(net7),
    .X(net809));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][10]$_DFFE_PP__2  (.LO(net166));
 sky130_fd_sc_hd__buf_1 place815 (.A(net4),
    .X(net815));
 sky130_fd_sc_hd__buf_12 place822 (.A(net13),
    .X(net822));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][18]$_DFFE_PP__9  (.LO(net173));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][17]$_DFFE_PP__8  (.LO(net172));
 sky130_fd_sc_hd__buf_12 place739 (.A(_1821_),
    .X(net739));
 sky130_fd_sc_hd__buf_12 place813 (.A(net812),
    .X(net813));
 sky130_fd_sc_hd__buf_6 place702 (.A(_2258_),
    .X(net702));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][23]$_DFFE_PP__14  (.LO(net178));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][24]$_DFFE_PP__15  (.LO(net179));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][25]$_DFFE_PP__16  (.LO(net180));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][27]$_DFFE_PP__17  (.LO(net181));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][28]$_DFFE_PP__18  (.LO(net182));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][29]$_DFFE_PP__19  (.LO(net183));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][30]$_DFFE_PP__20  (.LO(net184));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][31]$_DFFE_PP__21  (.LO(net185));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][3]$_DFFE_PP__22  (.LO(net186));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][4]$_DFFE_PP__23  (.LO(net187));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][5]$_DFFE_PP__24  (.LO(net188));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][6]$_DFFE_PP__25  (.LO(net189));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][7]$_DFFE_PP__26  (.LO(net190));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][8]$_DFFE_PP__27  (.LO(net191));
 sky130_fd_sc_hd__conb_1 \dp.rf.rf[0][9]$_DFFE_PP__28  (.LO(net192));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_150_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_159_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_162_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_169_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_189_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_192_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_193_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_193_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_194_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_195_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_196_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_198_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_199_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_200_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_201_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_202_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_202_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_203_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_203_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_204_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_204_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_205_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_205_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_206_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_206_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_207_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_207_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_208_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_208_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_209_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_209_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_210_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_210_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_211_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_211_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_212_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_212_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_213_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_213_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_214_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_214_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_215_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_215_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_216_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_216_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_217_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_217_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_218_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_218_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_219_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_219_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_220_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_220_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_221_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_221_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_222_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_222_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_223_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_223_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_224_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_224_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_225_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_225_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_226_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_226_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_227_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_227_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_228_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_228_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_229_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_229_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_230_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_230_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_231_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_231_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_232_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_232_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_233_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_233_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_234_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_234_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_235_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_235_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_236_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_236_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_237_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_237_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_238_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_238_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_239_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_239_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_240_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_240_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_241_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_241_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_242_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_242_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_243_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_243_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_244_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_244_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_245_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_245_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_246_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_246_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_247_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_247_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_248_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_248_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_249_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_249_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_250_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_250_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_251_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_251_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_254_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_254_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_255_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_255_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_256_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_256_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_257_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_257_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_258_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_258_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_259_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_259_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_260_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_260_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_262_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_262_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_263_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_263_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_264_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_264_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_265_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_265_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_266_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_266_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_267_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_267_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_268_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_268_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_269_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_269_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_270_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_270_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_271_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_271_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_272_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_272_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_273_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_273_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_274_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_274_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_275_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_275_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_276_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_276_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_277_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_277_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_278_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_278_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_279_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_279_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_280_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_280_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_281_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_281_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_282_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_282_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_283_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_283_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_284_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_284_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_285_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_285_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_286_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_286_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_287_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_287_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_288_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_288_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_289_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_289_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_290_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_290_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_291_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_291_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_292_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_292_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_293_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_293_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_294_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_294_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_295_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_295_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_296_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_296_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_297_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_297_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_298_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_298_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_299_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_299_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_300_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_300_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_301_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_301_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_302_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_302_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload0 (.A(clknet_5_0__leaf_clk));
 sky130_fd_sc_hd__clkinv_16 clkload1 (.A(clknet_5_5__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload2 (.A(clknet_5_6__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload3 (.A(clknet_5_9__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload4 (.A(clknet_5_11__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload5 (.A(clknet_5_13__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload6 (.A(clknet_5_19__leaf_clk));
 sky130_fd_sc_hd__inv_12 clkload7 (.A(clknet_5_20__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload8 (.A(clknet_5_23__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload9 (.A(clknet_5_25__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload10 (.A(clknet_5_27__leaf_clk));
 sky130_fd_sc_hd__inv_12 clkload11 (.A(clknet_5_29__leaf_clk));
 sky130_fd_sc_hd__inv_16 clkload12 (.A(clknet_5_30__leaf_clk));
 sky130_fd_sc_hd__clkinv_2 clkload13 (.A(clknet_leaf_286_clk));
 sky130_fd_sc_hd__clkinv_2 clkload14 (.A(clknet_leaf_292_clk));
 sky130_fd_sc_hd__clkinv_1 clkload15 (.A(clknet_leaf_293_clk));
 sky130_fd_sc_hd__clkinv_1 clkload16 (.A(clknet_leaf_294_clk));
 sky130_fd_sc_hd__bufinv_16 clkload17 (.A(clknet_leaf_270_clk));
 sky130_fd_sc_hd__bufinv_16 clkload18 (.A(clknet_leaf_276_clk));
 sky130_fd_sc_hd__clkinv_2 clkload19 (.A(clknet_leaf_277_clk));
 sky130_fd_sc_hd__clkinv_1 clkload20 (.A(clknet_leaf_278_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload21 (.A(clknet_leaf_279_clk));
 sky130_fd_sc_hd__clkinv_1 clkload22 (.A(clknet_leaf_285_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload23 (.A(clknet_leaf_296_clk));
 sky130_fd_sc_hd__clkinv_1 clkload24 (.A(clknet_leaf_235_clk));
 sky130_fd_sc_hd__clkinv_2 clkload25 (.A(clknet_leaf_237_clk));
 sky130_fd_sc_hd__clkinv_2 clkload26 (.A(clknet_leaf_283_clk));
 sky130_fd_sc_hd__clkinv_2 clkload27 (.A(clknet_leaf_284_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload28 (.A(clknet_leaf_288_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload29 (.A(clknet_leaf_289_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload30 (.A(clknet_leaf_242_clk));
 sky130_fd_sc_hd__clkinv_2 clkload31 (.A(clknet_leaf_254_clk));
 sky130_fd_sc_hd__clkinv_1 clkload32 (.A(clknet_leaf_255_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload33 (.A(clknet_leaf_268_clk));
 sky130_fd_sc_hd__clkinv_1 clkload34 (.A(clknet_leaf_280_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload35 (.A(clknet_leaf_281_clk));
 sky130_fd_sc_hd__clkinv_1 clkload36 (.A(clknet_leaf_282_clk));
 sky130_fd_sc_hd__bufinv_16 clkload37 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__bufinv_16 clkload38 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkinv_2 clkload39 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkinv_1 clkload40 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload41 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkinv_2 clkload42 (.A(clknet_leaf_297_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload43 (.A(clknet_leaf_298_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload44 (.A(clknet_leaf_299_clk));
 sky130_fd_sc_hd__clkinv_2 clkload45 (.A(clknet_leaf_300_clk));
 sky130_fd_sc_hd__clkinv_2 clkload46 (.A(clknet_leaf_301_clk));
 sky130_fd_sc_hd__clkinv_2 clkload47 (.A(clknet_leaf_302_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload48 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload49 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload50 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkinv_1 clkload51 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload52 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkinv_1 clkload53 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__bufinv_16 clkload54 (.A(clknet_leaf_256_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload55 (.A(clknet_leaf_265_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload56 (.A(clknet_leaf_267_clk));
 sky130_fd_sc_hd__bufinv_16 clkload57 (.A(clknet_leaf_271_clk));
 sky130_fd_sc_hd__clkinv_2 clkload58 (.A(clknet_leaf_272_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload59 (.A(clknet_leaf_273_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload60 (.A(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkinv_1 clkload61 (.A(clknet_leaf_259_clk));
 sky130_fd_sc_hd__clkinv_1 clkload62 (.A(clknet_leaf_260_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload63 (.A(clknet_leaf_262_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload64 (.A(clknet_leaf_263_clk));
 sky130_fd_sc_hd__clkinv_1 clkload65 (.A(clknet_leaf_266_clk));
 sky130_fd_sc_hd__clkinv_2 clkload66 (.A(clknet_leaf_225_clk));
 sky130_fd_sc_hd__clkinv_1 clkload67 (.A(clknet_leaf_226_clk));
 sky130_fd_sc_hd__clkinv_1 clkload68 (.A(clknet_leaf_228_clk));
 sky130_fd_sc_hd__clkinv_2 clkload69 (.A(clknet_leaf_229_clk));
 sky130_fd_sc_hd__bufinv_16 clkload70 (.A(clknet_leaf_230_clk));
 sky130_fd_sc_hd__clkinv_1 clkload71 (.A(clknet_leaf_231_clk));
 sky130_fd_sc_hd__clkinv_2 clkload72 (.A(clknet_leaf_232_clk));
 sky130_fd_sc_hd__clkinv_1 clkload73 (.A(clknet_leaf_233_clk));
 sky130_fd_sc_hd__bufinv_16 clkload74 (.A(clknet_leaf_234_clk));
 sky130_fd_sc_hd__clkinv_2 clkload75 (.A(clknet_leaf_236_clk));
 sky130_fd_sc_hd__clkinv_1 clkload76 (.A(clknet_leaf_238_clk));
 sky130_fd_sc_hd__bufinv_16 clkload77 (.A(clknet_leaf_239_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload78 (.A(clknet_leaf_222_clk));
 sky130_fd_sc_hd__clkinv_2 clkload79 (.A(clknet_leaf_223_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload80 (.A(clknet_leaf_240_clk));
 sky130_fd_sc_hd__bufinv_16 clkload81 (.A(clknet_leaf_243_clk));
 sky130_fd_sc_hd__clkinv_2 clkload82 (.A(clknet_leaf_244_clk));
 sky130_fd_sc_hd__clkinv_1 clkload83 (.A(clknet_leaf_245_clk));
 sky130_fd_sc_hd__clkinv_1 clkload84 (.A(clknet_leaf_247_clk));
 sky130_fd_sc_hd__clkinv_2 clkload85 (.A(clknet_leaf_248_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload86 (.A(clknet_leaf_249_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload87 (.A(clknet_leaf_206_clk));
 sky130_fd_sc_hd__clkinv_1 clkload88 (.A(clknet_leaf_207_clk));
 sky130_fd_sc_hd__clkinv_2 clkload89 (.A(clknet_leaf_208_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload90 (.A(clknet_leaf_209_clk));
 sky130_fd_sc_hd__clkinv_1 clkload91 (.A(clknet_leaf_210_clk));
 sky130_fd_sc_hd__clkinv_2 clkload92 (.A(clknet_leaf_211_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload93 (.A(clknet_leaf_213_clk));
 sky130_fd_sc_hd__clkinv_2 clkload94 (.A(clknet_leaf_214_clk));
 sky130_fd_sc_hd__clkinv_1 clkload95 (.A(clknet_leaf_216_clk));
 sky130_fd_sc_hd__clkinv_1 clkload96 (.A(clknet_leaf_217_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload97 (.A(clknet_leaf_218_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload98 (.A(clknet_leaf_196_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload99 (.A(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkinv_2 clkload100 (.A(clknet_leaf_198_clk));
 sky130_fd_sc_hd__bufinv_16 clkload101 (.A(clknet_leaf_200_clk));
 sky130_fd_sc_hd__bufinv_16 clkload102 (.A(clknet_leaf_201_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload103 (.A(clknet_leaf_202_clk));
 sky130_fd_sc_hd__clkinv_4 clkload104 (.A(clknet_leaf_203_clk));
 sky130_fd_sc_hd__clkinv_1 clkload105 (.A(clknet_leaf_204_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload106 (.A(clknet_leaf_205_clk));
 sky130_fd_sc_hd__clkinv_4 clkload107 (.A(clknet_leaf_220_clk));
 sky130_fd_sc_hd__clkinv_1 clkload108 (.A(clknet_leaf_221_clk));
 sky130_fd_sc_hd__clkinv_2 clkload109 (.A(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkinv_1 clkload110 (.A(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkinv_2 clkload111 (.A(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkinv_2 clkload112 (.A(clknet_leaf_193_clk));
 sky130_fd_sc_hd__clkinv_1 clkload113 (.A(clknet_leaf_258_clk));
 sky130_fd_sc_hd__clkinv_1 clkload114 (.A(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkinv_1 clkload115 (.A(clknet_leaf_169_clk));
 sky130_fd_sc_hd__clkinv_1 clkload116 (.A(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload117 (.A(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload118 (.A(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkinv_2 clkload119 (.A(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload120 (.A(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkinv_2 clkload121 (.A(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkinv_1 clkload122 (.A(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload123 (.A(clknet_leaf_195_clk));
 sky130_fd_sc_hd__clkinv_1 clkload124 (.A(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload125 (.A(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkinv_1 clkload126 (.A(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload127 (.A(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkinv_2 clkload128 (.A(clknet_leaf_189_clk));
 sky130_fd_sc_hd__clkinv_1 clkload129 (.A(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkinv_2 clkload130 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload131 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkinv_1 clkload132 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload133 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkinv_1 clkload134 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkinv_2 clkload135 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__bufinv_16 clkload136 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkinv_2 clkload137 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkinv_1 clkload138 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkinv_2 clkload139 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkinv_1 clkload140 (.A(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload141 (.A(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkinv_1 clkload142 (.A(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkinv_1 clkload143 (.A(clknet_leaf_65_clk));
 sky130_fd_sc_hd__bufinv_16 clkload144 (.A(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload145 (.A(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkinv_2 clkload146 (.A(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkinv_2 clkload147 (.A(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload148 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkinv_2 clkload149 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkinv_2 clkload150 (.A(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload151 (.A(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkinv_2 clkload152 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload153 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload154 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkinv_2 clkload155 (.A(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkinv_2 clkload156 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkinv_2 clkload157 (.A(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload158 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkinv_1 clkload159 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload160 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__bufinv_16 clkload161 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkinv_1 clkload162 (.A(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkinv_2 clkload163 (.A(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload164 (.A(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkinv_2 clkload165 (.A(clknet_leaf_58_clk));
 sky130_fd_sc_hd__bufinv_16 clkload166 (.A(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkinv_2 clkload167 (.A(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkinv_1 clkload168 (.A(clknet_leaf_74_clk));
 sky130_fd_sc_hd__bufinv_16 clkload169 (.A(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkinv_2 clkload170 (.A(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkinv_2 clkload171 (.A(clknet_leaf_79_clk));
 sky130_fd_sc_hd__bufinv_16 clkload172 (.A(clknet_leaf_90_clk));
 sky130_fd_sc_hd__bufinv_16 clkload173 (.A(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkinv_2 clkload174 (.A(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload175 (.A(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload176 (.A(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload177 (.A(clknet_leaf_95_clk));
 sky130_fd_sc_hd__bufinv_16 clkload178 (.A(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkinv_4 clkload179 (.A(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkinv_1 clkload180 (.A(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload181 (.A(clknet_leaf_99_clk));
 sky130_fd_sc_hd__bufinv_16 clkload182 (.A(clknet_leaf_100_clk));
 sky130_fd_sc_hd__bufinv_16 clkload183 (.A(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload184 (.A(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkinv_1 clkload185 (.A(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkinv_2 clkload186 (.A(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkinv_1 clkload187 (.A(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload188 (.A(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkinv_2 clkload189 (.A(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkinv_1 clkload190 (.A(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkinv_2 clkload191 (.A(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkinv_2 clkload192 (.A(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkinv_2 clkload193 (.A(clknet_leaf_86_clk));
 sky130_fd_sc_hd__bufinv_16 clkload194 (.A(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkinv_1 clkload195 (.A(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload196 (.A(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload197 (.A(clknet_leaf_109_clk));
 sky130_fd_sc_hd__bufinv_16 clkload198 (.A(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkinv_1 clkload199 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkinv_1 clkload200 (.A(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload201 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__bufinv_16 clkload202 (.A(clknet_leaf_40_clk));
 sky130_fd_sc_hd__bufinv_16 clkload203 (.A(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkinv_2 clkload204 (.A(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkinv_2 clkload205 (.A(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkinv_1 clkload206 (.A(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload207 (.A(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload208 (.A(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload209 (.A(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload210 (.A(clknet_leaf_135_clk));
 sky130_fd_sc_hd__bufinv_16 clkload211 (.A(clknet_leaf_111_clk));
 sky130_fd_sc_hd__bufinv_16 clkload212 (.A(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload213 (.A(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkinv_2 clkload214 (.A(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkinv_1 clkload215 (.A(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload216 (.A(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkinv_2 clkload217 (.A(clknet_leaf_117_clk));
 sky130_fd_sc_hd__bufinv_16 clkload218 (.A(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkinv_2 clkload219 (.A(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload220 (.A(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkinv_2 clkload221 (.A(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkinv_2 clkload222 (.A(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkinv_2 clkload223 (.A(clknet_leaf_107_clk));
 sky130_fd_sc_hd__bufinv_16 clkload224 (.A(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload225 (.A(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkinv_2 clkload226 (.A(clknet_leaf_126_clk));
 sky130_fd_sc_hd__bufinv_16 clkload227 (.A(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkinv_1 clkload228 (.A(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload229 (.A(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload230 (.A(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload231 (.A(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkinv_1 clkload232 (.A(clknet_leaf_162_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload233 (.A(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkinv_2 clkload234 (.A(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkinv_2 clkload235 (.A(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkinv_2 clkload236 (.A(clknet_leaf_166_clk));
 sky130_fd_sc_hd__buf_4 rebuffer1 (.A(_1752_),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_16 clone115 (.A(net309),
    .X(net308));
 sky130_fd_sc_hd__buf_1 rebuffer114 (.A(_1881_),
    .X(net307));
 sky130_fd_sc_hd__buf_1 rebuffer105 (.A(_2016_),
    .X(net298));
 sky130_fd_sc_hd__buf_6 rebuffer104 (.A(\dp.rf.rf[26][23] ),
    .X(net297));
 sky130_fd_sc_hd__buf_1 rebuffer99 (.A(_2381_),
    .X(net292));
 sky130_fd_sc_hd__buf_1 rebuffer96 (.A(net82),
    .X(net289));
 sky130_fd_sc_hd__buf_2 rebuffer93 (.A(net267),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_2 rebuffer92 (.A(_3254_[0]),
    .X(net285));
 sky130_fd_sc_hd__buf_1 rebuffer91 (.A(\dp.rf.rf[13][14] ),
    .X(net284));
 sky130_fd_sc_hd__buf_1 rebuffer90 (.A(\dp.rf.rf[12][14] ),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_2 rebuffer88 (.A(_3270_[0]),
    .X(net281));
 sky130_fd_sc_hd__buf_1 rebuffer78 (.A(_1628_),
    .X(net271));
 sky130_fd_sc_hd__buf_1 rebuffer70 (.A(_3237_[0]),
    .X(net270));
 sky130_fd_sc_hd__buf_1 rebuffer66 (.A(_1767_),
    .X(net262));
 sky130_fd_sc_hd__buf_1 rebuffer45 (.A(net66),
    .X(net256));
 sky130_fd_sc_hd__buf_2 rebuffer17 (.A(net210),
    .X(net209));
 sky130_fd_sc_hd__buf_2 rebuffer18 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__buf_2 rebuffer19 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__buf_2 rebuffer20 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__buf_2 rebuffer21 (.A(net214),
    .X(net213));
 sky130_fd_sc_hd__buf_2 rebuffer22 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__buf_2 rebuffer23 (.A(net216),
    .X(net215));
 sky130_fd_sc_hd__buf_2 rebuffer24 (.A(net217),
    .X(net216));
 sky130_fd_sc_hd__buf_2 rebuffer25 (.A(net218),
    .X(net217));
 sky130_fd_sc_hd__buf_6 rebuffer26 (.A(_1572_),
    .X(net218));
 sky130_fd_sc_hd__buf_4 rebuffer27 (.A(_2409_),
    .X(net219));
 sky130_fd_sc_hd__buf_1 rebuffer28 (.A(net219),
    .X(net220));
 sky130_fd_sc_hd__buf_1 rebuffer29 (.A(_2517_),
    .X(net221));
 sky130_fd_sc_hd__buf_1 rebuffer128 (.A(net74),
    .X(net321));
 sky130_fd_sc_hd__buf_6 rebuffer116 (.A(_1805_),
    .X(net309));
 sky130_fd_sc_hd__buf_1 rebuffer64 (.A(_1767_),
    .X(net258));
 sky130_fd_sc_hd__buf_6 rebuffer34 (.A(_2821_),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_16 clone33 (.A(_2821_),
    .X(net225));
 sky130_fd_sc_hd__buf_1 rebuffer31 (.A(net158),
    .X(net223));
 sky130_fd_sc_hd__buf_1 rebuffer30 (.A(net158),
    .X(net222));
 sky130_fd_sc_hd__buf_1 rebuffer190 (.A(net95),
    .X(net382));
 sky130_fd_sc_hd__buf_1 rebuffer121 (.A(_1964_),
    .X(net314));
 sky130_fd_sc_hd__buf_1 rebuffer120 (.A(_1964_),
    .X(net313));
 sky130_fd_sc_hd__buf_1 rebuffer119 (.A(net94),
    .X(net312));
 sky130_fd_sc_hd__buf_1 rebuffer41 (.A(net234),
    .X(net233));
 sky130_fd_sc_hd__buf_1 rebuffer42 (.A(net235),
    .X(net234));
 sky130_fd_sc_hd__buf_1 rebuffer43 (.A(net236),
    .X(net235));
 sky130_fd_sc_hd__buf_1 rebuffer44 (.A(_1744_),
    .X(net236));
 sky130_fd_sc_hd__buf_16 clone45 (.A(net226),
    .X(net237));
 sky130_fd_sc_hd__buf_1 rebuffer46 (.A(_1746_),
    .X(net238));
 sky130_fd_sc_hd__buf_1 rebuffer47 (.A(net155),
    .X(net239));
 sky130_fd_sc_hd__buf_2 rebuffer48 (.A(net155),
    .X(net240));
 sky130_fd_sc_hd__buf_6 rebuffer49 (.A(_2821_),
    .X(net241));
 sky130_fd_sc_hd__buf_1 rebuffer50 (.A(net241),
    .X(net242));
 sky130_fd_sc_hd__buf_1 rebuffer51 (.A(net241),
    .X(net243));
 sky130_fd_sc_hd__buf_1 rebuffer52 (.A(net256),
    .X(net244));
 sky130_fd_sc_hd__buf_1 rebuffer53 (.A(_1574_),
    .X(net245));
 sky130_fd_sc_hd__buf_1 rebuffer54 (.A(_3437_[0]),
    .X(net246));
 sky130_fd_sc_hd__buf_1 rebuffer55 (.A(net155),
    .X(net247));
 sky130_fd_sc_hd__buf_1 rebuffer56 (.A(net155),
    .X(net248));
 sky130_fd_sc_hd__buf_1 rebuffer57 (.A(_1672_),
    .X(net249));
 sky130_fd_sc_hd__buf_1 rebuffer58 (.A(\dp.rf.rf[29][1] ),
    .X(net250));
 sky130_fd_sc_hd__buf_1 rebuffer59 (.A(\dp.rf.rf[28][1] ),
    .X(net251));
 sky130_fd_sc_hd__buf_1 rebuffer61 (.A(_3237_[0]),
    .X(net253));
 sky130_fd_sc_hd__buf_1 rebuffer62 (.A(net81),
    .X(net254));
 sky130_fd_sc_hd__buf_1 rebuffer63 (.A(net83),
    .X(net255));
 sky130_fd_sc_hd__buf_12 rebuffer139 (.A(_1805_),
    .X(net331));
 sky130_fd_sc_hd__buf_1 rebuffer65 (.A(net289),
    .X(net257));
 sky130_fd_sc_hd__buf_1 rebuffer67 (.A(net80),
    .X(net259));
 sky130_fd_sc_hd__buf_1 rebuffer68 (.A(_2421_),
    .X(net260));
 sky130_fd_sc_hd__buf_2 rebuffer69 (.A(net89),
    .X(net261));
 sky130_fd_sc_hd__buf_1 rebuffer71 (.A(_3339_[0]),
    .X(net263));
 sky130_fd_sc_hd__buf_1 rebuffer72 (.A(_3341_[0]),
    .X(net264));
 sky130_fd_sc_hd__buf_1 rebuffer73 (.A(\dp.rf.rf[8][14] ),
    .X(net265));
 sky130_fd_sc_hd__buf_1 rebuffer74 (.A(\dp.rf.rf[9][14] ),
    .X(net266));
 sky130_fd_sc_hd__buf_2 rebuffer75 (.A(_2407_),
    .X(net267));
 sky130_fd_sc_hd__buf_1 rebuffer76 (.A(_1532_),
    .X(net268));
 sky130_fd_sc_hd__buf_1 rebuffer77 (.A(_1762_),
    .X(net269));
 sky130_fd_sc_hd__buf_1 rebuffer134 (.A(_1778_),
    .X(net326));
 sky130_fd_sc_hd__buf_1 rebuffer135 (.A(net86),
    .X(net327));
 sky130_fd_sc_hd__buf_1 rebuffer140 (.A(net71),
    .X(net332));
 sky130_fd_sc_hd__buf_1 rebuffer142 (.A(net79),
    .X(net334));
 sky130_fd_sc_hd__buf_1 rebuffer143 (.A(net325),
    .X(net335));
 sky130_fd_sc_hd__buf_12 rebuffer145 (.A(_0154_),
    .X(net337));
 sky130_fd_sc_hd__buf_1 rebuffer146 (.A(net337),
    .X(net338));
 sky130_fd_sc_hd__buf_1 rebuffer147 (.A(net337),
    .X(net339));
 sky130_fd_sc_hd__buf_1 rebuffer148 (.A(net329),
    .X(net340));
 sky130_fd_sc_hd__buf_1 rebuffer149 (.A(_2024_),
    .X(net341));
 sky130_fd_sc_hd__buf_1 rebuffer150 (.A(_2024_),
    .X(net342));
 sky130_fd_sc_hd__buf_1 rebuffer151 (.A(_1845_),
    .X(net343));
 sky130_fd_sc_hd__buf_1 rebuffer166 (.A(net321),
    .X(net358));
 sky130_fd_sc_hd__buf_1 rebuffer168 (.A(net96),
    .X(net360));
 sky130_fd_sc_hd__buf_1 rebuffer169 (.A(net70),
    .X(net361));
 sky130_fd_sc_hd__buf_1 rebuffer170 (.A(net702),
    .X(net362));
 sky130_fd_sc_hd__buf_1 rebuffer171 (.A(net702),
    .X(net363));
 sky130_fd_sc_hd__buf_1 rebuffer172 (.A(net292),
    .X(net364));
 sky130_fd_sc_hd__buf_1 rebuffer175 (.A(net69),
    .X(net367));
 sky130_fd_sc_hd__buf_1 rebuffer176 (.A(net72),
    .X(net368));
 sky130_fd_sc_hd__buf_1 rebuffer179 (.A(net97),
    .X(net371));
 sky130_fd_sc_hd__buf_1 rebuffer181 (.A(net67),
    .X(net373));
 sky130_fd_sc_hd__buf_1 rebuffer182 (.A(_2104_),
    .X(net374));
 sky130_fd_sc_hd__buf_1 rebuffer183 (.A(net68),
    .X(net375));
 sky130_fd_sc_hd__buf_1 rebuffer184 (.A(_2170_),
    .X(net376));
 sky130_fd_sc_hd__buf_1 rebuffer185 (.A(net93),
    .X(net377));
 sky130_fd_sc_hd__buf_1 rebuffer186 (.A(net88),
    .X(net378));
 sky130_fd_sc_hd__buf_1 rebuffer187 (.A(net308),
    .X(net379));
 sky130_fd_sc_hd__buf_1 rebuffer188 (.A(net77),
    .X(net380));
 sky130_fd_sc_hd__buf_1 rebuffer189 (.A(net92),
    .X(net381));
 sky130_fd_sc_hd__buf_1 rebuffer136 (.A(net91),
    .X(net329));
 sky130_fd_sc_hd__buf_1 rebuffer137 (.A(net159),
    .X(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(instr[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(instr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(instr[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(readdata[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(readdata[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(readdata[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(instr[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net735));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_0400_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(instr[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(instr[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(readdata[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(readdata[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(readdata[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(readdata[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(readdata[4]));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_777 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_653 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_714 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_777 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_606 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_777 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_484 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_777 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_452 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_570 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_387 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_534 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_400 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_777 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_583 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_614 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_750 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_548 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_240 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_168 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_572 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_653 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_550 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_782 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_540 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_771 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_524 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_770 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_733 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_594 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_520 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_710 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_272 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_392 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_242 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_554 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_666 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_196 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_747 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_464 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_733 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_620 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_584 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_668 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_732 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_498 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_136 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_552 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_774 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_782 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_730 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_380 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_460 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_498 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_630 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_417 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_732 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_762 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_520 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_514 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_744 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_337 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_594 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_709 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_620 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_717 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_734 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_117 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_766 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_384 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_486 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_498 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_726 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_782 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_640 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_516 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_720 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_216 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_653 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_516 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_540 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_692 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_704 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_709 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_87 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_488 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_576 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_768 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_638 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_766 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_572 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_640 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_246 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_470 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_540 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_730 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_777 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_711 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_450 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_683 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_709 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_668 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_774 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_782 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_709 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_740 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_420 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_777 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_548 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_670 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_650 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_773 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_201 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_443 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_584 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_141 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_330 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_512 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_756 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_708 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_612 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_698 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_417 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_537 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_717 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_604 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_234 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_534 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_452 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_495 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_740 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_460 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_488 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_756 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_462 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_644 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_261 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_426 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_614 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_714 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_614 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_678 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_704 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_734 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_86 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_417 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_740 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_444 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_704 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_420 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_668 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_501 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_550 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_150 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_384 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_687 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_766 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_660 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_444 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_640 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_774 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_674 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_777 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_462 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_432 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_747 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_484 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_708 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_636 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_801 ();
endmodule
