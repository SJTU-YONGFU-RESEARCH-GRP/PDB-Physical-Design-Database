module simple_spi_master (clk,
    rst_n,
    rx_valid,
    spi_clk,
    spi_cs_n,
    spi_miso,
    spi_mosi,
    tx_ready,
    tx_valid,
    rx_data,
    tx_data);
 input clk;
 input rst_n;
 output rx_valid;
 output spi_clk;
 output spi_cs_n;
 input spi_miso;
 output spi_mosi;
 output tx_ready;
 input tx_valid;
 output [7:0] rx_data;
 input [7:0] tx_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire \bit_count[0] ;
 wire \bit_count[1] ;
 wire \bit_count[2] ;
 wire \bit_count[3] ;
 wire \rx_shift_reg[0] ;
 wire \rx_shift_reg[1] ;
 wire \rx_shift_reg[2] ;
 wire \rx_shift_reg[3] ;
 wire \rx_shift_reg[4] ;
 wire \rx_shift_reg[5] ;
 wire \rx_shift_reg[6] ;
 wire \rx_shift_reg[7] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \tx_shift_reg[0] ;
 wire \tx_shift_reg[1] ;
 wire \tx_shift_reg[2] ;
 wire \tx_shift_reg[3] ;
 wire \tx_shift_reg[4] ;
 wire \tx_shift_reg[5] ;
 wire \tx_shift_reg[6] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net26;

 gf180mcu_fd_sc_mcu9t5v0__inv_3 _119_ (.I(\bit_count[3] ),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_2 _120_ (.A1(_100_),
    .A2(\bit_count[2] ),
    .A3(_098_),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _121_ (.I(_104_),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _122_ (.I(\bit_count[2] ),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _123_ (.I(\bit_count[0] ),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _124_ (.I(\bit_count[1] ),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu9t5v0__or3_2 _125_ (.A1(_096_),
    .A2(_097_),
    .A3(_034_),
    .Z(_101_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _126_ (.A1(\bit_count[3] ),
    .A2(_101_),
    .Z(_116_));
 gf180mcu_fd_sc_mcu9t5v0__inv_3 _127_ (.I(\state[0] ),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _128_ (.A1(_035_),
    .A2(net12),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _129_ (.A1(\bit_count[3] ),
    .A2(net22),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _130_ (.A1(\state[0] ),
    .A2(_037_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_4 _131_ (.A1(_036_),
    .A2(_038_),
    .B(\state[1] ),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_4 _132_ (.I(\state[1] ),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _133_ (.A1(\state[0] ),
    .A2(_040_),
    .A3(_037_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _134_ (.A1(_097_),
    .A2(_041_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _135_ (.A1(_097_),
    .A2(_039_),
    .B(_042_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _136_ (.A1(\state[0] ),
    .A2(_040_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu9t5v0__buf_4 _137_ (.I(_043_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _138_ (.A1(_037_),
    .A2(_044_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _139_ (.I(_099_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _140_ (.A1(_034_),
    .A2(_039_),
    .B1(_045_),
    .B2(_046_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_4 _141_ (.A1(\bit_count[2] ),
    .A2(_098_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _142_ (.A1(_096_),
    .A2(_039_),
    .B1(_045_),
    .B2(_047_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _143_ (.A1(_103_),
    .A2(_041_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _144_ (.A1(_100_),
    .A2(_039_),
    .B(_048_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_4 _145_ (.A1(_035_),
    .A2(\state[1] ),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _146_ (.I0(\rx_shift_reg[0] ),
    .I1(net13),
    .S(_049_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _147_ (.I0(\rx_shift_reg[1] ),
    .I1(net14),
    .S(_049_),
    .Z(_005_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _148_ (.I0(\rx_shift_reg[2] ),
    .I1(net15),
    .S(_049_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _149_ (.I0(\rx_shift_reg[3] ),
    .I1(net16),
    .S(_049_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _150_ (.I0(\rx_shift_reg[4] ),
    .I1(net17),
    .S(_049_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _151_ (.I0(\rx_shift_reg[5] ),
    .I1(net18),
    .S(_049_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _152_ (.I0(\rx_shift_reg[6] ),
    .I1(net19),
    .S(_049_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _153_ (.I0(\rx_shift_reg[7] ),
    .I1(net20),
    .S(_049_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _154_ (.A1(_114_),
    .A2(_112_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _155_ (.A1(\bit_count[0] ),
    .A2(_047_),
    .A3(_050_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _156_ (.A1(_102_),
    .A2(_117_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _157_ (.A1(_106_),
    .A2(_118_),
    .A3(_046_),
    .A4(_052_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _158_ (.A1(_103_),
    .A2(_041_),
    .A3(_051_),
    .A4(_053_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _159_ (.I0(\rx_shift_reg[0] ),
    .I1(net3),
    .S(_054_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _160_ (.A1(\bit_count[3] ),
    .A2(net22),
    .Z(_055_));
 gf180mcu_fd_sc_mcu9t5v0__nor4_4 _161_ (.A1(_035_),
    .A2(\state[1] ),
    .A3(_103_),
    .A4(_055_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _162_ (.A1(_099_),
    .A2(_056_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _163_ (.A1(_102_),
    .A2(_117_),
    .Z(_058_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _164_ (.A1(_106_),
    .A2(_118_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu9t5v0__and3_2 _165_ (.A1(_097_),
    .A2(net3),
    .A3(_050_),
    .Z(_060_));
 gf180mcu_fd_sc_mcu9t5v0__nand3_4 _166_ (.A1(_058_),
    .A2(_059_),
    .A3(_060_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu9t5v0__xor2_2 _167_ (.A1(\bit_count[2] ),
    .A2(_098_),
    .Z(_062_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _168_ (.A1(_100_),
    .A2(_097_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _169_ (.A1(_099_),
    .A2(_062_),
    .A3(_063_),
    .A4(_056_),
    .Z(_064_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _170_ (.I(\rx_shift_reg[1] ),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _171_ (.A1(_047_),
    .A2(_057_),
    .A3(_061_),
    .B1(_064_),
    .B2(_065_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _172_ (.A1(\bit_count[0] ),
    .A2(_050_),
    .A3(_058_),
    .A4(_059_),
    .Z(_066_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _173_ (.A1(_099_),
    .A2(_062_),
    .A3(_056_),
    .A4(_066_),
    .Z(_067_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _174_ (.I0(\rx_shift_reg[2] ),
    .I1(net3),
    .S(_067_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu9t5v0__or2_2 _175_ (.A1(_099_),
    .A2(_103_),
    .Z(_068_));
 gf180mcu_fd_sc_mcu9t5v0__or4_2 _176_ (.A1(_035_),
    .A2(\state[1] ),
    .A3(_055_),
    .A4(_068_),
    .Z(_069_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _177_ (.A1(\bit_count[0] ),
    .A2(_047_),
    .A3(_069_),
    .B(\rx_shift_reg[3] ),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _178_ (.A1(_047_),
    .A2(_061_),
    .A3(_069_),
    .B(_070_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _179_ (.A1(_046_),
    .A2(_062_),
    .A3(_056_),
    .A4(_066_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _180_ (.I0(\rx_shift_reg[4] ),
    .I1(net3),
    .S(_071_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _181_ (.A1(_099_),
    .A2(_047_),
    .A3(_063_),
    .A4(_056_),
    .Z(_072_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _182_ (.I(\rx_shift_reg[5] ),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu9t5v0__oai32_2 _183_ (.A1(_062_),
    .A2(_057_),
    .A3(_061_),
    .B1(_072_),
    .B2(_073_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu9t5v0__and4_2 _184_ (.A1(_099_),
    .A2(_047_),
    .A3(_056_),
    .A4(_066_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _185_ (.I0(\rx_shift_reg[6] ),
    .I1(net3),
    .S(_074_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _186_ (.A1(\bit_count[0] ),
    .A2(_062_),
    .A3(_069_),
    .B(\rx_shift_reg[7] ),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu9t5v0__oai31_2 _187_ (.A1(_062_),
    .A2(_061_),
    .A3(_069_),
    .B(_075_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _188_ (.I0(\state[1] ),
    .I1(net21),
    .S(\state[0] ),
    .Z(_020_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _189_ (.A1(_040_),
    .A2(_100_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu9t5v0__xnor2_2 _190_ (.A1(net22),
    .A2(_076_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu9t5v0__and2_2 _191_ (.A1(\state[0] ),
    .A2(_077_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _192_ (.A1(_040_),
    .A2(net12),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _193_ (.I0(net23),
    .I1(_078_),
    .S(_035_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _194_ (.I0(net11),
    .I1(\tx_shift_reg[6] ),
    .S(_044_),
    .Z(_079_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _195_ (.I(_110_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _196_ (.A1(\state[0] ),
    .A2(net22),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _197_ (.I(net12),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu9t5v0__oai22_2 _198_ (.A1(\state[0] ),
    .A2(_082_),
    .B1(_081_),
    .B2(\bit_count[3] ),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu9t5v0__oai211_2 _199_ (.A1(_080_),
    .A2(_081_),
    .B(_083_),
    .C(_040_),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _200_ (.I0(_079_),
    .I1(net24),
    .S(_084_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu9t5v0__oai21_2 _201_ (.A1(_107_),
    .A2(_055_),
    .B(\state[0] ),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu9t5v0__aoi21_2 _202_ (.A1(_036_),
    .A2(_085_),
    .B(\state[1] ),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _203_ (.A1(_107_),
    .A2(_045_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu9t5v0__nand2_2 _204_ (.A1(_035_),
    .A2(_040_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _205_ (.I0(_082_),
    .I1(net25),
    .S(_086_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_2 _206_ (.I(net4),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu9t5v0__nor2_2 _207_ (.A1(_087_),
    .A2(_044_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu9t5v0__and2_4 _208_ (.A1(_040_),
    .A2(_083_),
    .Z(_089_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _209_ (.I0(\tx_shift_reg[0] ),
    .I1(_088_),
    .S(_089_),
    .Z(_027_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _210_ (.I0(net5),
    .I1(\tx_shift_reg[0] ),
    .S(_044_),
    .Z(_090_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _211_ (.I0(\tx_shift_reg[1] ),
    .I1(_090_),
    .S(_089_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _212_ (.I0(net6),
    .I1(\tx_shift_reg[1] ),
    .S(_044_),
    .Z(_091_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _213_ (.I0(\tx_shift_reg[2] ),
    .I1(_091_),
    .S(_089_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _214_ (.I0(net7),
    .I1(\tx_shift_reg[2] ),
    .S(_044_),
    .Z(_092_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _215_ (.I0(\tx_shift_reg[3] ),
    .I1(_092_),
    .S(_089_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _216_ (.I0(net8),
    .I1(\tx_shift_reg[3] ),
    .S(_044_),
    .Z(_093_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _217_ (.I0(\tx_shift_reg[4] ),
    .I1(_093_),
    .S(_089_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _218_ (.I0(net9),
    .I1(\tx_shift_reg[4] ),
    .S(_044_),
    .Z(_094_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _219_ (.I0(\tx_shift_reg[5] ),
    .I1(_094_),
    .S(_089_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _220_ (.I0(net10),
    .I1(\tx_shift_reg[5] ),
    .S(_044_),
    .Z(_095_));
 gf180mcu_fd_sc_mcu9t5v0__mux2_2 _221_ (.I0(\tx_shift_reg[6] ),
    .I1(_095_),
    .S(_089_),
    .Z(_033_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _222_ (.A(\bit_count[0] ),
    .B(\bit_count[1] ),
    .CO(_098_),
    .S(_099_));
 gf180mcu_fd_sc_mcu9t5v0__addh_2 _223_ (.A(_100_),
    .B(_101_),
    .CO(_102_),
    .S(_103_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _224_ (.A(_100_),
    .B(_104_),
    .CO(_105_),
    .S(_106_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _225_ (.A(_100_),
    .B(_104_),
    .CO(_107_),
    .S(_108_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _226_ (.A(_100_),
    .B(_109_),
    .CO(_110_),
    .S(_111_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _227_ (.A(\bit_count[3] ),
    .B(_104_),
    .CO(_112_),
    .S(_113_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _228_ (.A(\bit_count[3] ),
    .B(_109_),
    .CO(_114_),
    .S(_115_));
 gf180mcu_fd_sc_mcu9t5v0__addh_1 _229_ (.A(_100_),
    .B(_116_),
    .CO(_117_),
    .S(_118_));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_count[0]$_DFFE_PN0P_  (.D(_000_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\bit_count[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_count[1]$_DFFE_PN0P_  (.D(_001_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\bit_count[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_count[2]$_DFFE_PN0P_  (.D(_002_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\bit_count[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \bit_count[3]$_DFFE_PN0P_  (.D(_003_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\bit_count[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[0]$_DFFE_PN0P_  (.D(_004_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net13));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[1]$_DFFE_PN0P_  (.D(_005_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net14));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[2]$_DFFE_PN0P_  (.D(_006_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net15));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[3]$_DFFE_PN0P_  (.D(_007_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net16));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[4]$_DFFE_PN0P_  (.D(_008_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net17));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[5]$_DFFE_PN0P_  (.D(_009_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[6]$_DFFE_PN0P_  (.D(_010_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_data[7]$_DFFE_PN0P_  (.D(_011_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[0]$_DFFE_PN0P_  (.D(_012_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\rx_shift_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[1]$_DFFE_PN0P_  (.D(_013_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\rx_shift_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[2]$_DFFE_PN0P_  (.D(_014_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\rx_shift_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[3]$_DFFE_PN0P_  (.D(_015_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\rx_shift_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[4]$_DFFE_PN0P_  (.D(_016_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\rx_shift_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[5]$_DFFE_PN0P_  (.D(_017_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\rx_shift_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[6]$_DFFE_PN0P_  (.D(_018_),
    .RN(net1),
    .CLK(clknet_2_1__leaf_clk),
    .Q(\rx_shift_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_shift_reg[7]$_DFFE_PN0P_  (.D(_019_),
    .RN(net1),
    .CLK(clknet_2_0__leaf_clk),
    .Q(\rx_shift_reg[7] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \rx_valid$_DFFE_PN0P_  (.D(_020_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \spi_clk$_DFFE_PN0P_  (.D(_021_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \spi_cs_n$_DFFE_PN1P_  (.D(_022_),
    .SETN(net2),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \spi_mosi$_DFFE_PN0P_  (.D(_023_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \state[0]$_DFFE_PN0P_  (.D(_024_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\state[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 \state[1]$_DFFE_PN0P_  (.D(_025_),
    .RN(net1),
    .CLK(clknet_2_2__leaf_clk),
    .Q(\state[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 \tx_ready$_DFFE_PN1P_  (.D(_026_),
    .SETN(net2),
    .CLK(clknet_2_2__leaf_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[0]$_DFFE_PN0P_  (.D(_027_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift_reg[0] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[1]$_DFFE_PN0P_  (.D(_028_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift_reg[1] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[2]$_DFFE_PN0P_  (.D(_029_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift_reg[2] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[3]$_DFFE_PN0P_  (.D(_030_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift_reg[3] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[4]$_DFFE_PN0P_  (.D(_031_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift_reg[4] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[5]$_DFFE_PN0P_  (.D(_032_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift_reg[5] ));
 gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 \tx_shift_reg[6]$_DFFE_PN0P_  (.D(_033_),
    .RN(net1),
    .CLK(clknet_2_3__leaf_clk),
    .Q(\tx_shift_reg[6] ));
 gf180mcu_fd_sc_mcu9t5v0__buf_12 hold1 (.I(net2),
    .Z(net1));
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_0_Left_26 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_1_Left_27 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_2_Left_28 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_3_Left_29 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_4_Left_30 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_5_Left_31 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_6_Left_32 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_7_Left_33 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_8_Left_34 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_9_Left_35 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_10_Left_36 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_11_Left_37 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_12_Left_38 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_13_Left_39 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_14_Left_40 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_15_Left_41 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_16_Left_42 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_17_Left_43 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_18_Left_44 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_19_Left_45 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_20_Left_46 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_21_Left_47 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_22_Left_48 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_23_Left_49 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_24_Left_50 ();
 gf180mcu_fd_sc_mcu9t5v0__endcap PHY_EDGE_ROW_25_Left_51 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_0_52 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_2_53 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_4_54 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_6_55 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_8_56 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_10_57 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_12_58 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_14_59 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_16_60 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_18_61 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_20_62 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_22_63 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_24_64 ();
 gf180mcu_fd_sc_mcu9t5v0__filltie TAP_TAPCELL_ROW_25_65 ();
 gf180mcu_fd_sc_mcu9t5v0__buf_2 input1 (.I(net26),
    .Z(net2));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input2 (.I(spi_miso),
    .Z(net3));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input3 (.I(tx_data[0]),
    .Z(net4));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input4 (.I(tx_data[1]),
    .Z(net5));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input5 (.I(tx_data[2]),
    .Z(net6));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input6 (.I(tx_data[3]),
    .Z(net7));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input7 (.I(tx_data[4]),
    .Z(net8));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input8 (.I(tx_data[5]),
    .Z(net9));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input9 (.I(tx_data[6]),
    .Z(net10));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 input10 (.I(tx_data[7]),
    .Z(net11));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 input11 (.I(tx_valid),
    .Z(net12));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output12 (.I(net13),
    .Z(rx_data[0]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output13 (.I(net14),
    .Z(rx_data[1]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output14 (.I(net15),
    .Z(rx_data[2]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output15 (.I(net16),
    .Z(rx_data[3]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output16 (.I(net17),
    .Z(rx_data[4]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output17 (.I(net18),
    .Z(rx_data[5]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output18 (.I(net19),
    .Z(rx_data[6]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output19 (.I(net20),
    .Z(rx_data[7]));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output20 (.I(net21),
    .Z(rx_valid));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output21 (.I(net22),
    .Z(spi_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output22 (.I(net23),
    .Z(spi_cs_n));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output23 (.I(net24),
    .Z(spi_mosi));
 gf180mcu_fd_sc_mcu9t5v0__dlyb_2 output24 (.I(net25),
    .Z(tx_ready));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_0__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_1__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_2__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 clkbuf_2_3__f_clk (.I(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload0 (.I(clknet_2_0__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__clkinv_3 clkload1 (.I(clknet_2_2__leaf_clk));
 gf180mcu_fd_sc_mcu9t5v0__dlyc_2 hold2 (.I(rst_n),
    .Z(net26));
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_85 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_101 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_0_129 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_0_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_0_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_0_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_0_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_0_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_87 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_89 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_1_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_1_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_1_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_1_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_1_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_2_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_166 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_2_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_2_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_2_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_2_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_3_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_127 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_3_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_3_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_134 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_4_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_4_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_4_212 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_4_228 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_4_236 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_4_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_103 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_5_135 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_5_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_5_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_203 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_5_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_5_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_6_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_90 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_6_111 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_151 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_6_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_6_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_6_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_6_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_84 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_7_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_192 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_7_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_7_213 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_7_221 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_7_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_8_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_116 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_139 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_8_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_8_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_8_211 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_9_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_46 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_113 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_9_169 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_9_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_88 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_95 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_125 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_157 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_10_161 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_10_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_10_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_10_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_80 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_96 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_11_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_11_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_11_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_204 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_11_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_11_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_12_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_82 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_86 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_12_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_12_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_143 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_12_175 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_12_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_12_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_13_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_108 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_13_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_13_155 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_13_171 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_13_206 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_13_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_14_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_107 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_14_123 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_14_142 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_174 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_14_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_14_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_14_238 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_22 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_109 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_117 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_15_121 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_15_140 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_15_172 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_15_188 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_15_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_15_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_4 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_39 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_47 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_51 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_98 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_102 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_16_152 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_16_168 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_16_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_16_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_16_186 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_21 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_17_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_92 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_94 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_17_106 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_122 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_17_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_17_182 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_17_233 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_17_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_42 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_71 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_75 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_110 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_118 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_148 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_150 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_18_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_18_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_198 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_18_229 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_18_237 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_18_241 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_19_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_44 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_60 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_19_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_19_163 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_19_179 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_19_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_19_225 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_18 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_26 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_28 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_63 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_67 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_69 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_93 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_97 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_104 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_20_120 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_124 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_20_126 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_20_144 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_20_180 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_196 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_20_219 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_21_99 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_131 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_21_147 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_21_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_21_184 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_21_200 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_21_223 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_62 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_22_100 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_22_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_170 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_22_197 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_22_232 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_22_240 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_187 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_189 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_23_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_23_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_50 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_58 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_16 FILLER_24_114 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_130 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_146 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_24_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_199 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_24_216 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_24_224 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_24_226 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_74 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_78 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_132 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_149 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_165 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_173 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_177 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_32 FILLER_25_195 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_8 FILLER_25_227 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_4 FILLER_25_235 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_2 FILLER_25_239 ();
 gf180mcu_fd_sc_mcu9t5v0__fill_1 FILLER_25_241 ();
endmodule
