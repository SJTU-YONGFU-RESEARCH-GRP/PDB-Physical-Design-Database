module parameterized_updown_counter (clk,
    enable,
    overflow,
    rst_n,
    up_down,
    count);
 input clk;
 input enable;
 output overflow;
 input rst_n;
 input up_down;
 output [3:0] count;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire _29_;
 wire _30_;
 wire _31_;
 wire _32_;
 wire _33_;
 wire _34_;
 wire _35_;
 wire _36_;
 wire _37_;
 wire _38_;
 wire _39_;
 wire _40_;
 wire _41_;
 wire _42_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 BUF_X1 _43_ (.A(rst_n),
    .Z(_05_));
 BUF_X2 _44_ (.A(enable),
    .Z(_06_));
 OAI21_X1 _45_ (.A(_05_),
    .B1(_06_),
    .B2(net1),
    .ZN(_07_));
 BUF_X4 _46_ (.A(net3),
    .Z(_08_));
 INV_X2 _47_ (.A(_08_),
    .ZN(_09_));
 INV_X1 _48_ (.A(net4),
    .ZN(_10_));
 INV_X1 _49_ (.A(_41_),
    .ZN(_11_));
 BUF_X4 _50_ (.A(up_down),
    .Z(_12_));
 INV_X2 _51_ (.A(_12_),
    .ZN(_13_));
 NOR4_X2 _52_ (.A1(_09_),
    .A2(_10_),
    .A3(_11_),
    .A4(_13_),
    .ZN(_14_));
 AOI21_X1 _53_ (.A(_07_),
    .B1(_14_),
    .B2(_06_),
    .ZN(_15_));
 NAND4_X1 _54_ (.A1(_09_),
    .A2(_10_),
    .A3(_39_),
    .A4(_13_),
    .ZN(_16_));
 NAND2_X1 _55_ (.A1(_06_),
    .A2(_16_),
    .ZN(_17_));
 OAI21_X1 _56_ (.A(_15_),
    .B1(_17_),
    .B2(_37_),
    .ZN(_18_));
 INV_X1 _57_ (.A(_18_),
    .ZN(_00_));
 XNOR2_X1 _58_ (.A(_12_),
    .B(_40_),
    .ZN(_19_));
 MUX2_X1 _59_ (.A(net2),
    .B(_19_),
    .S(_06_),
    .Z(_20_));
 AND2_X1 _60_ (.A1(_05_),
    .A2(_20_),
    .ZN(_01_));
 MUX2_X1 _61_ (.A(_39_),
    .B(_41_),
    .S(_12_),
    .Z(_21_));
 NAND2_X1 _62_ (.A1(_06_),
    .A2(_21_),
    .ZN(_22_));
 XNOR2_X1 _63_ (.A(_08_),
    .B(_22_),
    .ZN(_23_));
 AND2_X1 _64_ (.A1(_05_),
    .A2(_23_),
    .ZN(_02_));
 OAI21_X1 _65_ (.A(_05_),
    .B1(_06_),
    .B2(net4),
    .ZN(_24_));
 INV_X1 _66_ (.A(net2),
    .ZN(_25_));
 NOR4_X1 _67_ (.A1(_09_),
    .A2(net4),
    .A3(_37_),
    .A4(_25_),
    .ZN(_26_));
 OAI21_X1 _68_ (.A(_11_),
    .B1(_37_),
    .B2(_25_),
    .ZN(_27_));
 AOI21_X1 _69_ (.A(_10_),
    .B1(_27_),
    .B2(_08_),
    .ZN(_28_));
 OAI21_X1 _70_ (.A(_12_),
    .B1(_26_),
    .B2(_28_),
    .ZN(_29_));
 NOR3_X1 _71_ (.A1(_08_),
    .A2(net2),
    .A3(net1),
    .ZN(_30_));
 XNOR2_X1 _72_ (.A(_10_),
    .B(_30_),
    .ZN(_31_));
 AOI21_X1 _73_ (.A(_17_),
    .B1(_31_),
    .B2(_13_),
    .ZN(_32_));
 AOI21_X1 _74_ (.A(_24_),
    .B1(_29_),
    .B2(_32_),
    .ZN(_03_));
 OAI221_X1 _75_ (.A(_05_),
    .B1(_17_),
    .B2(_14_),
    .C1(net5),
    .C2(_06_),
    .ZN(_33_));
 INV_X1 _76_ (.A(_33_),
    .ZN(_04_));
 HA_X1 _77_ (.A(_37_),
    .B(_38_),
    .CO(_39_),
    .S(_40_));
 HA_X1 _78_ (.A(net1),
    .B(net2),
    .CO(_41_),
    .S(_42_));
 DFF_X2 \counter_reg[0]$_SDFFE_PN0P_  (.D(_00_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net1),
    .QN(_37_));
 DFF_X2 \counter_reg[1]$_SDFFE_PN0P_  (.D(_01_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net2),
    .QN(_38_));
 DFF_X1 \counter_reg[2]$_SDFFE_PN0P_  (.D(_02_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net3),
    .QN(_36_));
 DFF_X1 \counter_reg[3]$_SDFFE_PN0P_  (.D(_03_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net4),
    .QN(_35_));
 DFF_X1 \overflow_reg$_SDFFE_PN0P_  (.D(_04_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net5),
    .QN(_34_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_51 ();
 BUF_X1 output1 (.A(net1),
    .Z(count[0]));
 BUF_X1 output2 (.A(net2),
    .Z(count[1]));
 BUF_X1 output3 (.A(net3),
    .Z(count[2]));
 BUF_X1 output4 (.A(net4),
    .Z(count[3]));
 BUF_X1 output5 (.A(net5),
    .Z(overflow));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 CLKBUF_X1 clkload0 (.A(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X2 FILLER_0_193 ();
 FILLCELL_X1 FILLER_0_195 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X2 FILLER_1_193 ();
 FILLCELL_X1 FILLER_1_195 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X2 FILLER_2_193 ();
 FILLCELL_X1 FILLER_2_195 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X2 FILLER_3_193 ();
 FILLCELL_X1 FILLER_3_195 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X2 FILLER_4_193 ();
 FILLCELL_X1 FILLER_4_195 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X2 FILLER_5_193 ();
 FILLCELL_X1 FILLER_5_195 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X2 FILLER_6_193 ();
 FILLCELL_X1 FILLER_6_195 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X32 FILLER_7_161 ();
 FILLCELL_X2 FILLER_7_193 ();
 FILLCELL_X1 FILLER_7_195 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X32 FILLER_8_161 ();
 FILLCELL_X2 FILLER_8_193 ();
 FILLCELL_X1 FILLER_8_195 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X16 FILLER_9_65 ();
 FILLCELL_X4 FILLER_9_81 ();
 FILLCELL_X1 FILLER_9_85 ();
 FILLCELL_X32 FILLER_9_93 ();
 FILLCELL_X32 FILLER_9_125 ();
 FILLCELL_X32 FILLER_9_157 ();
 FILLCELL_X4 FILLER_9_189 ();
 FILLCELL_X2 FILLER_9_193 ();
 FILLCELL_X1 FILLER_9_195 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X32 FILLER_10_161 ();
 FILLCELL_X2 FILLER_10_193 ();
 FILLCELL_X1 FILLER_10_195 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X32 FILLER_11_129 ();
 FILLCELL_X32 FILLER_11_161 ();
 FILLCELL_X2 FILLER_11_193 ();
 FILLCELL_X1 FILLER_11_195 ();
 FILLCELL_X2 FILLER_12_1 ();
 FILLCELL_X16 FILLER_12_7 ();
 FILLCELL_X1 FILLER_12_23 ();
 FILLCELL_X4 FILLER_12_31 ();
 FILLCELL_X32 FILLER_12_41 ();
 FILLCELL_X32 FILLER_12_73 ();
 FILLCELL_X32 FILLER_12_105 ();
 FILLCELL_X32 FILLER_12_137 ();
 FILLCELL_X16 FILLER_12_169 ();
 FILLCELL_X8 FILLER_12_185 ();
 FILLCELL_X2 FILLER_12_193 ();
 FILLCELL_X1 FILLER_12_195 ();
 FILLCELL_X2 FILLER_13_1 ();
 FILLCELL_X4 FILLER_13_6 ();
 FILLCELL_X2 FILLER_13_13 ();
 FILLCELL_X1 FILLER_13_15 ();
 FILLCELL_X2 FILLER_13_35 ();
 FILLCELL_X8 FILLER_13_47 ();
 FILLCELL_X4 FILLER_13_65 ();
 FILLCELL_X2 FILLER_13_69 ();
 FILLCELL_X1 FILLER_13_73 ();
 FILLCELL_X32 FILLER_13_84 ();
 FILLCELL_X32 FILLER_13_116 ();
 FILLCELL_X32 FILLER_13_148 ();
 FILLCELL_X16 FILLER_13_180 ();
 FILLCELL_X8 FILLER_14_1 ();
 FILLCELL_X2 FILLER_14_9 ();
 FILLCELL_X1 FILLER_14_11 ();
 FILLCELL_X8 FILLER_14_39 ();
 FILLCELL_X4 FILLER_14_47 ();
 FILLCELL_X2 FILLER_14_51 ();
 FILLCELL_X1 FILLER_14_53 ();
 FILLCELL_X32 FILLER_14_91 ();
 FILLCELL_X32 FILLER_14_123 ();
 FILLCELL_X32 FILLER_14_155 ();
 FILLCELL_X8 FILLER_14_187 ();
 FILLCELL_X1 FILLER_14_195 ();
 FILLCELL_X8 FILLER_15_1 ();
 FILLCELL_X4 FILLER_15_9 ();
 FILLCELL_X2 FILLER_15_13 ();
 FILLCELL_X1 FILLER_15_15 ();
 FILLCELL_X1 FILLER_15_19 ();
 FILLCELL_X2 FILLER_15_22 ();
 FILLCELL_X16 FILLER_15_43 ();
 FILLCELL_X2 FILLER_15_59 ();
 FILLCELL_X32 FILLER_15_86 ();
 FILLCELL_X32 FILLER_15_118 ();
 FILLCELL_X32 FILLER_15_150 ();
 FILLCELL_X8 FILLER_15_182 ();
 FILLCELL_X4 FILLER_15_190 ();
 FILLCELL_X2 FILLER_15_194 ();
 FILLCELL_X4 FILLER_16_1 ();
 FILLCELL_X2 FILLER_16_8 ();
 FILLCELL_X32 FILLER_16_29 ();
 FILLCELL_X1 FILLER_16_61 ();
 FILLCELL_X2 FILLER_16_68 ();
 FILLCELL_X32 FILLER_16_74 ();
 FILLCELL_X32 FILLER_16_106 ();
 FILLCELL_X32 FILLER_16_138 ();
 FILLCELL_X16 FILLER_16_170 ();
 FILLCELL_X8 FILLER_16_186 ();
 FILLCELL_X2 FILLER_16_194 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X8 FILLER_17_33 ();
 FILLCELL_X4 FILLER_17_41 ();
 FILLCELL_X1 FILLER_17_45 ();
 FILLCELL_X8 FILLER_17_51 ();
 FILLCELL_X4 FILLER_17_59 ();
 FILLCELL_X32 FILLER_17_67 ();
 FILLCELL_X32 FILLER_17_99 ();
 FILLCELL_X32 FILLER_17_131 ();
 FILLCELL_X32 FILLER_17_163 ();
 FILLCELL_X1 FILLER_17_195 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_82 ();
 FILLCELL_X32 FILLER_18_114 ();
 FILLCELL_X32 FILLER_18_146 ();
 FILLCELL_X16 FILLER_18_178 ();
 FILLCELL_X2 FILLER_18_194 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X16 FILLER_19_33 ();
 FILLCELL_X8 FILLER_19_49 ();
 FILLCELL_X1 FILLER_19_57 ();
 FILLCELL_X32 FILLER_19_85 ();
 FILLCELL_X32 FILLER_19_117 ();
 FILLCELL_X32 FILLER_19_149 ();
 FILLCELL_X8 FILLER_19_181 ();
 FILLCELL_X4 FILLER_19_189 ();
 FILLCELL_X2 FILLER_19_193 ();
 FILLCELL_X1 FILLER_19_195 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X2 FILLER_20_65 ();
 FILLCELL_X1 FILLER_20_67 ();
 FILLCELL_X32 FILLER_20_73 ();
 FILLCELL_X32 FILLER_20_105 ();
 FILLCELL_X32 FILLER_20_137 ();
 FILLCELL_X16 FILLER_20_169 ();
 FILLCELL_X8 FILLER_20_185 ();
 FILLCELL_X2 FILLER_20_193 ();
 FILLCELL_X1 FILLER_20_195 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X2 FILLER_21_193 ();
 FILLCELL_X1 FILLER_21_195 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X2 FILLER_22_193 ();
 FILLCELL_X1 FILLER_22_195 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X2 FILLER_23_193 ();
 FILLCELL_X1 FILLER_23_195 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X2 FILLER_24_193 ();
 FILLCELL_X1 FILLER_24_195 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X8 FILLER_25_65 ();
 FILLCELL_X4 FILLER_25_73 ();
 FILLCELL_X1 FILLER_25_77 ();
 FILLCELL_X2 FILLER_25_81 ();
 FILLCELL_X32 FILLER_25_86 ();
 FILLCELL_X32 FILLER_25_118 ();
 FILLCELL_X32 FILLER_25_150 ();
 FILLCELL_X8 FILLER_25_182 ();
 FILLCELL_X4 FILLER_25_190 ();
 FILLCELL_X2 FILLER_25_194 ();
endmodule
