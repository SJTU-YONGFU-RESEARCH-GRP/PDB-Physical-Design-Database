module aes_cipher_top (clk,
    done,
    ld,
    rst,
    key,
    text_in,
    text_out);
 input clk;
 output done;
 input ld;
 input rst;
 input [127:0] key;
 input [127:0] text_in;
 output [127:0] text_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire net4044;
 wire net4041;
 wire net3996;
 wire net3986;
 wire net3988;
 wire clknet_leaf_36_clk;
 wire net4094;
 wire net4126;
 wire net3989;
 wire net3978;
 wire net3955;
 wire net3939;
 wire net3938;
 wire _00398_;
 wire net3952;
 wire net4078;
 wire net4134;
 wire net4076;
 wire net4062;
 wire net4115;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00832_;
 wire _00834_;
 wire _00836_;
 wire _00838_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00845_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00859_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00922_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00945_;
 wire _00946_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00960_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire net258;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire net257;
 wire _01018_;
 wire _01019_;
 wire net256;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire net255;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire net254;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire net253;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire net252;
 wire net251;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire net248;
 wire net247;
 wire net246;
 wire net243;
 wire net242;
 wire net241;
 wire net239;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire net238;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire net237;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire net236;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire net235;
 wire net234;
 wire net233;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire net232;
 wire net231;
 wire net230;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire net229;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire net228;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire net227;
 wire net226;
 wire net225;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire net224;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire net223;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire net222;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire net221;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire net220;
 wire _01470_;
 wire _01471_;
 wire net219;
 wire _01473_;
 wire net218;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire net217;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire net216;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire net215;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire net214;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire net213;
 wire _01514_;
 wire _01515_;
 wire net212;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire net211;
 wire _01521_;
 wire net210;
 wire _01523_;
 wire net209;
 wire _01525_;
 wire net208;
 wire _01527_;
 wire _01528_;
 wire net207;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire net206;
 wire net205;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire net203;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire net202;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire net201;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire net200;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire net199;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire net198;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire net197;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire net196;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire net195;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire net194;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire net193;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire net191;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire net189;
 wire net188;
 wire net186;
 wire net184;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire net182;
 wire net181;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire net180;
 wire _01923_;
 wire net179;
 wire net178;
 wire net177;
 wire net176;
 wire _01928_;
 wire _01929_;
 wire net175;
 wire net174;
 wire _01932_;
 wire _01933_;
 wire net173;
 wire _01935_;
 wire _01936_;
 wire net172;
 wire _01938_;
 wire net171;
 wire net170;
 wire _01941_;
 wire net169;
 wire _01943_;
 wire net168;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire net167;
 wire net166;
 wire _01953_;
 wire _01954_;
 wire net165;
 wire net164;
 wire net163;
 wire _01958_;
 wire _01959_;
 wire net162;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire net161;
 wire net160;
 wire net159;
 wire _01967_;
 wire _01968_;
 wire net158;
 wire net157;
 wire _01971_;
 wire net156;
 wire net155;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire net154;
 wire net153;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire net152;
 wire _01986_;
 wire _01987_;
 wire net151;
 wire net150;
 wire _01990_;
 wire _01991_;
 wire net149;
 wire net148;
 wire _01994_;
 wire net147;
 wire _01996_;
 wire _01997_;
 wire net146;
 wire net145;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire net144;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire net143;
 wire _02024_;
 wire _02025_;
 wire net142;
 wire _02027_;
 wire _02028_;
 wire net141;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire net140;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire net139;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire net138;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire net136;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire net135;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire net134;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire net133;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire net132;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire net131;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire net128;
 wire net125;
 wire net124;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire net122;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire net121;
 wire net120;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire net119;
 wire net118;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire net117;
 wire net116;
 wire net115;
 wire _02484_;
 wire net114;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire net113;
 wire net112;
 wire _02492_;
 wire net111;
 wire net110;
 wire _02495_;
 wire net109;
 wire net108;
 wire net107;
 wire _02499_;
 wire net106;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire net105;
 wire net104;
 wire _02507_;
 wire _02508_;
 wire net103;
 wire net102;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire net101;
 wire _02515_;
 wire _02516_;
 wire net100;
 wire net99;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire net98;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire net97;
 wire net96;
 wire net95;
 wire net94;
 wire net93;
 wire net92;
 wire _02532_;
 wire net91;
 wire net90;
 wire net89;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire net88;
 wire net87;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire net86;
 wire net85;
 wire net84;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire net83;
 wire net82;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire net81;
 wire net80;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire net79;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire net78;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire net77;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire net76;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire net75;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire net74;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire net73;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire net71;
 wire _02651_;
 wire net70;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire net69;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire net68;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire net67;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire net65;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire net63;
 wire net62;
 wire net60;
 wire net58;
 wire net57;
 wire net56;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire net54;
 wire net53;
 wire net52;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire net51;
 wire net50;
 wire net49;
 wire _03016_;
 wire _03017_;
 wire net48;
 wire net47;
 wire net46;
 wire _03021_;
 wire net45;
 wire net44;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire net43;
 wire net42;
 wire net41;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire net40;
 wire net38;
 wire net37;
 wire net36;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire net35;
 wire net34;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire net33;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire net32;
 wire net31;
 wire _03066_;
 wire net30;
 wire net29;
 wire _03069_;
 wire _03070_;
 wire net28;
 wire net27;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire net26;
 wire net25;
 wire net24;
 wire _03079_;
 wire _03080_;
 wire net23;
 wire net22;
 wire net21;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire net20;
 wire net19;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire net18;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire net17;
 wire _03101_;
 wire _03102_;
 wire net16;
 wire _03104_;
 wire net15;
 wire net14;
 wire net13;
 wire _03108_;
 wire _03109_;
 wire net12;
 wire net11;
 wire net10;
 wire net9;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire net8;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire net7;
 wire _03123_;
 wire net6;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire net5;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire net4;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire net3;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire net2;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire net1;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire net4145;
 wire net4144;
 wire net4143;
 wire net4142;
 wire _03574_;
 wire _03575_;
 wire clknet_leaf_34_clk;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire clknet_leaf_35_clk;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire clknet_leaf_33_clk;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_42_clk;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire net4128;
 wire net4129;
 wire net4123;
 wire net4130;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire net4107;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire net4110;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire net4091;
 wire net4090;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire net4093;
 wire _03639_;
 wire net4083;
 wire net4099;
 wire net4082;
 wire net4087;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire net4081;
 wire net4074;
 wire net4073;
 wire net4071;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire net4072;
 wire _03658_;
 wire net4127;
 wire net4067;
 wire net4064;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire net4077;
 wire net4066;
 wire net4063;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire net4118;
 wire net4102;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire net4116;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire net4069;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire net4150;
 wire net4207;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire net4117;
 wire _03704_;
 wire net4070;
 wire clknet_leaf_44_clk;
 wire net4121;
 wire net4059;
 wire net4056;
 wire net4057;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire net4055;
 wire net4048;
 wire net4035;
 wire net4037;
 wire net4038;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire net4032;
 wire net4034;
 wire net3999;
 wire net3995;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire net3994;
 wire net3997;
 wire net4002;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire net3985;
 wire net3981;
 wire net3980;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire net3983;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire net4012;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire net3982;
 wire net3974;
 wire _03787_;
 wire net3969;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire net3958;
 wire net3959;
 wire net3946;
 wire _03796_;
 wire net3947;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire net3948;
 wire net3943;
 wire net3944;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire net3945;
 wire net3937;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire net3932;
 wire _03826_;
 wire net3929;
 wire net3967;
 wire _03829_;
 wire clknet_leaf_57_clk;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire clknet_leaf_58_clk;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire net3927;
 wire _03851_;
 wire _03852_;
 wire net3928;
 wire net3930;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire clknet_leaf_59_clk;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire net3918;
 wire _03870_;
 wire _03871_;
 wire net3919;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire net3920;
 wire _03883_;
 wire _03884_;
 wire net3921;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire net3912;
 wire _03898_;
 wire _03899_;
 wire net3917;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire net3907;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire net3904;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire net3903;
 wire net3916;
 wire net3902;
 wire net3913;
 wire net3896;
 wire net3882;
 wire net388;
 wire net3885;
 wire net3893;
 wire net3891;
 wire _03942_;
 wire net3871;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire net3877;
 wire net3878;
 wire _03949_;
 wire _03950_;
 wire net3567;
 wire _03952_;
 wire _03953_;
 wire _03955_;
 wire net3573;
 wire _03957_;
 wire _03958_;
 wire _03960_;
 wire _03961_;
 wire net3572;
 wire _03964_;
 wire net3569;
 wire _03966_;
 wire _03967_;
 wire _03969_;
 wire net3706;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03977_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire net3744;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire net3824;
 wire net3820;
 wire _03991_;
 wire _03992_;
 wire _03995_;
 wire _03996_;
 wire clknet_leaf_19_clk;
 wire _03998_;
 wire clknet_leaf_20_clk;
 wire net4231;
 wire _04001_;
 wire _04002_;
 wire net4235;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire clknet_leaf_5_clk;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire net4225;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire net4224;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire net3560;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire net4218;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire net4222;
 wire _04068_;
 wire _04069_;
 wire clknet_leaf_21_clk;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire net4220;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire clknet_leaf_6_clk;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire clknet_leaf_8_clk;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire net4204;
 wire net4227;
 wire net4197;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04415_;
 wire _04416_;
 wire net4194;
 wire _04419_;
 wire clknet_leaf_9_clk;
 wire net4185;
 wire _04423_;
 wire net4181;
 wire net4182;
 wire net4180;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire net4178;
 wire _04432_;
 wire net4188;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire net4173;
 wire _04438_;
 wire net4172;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire net4164;
 wire _04447_;
 wire _04448_;
 wire net4175;
 wire _04450_;
 wire net4161;
 wire _04452_;
 wire _04453_;
 wire net4162;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire net4163;
 wire net4154;
 wire net4153;
 wire net4149;
 wire net4148;
 wire _04463_;
 wire _04464_;
 wire clknet_leaf_28_clk;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire net4139;
 wire net4141;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire net4152;
 wire _04480_;
 wire net4157;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire clknet_leaf_29_clk;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire clknet_leaf_25_clk;
 wire _04496_;
 wire _04497_;
 wire net4177;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire net4140;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire net4131;
 wire net4133;
 wire _04510_;
 wire clknet_leaf_30_clk;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire net4109;
 wire clknet_leaf_43_clk;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire net4135;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire net4113;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire net4106;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire net4124;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire net4104;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire net4179;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire net4103;
 wire net4097;
 wire net4105;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04904_;
 wire net4095;
 wire _04907_;
 wire _04908_;
 wire net4092;
 wire net4096;
 wire _04911_;
 wire _04912_;
 wire _04914_;
 wire _04915_;
 wire _04917_;
 wire net4098;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04928_;
 wire _04929_;
 wire _04931_;
 wire _04933_;
 wire net3703;
 wire _04935_;
 wire _04937_;
 wire net4089;
 wire _04939_;
 wire _04940_;
 wire net4086;
 wire _04942_;
 wire _04943_;
 wire net4084;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire net4228;
 wire net4079;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire net4088;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire net3702;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire net3578;
 wire _04999_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05024_;
 wire _05025_;
 wire net4080;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire net3579;
 wire _05055_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire net4229;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire net3582;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire net3698;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05107_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire net3581;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05388_;
 wire net3588;
 wire _05393_;
 wire _05394_;
 wire net3584;
 wire _05396_;
 wire _05398_;
 wire net3696;
 wire _05401_;
 wire net3580;
 wire _05404_;
 wire _05407_;
 wire net3587;
 wire _05409_;
 wire _05411_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05418_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire net3695;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire net3590;
 wire _05433_;
 wire _05437_;
 wire _05438_;
 wire net4238;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire net4239;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire net3591;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire net3592;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire net4240;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05874_;
 wire _05875_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire net3623;
 wire net3619;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05893_;
 wire _05895_;
 wire _05896_;
 wire net3594;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire net3595;
 wire net3617;
 wire net3614;
 wire net3597;
 wire net4075;
 wire _05911_;
 wire net3596;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05921_;
 wire net3599;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05927_;
 wire net3600;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05940_;
 wire net3605;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05947_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05953_;
 wire _05954_;
 wire net3604;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05960_;
 wire _05962_;
 wire _05963_;
 wire net3606;
 wire _05965_;
 wire _05966_;
 wire net3607;
 wire net3609;
 wire _05970_;
 wire _05971_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire net3611;
 wire _05982_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05991_;
 wire _05992_;
 wire _05994_;
 wire _05995_;
 wire _05997_;
 wire _05998_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire net3610;
 wire _06008_;
 wire _06009_;
 wire net3608;
 wire _06011_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06019_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06026_;
 wire _06028_;
 wire _06029_;
 wire net4119;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire clknet_leaf_14_clk;
 wire _06037_;
 wire _06038_;
 wire clknet_leaf_15_clk;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire net3612;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire net4058;
 wire _06053_;
 wire net4060;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire clknet_leaf_12_clk;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire clknet_leaf_16_clk;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire clknet_leaf_17_clk;
 wire _06072_;
 wire net4049;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire net4050;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire net4045;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire net4042;
 wire _06097_;
 wire _06098_;
 wire net4039;
 wire net4043;
 wire net4036;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire net4120;
 wire _06122_;
 wire net4033;
 wire _06124_;
 wire net4046;
 wire clknet_leaf_48_clk;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire net4017;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire net4021;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire net4013;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire net4014;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire net4011;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire net4005;
 wire net4001;
 wire _06477_;
 wire net4006;
 wire _06479_;
 wire net4009;
 wire _06481_;
 wire _06482_;
 wire net4051;
 wire net3998;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire net4000;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire net4010;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire net3991;
 wire _06505_;
 wire net3992;
 wire net4025;
 wire net3984;
 wire net4028;
 wire net3993;
 wire clknet_leaf_55_clk;
 wire _06512_;
 wire net3970;
 wire _06514_;
 wire net3962;
 wire net3976;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire net3960;
 wire net3957;
 wire net3956;
 wire net3953;
 wire net3954;
 wire net3940;
 wire _06527_;
 wire _06528_;
 wire net3935;
 wire _06530_;
 wire _06531_;
 wire net3941;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire net3966;
 wire net3964;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire net3931;
 wire net3933;
 wire net3951;
 wire net3910;
 wire net3922;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire net3905;
 wire net3914;
 wire _06553_;
 wire clknet_leaf_60_clk;
 wire net3899;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire clknet_leaf_61_clk;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire clknet_leaf_62_clk;
 wire _06564_;
 wire _06565_;
 wire net3895;
 wire net3894;
 wire _06568_;
 wire _06569_;
 wire net3900;
 wire net3890;
 wire net3886;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire net3883;
 wire net3906;
 wire net3924;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire net3879;
 wire _06583_;
 wire net3870;
 wire net3881;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire net3909;
 wire net3869;
 wire net3880;
 wire _06594_;
 wire clknet_leaf_66_clk;
 wire _06596_;
 wire net3865;
 wire net3867;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire net3868;
 wire _06605_;
 wire net3861;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire net3853;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire net3864;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire net3856;
 wire net3875;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire net3866;
 wire net3852;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire net3850;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire net3840;
 wire net3834;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire net3832;
 wire _06668_;
 wire net3835;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire net3827;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire net3836;
 wire _06731_;
 wire net3826;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire net3841;
 wire net3833;
 wire net3825;
 wire _06744_;
 wire net3805;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire net3828;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire net3830;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire net3807;
 wire net3803;
 wire _07074_;
 wire _07075_;
 wire net3804;
 wire net3814;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire net3799;
 wire _07084_;
 wire net3797;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire net3798;
 wire net3781;
 wire net3782;
 wire _07094_;
 wire net3765;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire net3771;
 wire net3772;
 wire net3755;
 wire net3752;
 wire net3745;
 wire net3746;
 wire clknet_3_7_0_clk;
 wire _07108_;
 wire net3741;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire net3732;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire net3742;
 wire net3729;
 wire _07126_;
 wire net3727;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire net3733;
 wire net3743;
 wire net3723;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire net3717;
 wire net3721;
 wire net3718;
 wire net3739;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire net3749;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire net3728;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire net3725;
 wire net389;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire net3751;
 wire net3750;
 wire net3748;
 wire _07173_;
 wire _07174_;
 wire net3756;
 wire net3757;
 wire net3758;
 wire _07178_;
 wire net3759;
 wire net3773;
 wire net3769;
 wire _07182_;
 wire clknet_leaf_89_clk;
 wire net3785;
 wire clknet_leaf_90_clk;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire net3777;
 wire net3783;
 wire _07193_;
 wire _07194_;
 wire clknet_leaf_83_clk;
 wire _07196_;
 wire _07197_;
 wire clknet_leaf_82_clk;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire net3784;
 wire net3806;
 wire clknet_leaf_70_clk;
 wire _07210_;
 wire net3844;
 wire _07212_;
 wire _07213_;
 wire net3872;
 wire _07215_;
 wire _07216_;
 wire net3714;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire net3837;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire net3838;
 wire _07230_;
 wire _07231_;
 wire net3842;
 wire net3854;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire net3843;
 wire _07239_;
 wire _07240_;
 wire net3858;
 wire clknet_leaf_67_clk;
 wire net3884;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire net3889;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire net3897;
 wire _07256_;
 wire net3898;
 wire clknet_leaf_64_clk;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire clknet_leaf_65_clk;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire clknet_leaf_63_clk;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire net3977;
 wire _07295_;
 wire _07296_;
 wire net3963;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire net3968;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire net4029;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire clknet_leaf_56_clk;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire net4019;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_51_clk;
 wire _07657_;
 wire net4024;
 wire net4007;
 wire _07660_;
 wire clknet_leaf_47_clk;
 wire net4015;
 wire net3715;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire net4018;
 wire _07670_;
 wire net4026;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire clknet_leaf_45_clk;
 wire _07678_;
 wire clknet_leaf_46_clk;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire net4040;
 wire net4047;
 wire net3613;
 wire _07692_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire net3625;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07712_;
 wire _07713_;
 wire net3694;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire net3693;
 wire _07723_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire net3692;
 wire net3626;
 wire _07732_;
 wire net3627;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire net3628;
 wire _07740_;
 wire net3629;
 wire net3630;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07749_;
 wire _07751_;
 wire net3686;
 wire net3673;
 wire _07754_;
 wire _07755_;
 wire net3672;
 wire _07758_;
 wire net3633;
 wire net3631;
 wire _07761_;
 wire net3632;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire net3639;
 wire _07768_;
 wire _07769_;
 wire _07771_;
 wire net3634;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire net3636;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire net3638;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire net3671;
 wire _07801_;
 wire _07803_;
 wire net3645;
 wire _07805_;
 wire net3648;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire net3654;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire net3651;
 wire _07843_;
 wire net3650;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire net3652;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire net3656;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire net3658;
 wire net3660;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08268_;
 wire _08270_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire net3661;
 wire _08289_;
 wire _08290_;
 wire net3662;
 wire _08293_;
 wire _08295_;
 wire net3665;
 wire _08298_;
 wire net3666;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08312_;
 wire _08314_;
 wire net3679;
 wire _08316_;
 wire net3682;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire net3680;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire net3681;
 wire _08338_;
 wire net405;
 wire net406;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire net3685;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire net3688;
 wire net3708;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08367_;
 wire _08368_;
 wire net3699;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08380_;
 wire _08381_;
 wire net3701;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire net3697;
 wire _08398_;
 wire _08400_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire net3691;
 wire _08415_;
 wire net3687;
 wire _08417_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08436_;
 wire _08437_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire net3683;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire net3677;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire net3678;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire net407;
 wire net3669;
 wire net3668;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08840_;
 wire net3670;
 wire _08842_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08851_;
 wire net3655;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire net3642;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08862_;
 wire _08863_;
 wire net3641;
 wire net3640;
 wire net3659;
 wire net3643;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire net3647;
 wire net3664;
 wire _08873_;
 wire _08874_;
 wire net3649;
 wire _08876_;
 wire net3663;
 wire _08878_;
 wire net3644;
 wire net3646;
 wire net3657;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08898_;
 wire _08899_;
 wire net3684;
 wire _08901_;
 wire _08902_;
 wire _08904_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire net3689;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08980_;
 wire _08981_;
 wire _08982_;
 wire _08983_;
 wire _08984_;
 wire _08985_;
 wire net3707;
 wire _08987_;
 wire net3768;
 wire net3794;
 wire net409;
 wire _08991_;
 wire _08992_;
 wire net3690;
 wire _08994_;
 wire _08995_;
 wire _08998_;
 wire net3700;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09004_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire _09035_;
 wire _09036_;
 wire _09037_;
 wire _09038_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire net3705;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire net3709;
 wire _09105_;
 wire _09106_;
 wire net3767;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire _09144_;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire net403;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire net3637;
 wire net402;
 wire net401;
 wire net3761;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire net399;
 wire _09408_;
 wire net398;
 wire _09410_;
 wire net396;
 wire _09412_;
 wire net397;
 wire net395;
 wire _09415_;
 wire net394;
 wire _09417_;
 wire _09418_;
 wire net393;
 wire _09420_;
 wire _09421_;
 wire net3722;
 wire net3735;
 wire _09424_;
 wire net3713;
 wire net3760;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire net3716;
 wire net3711;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire net3712;
 wire _09440_;
 wire net3720;
 wire net3719;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire net3730;
 wire _09448_;
 wire net3731;
 wire net3734;
 wire _09451_;
 wire _09452_;
 wire net3726;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire net391;
 wire _09459_;
 wire _09460_;
 wire net392;
 wire _09462_;
 wire net3740;
 wire net3753;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire net3724;
 wire net3754;
 wire _09470_;
 wire net3736;
 wire net3737;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire net390;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire net3747;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire clknet_3_4_0_clk;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire net3774;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire net3762;
 wire _09527_;
 wire net3766;
 wire net3775;
 wire net3776;
 wire _09531_;
 wire _09532_;
 wire net3770;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire clknet_leaf_91_clk;
 wire _09539_;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire clknet_3_1_0_clk;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire clknet_3_3_0_clk;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire clknet_leaf_88_clk;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire net3778;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire net3779;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire net3780;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire _09714_;
 wire _09715_;
 wire _09716_;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire _09720_;
 wire _09721_;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire _09737_;
 wire _09738_;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire _09883_;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire _09906_;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire clknet_leaf_85_clk;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire clknet_leaf_87_clk;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire net3787;
 wire clknet_leaf_80_clk;
 wire net3790;
 wire net3791;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire clknet_leaf_78_clk;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire net3815;
 wire _09952_;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire net3796;
 wire net3816;
 wire net3817;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire net3839;
 wire net3823;
 wire _09975_;
 wire net3822;
 wire _09977_;
 wire _09978_;
 wire net3942;
 wire net3800;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire net3801;
 wire _09992_;
 wire net3808;
 wire _09994_;
 wire net3809;
 wire net3810;
 wire _09997_;
 wire _09998_;
 wire net3811;
 wire net3812;
 wire net3949;
 wire _10002_;
 wire net3950;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire net3821;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire clknet_leaf_71_clk;
 wire _10012_;
 wire clknet_leaf_72_clk;
 wire _10014_;
 wire clknet_leaf_77_clk;
 wire _10016_;
 wire _10017_;
 wire net3829;
 wire _10019_;
 wire _10020_;
 wire net3831;
 wire _10023_;
 wire net3845;
 wire _10026_;
 wire net3624;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10036_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10043_;
 wire _10045_;
 wire _10046_;
 wire net3616;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10053_;
 wire _10054_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire net3601;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10076_;
 wire _10077_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire net3598;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire _10433_;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire _10440_;
 wire _10441_;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire _10474_;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10509_;
 wire net3615;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire net3620;
 wire net3618;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire net3622;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire net3621;
 wire _10552_;
 wire _10554_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire net3936;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire net3846;
 wire _10567_;
 wire net3847;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire net3873;
 wire net3862;
 wire net3926;
 wire net3934;
 wire _10579_;
 wire _10580_;
 wire net3848;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire net3874;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire net3851;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire net3849;
 wire net3876;
 wire net3855;
 wire _10602_;
 wire net3859;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire _10608_;
 wire _10609_;
 wire net3589;
 wire _10611_;
 wire net3925;
 wire _10614_;
 wire net3586;
 wire net3863;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire net3585;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire net3583;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10667_;
 wire _10668_;
 wire net3577;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10703_;
 wire clknet_leaf_68_clk;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire clknet_leaf_69_clk;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire net3575;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire net3795;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire net3565;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire net3819;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire net3704;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire net3571;
 wire net3566;
 wire net3563;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire net3818;
 wire net4138;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire net4137;
 wire _11105_;
 wire clknet_leaf_10_clk;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire net4136;
 wire net4114;
 wire _11112_;
 wire net4125;
 wire _11114_;
 wire _11115_;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire clknet_leaf_31_clk;
 wire _11124_;
 wire _11125_;
 wire net4132;
 wire _11127_;
 wire _11128_;
 wire net4108;
 wire _11130_;
 wire _11131_;
 wire net3574;
 wire net4101;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire net3576;
 wire _11144_;
 wire _11145_;
 wire clknet_leaf_11_clk;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_53_clk;
 wire _11152_;
 wire _11153_;
 wire net4016;
 wire net4004;
 wire _11156_;
 wire net4023;
 wire net3990;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire _11166_;
 wire _11167_;
 wire net3975;
 wire _11169_;
 wire _11170_;
 wire net3961;
 wire _11172_;
 wire net4030;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire net3915;
 wire net3892;
 wire net3923;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire net3857;
 wire _11188_;
 wire net3813;
 wire _11190_;
 wire _11191_;
 wire clknet_leaf_81_clk;
 wire _11193_;
 wire _11194_;
 wire net3793;
 wire clknet_3_6_0_clk;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire net3738;
 wire _11201_;
 wire _11202_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11673_;
 wire _11676_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11684_;
 wire _11686_;
 wire _11688_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11696_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11719_;
 wire _11723_;
 wire _11726_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11740_;
 wire _11743_;
 wire _11744_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11761_;
 wire _11762_;
 wire _11765_;
 wire _11766_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11789_;
 wire _11790_;
 wire _11792_;
 wire _11793_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire net3908;
 wire net3901;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire net3911;
 wire net4112;
 wire net4209;
 wire net4068;
 wire net4065;
 wire net4208;
 wire net4061;
 wire net4111;
 wire net4122;
 wire net4100;
 wire net4085;
 wire net3979;
 wire net3973;
 wire net3971;
 wire net3593;
 wire net4054;
 wire net3603;
 wire net3987;
 wire net3888;
 wire net4003;
 wire net4008;
 wire net3972;
 wire net4022;
 wire net3764;
 wire net3965;
 wire net3802;
 wire net3788;
 wire clknet_3_5_0_clk;
 wire net3763;
 wire net3653;
 wire net4020;
 wire net4027;
 wire net3676;
 wire net410;
 wire net3675;
 wire net3674;
 wire net3667;
 wire net408;
 wire net3635;
 wire clknet_3_2_0_clk;
 wire net3710;
 wire net404;
 wire clknet_leaf_79_clk;
 wire net3602;
 wire clknet_leaf_86_clk;
 wire net3786;
 wire net3792;
 wire net3789;
 wire net3860;
 wire net3568;
 wire net3570;
 wire net3564;
 wire net244;
 wire net204;
 wire net250;
 wire net249;
 wire net240;
 wire net245;
 wire net185;
 wire net137;
 wire net192;
 wire net190;
 wire net183;
 wire net187;
 wire net126;
 wire net72;
 wire net130;
 wire net129;
 wire net123;
 wire net127;
 wire net59;
 wire net39;
 wire net66;
 wire net64;
 wire net55;
 wire net61;
 wire \dcnt[0] ;
 wire \dcnt[1] ;
 wire \dcnt[2] ;
 wire \dcnt[3] ;
 wire net259;
 wire ld_r;
 wire \sa00_sr[0] ;
 wire \sa00_sr[1] ;
 wire \sa00_sr[2] ;
 wire \sa00_sr[3] ;
 wire \sa00_sr[4] ;
 wire \sa00_sr[5] ;
 wire \sa00_sr[6] ;
 wire \sa00_sr[7] ;
 wire \sa01_sr[0] ;
 wire \sa01_sr[1] ;
 wire \sa01_sr[2] ;
 wire \sa01_sr[3] ;
 wire \sa01_sr[4] ;
 wire \sa01_sr[5] ;
 wire \sa01_sr[6] ;
 wire \sa01_sr[7] ;
 wire \sa02_sr[0] ;
 wire \sa02_sr[1] ;
 wire \sa02_sr[2] ;
 wire \sa02_sr[3] ;
 wire \sa02_sr[4] ;
 wire \sa02_sr[5] ;
 wire \sa02_sr[6] ;
 wire \sa02_sr[7] ;
 wire \sa03_sr[0] ;
 wire \sa03_sr[1] ;
 wire \sa03_sr[2] ;
 wire \sa03_sr[3] ;
 wire \sa03_sr[4] ;
 wire \sa03_sr[5] ;
 wire \sa03_sr[6] ;
 wire \sa03_sr[7] ;
 wire \sa10_sr[0] ;
 wire \sa10_sr[1] ;
 wire \sa10_sr[2] ;
 wire \sa10_sr[3] ;
 wire \sa10_sr[4] ;
 wire \sa10_sr[5] ;
 wire \sa10_sr[6] ;
 wire \sa10_sr[7] ;
 wire \sa10_sub[0] ;
 wire \sa10_sub[1] ;
 wire \sa10_sub[2] ;
 wire \sa10_sub[3] ;
 wire \sa10_sub[4] ;
 wire \sa10_sub[5] ;
 wire \sa10_sub[6] ;
 wire \sa10_sub[7] ;
 wire \sa11_sr[0] ;
 wire \sa11_sr[1] ;
 wire \sa11_sr[2] ;
 wire \sa11_sr[3] ;
 wire \sa11_sr[4] ;
 wire \sa11_sr[5] ;
 wire \sa11_sr[6] ;
 wire \sa11_sr[7] ;
 wire \sa12_sr[0] ;
 wire \sa12_sr[1] ;
 wire \sa12_sr[2] ;
 wire \sa12_sr[3] ;
 wire \sa12_sr[4] ;
 wire \sa12_sr[5] ;
 wire \sa12_sr[6] ;
 wire \sa12_sr[7] ;
 wire \sa20_sr[0] ;
 wire \sa20_sr[1] ;
 wire \sa20_sr[2] ;
 wire \sa20_sr[3] ;
 wire \sa20_sr[4] ;
 wire \sa20_sr[5] ;
 wire \sa20_sr[6] ;
 wire \sa20_sr[7] ;
 wire \sa20_sub[0] ;
 wire \sa20_sub[1] ;
 wire \sa20_sub[2] ;
 wire \sa20_sub[3] ;
 wire \sa20_sub[4] ;
 wire \sa20_sub[5] ;
 wire \sa20_sub[6] ;
 wire \sa20_sub[7] ;
 wire \sa21_sr[0] ;
 wire \sa21_sr[1] ;
 wire \sa21_sr[2] ;
 wire \sa21_sr[3] ;
 wire \sa21_sr[4] ;
 wire \sa21_sr[5] ;
 wire \sa21_sr[6] ;
 wire \sa21_sr[7] ;
 wire \sa21_sub[0] ;
 wire \sa21_sub[1] ;
 wire \sa21_sub[2] ;
 wire \sa21_sub[3] ;
 wire \sa21_sub[4] ;
 wire \sa21_sub[5] ;
 wire \sa21_sub[6] ;
 wire \sa21_sub[7] ;
 wire \sa30_sr[0] ;
 wire \sa30_sr[1] ;
 wire \sa30_sr[2] ;
 wire \sa30_sr[3] ;
 wire \sa30_sr[4] ;
 wire \sa30_sr[5] ;
 wire \sa30_sr[6] ;
 wire \sa30_sr[7] ;
 wire \sa30_sub[0] ;
 wire \sa30_sub[1] ;
 wire \sa30_sub[2] ;
 wire \sa30_sub[3] ;
 wire \sa30_sub[4] ;
 wire \sa30_sub[5] ;
 wire \sa30_sub[6] ;
 wire \sa30_sub[7] ;
 wire \sa31_sub[0] ;
 wire \sa31_sub[1] ;
 wire \sa31_sub[2] ;
 wire \sa31_sub[3] ;
 wire \sa31_sub[4] ;
 wire \sa31_sub[5] ;
 wire \sa31_sub[6] ;
 wire \sa31_sub[7] ;
 wire \sa32_sub[0] ;
 wire \sa32_sub[1] ;
 wire \sa32_sub[2] ;
 wire \sa32_sub[3] ;
 wire \sa32_sub[4] ;
 wire \sa32_sub[5] ;
 wire \sa32_sub[6] ;
 wire \sa32_sub[7] ;
 wire \text_in_r[0] ;
 wire \text_in_r[100] ;
 wire \text_in_r[101] ;
 wire \text_in_r[102] ;
 wire \text_in_r[103] ;
 wire \text_in_r[104] ;
 wire \text_in_r[105] ;
 wire \text_in_r[106] ;
 wire \text_in_r[107] ;
 wire \text_in_r[108] ;
 wire \text_in_r[109] ;
 wire \text_in_r[10] ;
 wire \text_in_r[110] ;
 wire \text_in_r[111] ;
 wire \text_in_r[112] ;
 wire \text_in_r[113] ;
 wire \text_in_r[114] ;
 wire \text_in_r[115] ;
 wire \text_in_r[116] ;
 wire \text_in_r[117] ;
 wire \text_in_r[118] ;
 wire \text_in_r[119] ;
 wire \text_in_r[11] ;
 wire \text_in_r[120] ;
 wire \text_in_r[121] ;
 wire \text_in_r[122] ;
 wire \text_in_r[123] ;
 wire \text_in_r[124] ;
 wire \text_in_r[125] ;
 wire \text_in_r[126] ;
 wire \text_in_r[127] ;
 wire \text_in_r[12] ;
 wire \text_in_r[13] ;
 wire \text_in_r[14] ;
 wire \text_in_r[15] ;
 wire \text_in_r[16] ;
 wire \text_in_r[17] ;
 wire \text_in_r[18] ;
 wire \text_in_r[19] ;
 wire \text_in_r[1] ;
 wire \text_in_r[20] ;
 wire \text_in_r[21] ;
 wire \text_in_r[22] ;
 wire \text_in_r[23] ;
 wire \text_in_r[24] ;
 wire \text_in_r[25] ;
 wire \text_in_r[26] ;
 wire \text_in_r[27] ;
 wire \text_in_r[28] ;
 wire \text_in_r[29] ;
 wire \text_in_r[2] ;
 wire \text_in_r[30] ;
 wire \text_in_r[31] ;
 wire \text_in_r[32] ;
 wire \text_in_r[33] ;
 wire \text_in_r[34] ;
 wire \text_in_r[35] ;
 wire \text_in_r[36] ;
 wire \text_in_r[37] ;
 wire \text_in_r[38] ;
 wire \text_in_r[39] ;
 wire \text_in_r[3] ;
 wire \text_in_r[40] ;
 wire \text_in_r[41] ;
 wire \text_in_r[42] ;
 wire \text_in_r[43] ;
 wire \text_in_r[44] ;
 wire \text_in_r[45] ;
 wire \text_in_r[46] ;
 wire \text_in_r[47] ;
 wire \text_in_r[48] ;
 wire \text_in_r[49] ;
 wire \text_in_r[4] ;
 wire \text_in_r[50] ;
 wire \text_in_r[51] ;
 wire \text_in_r[52] ;
 wire \text_in_r[53] ;
 wire \text_in_r[54] ;
 wire \text_in_r[55] ;
 wire \text_in_r[56] ;
 wire \text_in_r[57] ;
 wire \text_in_r[58] ;
 wire \text_in_r[59] ;
 wire \text_in_r[5] ;
 wire \text_in_r[60] ;
 wire \text_in_r[61] ;
 wire \text_in_r[62] ;
 wire \text_in_r[63] ;
 wire \text_in_r[64] ;
 wire \text_in_r[65] ;
 wire \text_in_r[66] ;
 wire \text_in_r[67] ;
 wire \text_in_r[68] ;
 wire \text_in_r[69] ;
 wire \text_in_r[6] ;
 wire \text_in_r[70] ;
 wire \text_in_r[71] ;
 wire \text_in_r[72] ;
 wire \text_in_r[73] ;
 wire \text_in_r[74] ;
 wire \text_in_r[75] ;
 wire \text_in_r[76] ;
 wire \text_in_r[77] ;
 wire \text_in_r[78] ;
 wire \text_in_r[79] ;
 wire \text_in_r[7] ;
 wire \text_in_r[80] ;
 wire \text_in_r[81] ;
 wire \text_in_r[82] ;
 wire \text_in_r[83] ;
 wire \text_in_r[84] ;
 wire \text_in_r[85] ;
 wire \text_in_r[86] ;
 wire \text_in_r[87] ;
 wire \text_in_r[88] ;
 wire \text_in_r[89] ;
 wire \text_in_r[8] ;
 wire \text_in_r[90] ;
 wire \text_in_r[91] ;
 wire \text_in_r[92] ;
 wire \text_in_r[93] ;
 wire \text_in_r[94] ;
 wire \text_in_r[95] ;
 wire \text_in_r[96] ;
 wire \text_in_r[97] ;
 wire \text_in_r[98] ;
 wire \text_in_r[99] ;
 wire \text_in_r[9] ;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire \u0.r0.out[24] ;
 wire \u0.r0.out[25] ;
 wire \u0.r0.out[26] ;
 wire \u0.r0.out[27] ;
 wire \u0.r0.out[28] ;
 wire \u0.r0.out[29] ;
 wire \u0.r0.out[30] ;
 wire \u0.r0.out[31] ;
 wire \u0.r0.rcnt[0] ;
 wire \u0.r0.rcnt[1] ;
 wire \u0.r0.rcnt[2] ;
 wire \u0.r0.rcnt[3] ;
 wire \u0.r0.rcnt_next[0] ;
 wire \u0.r0.rcnt_next[1] ;
 wire \u0.subword[0] ;
 wire \u0.subword[10] ;
 wire \u0.subword[11] ;
 wire \u0.subword[12] ;
 wire \u0.subword[13] ;
 wire \u0.subword[14] ;
 wire \u0.subword[15] ;
 wire \u0.subword[16] ;
 wire \u0.subword[17] ;
 wire \u0.subword[18] ;
 wire \u0.subword[19] ;
 wire \u0.subword[1] ;
 wire \u0.subword[20] ;
 wire \u0.subword[21] ;
 wire \u0.subword[22] ;
 wire \u0.subword[23] ;
 wire \u0.subword[24] ;
 wire \u0.subword[25] ;
 wire \u0.subword[26] ;
 wire \u0.subword[27] ;
 wire \u0.subword[28] ;
 wire \u0.subword[29] ;
 wire \u0.subword[2] ;
 wire \u0.subword[30] ;
 wire \u0.subword[31] ;
 wire \u0.subword[3] ;
 wire \u0.subword[4] ;
 wire \u0.subword[5] ;
 wire \u0.subword[6] ;
 wire \u0.subword[7] ;
 wire \u0.subword[8] ;
 wire \u0.subword[9] ;
 wire \u0.tmp_w[0] ;
 wire \u0.tmp_w[10] ;
 wire \u0.tmp_w[11] ;
 wire \u0.tmp_w[12] ;
 wire \u0.tmp_w[13] ;
 wire \u0.tmp_w[14] ;
 wire \u0.tmp_w[15] ;
 wire \u0.tmp_w[16] ;
 wire \u0.tmp_w[17] ;
 wire \u0.tmp_w[18] ;
 wire \u0.tmp_w[19] ;
 wire \u0.tmp_w[1] ;
 wire \u0.tmp_w[20] ;
 wire \u0.tmp_w[21] ;
 wire \u0.tmp_w[22] ;
 wire \u0.tmp_w[23] ;
 wire \u0.tmp_w[24] ;
 wire \u0.tmp_w[25] ;
 wire \u0.tmp_w[26] ;
 wire \u0.tmp_w[27] ;
 wire \u0.tmp_w[28] ;
 wire \u0.tmp_w[29] ;
 wire \u0.tmp_w[2] ;
 wire \u0.tmp_w[30] ;
 wire \u0.tmp_w[31] ;
 wire \u0.tmp_w[3] ;
 wire \u0.tmp_w[4] ;
 wire \u0.tmp_w[5] ;
 wire \u0.tmp_w[6] ;
 wire \u0.tmp_w[7] ;
 wire \u0.tmp_w[8] ;
 wire \u0.tmp_w[9] ;
 wire \u0.w[0][0] ;
 wire \u0.w[0][10] ;
 wire \u0.w[0][11] ;
 wire \u0.w[0][12] ;
 wire \u0.w[0][13] ;
 wire \u0.w[0][14] ;
 wire \u0.w[0][15] ;
 wire \u0.w[0][16] ;
 wire \u0.w[0][17] ;
 wire \u0.w[0][18] ;
 wire \u0.w[0][19] ;
 wire \u0.w[0][1] ;
 wire \u0.w[0][20] ;
 wire \u0.w[0][21] ;
 wire \u0.w[0][22] ;
 wire \u0.w[0][23] ;
 wire \u0.w[0][24] ;
 wire \u0.w[0][25] ;
 wire \u0.w[0][26] ;
 wire \u0.w[0][27] ;
 wire \u0.w[0][28] ;
 wire \u0.w[0][29] ;
 wire \u0.w[0][2] ;
 wire \u0.w[0][30] ;
 wire \u0.w[0][31] ;
 wire \u0.w[0][3] ;
 wire \u0.w[0][4] ;
 wire \u0.w[0][5] ;
 wire \u0.w[0][6] ;
 wire \u0.w[0][7] ;
 wire \u0.w[0][8] ;
 wire \u0.w[0][9] ;
 wire \u0.w[1][0] ;
 wire \u0.w[1][10] ;
 wire \u0.w[1][11] ;
 wire \u0.w[1][12] ;
 wire \u0.w[1][13] ;
 wire \u0.w[1][14] ;
 wire \u0.w[1][15] ;
 wire \u0.w[1][16] ;
 wire \u0.w[1][17] ;
 wire \u0.w[1][18] ;
 wire \u0.w[1][19] ;
 wire \u0.w[1][1] ;
 wire \u0.w[1][20] ;
 wire \u0.w[1][21] ;
 wire \u0.w[1][22] ;
 wire \u0.w[1][23] ;
 wire \u0.w[1][24] ;
 wire \u0.w[1][25] ;
 wire \u0.w[1][26] ;
 wire \u0.w[1][27] ;
 wire \u0.w[1][28] ;
 wire \u0.w[1][29] ;
 wire \u0.w[1][2] ;
 wire \u0.w[1][30] ;
 wire \u0.w[1][31] ;
 wire \u0.w[1][3] ;
 wire \u0.w[1][4] ;
 wire \u0.w[1][5] ;
 wire \u0.w[1][6] ;
 wire \u0.w[1][7] ;
 wire \u0.w[1][8] ;
 wire \u0.w[1][9] ;
 wire \u0.w[2][0] ;
 wire \u0.w[2][10] ;
 wire \u0.w[2][11] ;
 wire \u0.w[2][12] ;
 wire \u0.w[2][13] ;
 wire \u0.w[2][14] ;
 wire \u0.w[2][15] ;
 wire \u0.w[2][16] ;
 wire \u0.w[2][17] ;
 wire \u0.w[2][18] ;
 wire \u0.w[2][19] ;
 wire \u0.w[2][1] ;
 wire \u0.w[2][20] ;
 wire \u0.w[2][21] ;
 wire \u0.w[2][22] ;
 wire \u0.w[2][23] ;
 wire \u0.w[2][24] ;
 wire \u0.w[2][25] ;
 wire \u0.w[2][26] ;
 wire \u0.w[2][27] ;
 wire \u0.w[2][28] ;
 wire \u0.w[2][29] ;
 wire \u0.w[2][2] ;
 wire \u0.w[2][30] ;
 wire \u0.w[2][31] ;
 wire \u0.w[2][3] ;
 wire \u0.w[2][4] ;
 wire \u0.w[2][5] ;
 wire \u0.w[2][6] ;
 wire \u0.w[2][7] ;
 wire \u0.w[2][8] ;
 wire \u0.w[2][9] ;
 wire clknet_leaf_26_clk;
 wire net4146;
 wire net4147;
 wire net4191;
 wire net4151;
 wire net4206;
 wire net4155;
 wire net4156;
 wire net4158;
 wire net4159;
 wire net4160;
 wire net4165;
 wire net4166;
 wire net4167;
 wire net4168;
 wire net4169;
 wire net4170;
 wire net4171;
 wire net4174;
 wire clknet_leaf_24_clk;
 wire net4183;
 wire net4176;
 wire net4184;
 wire net4186;
 wire net4187;
 wire net4189;
 wire clknet_leaf_4_clk;
 wire net4190;
 wire net4192;
 wire net4193;
 wire net4195;
 wire net4196;
 wire net4200;
 wire net4199;
 wire net4198;
 wire net4201;
 wire clknet_leaf_3_clk;
 wire net4202;
 wire net4203;
 wire net4205;
 wire net4210;
 wire net4211;
 wire net4212;
 wire net4214;
 wire net4219;
 wire net4213;
 wire net4216;
 wire net4215;
 wire net4217;
 wire clknet_leaf_2_clk;
 wire net4234;
 wire net4221;
 wire net4233;
 wire net4223;
 wire net4226;
 wire net4232;
 wire net4236;
 wire net4230;
 wire net4237;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_18_clk;
 wire net4053;
 wire net4052;
 wire net4031;
 wire net3562;
 wire net3561;
 wire [0:0] _11828_;
 wire [0:0] _11829_;
 wire [0:0] _11830_;
 wire [0:0] _11831_;
 wire [0:0] _11833_;
 wire [0:0] _11834_;
 wire [0:0] _11835_;
 wire [0:0] _11836_;
 wire [0:0] _11838_;
 wire [0:0] _11839_;
 wire [0:0] _11840_;
 wire [0:0] _11841_;
 wire [0:0] _11842_;
 wire [0:0] _11843_;
 wire [0:0] _11844_;
 wire [0:0] _11845_;
 wire [0:0] _11847_;
 wire [0:0] _11848_;
 wire [0:0] _11849_;
 wire [0:0] _11850_;
 wire [0:0] _11852_;
 wire [0:0] _11853_;
 wire [0:0] _11854_;
 wire [0:0] _11855_;
 wire [0:0] _11856_;
 wire [0:0] _11857_;
 wire [0:0] _11858_;
 wire [0:0] _11859_;
 wire [0:0] _11860_;
 wire [0:0] _11862_;
 wire [0:0] _11863_;
 wire [0:0] _11864_;
 wire [0:0] _11865_;
 wire [0:0] _11867_;
 wire [0:0] _11868_;
 wire [0:0] _11869_;
 wire [0:0] _11870_;
 wire [0:0] _11872_;
 wire [0:0] _11873_;
 wire [0:0] _11874_;
 wire [0:0] _11875_;
 wire [0:0] _11876_;
 wire [0:0] _11877_;
 wire [0:0] _11878_;
 wire [0:0] _11879_;
 wire [0:0] _11881_;
 wire [0:0] _11882_;
 wire [0:0] _11883_;
 wire [0:0] _11884_;
 wire [0:0] _11886_;
 wire [0:0] _11887_;
 wire [0:0] _11888_;
 wire [0:0] _11889_;
 wire [0:0] _11890_;
 wire [0:0] _11891_;
 wire [0:0] _11892_;
 wire [0:0] _11893_;
 wire [0:0] _11896_;
 wire [0:0] _11897_;
 wire [0:0] _11898_;
 wire [0:0] _11899_;
 wire [0:0] _11901_;
 wire [0:0] _11902_;
 wire [0:0] _11903_;
 wire [0:0] _11904_;
 wire [0:0] _11906_;
 wire [0:0] _11907_;
 wire [0:0] _11908_;
 wire [0:0] _11909_;
 wire [0:0] _11910_;
 wire [0:0] _11911_;
 wire [0:0] _11912_;
 wire [0:0] _11913_;
 wire [0:0] _11915_;
 wire [0:0] _11916_;
 wire [0:0] _11917_;
 wire [0:0] _11918_;
 wire [0:0] _11920_;
 wire [0:0] _11921_;
 wire [0:0] _11922_;
 wire [0:0] _11923_;
 wire [0:0] _11924_;
 wire [0:0] _11925_;
 wire [0:0] _11926_;
 wire [0:0] _11927_;
 wire [0:0] _11930_;
 wire [0:0] _11931_;
 wire [0:0] _11932_;
 wire [0:0] _11933_;
 wire [0:0] _11935_;
 wire [0:0] _11936_;
 wire [0:0] _11937_;
 wire [0:0] _11938_;
 wire [0:0] _11940_;
 wire [0:0] _11941_;
 wire [0:0] _11942_;
 wire [0:0] _11943_;
 wire [0:0] _11944_;
 wire [0:0] _11945_;
 wire [0:0] _11946_;
 wire [0:0] _11947_;
 wire [0:0] _11949_;
 wire [0:0] _11950_;
 wire [0:0] _11951_;
 wire [0:0] _11952_;
 wire [0:0] _11954_;
 wire [0:0] _11955_;
 wire [0:0] _11956_;
 wire [0:0] _11957_;
 wire [0:0] _11958_;
 wire [0:0] _11959_;
 wire [0:0] _11960_;
 wire [0:0] _11961_;
 wire [0:0] _11964_;
 wire [0:0] _11965_;
 wire [0:0] _11966_;
 wire [0:0] _11967_;
 wire [0:0] _11969_;
 wire [0:0] _11970_;
 wire [0:0] _11972_;
 wire [0:0] _11973_;
 wire [0:0] _11974_;
 wire [0:0] _11975_;
 wire [0:0] _11976_;
 wire [0:0] _11977_;
 wire [0:0] _11978_;
 wire [0:0] _11979_;
 wire [0:0] _11981_;
 wire [0:0] _11982_;
 wire [0:0] _11983_;
 wire [0:0] _11984_;
 wire [0:0] _11985_;
 wire [0:0] _11986_;
 wire [0:0] _11988_;
 wire [0:0] _11989_;
 wire [0:0] _11990_;
 wire [0:0] _11991_;
 wire [0:0] _11992_;
 wire [0:0] _11993_;
 wire [0:0] _11996_;
 wire [0:0] _11997_;
 wire [0:0] _11998_;
 wire [0:0] _11999_;
 wire [0:0] _12001_;
 wire [0:0] _12002_;
 wire [0:0] _12004_;
 wire [0:0] _12005_;
 wire [0:0] _12006_;
 wire [0:0] _12007_;
 wire [0:0] _12008_;
 wire [0:0] _12009_;
 wire [0:0] _12010_;
 wire [0:0] _12011_;
 wire [0:0] _12013_;
 wire [0:0] _12014_;
 wire [0:0] _12015_;
 wire [0:0] _12016_;
 wire [0:0] _12017_;
 wire [0:0] _12018_;
 wire [0:0] _12020_;
 wire [0:0] _12021_;
 wire [0:0] _12022_;
 wire [0:0] _12023_;
 wire [0:0] _12024_;
 wire [0:0] _12025_;
 wire [0:0] _12028_;
 wire [0:0] _12029_;
 wire [0:0] _12030_;
 wire [0:0] _12031_;
 wire [0:0] _12033_;
 wire [0:0] _12034_;
 wire [0:0] _12036_;
 wire [0:0] _12037_;
 wire [0:0] _12038_;
 wire [0:0] _12039_;
 wire [0:0] _12040_;
 wire [0:0] _12041_;
 wire [0:0] _12042_;
 wire [0:0] _12043_;
 wire [0:0] _12045_;
 wire [0:0] _12046_;
 wire [0:0] _12047_;
 wire [0:0] _12048_;
 wire [0:0] _12049_;
 wire [0:0] _12050_;
 wire [0:0] _12052_;
 wire [0:0] _12053_;
 wire [0:0] _12054_;
 wire [0:0] _12055_;
 wire [0:0] _12056_;
 wire [0:0] _12057_;
 wire [0:0] _12060_;
 wire [0:0] _12061_;
 wire [0:0] _12062_;
 wire [0:0] _12063_;
 wire [0:0] _12065_;
 wire [0:0] _12066_;
 wire [0:0] _12068_;
 wire [0:0] _12069_;
 wire [0:0] _12070_;
 wire [0:0] _12071_;
 wire [0:0] _12072_;
 wire [0:0] _12073_;
 wire [0:0] _12074_;
 wire [0:0] _12075_;
 wire [0:0] _12077_;
 wire [0:0] _12078_;
 wire [0:0] _12079_;
 wire [0:0] _12080_;
 wire [0:0] _12081_;
 wire [0:0] _12082_;
 wire [0:0] _12084_;
 wire [0:0] _12085_;
 wire [0:0] _12086_;
 wire [0:0] _12087_;
 wire [0:0] _12088_;
 wire [0:0] _12089_;
 wire [0:0] _12092_;
 wire [0:0] _12093_;
 wire [0:0] _12094_;
 wire [0:0] _12095_;
 wire [0:0] _12097_;
 wire [0:0] _12098_;
 wire [0:0] _12100_;
 wire [0:0] _12101_;
 wire [0:0] _12102_;
 wire [0:0] _12103_;
 wire [0:0] _12104_;
 wire [0:0] _12105_;
 wire [0:0] _12106_;
 wire [0:0] _12107_;
 wire [0:0] _12109_;
 wire [0:0] _12110_;
 wire [0:0] _12111_;
 wire [0:0] _12112_;
 wire [0:0] _12113_;
 wire [0:0] _12114_;
 wire [0:0] _12116_;
 wire [0:0] _12117_;
 wire [0:0] _12118_;
 wire [0:0] _12119_;
 wire [0:0] _12120_;
 wire [0:0] _12121_;
 wire [0:0] _12124_;
 wire [0:0] _12125_;
 wire [0:0] _12126_;
 wire [0:0] _12127_;
 wire [0:0] _12129_;
 wire [0:0] _12130_;
 wire [0:0] _12132_;
 wire [0:0] _12133_;
 wire [0:0] _12134_;
 wire [0:0] _12135_;
 wire [0:0] _12136_;
 wire [0:0] _12137_;
 wire [0:0] _12138_;
 wire [0:0] _12139_;
 wire [0:0] _12141_;
 wire [0:0] _12142_;
 wire [0:0] _12143_;
 wire [0:0] _12144_;
 wire [0:0] _12145_;
 wire [0:0] _12146_;
 wire [0:0] _12148_;
 wire [0:0] _12149_;
 wire [0:0] _12150_;
 wire [0:0] _12151_;
 wire [0:0] _12152_;
 wire [0:0] _12153_;
 wire [0:0] _12156_;
 wire [0:0] _12157_;
 wire [0:0] _12158_;
 wire [0:0] _12159_;
 wire [0:0] _12161_;
 wire [0:0] _12162_;
 wire [0:0] _12164_;
 wire [0:0] _12165_;
 wire [0:0] _12166_;
 wire [0:0] _12167_;
 wire [0:0] _12168_;
 wire [0:0] _12169_;
 wire [0:0] _12170_;
 wire [0:0] _12171_;
 wire [0:0] _12173_;
 wire [0:0] _12174_;
 wire [0:0] _12175_;
 wire [0:0] _12176_;
 wire [0:0] _12177_;
 wire [0:0] _12178_;
 wire [0:0] _12180_;
 wire [0:0] _12181_;
 wire [0:0] _12182_;
 wire [0:0] _12183_;
 wire [0:0] _12184_;
 wire [0:0] _12185_;
 wire [0:0] _12188_;
 wire [0:0] _12189_;
 wire [0:0] _12190_;
 wire [0:0] _12191_;
 wire [0:0] _12193_;
 wire [0:0] _12194_;
 wire [0:0] _12196_;
 wire [0:0] _12197_;
 wire [0:0] _12198_;
 wire [0:0] _12199_;
 wire [0:0] _12200_;
 wire [0:0] _12201_;
 wire [0:0] _12202_;
 wire [0:0] _12203_;
 wire [0:0] _12205_;
 wire [0:0] _12206_;
 wire [0:0] _12207_;
 wire [0:0] _12208_;
 wire [0:0] _12209_;
 wire [0:0] _12210_;
 wire [0:0] _12212_;
 wire [0:0] _12213_;
 wire [0:0] _12214_;
 wire [0:0] _12215_;
 wire [0:0] _12216_;
 wire [0:0] _12217_;
 wire [0:0] _12220_;
 wire [0:0] _12221_;
 wire [0:0] _12222_;
 wire [0:0] _12223_;
 wire [0:0] _12225_;
 wire [0:0] _12226_;
 wire [0:0] _12227_;
 wire [0:0] _12228_;
 wire [0:0] _12230_;
 wire [0:0] _12231_;
 wire [0:0] _12232_;
 wire [0:0] _12233_;
 wire [0:0] _12234_;
 wire [0:0] _12235_;
 wire [0:0] _12236_;
 wire [0:0] _12237_;
 wire [0:0] _12239_;
 wire [0:0] _12240_;
 wire [0:0] _12241_;
 wire [0:0] _12242_;
 wire [0:0] _12243_;
 wire [0:0] _12244_;
 wire [0:0] _12246_;
 wire [0:0] _12247_;
 wire [0:0] _12248_;
 wire [0:0] _12249_;
 wire [0:0] _12250_;
 wire [0:0] _12251_;
 wire [0:0] _12252_;
 wire [0:0] _12253_;
 wire [0:0] _12256_;
 wire [0:0] _12257_;
 wire [0:0] _12258_;
 wire [0:0] _12259_;
 wire [0:0] _12261_;
 wire [0:0] _12262_;
 wire [0:0] _12263_;
 wire [0:0] _12264_;
 wire [0:0] _12266_;
 wire [0:0] _12267_;
 wire [0:0] _12268_;
 wire [0:0] _12269_;
 wire [0:0] _12270_;
 wire [0:0] _12271_;
 wire [0:0] _12272_;
 wire [0:0] _12273_;
 wire [0:0] _12275_;
 wire [0:0] _12276_;
 wire [0:0] _12277_;
 wire [0:0] _12278_;
 wire [0:0] _12279_;
 wire [0:0] _12280_;
 wire [0:0] _12282_;
 wire [0:0] _12283_;
 wire [0:0] _12284_;
 wire [0:0] _12285_;
 wire [0:0] _12286_;
 wire [0:0] _12287_;
 wire [0:0] _12288_;
 wire [0:0] _12289_;
 wire [0:0] _12292_;
 wire [0:0] _12293_;
 wire [0:0] _12294_;
 wire [0:0] _12295_;
 wire [0:0] _12297_;
 wire [0:0] _12298_;
 wire [0:0] _12299_;
 wire [0:0] _12300_;
 wire [0:0] _12302_;
 wire [0:0] _12303_;
 wire [0:0] _12304_;
 wire [0:0] _12305_;
 wire [0:0] _12306_;
 wire [0:0] _12307_;
 wire [0:0] _12308_;
 wire [0:0] _12309_;
 wire [0:0] _12311_;
 wire [0:0] _12312_;
 wire [0:0] _12313_;
 wire [0:0] _12314_;
 wire [0:0] _12315_;
 wire [0:0] _12316_;
 wire [0:0] _12318_;
 wire [0:0] _12319_;
 wire [0:0] _12320_;
 wire [0:0] _12321_;
 wire [0:0] _12322_;
 wire [0:0] _12323_;
 wire [0:0] _12324_;
 wire [0:0] _12325_;
 wire [0:0] _12328_;
 wire [0:0] _12329_;
 wire [0:0] _12330_;
 wire [0:0] _12331_;
 wire [0:0] _12333_;
 wire [0:0] _12334_;
 wire [0:0] _12335_;
 wire [0:0] _12336_;
 wire [0:0] _12338_;
 wire [0:0] _12339_;
 wire [0:0] _12340_;
 wire [0:0] _12341_;
 wire [0:0] _12342_;
 wire [0:0] _12343_;
 wire [0:0] _12344_;
 wire [0:0] _12345_;
 wire [0:0] _12347_;
 wire [0:0] _12348_;
 wire [0:0] _12349_;
 wire [0:0] _12350_;
 wire [0:0] _12351_;
 wire [0:0] _12352_;
 wire [0:0] _12354_;
 wire [0:0] _12355_;
 wire [0:0] _12356_;
 wire [0:0] _12357_;
 wire [0:0] _12358_;
 wire [0:0] _12359_;
 wire [0:0] _12360_;
 wire [0:0] _12361_;
 wire [0:0] _12364_;
 wire [0:0] _12365_;
 wire [0:0] _12366_;
 wire [0:0] _12367_;
 wire [0:0] _12369_;
 wire [0:0] _12370_;
 wire [0:0] _12372_;
 wire [0:0] _12373_;
 wire [0:0] _12374_;
 wire [0:0] _12375_;
 wire [0:0] _12376_;
 wire [0:0] _12377_;
 wire [0:0] _12378_;
 wire [0:0] _12379_;
 wire [0:0] _12381_;
 wire [0:0] _12382_;
 wire [0:0] _12383_;
 wire [0:0] _12384_;
 wire [0:0] _12385_;
 wire [0:0] _12386_;
 wire [0:0] _12388_;
 wire [0:0] _12389_;
 wire [0:0] _12390_;
 wire [0:0] _12391_;
 wire [0:0] _12392_;
 wire [0:0] _12393_;
 wire [0:0] _12396_;
 wire [0:0] _12397_;
 wire [0:0] _12398_;
 wire [0:0] _12399_;
 wire [0:0] _12401_;
 wire [0:0] _12402_;
 wire [0:0] _12404_;
 wire [0:0] _12405_;
 wire [0:0] _12406_;
 wire [0:0] _12407_;
 wire [0:0] _12408_;
 wire [0:0] _12409_;
 wire [0:0] _12410_;
 wire [0:0] _12411_;
 wire [0:0] _12413_;
 wire [0:0] _12414_;
 wire [0:0] _12415_;
 wire [0:0] _12416_;
 wire [0:0] _12417_;
 wire [0:0] _12418_;
 wire [0:0] _12420_;
 wire [0:0] _12421_;
 wire [0:0] _12422_;
 wire [0:0] _12423_;
 wire [0:0] _12424_;
 wire [0:0] _12425_;
 wire [0:0] _12428_;
 wire [0:0] _12429_;
 wire [0:0] _12430_;
 wire [0:0] _12431_;
 wire [0:0] _12433_;
 wire [0:0] _12434_;
 wire [0:0] _12436_;
 wire [0:0] _12437_;
 wire [0:0] _12438_;
 wire [0:0] _12439_;
 wire [0:0] _12440_;
 wire [0:0] _12441_;
 wire [0:0] _12442_;
 wire [0:0] _12443_;
 wire [0:0] _12445_;
 wire [0:0] _12446_;
 wire [0:0] _12447_;
 wire [0:0] _12448_;
 wire [0:0] _12449_;
 wire [0:0] _12450_;
 wire [0:0] _12452_;
 wire [0:0] _12453_;
 wire [0:0] _12454_;
 wire [0:0] _12455_;
 wire [0:0] _12456_;
 wire [0:0] _12457_;
 wire [0:0] _12460_;
 wire [0:0] _12461_;
 wire [0:0] _12462_;
 wire [0:0] _12463_;
 wire [0:0] _12465_;
 wire [0:0] _12466_;
 wire [0:0] _12468_;
 wire [0:0] _12469_;
 wire [0:0] _12470_;
 wire [0:0] _12471_;
 wire [0:0] _12472_;
 wire [0:0] _12473_;
 wire [0:0] _12474_;
 wire [0:0] _12475_;
 wire [0:0] _12477_;
 wire [0:0] _12478_;
 wire [0:0] _12479_;
 wire [0:0] _12480_;
 wire [0:0] _12481_;
 wire [0:0] _12482_;
 wire [0:0] _12484_;
 wire [0:0] _12485_;
 wire [0:0] _12486_;
 wire [0:0] _12487_;
 wire [0:0] _12488_;
 wire [0:0] _12489_;
 wire [0:0] _12490_;
 wire [0:0] _12491_;
 wire [0:0] _12492_;
 wire [0:0] _12493_;
 wire [0:0] _12494_;
 wire [0:0] _12495_;
 wire [0:0] _12496_;
 wire [0:0] _12497_;
 wire [0:0] _12498_;
 wire [0:0] _12499_;

 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1400 ();
 sky130_fd_sc_hd__xor3_1 _12504_ (.A(\u0.w[0][19] ),
    .B(\u0.w[1][19] ),
    .C(\u0.subword[19] ),
    .X(_03574_));
 sky130_fd_sc_hd__xnor3_1 _12505_ (.A(\u0.tmp_w[19] ),
    .B(\u0.w[2][19] ),
    .C(_03574_),
    .X(_03575_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1399 ();
 sky130_fd_sc_hd__nand2_1 _12507_ (.A(net4234),
    .B(net39),
    .Y(_03577_));
 sky130_fd_sc_hd__o21a_4 _12508_ (.A1(net4234),
    .A2(_03575_),
    .B1(_03577_),
    .X(_03578_));
 sky130_fd_sc_hd__clkinv_16 _12509_ (.A(_03578_),
    .Y(_03579_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1397 ();
 sky130_fd_sc_hd__xor2_2 _12512_ (.A(\u0.w[0][16] ),
    .B(\u0.subword[16] ),
    .X(_03581_));
 sky130_fd_sc_hd__xor2_2 _12513_ (.A(\u0.w[2][16] ),
    .B(\u0.w[1][16] ),
    .X(_03582_));
 sky130_fd_sc_hd__xnor3_1 _12514_ (.A(\u0.tmp_w[16] ),
    .B(_03581_),
    .C(_03582_),
    .X(_03583_));
 sky130_fd_sc_hd__nand2_2 _12515_ (.A(net129),
    .B(net36),
    .Y(_03584_));
 sky130_fd_sc_hd__o21ai_4 _12516_ (.A1(net129),
    .A2(_03583_),
    .B1(_03584_),
    .Y(_03585_));
 sky130_fd_sc_hd__inv_16 _12517_ (.A(net4106),
    .Y(_03586_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1396 ();
 sky130_fd_sc_hd__xor2_2 _12519_ (.A(\u0.w[0][17] ),
    .B(\u0.subword[17] ),
    .X(_03587_));
 sky130_fd_sc_hd__xor2_2 _12520_ (.A(\u0.w[2][17] ),
    .B(\u0.w[1][17] ),
    .X(_03588_));
 sky130_fd_sc_hd__xnor3_1 _12521_ (.A(\u0.tmp_w[17] ),
    .B(_03587_),
    .C(_03588_),
    .X(_03589_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1395 ();
 sky130_fd_sc_hd__nand2_2 _12523_ (.A(net129),
    .B(net37),
    .Y(_03591_));
 sky130_fd_sc_hd__o21ai_4 _12524_ (.A1(net129),
    .A2(_03589_),
    .B1(_03591_),
    .Y(_03592_));
 sky130_fd_sc_hd__inv_16 _12525_ (.A(net4104),
    .Y(_03593_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1390 ();
 sky130_fd_sc_hd__xnor3_1 _12531_ (.A(\u0.w[0][21] ),
    .B(\u0.w[1][21] ),
    .C(\u0.subword[21] ),
    .X(_03598_));
 sky130_fd_sc_hd__xor3_1 _12532_ (.A(\u0.tmp_w[21] ),
    .B(\u0.w[2][21] ),
    .C(_03598_),
    .X(_03599_));
 sky130_fd_sc_hd__nor2_2 _12533_ (.A(net4234),
    .B(_03599_),
    .Y(_03600_));
 sky130_fd_sc_hd__a21oi_4 _12534_ (.A1(net4234),
    .A2(net42),
    .B1(_03600_),
    .Y(_03601_));
 sky130_fd_sc_hd__inv_16 _12535_ (.A(_03601_),
    .Y(_03602_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1385 ();
 sky130_fd_sc_hd__xnor3_1 _12541_ (.A(\u0.w[0][20] ),
    .B(\u0.w[1][20] ),
    .C(\u0.subword[20] ),
    .X(_03607_));
 sky130_fd_sc_hd__xor3_1 _12542_ (.A(\u0.tmp_w[20] ),
    .B(\u0.w[2][20] ),
    .C(_03607_),
    .X(_03608_));
 sky130_fd_sc_hd__nand2_1 _12543_ (.A(net4233),
    .B(net41),
    .Y(_03609_));
 sky130_fd_sc_hd__o21a_4 _12544_ (.A1(net4233),
    .A2(_03608_),
    .B1(_03609_),
    .X(_03610_));
 sky130_fd_sc_hd__clkinv_16 _12545_ (.A(_03610_),
    .Y(_03611_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1383 ();
 sky130_fd_sc_hd__xor2_4 _12548_ (.A(\u0.subword[18] ),
    .B(\u0.w[0][18] ),
    .X(_03613_));
 sky130_fd_sc_hd__xor2_2 _12549_ (.A(\u0.w[2][18] ),
    .B(\u0.w[1][18] ),
    .X(_03614_));
 sky130_fd_sc_hd__xnor3_1 _12550_ (.A(\u0.tmp_w[18] ),
    .B(_03613_),
    .C(_03614_),
    .X(_03615_));
 sky130_fd_sc_hd__nand2_1 _12551_ (.A(net4234),
    .B(net38),
    .Y(_03616_));
 sky130_fd_sc_hd__o21a_4 _12552_ (.A1(net4234),
    .A2(_03615_),
    .B1(_03616_),
    .X(_03617_));
 sky130_fd_sc_hd__clkinv_16 _12553_ (.A(_03617_),
    .Y(_03618_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1381 ();
 sky130_fd_sc_hd__xor2_2 _12556_ (.A(\u0.w[0][0] ),
    .B(\u0.subword[0] ),
    .X(_03620_));
 sky130_fd_sc_hd__xor2_1 _12557_ (.A(\u0.w[2][0] ),
    .B(\u0.w[1][0] ),
    .X(_03621_));
 sky130_fd_sc_hd__xnor3_1 _12558_ (.A(\u0.tmp_w[0] ),
    .B(_03620_),
    .C(_03621_),
    .X(_03622_));
 sky130_fd_sc_hd__nand2_2 _12559_ (.A(net129),
    .B(net1),
    .Y(_03623_));
 sky130_fd_sc_hd__o21ai_4 _12560_ (.A1(net129),
    .A2(_03622_),
    .B1(_03623_),
    .Y(_03624_));
 sky130_fd_sc_hd__inv_12 _12561_ (.A(_03624_),
    .Y(_03625_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1380 ();
 sky130_fd_sc_hd__xor2_2 _12563_ (.A(\u0.w[0][1] ),
    .B(\u0.subword[1] ),
    .X(_03626_));
 sky130_fd_sc_hd__xor2_1 _12564_ (.A(\u0.w[2][1] ),
    .B(\u0.w[1][1] ),
    .X(_03627_));
 sky130_fd_sc_hd__xnor3_1 _12565_ (.A(\u0.tmp_w[1] ),
    .B(_03626_),
    .C(_03627_),
    .X(_03628_));
 sky130_fd_sc_hd__nand2_1 _12566_ (.A(net129),
    .B(net40),
    .Y(_03629_));
 sky130_fd_sc_hd__o21ai_4 _12567_ (.A1(net129),
    .A2(_03628_),
    .B1(_03629_),
    .Y(_03630_));
 sky130_fd_sc_hd__inv_16 _12568_ (.A(_03630_),
    .Y(_03631_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1377 ();
 sky130_fd_sc_hd__xnor3_1 _12572_ (.A(\u0.subword[2] ),
    .B(\u0.w[0][2] ),
    .C(\u0.w[1][2] ),
    .X(_03634_));
 sky130_fd_sc_hd__xor3_1 _12573_ (.A(\u0.tmp_w[2] ),
    .B(\u0.w[2][2] ),
    .C(_03634_),
    .X(_03635_));
 sky130_fd_sc_hd__nand2_1 _12574_ (.A(net129),
    .B(net51),
    .Y(_03636_));
 sky130_fd_sc_hd__o21a_4 _12575_ (.A1(net129),
    .A2(_03635_),
    .B1(_03636_),
    .X(_03637_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1376 ();
 sky130_fd_sc_hd__clkinv_16 _12577_ (.A(_03637_),
    .Y(_03639_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1371 ();
 sky130_fd_sc_hd__xnor3_1 _12583_ (.A(\u0.w[0][3] ),
    .B(\u0.w[1][3] ),
    .C(\u0.subword[3] ),
    .X(_03644_));
 sky130_fd_sc_hd__xnor3_1 _12584_ (.A(\u0.tmp_w[3] ),
    .B(\u0.w[2][3] ),
    .C(_03644_),
    .X(_03645_));
 sky130_fd_sc_hd__nand2b_2 _12585_ (.A_N(net62),
    .B(net129),
    .Y(_03646_));
 sky130_fd_sc_hd__o21ai_4 _12586_ (.A1(net129),
    .A2(_03645_),
    .B1(_03646_),
    .Y(_03647_));
 sky130_fd_sc_hd__clkinv_16 _12587_ (.A(_03647_),
    .Y(_03648_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1366 ();
 sky130_fd_sc_hd__xnor3_1 _12593_ (.A(\u0.w[0][4] ),
    .B(\u0.w[1][4] ),
    .C(\u0.subword[4] ),
    .X(_03653_));
 sky130_fd_sc_hd__xor3_1 _12594_ (.A(\u0.tmp_w[4] ),
    .B(\u0.w[2][4] ),
    .C(_03653_),
    .X(_03654_));
 sky130_fd_sc_hd__nand2_1 _12595_ (.A(net4233),
    .B(net73),
    .Y(_03655_));
 sky130_fd_sc_hd__o21a_4 _12596_ (.A1(net4233),
    .A2(_03654_),
    .B1(_03655_),
    .X(_03656_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1365 ();
 sky130_fd_sc_hd__inv_16 _12598_ (.A(_03656_),
    .Y(_03658_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1361 ();
 sky130_fd_sc_hd__xnor3_1 _12603_ (.A(\u0.w[0][5] ),
    .B(\u0.w[1][5] ),
    .C(\u0.subword[5] ),
    .X(_03662_));
 sky130_fd_sc_hd__xor2_2 _12604_ (.A(\u0.w[2][5] ),
    .B(_03662_),
    .X(_03663_));
 sky130_fd_sc_hd__xor2_2 _12605_ (.A(\u0.tmp_w[5] ),
    .B(_03663_),
    .X(_03664_));
 sky130_fd_sc_hd__nand2_1 _12606_ (.A(net129),
    .B(net84),
    .Y(_03665_));
 sky130_fd_sc_hd__o21a_4 _12607_ (.A1(net129),
    .A2(_03664_),
    .B1(_03665_),
    .X(_03666_));
 sky130_fd_sc_hd__clkinv_16 _12608_ (.A(_03666_),
    .Y(_03667_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1357 ();
 sky130_fd_sc_hd__xnor3_1 _12613_ (.A(\u0.w[0][6] ),
    .B(\u0.w[1][6] ),
    .C(\u0.subword[6] ),
    .X(_03671_));
 sky130_fd_sc_hd__xor2_2 _12614_ (.A(\u0.w[2][6] ),
    .B(_03671_),
    .X(_03672_));
 sky130_fd_sc_hd__xor2_1 _12615_ (.A(\u0.tmp_w[6] ),
    .B(_03672_),
    .X(_03673_));
 sky130_fd_sc_hd__nand2_1 _12616_ (.A(net4233),
    .B(net95),
    .Y(_03674_));
 sky130_fd_sc_hd__o21a_4 _12617_ (.A1(net4233),
    .A2(_03673_),
    .B1(_03674_),
    .X(_03675_));
 sky130_fd_sc_hd__clkinv_16 _12618_ (.A(_03675_),
    .Y(_03676_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1354 ();
 sky130_fd_sc_hd__xor2_1 _12622_ (.A(\u0.w[0][7] ),
    .B(\u0.subword[7] ),
    .X(_03679_));
 sky130_fd_sc_hd__xnor2_2 _12623_ (.A(\u0.w[1][7] ),
    .B(_03679_),
    .Y(_03680_));
 sky130_fd_sc_hd__xnor2_1 _12624_ (.A(\u0.w[2][7] ),
    .B(_03680_),
    .Y(_03681_));
 sky130_fd_sc_hd__xnor2_1 _12625_ (.A(\u0.tmp_w[7] ),
    .B(_03681_),
    .Y(_03682_));
 sky130_fd_sc_hd__nor2_2 _12626_ (.A(net4233),
    .B(_03682_),
    .Y(_03683_));
 sky130_fd_sc_hd__a21oi_4 _12627_ (.A1(net4233),
    .A2(net106),
    .B1(_03683_),
    .Y(_03684_));
 sky130_fd_sc_hd__inv_12 _12628_ (.A(_03684_),
    .Y(_03685_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1352 ();
 sky130_fd_sc_hd__xnor3_1 _12631_ (.A(\u0.w[0][8] ),
    .B(\u0.w[1][8] ),
    .C(\u0.subword[8] ),
    .X(_03687_));
 sky130_fd_sc_hd__xor3_1 _12632_ (.A(\u0.tmp_w[8] ),
    .B(\u0.w[2][8] ),
    .C(_03687_),
    .X(_03688_));
 sky130_fd_sc_hd__nand2_2 _12633_ (.A(net129),
    .B(net117),
    .Y(_03689_));
 sky130_fd_sc_hd__o21ai_4 _12634_ (.A1(net129),
    .A2(_03688_),
    .B1(_03689_),
    .Y(_03690_));
 sky130_fd_sc_hd__clkinvlp_4 _12635_ (.A(_03690_),
    .Y(_03691_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1350 ();
 sky130_fd_sc_hd__xnor3_1 _12638_ (.A(\u0.w[0][9] ),
    .B(\u0.w[1][9] ),
    .C(\u0.subword[9] ),
    .X(_03693_));
 sky130_fd_sc_hd__xor3_1 _12639_ (.A(\u0.tmp_w[9] ),
    .B(\u0.w[2][9] ),
    .C(_03693_),
    .X(_03694_));
 sky130_fd_sc_hd__nand2_2 _12640_ (.A(net129),
    .B(net128),
    .Y(_03695_));
 sky130_fd_sc_hd__o21ai_4 _12641_ (.A1(net129),
    .A2(_03694_),
    .B1(_03695_),
    .Y(_11860_[0]));
 sky130_fd_sc_hd__clkinv_16 _12642_ (.A(_11860_[0]),
    .Y(_03696_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1347 ();
 sky130_fd_sc_hd__xor3_1 _12646_ (.A(\u0.subword[10] ),
    .B(\u0.w[0][10] ),
    .C(\u0.w[1][10] ),
    .X(_03699_));
 sky130_fd_sc_hd__xnor3_1 _12647_ (.A(\u0.tmp_w[10] ),
    .B(\u0.w[2][10] ),
    .C(_03699_),
    .X(_03700_));
 sky130_fd_sc_hd__nand2_1 _12648_ (.A(net4237),
    .B(net12),
    .Y(_03701_));
 sky130_fd_sc_hd__o21a_4 _12649_ (.A1(net4237),
    .A2(_03700_),
    .B1(_03701_),
    .X(_03702_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1346 ();
 sky130_fd_sc_hd__clkinv_16 _12651_ (.A(_03702_),
    .Y(_03704_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1339 ();
 sky130_fd_sc_hd__xor3_1 _12659_ (.A(\u0.w[0][11] ),
    .B(\u0.w[1][11] ),
    .C(\u0.subword[11] ),
    .X(_03711_));
 sky130_fd_sc_hd__xnor3_1 _12660_ (.A(\u0.tmp_w[11] ),
    .B(\u0.w[2][11] ),
    .C(_03711_),
    .X(_03712_));
 sky130_fd_sc_hd__nand2_1 _12661_ (.A(net4237),
    .B(net23),
    .Y(_03713_));
 sky130_fd_sc_hd__o21a_4 _12662_ (.A1(net4237),
    .A2(_03712_),
    .B1(_03713_),
    .X(_03714_));
 sky130_fd_sc_hd__clkinv_16 _12663_ (.A(_03714_),
    .Y(_03715_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1333 ();
 sky130_fd_sc_hd__xnor3_1 _12670_ (.A(\u0.w[0][12] ),
    .B(\u0.w[1][12] ),
    .C(\u0.subword[12] ),
    .X(_03721_));
 sky130_fd_sc_hd__xor3_1 _12671_ (.A(\u0.tmp_w[12] ),
    .B(\u0.w[2][12] ),
    .C(_03721_),
    .X(_03722_));
 sky130_fd_sc_hd__nor2_1 _12672_ (.A(net4237),
    .B(_03722_),
    .Y(_03723_));
 sky130_fd_sc_hd__a21oi_4 _12673_ (.A1(net4237),
    .A2(net32),
    .B1(_03723_),
    .Y(_03724_));
 sky130_fd_sc_hd__clkinv_16 _12674_ (.A(_03724_),
    .Y(_03725_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1328 ();
 sky130_fd_sc_hd__xnor3_1 _12680_ (.A(\u0.w[0][13] ),
    .B(\u0.w[1][13] ),
    .C(\u0.subword[13] ),
    .X(_03730_));
 sky130_fd_sc_hd__xnor2_2 _12681_ (.A(\u0.w[2][13] ),
    .B(_03730_),
    .Y(_03731_));
 sky130_fd_sc_hd__xnor2_1 _12682_ (.A(\u0.tmp_w[13] ),
    .B(_03731_),
    .Y(_03732_));
 sky130_fd_sc_hd__nand2_1 _12683_ (.A(net4237),
    .B(net33),
    .Y(_03733_));
 sky130_fd_sc_hd__o21a_4 _12684_ (.A1(net4237),
    .A2(_03732_),
    .B1(_03733_),
    .X(_03734_));
 sky130_fd_sc_hd__clkinv_16 _12685_ (.A(_03734_),
    .Y(_03735_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1324 ();
 sky130_fd_sc_hd__xnor3_1 _12690_ (.A(\u0.w[0][14] ),
    .B(\u0.w[1][14] ),
    .C(\u0.subword[14] ),
    .X(_03739_));
 sky130_fd_sc_hd__xor2_1 _12691_ (.A(\u0.w[2][14] ),
    .B(_03739_),
    .X(_03740_));
 sky130_fd_sc_hd__xor2_1 _12692_ (.A(\u0.tmp_w[14] ),
    .B(_03740_),
    .X(_03741_));
 sky130_fd_sc_hd__nor2_1 _12693_ (.A(net4237),
    .B(_03741_),
    .Y(_03742_));
 sky130_fd_sc_hd__a21oi_4 _12694_ (.A1(net4237),
    .A2(net34),
    .B1(_03742_),
    .Y(_03743_));
 sky130_fd_sc_hd__inv_12 _12695_ (.A(_03743_),
    .Y(_03744_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1323 ();
 sky130_fd_sc_hd__xor2_1 _12697_ (.A(\u0.w[0][15] ),
    .B(\u0.subword[15] ),
    .X(_03745_));
 sky130_fd_sc_hd__xnor2_1 _12698_ (.A(\u0.w[1][15] ),
    .B(_03745_),
    .Y(_03746_));
 sky130_fd_sc_hd__xnor2_2 _12699_ (.A(\u0.w[2][15] ),
    .B(_03746_),
    .Y(_03747_));
 sky130_fd_sc_hd__xnor2_1 _12700_ (.A(\u0.tmp_w[15] ),
    .B(_03747_),
    .Y(_03748_));
 sky130_fd_sc_hd__nor2_2 _12701_ (.A(net4237),
    .B(_03748_),
    .Y(_03749_));
 sky130_fd_sc_hd__a21oi_4 _12702_ (.A1(net4237),
    .A2(net35),
    .B1(_03749_),
    .Y(_03750_));
 sky130_fd_sc_hd__inv_12 _12703_ (.A(_03750_),
    .Y(_03751_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1319 ();
 sky130_fd_sc_hd__xnor3_1 _12708_ (.A(\u0.w[0][22] ),
    .B(\u0.w[1][22] ),
    .C(\u0.subword[22] ),
    .X(_03755_));
 sky130_fd_sc_hd__xor3_1 _12709_ (.A(\u0.tmp_w[22] ),
    .B(\u0.w[2][22] ),
    .C(_03755_),
    .X(_03756_));
 sky130_fd_sc_hd__nand2_1 _12710_ (.A(net4234),
    .B(net43),
    .Y(_03757_));
 sky130_fd_sc_hd__o21a_4 _12711_ (.A1(net4234),
    .A2(_03756_),
    .B1(_03757_),
    .X(_03758_));
 sky130_fd_sc_hd__clkinv_16 _12712_ (.A(_03758_),
    .Y(_03759_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1317 ();
 sky130_fd_sc_hd__xor2_2 _12715_ (.A(\u0.w[0][23] ),
    .B(\u0.subword[23] ),
    .X(_03761_));
 sky130_fd_sc_hd__xnor2_4 _12716_ (.A(\u0.w[1][23] ),
    .B(_03761_),
    .Y(_03762_));
 sky130_fd_sc_hd__xnor2_1 _12717_ (.A(\u0.w[2][23] ),
    .B(_03762_),
    .Y(_03763_));
 sky130_fd_sc_hd__xnor2_1 _12718_ (.A(\u0.tmp_w[23] ),
    .B(_03763_),
    .Y(_03764_));
 sky130_fd_sc_hd__nor2_1 _12719_ (.A(net4233),
    .B(_03764_),
    .Y(_03765_));
 sky130_fd_sc_hd__a21oi_4 _12720_ (.A1(net4233),
    .A2(net44),
    .B1(_03765_),
    .Y(_03766_));
 sky130_fd_sc_hd__inv_12 _12721_ (.A(_03766_),
    .Y(_03767_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1315 ();
 sky130_fd_sc_hd__xnor3_1 _12724_ (.A(\u0.w[0][24] ),
    .B(\u0.subword[24] ),
    .C(\u0.r0.out[24] ),
    .X(_03769_));
 sky130_fd_sc_hd__xor2_1 _12725_ (.A(\u0.tmp_w[24] ),
    .B(\u0.w[2][24] ),
    .X(_03770_));
 sky130_fd_sc_hd__xnor3_1 _12726_ (.A(\u0.w[1][24] ),
    .B(_03769_),
    .C(_03770_),
    .X(_03771_));
 sky130_fd_sc_hd__mux2_8 _12727_ (.A0(_03771_),
    .A1(net45),
    .S(net129),
    .X(_03772_));
 sky130_fd_sc_hd__clkinv_16 _12728_ (.A(_03772_),
    .Y(_03773_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1314 ();
 sky130_fd_sc_hd__xnor3_1 _12730_ (.A(\u0.w[0][25] ),
    .B(\u0.subword[25] ),
    .C(\u0.r0.out[25] ),
    .X(_03774_));
 sky130_fd_sc_hd__xor2_1 _12731_ (.A(\u0.tmp_w[25] ),
    .B(\u0.w[2][25] ),
    .X(_03775_));
 sky130_fd_sc_hd__xnor3_1 _12732_ (.A(\u0.w[1][25] ),
    .B(_03774_),
    .C(_03775_),
    .X(_03776_));
 sky130_fd_sc_hd__mux2_8 _12733_ (.A0(_03776_),
    .A1(net46),
    .S(net129),
    .X(_03777_));
 sky130_fd_sc_hd__clkinv_16 _12734_ (.A(_03777_),
    .Y(_03778_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1313 ();
 sky130_fd_sc_hd__xnor3_1 _12736_ (.A(\u0.w[0][26] ),
    .B(\u0.subword[26] ),
    .C(\u0.r0.out[26] ),
    .X(_03779_));
 sky130_fd_sc_hd__xnor2_1 _12737_ (.A(\u0.tmp_w[26] ),
    .B(\u0.w[2][26] ),
    .Y(_03780_));
 sky130_fd_sc_hd__xnor3_1 _12738_ (.A(\u0.w[1][26] ),
    .B(_03779_),
    .C(_03780_),
    .X(_03781_));
 sky130_fd_sc_hd__inv_1 _12739_ (.A(net47),
    .Y(_03782_));
 sky130_fd_sc_hd__mux2i_1 _12740_ (.A0(_03781_),
    .A1(_03782_),
    .S(net129),
    .Y(_03783_));
 sky130_fd_sc_hd__clkinv_16 _12741_ (.A(net4078),
    .Y(_03784_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1310 ();
 sky130_fd_sc_hd__xnor3_1 _12745_ (.A(\u0.w[0][27] ),
    .B(\u0.subword[27] ),
    .C(\u0.r0.out[27] ),
    .X(_03787_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1309 ();
 sky130_fd_sc_hd__xor2_1 _12747_ (.A(\u0.tmp_w[27] ),
    .B(\u0.w[2][27] ),
    .X(_03789_));
 sky130_fd_sc_hd__xnor3_1 _12748_ (.A(\u0.w[1][27] ),
    .B(_03787_),
    .C(_03789_),
    .X(_03790_));
 sky130_fd_sc_hd__mux2i_4 _12749_ (.A0(_03790_),
    .A1(net48),
    .S(net129),
    .Y(_03791_));
 sky130_fd_sc_hd__inv_16 _12750_ (.A(_03791_),
    .Y(_03792_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1305 ();
 sky130_fd_sc_hd__xnor3_1 _12755_ (.A(\u0.w[0][28] ),
    .B(\u0.subword[28] ),
    .C(\u0.r0.out[28] ),
    .X(_03796_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1304 ();
 sky130_fd_sc_hd__xor2_1 _12757_ (.A(\u0.tmp_w[28] ),
    .B(\u0.w[2][28] ),
    .X(_03798_));
 sky130_fd_sc_hd__xnor3_1 _12758_ (.A(\u0.w[1][28] ),
    .B(_03796_),
    .C(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__mux2i_4 _12759_ (.A0(_03799_),
    .A1(net49),
    .S(net129),
    .Y(_03800_));
 sky130_fd_sc_hd__inv_16 _12760_ (.A(_03800_),
    .Y(_03801_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1300 ();
 sky130_fd_sc_hd__xnor2_1 _12765_ (.A(\u0.w[0][29] ),
    .B(\u0.subword[29] ),
    .Y(_03805_));
 sky130_fd_sc_hd__xnor3_1 _12766_ (.A(\u0.w[1][29] ),
    .B(\u0.r0.out[29] ),
    .C(_03805_),
    .X(_03806_));
 sky130_fd_sc_hd__xnor3_1 _12767_ (.A(\u0.tmp_w[29] ),
    .B(\u0.w[2][29] ),
    .C(_03806_),
    .X(_03807_));
 sky130_fd_sc_hd__nand2_1 _12768_ (.A(net129),
    .B(net50),
    .Y(_03808_));
 sky130_fd_sc_hd__o21a_4 _12769_ (.A1(net129),
    .A2(_03807_),
    .B1(_03808_),
    .X(_03809_));
 sky130_fd_sc_hd__inv_16 _12770_ (.A(_03809_),
    .Y(_03810_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1297 ();
 sky130_fd_sc_hd__xnor3_1 _12774_ (.A(\u0.w[0][30] ),
    .B(\u0.subword[30] ),
    .C(\u0.r0.out[30] ),
    .X(_03813_));
 sky130_fd_sc_hd__xnor3_1 _12775_ (.A(\u0.w[2][30] ),
    .B(\u0.w[1][30] ),
    .C(_03813_),
    .X(_03814_));
 sky130_fd_sc_hd__xnor2_1 _12776_ (.A(\u0.tmp_w[30] ),
    .B(_03814_),
    .Y(_03815_));
 sky130_fd_sc_hd__nand2_1 _12777_ (.A(net129),
    .B(net52),
    .Y(_03816_));
 sky130_fd_sc_hd__o21a_4 _12778_ (.A1(net129),
    .A2(_03815_),
    .B1(_03816_),
    .X(_03817_));
 sky130_fd_sc_hd__inv_12 _12779_ (.A(_03817_),
    .Y(_00398_));
 sky130_fd_sc_hd__xor2_1 _12780_ (.A(\u0.subword[31] ),
    .B(\u0.r0.out[31] ),
    .X(_03818_));
 sky130_fd_sc_hd__xnor2_1 _12781_ (.A(\u0.w[0][31] ),
    .B(_03818_),
    .Y(_03819_));
 sky130_fd_sc_hd__xnor2_2 _12782_ (.A(\u0.w[1][31] ),
    .B(_03819_),
    .Y(_03820_));
 sky130_fd_sc_hd__xnor2_1 _12783_ (.A(\u0.w[2][31] ),
    .B(_03820_),
    .Y(_03821_));
 sky130_fd_sc_hd__xor2_1 _12784_ (.A(\u0.tmp_w[31] ),
    .B(_03821_),
    .X(_03822_));
 sky130_fd_sc_hd__nand2_2 _12785_ (.A(net4232),
    .B(net53),
    .Y(_03823_));
 sky130_fd_sc_hd__o21ai_4 _12786_ (.A1(net4232),
    .A2(_03822_),
    .B1(_03823_),
    .Y(_03824_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1295 ();
 sky130_fd_sc_hd__xor2_1 _12789_ (.A(_03620_),
    .B(_03621_),
    .X(_03826_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1293 ();
 sky130_fd_sc_hd__mux2_1 _12792_ (.A0(_03826_),
    .A1(net54),
    .S(net4235),
    .X(_00353_));
 sky130_fd_sc_hd__xor2_1 _12793_ (.A(_03626_),
    .B(_03627_),
    .X(_03829_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1292 ();
 sky130_fd_sc_hd__mux2_1 _12795_ (.A0(_03829_),
    .A1(net55),
    .S(net129),
    .X(_00364_));
 sky130_fd_sc_hd__xnor2_1 _12796_ (.A(\u0.w[2][2] ),
    .B(_03634_),
    .Y(_03831_));
 sky130_fd_sc_hd__mux2_1 _12797_ (.A0(_03831_),
    .A1(net56),
    .S(net129),
    .X(_00375_));
 sky130_fd_sc_hd__xnor2_1 _12798_ (.A(\u0.w[2][3] ),
    .B(_03644_),
    .Y(_03832_));
 sky130_fd_sc_hd__mux2_1 _12799_ (.A0(_03832_),
    .A1(net57),
    .S(net129),
    .X(_00378_));
 sky130_fd_sc_hd__xnor2_1 _12800_ (.A(\u0.w[2][4] ),
    .B(_03653_),
    .Y(_03833_));
 sky130_fd_sc_hd__mux2_1 _12801_ (.A0(_03833_),
    .A1(net58),
    .S(net129),
    .X(_00379_));
 sky130_fd_sc_hd__inv_1 _12802_ (.A(net59),
    .Y(_03834_));
 sky130_fd_sc_hd__mux2i_1 _12803_ (.A0(_03663_),
    .A1(_03834_),
    .S(net129),
    .Y(_00380_));
 sky130_fd_sc_hd__inv_1 _12804_ (.A(net60),
    .Y(_03835_));
 sky130_fd_sc_hd__mux2i_1 _12805_ (.A0(_03672_),
    .A1(_03835_),
    .S(net4232),
    .Y(_00381_));
 sky130_fd_sc_hd__mux2_1 _12806_ (.A0(_03681_),
    .A1(net61),
    .S(net129),
    .X(_00382_));
 sky130_fd_sc_hd__xnor2_1 _12807_ (.A(\u0.w[2][8] ),
    .B(_03687_),
    .Y(_03836_));
 sky130_fd_sc_hd__mux2_1 _12808_ (.A0(_03836_),
    .A1(net63),
    .S(net4237),
    .X(_00383_));
 sky130_fd_sc_hd__xnor2_1 _12809_ (.A(\u0.w[2][9] ),
    .B(_03693_),
    .Y(_03837_));
 sky130_fd_sc_hd__mux2_1 _12810_ (.A0(_03837_),
    .A1(net64),
    .S(net4236),
    .X(_00384_));
 sky130_fd_sc_hd__xor2_1 _12811_ (.A(\u0.w[2][10] ),
    .B(_03699_),
    .X(_03838_));
 sky130_fd_sc_hd__mux2_1 _12812_ (.A0(_03838_),
    .A1(net65),
    .S(net4237),
    .X(_00354_));
 sky130_fd_sc_hd__xor2_1 _12813_ (.A(net4141),
    .B(_03711_),
    .X(_03839_));
 sky130_fd_sc_hd__mux2_1 _12814_ (.A0(_03839_),
    .A1(net66),
    .S(net4238),
    .X(_00355_));
 sky130_fd_sc_hd__xnor2_1 _12815_ (.A(net4140),
    .B(_03721_),
    .Y(_03840_));
 sky130_fd_sc_hd__mux2_1 _12816_ (.A0(_03840_),
    .A1(net67),
    .S(net4238),
    .X(_00356_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1291 ();
 sky130_fd_sc_hd__mux2_1 _12818_ (.A0(_03731_),
    .A1(net68),
    .S(net4237),
    .X(_00357_));
 sky130_fd_sc_hd__inv_1 _12819_ (.A(net69),
    .Y(_03842_));
 sky130_fd_sc_hd__mux2i_1 _12820_ (.A0(_03740_),
    .A1(_03842_),
    .S(net4237),
    .Y(_00358_));
 sky130_fd_sc_hd__mux2_1 _12821_ (.A0(_03747_),
    .A1(net70),
    .S(net4239),
    .X(_00359_));
 sky130_fd_sc_hd__xor2_1 _12822_ (.A(net4124),
    .B(_03582_),
    .X(_03843_));
 sky130_fd_sc_hd__mux2_1 _12823_ (.A0(_03843_),
    .A1(net71),
    .S(net4235),
    .X(_00360_));
 sky130_fd_sc_hd__xor2_1 _12824_ (.A(net4123),
    .B(_03588_),
    .X(_03844_));
 sky130_fd_sc_hd__mux2_1 _12825_ (.A0(_03844_),
    .A1(net72),
    .S(net4236),
    .X(_00361_));
 sky130_fd_sc_hd__xor2_1 _12826_ (.A(_03613_),
    .B(_03614_),
    .X(_03845_));
 sky130_fd_sc_hd__mux2_1 _12827_ (.A0(_03845_),
    .A1(net74),
    .S(net4235),
    .X(_00362_));
 sky130_fd_sc_hd__xor2_1 _12828_ (.A(\u0.w[2][19] ),
    .B(net4125),
    .X(_03846_));
 sky130_fd_sc_hd__mux2_1 _12829_ (.A0(_03846_),
    .A1(net75),
    .S(net4235),
    .X(_00363_));
 sky130_fd_sc_hd__xnor2_1 _12830_ (.A(net4138),
    .B(_03607_),
    .Y(_03847_));
 sky130_fd_sc_hd__mux2_1 _12831_ (.A0(_03847_),
    .A1(net76),
    .S(net4233),
    .X(_00365_));
 sky130_fd_sc_hd__xnor2_1 _12832_ (.A(\u0.w[2][21] ),
    .B(_03598_),
    .Y(_03848_));
 sky130_fd_sc_hd__mux2_1 _12833_ (.A0(_03848_),
    .A1(net77),
    .S(net4235),
    .X(_00366_));
 sky130_fd_sc_hd__xnor2_1 _12834_ (.A(\u0.w[2][22] ),
    .B(_03755_),
    .Y(_03849_));
 sky130_fd_sc_hd__mux2_1 _12835_ (.A0(_03849_),
    .A1(net78),
    .S(net4235),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_1 _12836_ (.A0(_03763_),
    .A1(net79),
    .S(net4233),
    .X(_00368_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1290 ();
 sky130_fd_sc_hd__xnor2_1 _12838_ (.A(net4151),
    .B(_03769_),
    .Y(_03851_));
 sky130_fd_sc_hd__xnor2_1 _12839_ (.A(\u0.w[2][24] ),
    .B(_03851_),
    .Y(_03852_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1288 ();
 sky130_fd_sc_hd__nand2_1 _12842_ (.A(net4235),
    .B(net80),
    .Y(_03855_));
 sky130_fd_sc_hd__o21ai_0 _12843_ (.A1(net4235),
    .A2(_03852_),
    .B1(_03855_),
    .Y(_00369_));
 sky130_fd_sc_hd__xnor2_1 _12844_ (.A(\u0.w[1][25] ),
    .B(_03774_),
    .Y(_03856_));
 sky130_fd_sc_hd__xnor2_1 _12845_ (.A(net4137),
    .B(_03856_),
    .Y(_03857_));
 sky130_fd_sc_hd__nand2_1 _12846_ (.A(net129),
    .B(net81),
    .Y(_03858_));
 sky130_fd_sc_hd__o21ai_0 _12847_ (.A1(net129),
    .A2(_03857_),
    .B1(_03858_),
    .Y(_00370_));
 sky130_fd_sc_hd__xnor2_1 _12848_ (.A(net4149),
    .B(_03779_),
    .Y(_03859_));
 sky130_fd_sc_hd__xnor2_1 _12849_ (.A(\u0.w[2][26] ),
    .B(_03859_),
    .Y(_03860_));
 sky130_fd_sc_hd__nand2_1 _12850_ (.A(net4232),
    .B(net82),
    .Y(_03861_));
 sky130_fd_sc_hd__o21ai_0 _12851_ (.A1(net129),
    .A2(_03860_),
    .B1(_03861_),
    .Y(_00371_));
 sky130_fd_sc_hd__xnor2_1 _12852_ (.A(\u0.w[1][27] ),
    .B(_03787_),
    .Y(_03862_));
 sky130_fd_sc_hd__xnor2_1 _12853_ (.A(\u0.w[2][27] ),
    .B(_03862_),
    .Y(_03863_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1287 ();
 sky130_fd_sc_hd__nand2_1 _12855_ (.A(net129),
    .B(net83),
    .Y(_03865_));
 sky130_fd_sc_hd__o21ai_0 _12856_ (.A1(net4232),
    .A2(_03863_),
    .B1(_03865_),
    .Y(_00372_));
 sky130_fd_sc_hd__xnor2_1 _12857_ (.A(\u0.w[1][28] ),
    .B(_03796_),
    .Y(_03866_));
 sky130_fd_sc_hd__xnor2_1 _12858_ (.A(\u0.w[2][28] ),
    .B(_03866_),
    .Y(_03867_));
 sky130_fd_sc_hd__nand2_1 _12859_ (.A(net4232),
    .B(net85),
    .Y(_03868_));
 sky130_fd_sc_hd__o21ai_0 _12860_ (.A1(net4232),
    .A2(_03867_),
    .B1(_03868_),
    .Y(_00373_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1286 ();
 sky130_fd_sc_hd__xnor2_1 _12862_ (.A(\u0.w[2][29] ),
    .B(_03806_),
    .Y(_03870_));
 sky130_fd_sc_hd__nand2_1 _12863_ (.A(net4232),
    .B(net86),
    .Y(_03871_));
 sky130_fd_sc_hd__o21ai_0 _12864_ (.A1(net4232),
    .A2(_03870_),
    .B1(_03871_),
    .Y(_00374_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1285 ();
 sky130_fd_sc_hd__mux2_1 _12866_ (.A0(_03814_),
    .A1(net87),
    .S(net4232),
    .X(_00376_));
 sky130_fd_sc_hd__nand2_1 _12867_ (.A(net4232),
    .B(net88),
    .Y(_03873_));
 sky130_fd_sc_hd__o21ai_0 _12868_ (.A1(net4232),
    .A2(_03821_),
    .B1(_03873_),
    .Y(_00377_));
 sky130_fd_sc_hd__xnor2_1 _12869_ (.A(net4157),
    .B(_03620_),
    .Y(_03874_));
 sky130_fd_sc_hd__nand2_1 _12870_ (.A(net4235),
    .B(net89),
    .Y(_03875_));
 sky130_fd_sc_hd__o21ai_0 _12871_ (.A1(net129),
    .A2(_03874_),
    .B1(_03875_),
    .Y(_00321_));
 sky130_fd_sc_hd__xnor2_1 _12872_ (.A(net4153),
    .B(_03626_),
    .Y(_03876_));
 sky130_fd_sc_hd__nand2_1 _12873_ (.A(net129),
    .B(net90),
    .Y(_03877_));
 sky130_fd_sc_hd__o21ai_0 _12874_ (.A1(net129),
    .A2(_03876_),
    .B1(_03877_),
    .Y(_00332_));
 sky130_fd_sc_hd__nand2_1 _12875_ (.A(net4236),
    .B(net91),
    .Y(_03878_));
 sky130_fd_sc_hd__o21ai_0 _12876_ (.A1(net4236),
    .A2(_03634_),
    .B1(_03878_),
    .Y(_00343_));
 sky130_fd_sc_hd__nand2_1 _12877_ (.A(net4235),
    .B(net92),
    .Y(_03879_));
 sky130_fd_sc_hd__o21ai_0 _12878_ (.A1(net4235),
    .A2(_03644_),
    .B1(_03879_),
    .Y(_00346_));
 sky130_fd_sc_hd__nand2_1 _12879_ (.A(net4235),
    .B(net93),
    .Y(_03880_));
 sky130_fd_sc_hd__o21ai_0 _12880_ (.A1(net4235),
    .A2(_03653_),
    .B1(_03880_),
    .Y(_00347_));
 sky130_fd_sc_hd__nand2_1 _12881_ (.A(net4236),
    .B(net94),
    .Y(_03881_));
 sky130_fd_sc_hd__o21ai_0 _12882_ (.A1(net4236),
    .A2(_03662_),
    .B1(_03881_),
    .Y(_00348_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1284 ();
 sky130_fd_sc_hd__nand2_1 _12884_ (.A(net4236),
    .B(net96),
    .Y(_03883_));
 sky130_fd_sc_hd__o21ai_0 _12885_ (.A1(net4236),
    .A2(_03671_),
    .B1(_03883_),
    .Y(_00349_));
 sky130_fd_sc_hd__nand2_1 _12886_ (.A(net4235),
    .B(net97),
    .Y(_03884_));
 sky130_fd_sc_hd__o21ai_0 _12887_ (.A1(net4235),
    .A2(_03680_),
    .B1(_03884_),
    .Y(_00350_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1283 ();
 sky130_fd_sc_hd__nand2_1 _12889_ (.A(net4237),
    .B(net98),
    .Y(_03886_));
 sky130_fd_sc_hd__o21ai_0 _12890_ (.A1(net4237),
    .A2(_03687_),
    .B1(_03886_),
    .Y(_00351_));
 sky130_fd_sc_hd__nand2_1 _12891_ (.A(net4236),
    .B(net99),
    .Y(_03887_));
 sky130_fd_sc_hd__o21ai_0 _12892_ (.A1(net4236),
    .A2(_03693_),
    .B1(_03887_),
    .Y(_00352_));
 sky130_fd_sc_hd__mux2_1 _12893_ (.A0(_03699_),
    .A1(net100),
    .S(net4237),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _12894_ (.A0(_03711_),
    .A1(net101),
    .S(net4238),
    .X(_00323_));
 sky130_fd_sc_hd__nand2_1 _12895_ (.A(net4238),
    .B(net102),
    .Y(_03888_));
 sky130_fd_sc_hd__o21ai_0 _12896_ (.A1(net4238),
    .A2(_03721_),
    .B1(_03888_),
    .Y(_00324_));
 sky130_fd_sc_hd__nand2_1 _12897_ (.A(net4237),
    .B(net103),
    .Y(_03889_));
 sky130_fd_sc_hd__o21ai_0 _12898_ (.A1(net4237),
    .A2(_03730_),
    .B1(_03889_),
    .Y(_00325_));
 sky130_fd_sc_hd__nand2_1 _12899_ (.A(net4237),
    .B(net104),
    .Y(_03890_));
 sky130_fd_sc_hd__o21ai_0 _12900_ (.A1(net4237),
    .A2(_03739_),
    .B1(_03890_),
    .Y(_00326_));
 sky130_fd_sc_hd__nand2_1 _12901_ (.A(net4239),
    .B(net105),
    .Y(_03891_));
 sky130_fd_sc_hd__o21ai_0 _12902_ (.A1(net4239),
    .A2(_03746_),
    .B1(_03891_),
    .Y(_00327_));
 sky130_fd_sc_hd__xnor2_1 _12903_ (.A(net4155),
    .B(net4124),
    .Y(_03892_));
 sky130_fd_sc_hd__nand2_1 _12904_ (.A(net4235),
    .B(net107),
    .Y(_03893_));
 sky130_fd_sc_hd__o21ai_0 _12905_ (.A1(net4235),
    .A2(_03892_),
    .B1(_03893_),
    .Y(_00328_));
 sky130_fd_sc_hd__xnor2_1 _12906_ (.A(net4154),
    .B(net4123),
    .Y(_03894_));
 sky130_fd_sc_hd__nand2_1 _12907_ (.A(net4236),
    .B(net108),
    .Y(_03895_));
 sky130_fd_sc_hd__o21ai_0 _12908_ (.A1(net4236),
    .A2(_03894_),
    .B1(_03895_),
    .Y(_00329_));
 sky130_fd_sc_hd__xnor2_1 _12909_ (.A(\u0.w[1][18] ),
    .B(_03613_),
    .Y(_03896_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1282 ();
 sky130_fd_sc_hd__nand2_1 _12911_ (.A(net4236),
    .B(net109),
    .Y(_03898_));
 sky130_fd_sc_hd__o21ai_0 _12912_ (.A1(net4236),
    .A2(_03896_),
    .B1(_03898_),
    .Y(_00330_));
 sky130_fd_sc_hd__mux2_1 _12913_ (.A0(net4125),
    .A1(net110),
    .S(net4236),
    .X(_00331_));
 sky130_fd_sc_hd__nand2_1 _12914_ (.A(net4239),
    .B(net111),
    .Y(_03899_));
 sky130_fd_sc_hd__o21ai_0 _12915_ (.A1(net4239),
    .A2(_03607_),
    .B1(_03899_),
    .Y(_00333_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1281 ();
 sky130_fd_sc_hd__nand2_1 _12917_ (.A(net4240),
    .B(net112),
    .Y(_03901_));
 sky130_fd_sc_hd__o21ai_0 _12918_ (.A1(net4240),
    .A2(_03598_),
    .B1(_03901_),
    .Y(_00334_));
 sky130_fd_sc_hd__nand2_1 _12919_ (.A(net4240),
    .B(net113),
    .Y(_03902_));
 sky130_fd_sc_hd__o21ai_0 _12920_ (.A1(net4240),
    .A2(_03755_),
    .B1(_03902_),
    .Y(_00335_));
 sky130_fd_sc_hd__nand2_1 _12921_ (.A(net4240),
    .B(net114),
    .Y(_03903_));
 sky130_fd_sc_hd__o21ai_0 _12922_ (.A1(net4240),
    .A2(_03762_),
    .B1(_03903_),
    .Y(_00336_));
 sky130_fd_sc_hd__mux2_1 _12923_ (.A0(_03851_),
    .A1(net115),
    .S(net4235),
    .X(_00337_));
 sky130_fd_sc_hd__mux2_1 _12924_ (.A0(_03856_),
    .A1(net116),
    .S(net129),
    .X(_00338_));
 sky130_fd_sc_hd__mux2_1 _12925_ (.A0(_03859_),
    .A1(net118),
    .S(net129),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _12926_ (.A0(_03862_),
    .A1(net119),
    .S(net129),
    .X(_00340_));
 sky130_fd_sc_hd__mux2_1 _12927_ (.A0(_03866_),
    .A1(net120),
    .S(net4232),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_1 _12928_ (.A0(_03806_),
    .A1(net121),
    .S(net4236),
    .X(_00342_));
 sky130_fd_sc_hd__xnor2_1 _12929_ (.A(\u0.w[1][30] ),
    .B(_03813_),
    .Y(_03904_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1280 ();
 sky130_fd_sc_hd__mux2_1 _12931_ (.A0(_03904_),
    .A1(net122),
    .S(net4235),
    .X(_00344_));
 sky130_fd_sc_hd__mux2_1 _12932_ (.A0(_03820_),
    .A1(net123),
    .S(net4236),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _12933_ (.A0(_03620_),
    .A1(net124),
    .S(net4235),
    .X(_00289_));
 sky130_fd_sc_hd__mux2_1 _12934_ (.A0(_03626_),
    .A1(net125),
    .S(net129),
    .X(_00300_));
 sky130_fd_sc_hd__xor2_1 _12935_ (.A(\u0.subword[2] ),
    .B(\u0.w[0][2] ),
    .X(_03906_));
 sky130_fd_sc_hd__mux2_1 _12936_ (.A0(_03906_),
    .A1(net126),
    .S(net4236),
    .X(_00311_));
 sky130_fd_sc_hd__xor2_1 _12937_ (.A(net4163),
    .B(\u0.subword[3] ),
    .X(_03907_));
 sky130_fd_sc_hd__mux2_1 _12938_ (.A0(_03907_),
    .A1(net127),
    .S(net4235),
    .X(_00314_));
 sky130_fd_sc_hd__xor2_1 _12939_ (.A(\u0.w[0][4] ),
    .B(\u0.subword[4] ),
    .X(_03908_));
 sky130_fd_sc_hd__mux2_1 _12940_ (.A0(_03908_),
    .A1(net2),
    .S(net4235),
    .X(_00315_));
 sky130_fd_sc_hd__xor2_1 _12941_ (.A(net4161),
    .B(\u0.subword[5] ),
    .X(_03909_));
 sky130_fd_sc_hd__mux2_1 _12942_ (.A0(_03909_),
    .A1(net3),
    .S(net4236),
    .X(_00316_));
 sky130_fd_sc_hd__xor2_1 _12943_ (.A(net4160),
    .B(\u0.subword[6] ),
    .X(_03910_));
 sky130_fd_sc_hd__mux2_1 _12944_ (.A0(_03910_),
    .A1(net4),
    .S(net4236),
    .X(_00317_));
 sky130_fd_sc_hd__mux2_1 _12945_ (.A0(_03679_),
    .A1(net5),
    .S(net4235),
    .X(_00318_));
 sky130_fd_sc_hd__xor2_1 _12946_ (.A(\u0.w[0][8] ),
    .B(\u0.subword[8] ),
    .X(_03911_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1279 ();
 sky130_fd_sc_hd__mux2_1 _12948_ (.A0(_03911_),
    .A1(net6),
    .S(net4240),
    .X(_00319_));
 sky130_fd_sc_hd__xor2_1 _12949_ (.A(net4158),
    .B(\u0.subword[9] ),
    .X(_03913_));
 sky130_fd_sc_hd__mux2_1 _12950_ (.A0(_03913_),
    .A1(net7),
    .S(net4236),
    .X(_00320_));
 sky130_fd_sc_hd__xor2_1 _12951_ (.A(\u0.subword[10] ),
    .B(\u0.w[0][10] ),
    .X(_03914_));
 sky130_fd_sc_hd__mux2_1 _12952_ (.A0(_03914_),
    .A1(net8),
    .S(net4237),
    .X(_00290_));
 sky130_fd_sc_hd__xor2_1 _12953_ (.A(net4177),
    .B(\u0.subword[11] ),
    .X(_03915_));
 sky130_fd_sc_hd__mux2_1 _12954_ (.A0(_03915_),
    .A1(net9),
    .S(net4238),
    .X(_00291_));
 sky130_fd_sc_hd__xor2_1 _12955_ (.A(net4176),
    .B(\u0.subword[12] ),
    .X(_03916_));
 sky130_fd_sc_hd__mux2_1 _12956_ (.A0(_03916_),
    .A1(net10),
    .S(net4238),
    .X(_00292_));
 sky130_fd_sc_hd__xor2_1 _12957_ (.A(net4175),
    .B(\u0.subword[13] ),
    .X(_03917_));
 sky130_fd_sc_hd__mux2_1 _12958_ (.A0(_03917_),
    .A1(net11),
    .S(net4237),
    .X(_00293_));
 sky130_fd_sc_hd__xor2_1 _12959_ (.A(net4174),
    .B(\u0.subword[14] ),
    .X(_03918_));
 sky130_fd_sc_hd__mux2_1 _12960_ (.A0(_03918_),
    .A1(net13),
    .S(net4237),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _12961_ (.A0(_03745_),
    .A1(net14),
    .S(net4239),
    .X(_00295_));
 sky130_fd_sc_hd__mux2_1 _12962_ (.A0(net4124),
    .A1(net15),
    .S(net4237),
    .X(_00296_));
 sky130_fd_sc_hd__mux2_1 _12963_ (.A0(net4123),
    .A1(net16),
    .S(net4238),
    .X(_00297_));
 sky130_fd_sc_hd__mux2_1 _12964_ (.A0(_03613_),
    .A1(net17),
    .S(net4239),
    .X(_00298_));
 sky130_fd_sc_hd__xor2_1 _12965_ (.A(\u0.w[0][19] ),
    .B(\u0.subword[19] ),
    .X(_03919_));
 sky130_fd_sc_hd__mux2_1 _12966_ (.A0(_03919_),
    .A1(net18),
    .S(net4236),
    .X(_00299_));
 sky130_fd_sc_hd__xor2_1 _12967_ (.A(\u0.w[0][20] ),
    .B(\u0.subword[20] ),
    .X(_03920_));
 sky130_fd_sc_hd__mux2_1 _12968_ (.A0(_03920_),
    .A1(net19),
    .S(net4239),
    .X(_00301_));
 sky130_fd_sc_hd__xor2_1 _12969_ (.A(net4172),
    .B(\u0.subword[21] ),
    .X(_03921_));
 sky130_fd_sc_hd__mux2_1 _12970_ (.A0(_03921_),
    .A1(net20),
    .S(net4240),
    .X(_00302_));
 sky130_fd_sc_hd__xor2_1 _12971_ (.A(net4171),
    .B(\u0.subword[22] ),
    .X(_03922_));
 sky130_fd_sc_hd__mux2_1 _12972_ (.A0(_03922_),
    .A1(net21),
    .S(net4240),
    .X(_00303_));
 sky130_fd_sc_hd__mux2_1 _12973_ (.A0(_03761_),
    .A1(net22),
    .S(net4240),
    .X(_00304_));
 sky130_fd_sc_hd__nand2_1 _12974_ (.A(net4235),
    .B(net24),
    .Y(_03923_));
 sky130_fd_sc_hd__o21ai_0 _12975_ (.A1(net4235),
    .A2(_03769_),
    .B1(_03923_),
    .Y(_00305_));
 sky130_fd_sc_hd__nand2_1 _12976_ (.A(net129),
    .B(net25),
    .Y(_03924_));
 sky130_fd_sc_hd__o21ai_0 _12977_ (.A1(net129),
    .A2(_03774_),
    .B1(_03924_),
    .Y(_00306_));
 sky130_fd_sc_hd__nand2_1 _12978_ (.A(net4235),
    .B(net26),
    .Y(_03925_));
 sky130_fd_sc_hd__o21ai_0 _12979_ (.A1(net4235),
    .A2(_03779_),
    .B1(_03925_),
    .Y(_00307_));
 sky130_fd_sc_hd__nand2_1 _12980_ (.A(net4235),
    .B(net27),
    .Y(_03926_));
 sky130_fd_sc_hd__o21ai_0 _12981_ (.A1(net4235),
    .A2(_03787_),
    .B1(_03926_),
    .Y(_00308_));
 sky130_fd_sc_hd__nand2_1 _12982_ (.A(net4235),
    .B(net28),
    .Y(_03927_));
 sky130_fd_sc_hd__o21ai_0 _12983_ (.A1(net4235),
    .A2(_03796_),
    .B1(_03927_),
    .Y(_00309_));
 sky130_fd_sc_hd__xor2_1 _12984_ (.A(\u0.r0.out[29] ),
    .B(_03805_),
    .X(_03928_));
 sky130_fd_sc_hd__nand2_1 _12985_ (.A(net4236),
    .B(net29),
    .Y(_03929_));
 sky130_fd_sc_hd__o21ai_0 _12986_ (.A1(net4236),
    .A2(_03928_),
    .B1(_03929_),
    .Y(_00310_));
 sky130_fd_sc_hd__nand2_1 _12987_ (.A(net4235),
    .B(net30),
    .Y(_03930_));
 sky130_fd_sc_hd__o21ai_0 _12988_ (.A1(net4235),
    .A2(_03813_),
    .B1(_03930_),
    .Y(_00312_));
 sky130_fd_sc_hd__nand2_1 _12989_ (.A(net4236),
    .B(net31),
    .Y(_03931_));
 sky130_fd_sc_hd__o21ai_0 _12990_ (.A1(net4236),
    .A2(_03819_),
    .B1(_03931_),
    .Y(_00313_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1266 ();
 sky130_fd_sc_hd__nand2_4 _13004_ (.A(_03593_),
    .B(net4101),
    .Y(_03942_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1265 ();
 sky130_fd_sc_hd__clkinvlp_4 _13006_ (.A(_11829_[0]),
    .Y(_03944_));
 sky130_fd_sc_hd__nand2_8 _13007_ (.A(_03944_),
    .B(net4102),
    .Y(_03945_));
 sky130_fd_sc_hd__a21oi_1 _13008_ (.A1(net4107),
    .A2(_03593_),
    .B1(_03945_),
    .Y(_03946_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1263 ();
 sky130_fd_sc_hd__a311oi_1 _13011_ (.A1(_11829_[0]),
    .A2(net4107),
    .A3(_03942_),
    .B1(_03946_),
    .C1(_03610_),
    .Y(_03949_));
 sky130_fd_sc_hd__nor2_4 _13012_ (.A(net4108),
    .B(net4102),
    .Y(_03950_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1262 ();
 sky130_fd_sc_hd__nand2_4 _13014_ (.A(net4107),
    .B(_03617_),
    .Y(_03952_));
 sky130_fd_sc_hd__nor2_2 _13015_ (.A(_11838_[0]),
    .B(_03952_),
    .Y(_03953_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1261 ();
 sky130_fd_sc_hd__nor2_4 _13017_ (.A(_03579_),
    .B(net4101),
    .Y(_03955_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1260 ();
 sky130_fd_sc_hd__nor2_4 _13019_ (.A(_03578_),
    .B(_03618_),
    .Y(_03957_));
 sky130_fd_sc_hd__nor2_2 _13020_ (.A(_03955_),
    .B(_03957_),
    .Y(_03958_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1259 ();
 sky130_fd_sc_hd__o21ai_0 _13022_ (.A1(_11842_[0]),
    .A2(_03958_),
    .B1(net4103),
    .Y(_03960_));
 sky130_fd_sc_hd__a211oi_1 _13023_ (.A1(_11829_[0]),
    .A2(_03950_),
    .B1(_03953_),
    .C1(_03960_),
    .Y(_03961_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1257 ();
 sky130_fd_sc_hd__o21ai_0 _13026_ (.A1(_03949_),
    .A2(_03961_),
    .B1(_03758_),
    .Y(_03964_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1256 ();
 sky130_fd_sc_hd__nand2_8 _13028_ (.A(_11833_[0]),
    .B(net4100),
    .Y(_03966_));
 sky130_fd_sc_hd__nand2_4 _13029_ (.A(_03593_),
    .B(_03618_),
    .Y(_03967_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1255 ();
 sky130_fd_sc_hd__nor2_4 _13031_ (.A(net4106),
    .B(_03618_),
    .Y(_03969_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1253 ();
 sky130_fd_sc_hd__nor2_2 _13034_ (.A(_11830_[0]),
    .B(net4101),
    .Y(_03972_));
 sky130_fd_sc_hd__nor3_1 _13035_ (.A(net4108),
    .B(_03969_),
    .C(_03972_),
    .Y(_03973_));
 sky130_fd_sc_hd__a311oi_2 _13036_ (.A1(net4108),
    .A2(_03966_),
    .A3(_03967_),
    .B1(_03973_),
    .C1(net4103),
    .Y(_03974_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1251 ();
 sky130_fd_sc_hd__nand2_8 _13039_ (.A(_03586_),
    .B(net4101),
    .Y(_03977_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1249 ();
 sky130_fd_sc_hd__nand2_8 _13042_ (.A(_11828_[0]),
    .B(_03618_),
    .Y(_03980_));
 sky130_fd_sc_hd__nand3_1 _13043_ (.A(_03579_),
    .B(_03977_),
    .C(_03980_),
    .Y(_03981_));
 sky130_fd_sc_hd__nand2_4 _13044_ (.A(_03610_),
    .B(_03981_),
    .Y(_03982_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1248 ();
 sky130_fd_sc_hd__nand2_1 _13046_ (.A(_11844_[0]),
    .B(_03618_),
    .Y(_03984_));
 sky130_fd_sc_hd__a21oi_1 _13047_ (.A1(_03942_),
    .A2(_03984_),
    .B1(_03579_),
    .Y(_03985_));
 sky130_fd_sc_hd__nor2_1 _13048_ (.A(_03982_),
    .B(_03985_),
    .Y(_03986_));
 sky130_fd_sc_hd__o21ai_0 _13049_ (.A1(_03974_),
    .A2(_03986_),
    .B1(_03759_),
    .Y(_03987_));
 sky130_fd_sc_hd__nand3_1 _13050_ (.A(_03766_),
    .B(_03964_),
    .C(_03987_),
    .Y(_03988_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1246 ();
 sky130_fd_sc_hd__nor2_1 _13053_ (.A(net4069),
    .B(_03759_),
    .Y(_03991_));
 sky130_fd_sc_hd__a21oi_1 _13054_ (.A1(_03759_),
    .A2(_03950_),
    .B1(_03991_),
    .Y(_03992_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1244 ();
 sky130_fd_sc_hd__nand2_1 _13057_ (.A(net4069),
    .B(_03758_),
    .Y(_03995_));
 sky130_fd_sc_hd__nand2_8 _13058_ (.A(_11840_[0]),
    .B(_03618_),
    .Y(_03996_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1243 ();
 sky130_fd_sc_hd__o21ai_0 _13060_ (.A1(_11835_[0]),
    .A2(_03758_),
    .B1(net4101),
    .Y(_03998_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1241 ();
 sky130_fd_sc_hd__o211ai_1 _13063_ (.A1(_03758_),
    .A2(_03996_),
    .B1(_03998_),
    .C1(net4108),
    .Y(_04001_));
 sky130_fd_sc_hd__o221ai_1 _13064_ (.A1(_11829_[0]),
    .A2(_03992_),
    .B1(_03995_),
    .B2(_11854_[0]),
    .C1(_04001_),
    .Y(_04002_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1240 ();
 sky130_fd_sc_hd__nand2_8 _13066_ (.A(_11842_[0]),
    .B(_03618_),
    .Y(_04004_));
 sky130_fd_sc_hd__nor2_1 _13067_ (.A(_11833_[0]),
    .B(net4101),
    .Y(_04005_));
 sky130_fd_sc_hd__nor2_1 _13068_ (.A(_03969_),
    .B(_04005_),
    .Y(_04006_));
 sky130_fd_sc_hd__nor2_1 _13069_ (.A(net4069),
    .B(_04006_),
    .Y(_04007_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1239 ();
 sky130_fd_sc_hd__a311oi_1 _13071_ (.A1(net4069),
    .A2(_03977_),
    .A3(_04004_),
    .B1(_04007_),
    .C1(_03611_),
    .Y(_04009_));
 sky130_fd_sc_hd__a311oi_1 _13072_ (.A1(_11835_[0]),
    .A2(net4108),
    .A3(net4101),
    .B1(_03758_),
    .C1(_03982_),
    .Y(_04010_));
 sky130_fd_sc_hd__a221oi_1 _13073_ (.A1(_03611_),
    .A2(_04002_),
    .B1(_04009_),
    .B2(_03758_),
    .C1(_04010_),
    .Y(_04011_));
 sky130_fd_sc_hd__nand2_1 _13074_ (.A(_03767_),
    .B(_04011_),
    .Y(_04012_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1238 ();
 sky130_fd_sc_hd__o211ai_1 _13076_ (.A1(_11835_[0]),
    .A2(net4100),
    .B1(_03966_),
    .C1(net4067),
    .Y(_04014_));
 sky130_fd_sc_hd__nand2_1 _13077_ (.A(_03578_),
    .B(_03977_),
    .Y(_04015_));
 sky130_fd_sc_hd__nor2_4 _13078_ (.A(_03944_),
    .B(net4101),
    .Y(_04016_));
 sky130_fd_sc_hd__nor2_2 _13079_ (.A(_11828_[0]),
    .B(_03618_),
    .Y(_04017_));
 sky130_fd_sc_hd__or3_1 _13080_ (.A(_03579_),
    .B(_04016_),
    .C(_04017_),
    .X(_04018_));
 sky130_fd_sc_hd__nand2b_4 _13081_ (.A_N(_11842_[0]),
    .B(_03617_),
    .Y(_04019_));
 sky130_fd_sc_hd__o211ai_1 _13082_ (.A1(_11838_[0]),
    .A2(net4100),
    .B1(_04019_),
    .C1(_03579_),
    .Y(_04020_));
 sky130_fd_sc_hd__a21oi_1 _13083_ (.A1(_04018_),
    .A2(_04020_),
    .B1(_03759_),
    .Y(_04021_));
 sky130_fd_sc_hd__a311o_1 _13084_ (.A1(_03759_),
    .A2(_04014_),
    .A3(_04015_),
    .B1(_04021_),
    .C1(_03611_),
    .X(_04022_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1237 ();
 sky130_fd_sc_hd__nand2_8 _13086_ (.A(_03944_),
    .B(_03618_),
    .Y(_04024_));
 sky130_fd_sc_hd__clkinv_2 _13087_ (.A(_11830_[0]),
    .Y(_04025_));
 sky130_fd_sc_hd__nand2_4 _13088_ (.A(_04025_),
    .B(net4100),
    .Y(_04026_));
 sky130_fd_sc_hd__nand2_1 _13089_ (.A(_04024_),
    .B(_04026_),
    .Y(_04027_));
 sky130_fd_sc_hd__nand2_8 _13090_ (.A(_03586_),
    .B(_03618_),
    .Y(_04028_));
 sky130_fd_sc_hd__a21oi_1 _13091_ (.A1(_03966_),
    .A2(_04028_),
    .B1(net4069),
    .Y(_04029_));
 sky130_fd_sc_hd__a211oi_1 _13092_ (.A1(net4068),
    .A2(_04027_),
    .B1(_04029_),
    .C1(_03758_),
    .Y(_04030_));
 sky130_fd_sc_hd__nand2_2 _13093_ (.A(net4106),
    .B(net4100),
    .Y(_04031_));
 sky130_fd_sc_hd__nand2_4 _13094_ (.A(_03586_),
    .B(net4105),
    .Y(_04032_));
 sky130_fd_sc_hd__a21o_1 _13095_ (.A1(_04031_),
    .A2(_04032_),
    .B1(net4068),
    .X(_04033_));
 sky130_fd_sc_hd__nand3_1 _13096_ (.A(net4068),
    .B(_04031_),
    .C(_04032_),
    .Y(_04034_));
 sky130_fd_sc_hd__a21oi_1 _13097_ (.A1(_04033_),
    .A2(_04034_),
    .B1(_03759_),
    .Y(_04035_));
 sky130_fd_sc_hd__o21ai_0 _13098_ (.A1(_04030_),
    .A2(_04035_),
    .B1(_03611_),
    .Y(_04036_));
 sky130_fd_sc_hd__a21oi_1 _13099_ (.A1(_04022_),
    .A2(_04036_),
    .B1(_03767_),
    .Y(_04037_));
 sky130_fd_sc_hd__nor2_4 _13100_ (.A(_11829_[0]),
    .B(_03618_),
    .Y(_04038_));
 sky130_fd_sc_hd__nor2_4 _13101_ (.A(net4105),
    .B(net4100),
    .Y(_04039_));
 sky130_fd_sc_hd__o21ai_2 _13102_ (.A1(_04038_),
    .A2(_04039_),
    .B1(net4108),
    .Y(_04040_));
 sky130_fd_sc_hd__nor2_4 _13103_ (.A(_03586_),
    .B(_03617_),
    .Y(_04041_));
 sky130_fd_sc_hd__nor2_1 _13104_ (.A(_11838_[0]),
    .B(_03618_),
    .Y(_04042_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1236 ();
 sky130_fd_sc_hd__o21ai_0 _13106_ (.A1(_04041_),
    .A2(_04042_),
    .B1(net4069),
    .Y(_04044_));
 sky130_fd_sc_hd__and2_4 _13107_ (.A(_11833_[0]),
    .B(_03618_),
    .X(_04045_));
 sky130_fd_sc_hd__nor2_4 _13108_ (.A(_11840_[0]),
    .B(_03618_),
    .Y(_04046_));
 sky130_fd_sc_hd__nor3_1 _13109_ (.A(net4108),
    .B(_04045_),
    .C(_04046_),
    .Y(_04047_));
 sky130_fd_sc_hd__a211oi_1 _13110_ (.A1(_11844_[0]),
    .A2(_03955_),
    .B1(_04047_),
    .C1(_03759_),
    .Y(_04048_));
 sky130_fd_sc_hd__a311oi_1 _13111_ (.A1(_03759_),
    .A2(_04040_),
    .A3(_04044_),
    .B1(_04048_),
    .C1(_03611_),
    .Y(_04049_));
 sky130_fd_sc_hd__o21ai_0 _13112_ (.A1(_04005_),
    .A2(_04042_),
    .B1(net4108),
    .Y(_04050_));
 sky130_fd_sc_hd__a21oi_1 _13113_ (.A1(_11844_[0]),
    .A2(_03950_),
    .B1(_03759_),
    .Y(_04051_));
 sky130_fd_sc_hd__nand2_2 _13114_ (.A(_03579_),
    .B(_03618_),
    .Y(_04052_));
 sky130_fd_sc_hd__nor2_1 _13115_ (.A(_11844_[0]),
    .B(net4101),
    .Y(_04053_));
 sky130_fd_sc_hd__a21oi_1 _13116_ (.A1(_11842_[0]),
    .A2(net4101),
    .B1(_04053_),
    .Y(_04054_));
 sky130_fd_sc_hd__o22ai_1 _13117_ (.A1(_11835_[0]),
    .A2(_04052_),
    .B1(_04054_),
    .B2(_03579_),
    .Y(_04055_));
 sky130_fd_sc_hd__a221oi_1 _13118_ (.A1(_04050_),
    .A2(_04051_),
    .B1(_04055_),
    .B2(_03759_),
    .C1(_03610_),
    .Y(_04056_));
 sky130_fd_sc_hd__o21a_1 _13119_ (.A1(_04049_),
    .A2(_04056_),
    .B1(_03767_),
    .X(_04057_));
 sky130_fd_sc_hd__nor3_1 _13120_ (.A(net4066),
    .B(_04037_),
    .C(_04057_),
    .Y(_04058_));
 sky130_fd_sc_hd__a31oi_1 _13121_ (.A1(net4066),
    .A2(_03988_),
    .A3(_04012_),
    .B1(_04058_),
    .Y(_00000_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1235 ();
 sky130_fd_sc_hd__nand2_8 _13123_ (.A(_11829_[0]),
    .B(_03618_),
    .Y(_04060_));
 sky130_fd_sc_hd__nand2b_4 _13124_ (.A_N(_11835_[0]),
    .B(net4101),
    .Y(_04061_));
 sky130_fd_sc_hd__and3_1 _13125_ (.A(net4108),
    .B(_03977_),
    .C(_04004_),
    .X(_04062_));
 sky130_fd_sc_hd__a311oi_1 _13126_ (.A1(_03579_),
    .A2(_04060_),
    .A3(_04061_),
    .B1(_04062_),
    .C1(_03758_),
    .Y(_04063_));
 sky130_fd_sc_hd__nand2_1 _13127_ (.A(_11847_[0]),
    .B(net4069),
    .Y(_04064_));
 sky130_fd_sc_hd__nand2_4 _13128_ (.A(_11835_[0]),
    .B(net4100),
    .Y(_04065_));
 sky130_fd_sc_hd__nand3_1 _13129_ (.A(net4108),
    .B(_03967_),
    .C(_04065_),
    .Y(_04066_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1234 ();
 sky130_fd_sc_hd__a21oi_1 _13131_ (.A1(_04064_),
    .A2(_04066_),
    .B1(_03759_),
    .Y(_04068_));
 sky130_fd_sc_hd__o21ai_0 _13132_ (.A1(_04063_),
    .A2(_04068_),
    .B1(_03611_),
    .Y(_04069_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1233 ();
 sky130_fd_sc_hd__nand2_1 _13134_ (.A(net4106),
    .B(net4105),
    .Y(_04071_));
 sky130_fd_sc_hd__nand3_1 _13135_ (.A(_03579_),
    .B(_04028_),
    .C(_04071_),
    .Y(_04072_));
 sky130_fd_sc_hd__o31ai_1 _13136_ (.A1(_03579_),
    .A2(_04041_),
    .A3(_04038_),
    .B1(_04072_),
    .Y(_04073_));
 sky130_fd_sc_hd__nand2_4 _13137_ (.A(_04025_),
    .B(_03618_),
    .Y(_04074_));
 sky130_fd_sc_hd__a31oi_1 _13138_ (.A1(_03579_),
    .A2(_03945_),
    .A3(_04074_),
    .B1(_03759_),
    .Y(_04075_));
 sky130_fd_sc_hd__nand2_4 _13139_ (.A(_11833_[0]),
    .B(_03618_),
    .Y(_04076_));
 sky130_fd_sc_hd__a31oi_2 _13140_ (.A1(net4108),
    .A2(_04076_),
    .A3(_04061_),
    .B1(_03611_),
    .Y(_04077_));
 sky130_fd_sc_hd__a32oi_1 _13141_ (.A1(_03610_),
    .A2(_03759_),
    .A3(_04073_),
    .B1(_04075_),
    .B2(_04077_),
    .Y(_04078_));
 sky130_fd_sc_hd__nand2_4 _13142_ (.A(_11835_[0]),
    .B(_03618_),
    .Y(_04079_));
 sky130_fd_sc_hd__a21oi_1 _13143_ (.A1(_03977_),
    .A2(_04024_),
    .B1(net4108),
    .Y(_04080_));
 sky130_fd_sc_hd__a31oi_1 _13144_ (.A1(net4108),
    .A2(_03977_),
    .A3(_04079_),
    .B1(_04080_),
    .Y(_04081_));
 sky130_fd_sc_hd__nand2_2 _13145_ (.A(_03578_),
    .B(_03618_),
    .Y(_04082_));
 sky130_fd_sc_hd__nand3_1 _13146_ (.A(net4069),
    .B(_04026_),
    .C(_03967_),
    .Y(_04083_));
 sky130_fd_sc_hd__o211ai_1 _13147_ (.A1(_11828_[0]),
    .A2(_04082_),
    .B1(_04083_),
    .C1(_03759_),
    .Y(_04084_));
 sky130_fd_sc_hd__o21ai_0 _13148_ (.A1(_03759_),
    .A2(_04081_),
    .B1(_04084_),
    .Y(_04085_));
 sky130_fd_sc_hd__nand2_1 _13149_ (.A(_11835_[0]),
    .B(_03955_),
    .Y(_04086_));
 sky130_fd_sc_hd__nand2_4 _13150_ (.A(_11828_[0]),
    .B(net4101),
    .Y(_04087_));
 sky130_fd_sc_hd__nand3_1 _13151_ (.A(_03579_),
    .B(_04060_),
    .C(_04087_),
    .Y(_04088_));
 sky130_fd_sc_hd__nand3_1 _13152_ (.A(_03759_),
    .B(_04086_),
    .C(_04088_),
    .Y(_04089_));
 sky130_fd_sc_hd__nand2_4 _13153_ (.A(net4067),
    .B(net4100),
    .Y(_04090_));
 sky130_fd_sc_hd__nor2_2 _13154_ (.A(_03593_),
    .B(_03618_),
    .Y(_04091_));
 sky130_fd_sc_hd__nor2_1 _13155_ (.A(_03586_),
    .B(net4105),
    .Y(_04092_));
 sky130_fd_sc_hd__o21ai_2 _13156_ (.A1(_04091_),
    .A2(_04092_),
    .B1(net4107),
    .Y(_04093_));
 sky130_fd_sc_hd__o211ai_1 _13157_ (.A1(_11833_[0]),
    .A2(_04090_),
    .B1(_04093_),
    .C1(_03758_),
    .Y(_04094_));
 sky130_fd_sc_hd__a21oi_1 _13158_ (.A1(_04089_),
    .A2(_04094_),
    .B1(_03611_),
    .Y(_04095_));
 sky130_fd_sc_hd__a211oi_1 _13159_ (.A1(_03611_),
    .A2(_04085_),
    .B1(_04095_),
    .C1(net4066),
    .Y(_04096_));
 sky130_fd_sc_hd__a31oi_2 _13160_ (.A1(net4066),
    .A2(_04069_),
    .A3(_04078_),
    .B1(_04096_),
    .Y(_04097_));
 sky130_fd_sc_hd__nand2_4 _13161_ (.A(net4105),
    .B(_03617_),
    .Y(_04098_));
 sky130_fd_sc_hd__and3_4 _13162_ (.A(_03579_),
    .B(_04098_),
    .C(_04079_),
    .X(_04099_));
 sky130_fd_sc_hd__a31oi_1 _13163_ (.A1(_03578_),
    .A2(_04019_),
    .A3(_04028_),
    .B1(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__nand3_1 _13164_ (.A(_03579_),
    .B(_03945_),
    .C(_04004_),
    .Y(_04101_));
 sky130_fd_sc_hd__o311ai_0 _13165_ (.A1(_03579_),
    .A2(_03969_),
    .A3(_04053_),
    .B1(_04101_),
    .C1(_03611_),
    .Y(_04102_));
 sky130_fd_sc_hd__o21ai_0 _13166_ (.A1(_03611_),
    .A2(_04100_),
    .B1(_04102_),
    .Y(_04103_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1232 ();
 sky130_fd_sc_hd__nand2_1 _13168_ (.A(_03977_),
    .B(_03980_),
    .Y(_04105_));
 sky130_fd_sc_hd__nand2_1 _13169_ (.A(net4108),
    .B(_04105_),
    .Y(_04106_));
 sky130_fd_sc_hd__a21oi_1 _13170_ (.A1(_03944_),
    .A2(_03950_),
    .B1(_03611_),
    .Y(_04107_));
 sky130_fd_sc_hd__o211ai_1 _13171_ (.A1(_11844_[0]),
    .A2(_03618_),
    .B1(_04074_),
    .C1(net4108),
    .Y(_04108_));
 sky130_fd_sc_hd__a21oi_1 _13172_ (.A1(_04088_),
    .A2(_04108_),
    .B1(_03610_),
    .Y(_04109_));
 sky130_fd_sc_hd__a211oi_1 _13173_ (.A1(_04106_),
    .A2(_04107_),
    .B1(_04109_),
    .C1(_03602_),
    .Y(_04110_));
 sky130_fd_sc_hd__a211oi_1 _13174_ (.A1(_03602_),
    .A2(_04103_),
    .B1(_04110_),
    .C1(_03758_),
    .Y(_04111_));
 sky130_fd_sc_hd__nor2_1 _13175_ (.A(_11842_[0]),
    .B(_03618_),
    .Y(_04112_));
 sky130_fd_sc_hd__nor3_1 _13176_ (.A(_03579_),
    .B(_04112_),
    .C(_04041_),
    .Y(_04113_));
 sky130_fd_sc_hd__nor2_2 _13177_ (.A(_11833_[0]),
    .B(_03618_),
    .Y(_04114_));
 sky130_fd_sc_hd__nor2_1 _13178_ (.A(_11828_[0]),
    .B(net4100),
    .Y(_04115_));
 sky130_fd_sc_hd__nor3_1 _13179_ (.A(net4107),
    .B(_04114_),
    .C(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__o21ai_1 _13180_ (.A1(_04113_),
    .A2(_04116_),
    .B1(_03602_),
    .Y(_04117_));
 sky130_fd_sc_hd__nand2_8 _13181_ (.A(net4106),
    .B(_03618_),
    .Y(_04118_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1231 ();
 sky130_fd_sc_hd__a21oi_1 _13183_ (.A1(_04118_),
    .A2(_04098_),
    .B1(_03579_),
    .Y(_04120_));
 sky130_fd_sc_hd__o21ai_0 _13184_ (.A1(_04099_),
    .A2(_04120_),
    .B1(_03601_),
    .Y(_04121_));
 sky130_fd_sc_hd__nand2_4 _13185_ (.A(_11838_[0]),
    .B(_03617_),
    .Y(_04122_));
 sky130_fd_sc_hd__nor2_1 _13186_ (.A(_11856_[0]),
    .B(net4107),
    .Y(_04123_));
 sky130_fd_sc_hd__a32oi_1 _13187_ (.A1(net4107),
    .A2(_04122_),
    .A3(_03980_),
    .B1(_04123_),
    .B2(_03601_),
    .Y(_04124_));
 sky130_fd_sc_hd__nor2_1 _13188_ (.A(_03611_),
    .B(_04124_),
    .Y(_04125_));
 sky130_fd_sc_hd__a31oi_1 _13189_ (.A1(_03611_),
    .A2(_04117_),
    .A3(_04121_),
    .B1(_04125_),
    .Y(_04126_));
 sky130_fd_sc_hd__nor2_1 _13190_ (.A(_03759_),
    .B(_04126_),
    .Y(_04127_));
 sky130_fd_sc_hd__nor3_1 _13191_ (.A(_03767_),
    .B(_04111_),
    .C(_04127_),
    .Y(_04128_));
 sky130_fd_sc_hd__a21oi_1 _13192_ (.A1(_03767_),
    .A2(_04097_),
    .B1(_04128_),
    .Y(_00001_));
 sky130_fd_sc_hd__nor2_4 _13193_ (.A(_03593_),
    .B(_03617_),
    .Y(_04129_));
 sky130_fd_sc_hd__nand2_2 _13194_ (.A(_11829_[0]),
    .B(_03617_),
    .Y(_04130_));
 sky130_fd_sc_hd__o211ai_1 _13195_ (.A1(_11838_[0]),
    .A2(_03617_),
    .B1(_04130_),
    .C1(_03579_),
    .Y(_04131_));
 sky130_fd_sc_hd__o311ai_0 _13196_ (.A1(_03579_),
    .A2(_04112_),
    .A3(_04129_),
    .B1(_04131_),
    .C1(_03759_),
    .Y(_04132_));
 sky130_fd_sc_hd__or3_4 _13197_ (.A(net4107),
    .B(_04114_),
    .C(_04039_),
    .X(_04133_));
 sky130_fd_sc_hd__o211ai_1 _13198_ (.A1(_11849_[0]),
    .A2(_03579_),
    .B1(_03758_),
    .C1(_04133_),
    .Y(_04134_));
 sky130_fd_sc_hd__nand2_1 _13199_ (.A(_11856_[0]),
    .B(net4107),
    .Y(_04135_));
 sky130_fd_sc_hd__or3_1 _13200_ (.A(net4107),
    .B(_04091_),
    .C(_04092_),
    .X(_04136_));
 sky130_fd_sc_hd__nor2_2 _13201_ (.A(_03579_),
    .B(_03966_),
    .Y(_04137_));
 sky130_fd_sc_hd__a211oi_1 _13202_ (.A1(_11852_[0]),
    .A2(_03579_),
    .B1(_03759_),
    .C1(_04137_),
    .Y(_04138_));
 sky130_fd_sc_hd__a311oi_1 _13203_ (.A1(_03759_),
    .A2(_04135_),
    .A3(_04136_),
    .B1(_04138_),
    .C1(_03611_),
    .Y(_04139_));
 sky130_fd_sc_hd__a31oi_1 _13204_ (.A1(_03611_),
    .A2(_04132_),
    .A3(_04134_),
    .B1(_04139_),
    .Y(_04140_));
 sky130_fd_sc_hd__nand2_1 _13205_ (.A(_03579_),
    .B(_04129_),
    .Y(_04141_));
 sky130_fd_sc_hd__nor2_4 _13206_ (.A(_03579_),
    .B(_03618_),
    .Y(_04142_));
 sky130_fd_sc_hd__a21oi_1 _13207_ (.A1(_04118_),
    .A2(_04065_),
    .B1(net4107),
    .Y(_04143_));
 sky130_fd_sc_hd__a211oi_1 _13208_ (.A1(_11830_[0]),
    .A2(_04142_),
    .B1(_04143_),
    .C1(_03610_),
    .Y(_04144_));
 sky130_fd_sc_hd__a31oi_1 _13209_ (.A1(_03610_),
    .A2(_04065_),
    .A3(_04141_),
    .B1(_04144_),
    .Y(_04145_));
 sky130_fd_sc_hd__o21ai_0 _13210_ (.A1(_03579_),
    .A2(_03996_),
    .B1(_03759_),
    .Y(_04146_));
 sky130_fd_sc_hd__o21ai_2 _13211_ (.A1(_11835_[0]),
    .A2(_03617_),
    .B1(_04026_),
    .Y(_04147_));
 sky130_fd_sc_hd__nand2_1 _13212_ (.A(net4107),
    .B(_04147_),
    .Y(_04148_));
 sky130_fd_sc_hd__a21oi_1 _13213_ (.A1(_04076_),
    .A2(_04061_),
    .B1(_03578_),
    .Y(_04149_));
 sky130_fd_sc_hd__nor2_1 _13214_ (.A(_03611_),
    .B(_04149_),
    .Y(_04150_));
 sky130_fd_sc_hd__a32o_1 _13215_ (.A1(_03611_),
    .A2(_04133_),
    .A3(_04148_),
    .B1(_04150_),
    .B2(_04040_),
    .X(_04151_));
 sky130_fd_sc_hd__o221a_1 _13216_ (.A1(_04145_),
    .A2(_04146_),
    .B1(_04151_),
    .B2(_03759_),
    .C1(_03766_),
    .X(_04152_));
 sky130_fd_sc_hd__a21oi_1 _13217_ (.A1(_03767_),
    .A2(_04140_),
    .B1(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__nand2_1 _13218_ (.A(_11840_[0]),
    .B(_03617_),
    .Y(_04154_));
 sky130_fd_sc_hd__nor3_2 _13219_ (.A(net4108),
    .B(_04016_),
    .C(_04038_),
    .Y(_04155_));
 sky130_fd_sc_hd__a31oi_1 _13220_ (.A1(net4107),
    .A2(_04118_),
    .A3(_04154_),
    .B1(_04155_),
    .Y(_04156_));
 sky130_fd_sc_hd__a21oi_1 _13221_ (.A1(_04074_),
    .A2(_04087_),
    .B1(_03578_),
    .Y(_04157_));
 sky130_fd_sc_hd__o21ai_0 _13222_ (.A1(_04137_),
    .A2(_04157_),
    .B1(_03758_),
    .Y(_04158_));
 sky130_fd_sc_hd__o21ai_0 _13223_ (.A1(_03758_),
    .A2(_04156_),
    .B1(_04158_),
    .Y(_04159_));
 sky130_fd_sc_hd__a21oi_1 _13224_ (.A1(_04060_),
    .A2(_03942_),
    .B1(net4069),
    .Y(_04160_));
 sky130_fd_sc_hd__nand2_4 _13225_ (.A(_11844_[0]),
    .B(net4101),
    .Y(_04161_));
 sky130_fd_sc_hd__a21oi_1 _13226_ (.A1(_04118_),
    .A2(_04161_),
    .B1(_03578_),
    .Y(_04162_));
 sky130_fd_sc_hd__a21oi_1 _13227_ (.A1(_04028_),
    .A2(_04026_),
    .B1(_03579_),
    .Y(_04163_));
 sky130_fd_sc_hd__a21oi_2 _13228_ (.A1(_03593_),
    .A2(net4101),
    .B1(net4108),
    .Y(_04164_));
 sky130_fd_sc_hd__and2_0 _13229_ (.A(_03996_),
    .B(_04164_),
    .X(_04165_));
 sky130_fd_sc_hd__o21ai_0 _13230_ (.A1(_04163_),
    .A2(_04165_),
    .B1(_03759_),
    .Y(_04166_));
 sky130_fd_sc_hd__o311ai_0 _13231_ (.A1(_03759_),
    .A2(_04160_),
    .A3(_04162_),
    .B1(_04166_),
    .C1(_03611_),
    .Y(_04167_));
 sky130_fd_sc_hd__o21ai_0 _13232_ (.A1(_03611_),
    .A2(_04159_),
    .B1(_04167_),
    .Y(_04168_));
 sky130_fd_sc_hd__o21ai_0 _13233_ (.A1(_11849_[0]),
    .A2(_04041_),
    .B1(_03579_),
    .Y(_04169_));
 sky130_fd_sc_hd__nor2_1 _13234_ (.A(_03578_),
    .B(_04028_),
    .Y(_04170_));
 sky130_fd_sc_hd__nor2_1 _13235_ (.A(_11828_[0]),
    .B(_03958_),
    .Y(_04171_));
 sky130_fd_sc_hd__nor4_1 _13236_ (.A(_03759_),
    .B(_03953_),
    .C(_04170_),
    .D(_04171_),
    .Y(_04172_));
 sky130_fd_sc_hd__a311oi_1 _13237_ (.A1(_03759_),
    .A2(_04040_),
    .A3(_04169_),
    .B1(_04172_),
    .C1(net4103),
    .Y(_04173_));
 sky130_fd_sc_hd__a21oi_1 _13238_ (.A1(_04060_),
    .A2(_04065_),
    .B1(net4108),
    .Y(_04174_));
 sky130_fd_sc_hd__nor2_1 _13239_ (.A(_11842_[0]),
    .B(_04082_),
    .Y(_04175_));
 sky130_fd_sc_hd__nand2_1 _13240_ (.A(_11854_[0]),
    .B(net4108),
    .Y(_04176_));
 sky130_fd_sc_hd__o311ai_0 _13241_ (.A1(net4108),
    .A2(_04045_),
    .A3(_04038_),
    .B1(_04176_),
    .C1(_03759_),
    .Y(_04177_));
 sky130_fd_sc_hd__o311ai_0 _13242_ (.A1(_03759_),
    .A2(_04174_),
    .A3(_04175_),
    .B1(_04177_),
    .C1(net4103),
    .Y(_04178_));
 sky130_fd_sc_hd__nand2_2 _13243_ (.A(_03767_),
    .B(_04178_),
    .Y(_04179_));
 sky130_fd_sc_hd__o221ai_1 _13244_ (.A1(_03767_),
    .A2(_04168_),
    .B1(_04173_),
    .B2(_04179_),
    .C1(_03602_),
    .Y(_04180_));
 sky130_fd_sc_hd__o21ai_1 _13245_ (.A1(_03602_),
    .A2(_04153_),
    .B1(_04180_),
    .Y(_00002_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1230 ();
 sky130_fd_sc_hd__a22oi_1 _13247_ (.A1(_03578_),
    .A2(_04041_),
    .B1(_03958_),
    .B2(_11840_[0]),
    .Y(_04182_));
 sky130_fd_sc_hd__a21oi_1 _13248_ (.A1(_04060_),
    .A2(_04031_),
    .B1(net4068),
    .Y(_04183_));
 sky130_fd_sc_hd__and3_1 _13249_ (.A(net4068),
    .B(_04118_),
    .C(_04026_),
    .X(_04184_));
 sky130_fd_sc_hd__o21ai_0 _13250_ (.A1(_04183_),
    .A2(_04184_),
    .B1(net4066),
    .Y(_04185_));
 sky130_fd_sc_hd__o211ai_1 _13251_ (.A1(net4066),
    .A2(_04182_),
    .B1(_04185_),
    .C1(net4103),
    .Y(_04186_));
 sky130_fd_sc_hd__nor2_1 _13252_ (.A(_03602_),
    .B(_04090_),
    .Y(_04187_));
 sky130_fd_sc_hd__a21oi_1 _13253_ (.A1(_03602_),
    .A2(_03955_),
    .B1(_04187_),
    .Y(_04188_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1229 ();
 sky130_fd_sc_hd__o211ai_1 _13255_ (.A1(_04039_),
    .A2(_04042_),
    .B1(net4108),
    .C1(net4066),
    .Y(_04190_));
 sky130_fd_sc_hd__nand2_1 _13256_ (.A(_11844_[0]),
    .B(_03950_),
    .Y(_04191_));
 sky130_fd_sc_hd__o2111ai_1 _13257_ (.A1(_11829_[0]),
    .A2(_04188_),
    .B1(_04190_),
    .C1(_04191_),
    .D1(_03611_),
    .Y(_04192_));
 sky130_fd_sc_hd__o32a_1 _13258_ (.A1(_11849_[0]),
    .A2(_03579_),
    .A3(_04041_),
    .B1(_04090_),
    .B2(_11829_[0]),
    .X(_04193_));
 sky130_fd_sc_hd__a21oi_1 _13259_ (.A1(_04118_),
    .A2(_04032_),
    .B1(net4068),
    .Y(_04194_));
 sky130_fd_sc_hd__a311oi_1 _13260_ (.A1(net4068),
    .A2(_04060_),
    .A3(_04098_),
    .B1(_04194_),
    .C1(_03611_),
    .Y(_04195_));
 sky130_fd_sc_hd__a21oi_1 _13261_ (.A1(_03611_),
    .A2(_04193_),
    .B1(_04195_),
    .Y(_04196_));
 sky130_fd_sc_hd__nand2_1 _13262_ (.A(_11838_[0]),
    .B(_03618_),
    .Y(_04197_));
 sky130_fd_sc_hd__and3_1 _13263_ (.A(_03578_),
    .B(_03977_),
    .C(_04197_),
    .X(_04198_));
 sky130_fd_sc_hd__a311o_1 _13264_ (.A1(net4069),
    .A2(_04004_),
    .A3(_04130_),
    .B1(_04198_),
    .C1(net4103),
    .X(_04199_));
 sky130_fd_sc_hd__a21oi_1 _13265_ (.A1(_04074_),
    .A2(_04061_),
    .B1(_03578_),
    .Y(_04200_));
 sky130_fd_sc_hd__o21ai_0 _13266_ (.A1(_04160_),
    .A2(_04200_),
    .B1(net4103),
    .Y(_04201_));
 sky130_fd_sc_hd__a21oi_1 _13267_ (.A1(_04199_),
    .A2(_04201_),
    .B1(net4066),
    .Y(_04202_));
 sky130_fd_sc_hd__a211oi_1 _13268_ (.A1(net4066),
    .A2(_04196_),
    .B1(_04202_),
    .C1(net3627),
    .Y(_04203_));
 sky130_fd_sc_hd__a31oi_1 _13269_ (.A1(net3627),
    .A2(_04186_),
    .A3(_04192_),
    .B1(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__and3_1 _13270_ (.A(_03579_),
    .B(_04028_),
    .C(_04154_),
    .X(_04205_));
 sky130_fd_sc_hd__a21oi_1 _13271_ (.A1(_04122_),
    .A2(_03980_),
    .B1(_03579_),
    .Y(_04206_));
 sky130_fd_sc_hd__o21a_1 _13272_ (.A1(_04205_),
    .A2(_04206_),
    .B1(net4103),
    .X(_04207_));
 sky130_fd_sc_hd__a211oi_1 _13273_ (.A1(_03611_),
    .A2(_04163_),
    .B1(_04207_),
    .C1(_03602_),
    .Y(_04208_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1228 ();
 sky130_fd_sc_hd__a21oi_1 _13275_ (.A1(_04024_),
    .A2(_04026_),
    .B1(net4069),
    .Y(_04210_));
 sky130_fd_sc_hd__a31oi_1 _13276_ (.A1(net4069),
    .A2(_03977_),
    .A3(_03996_),
    .B1(_04210_),
    .Y(_04211_));
 sky130_fd_sc_hd__o2111ai_1 _13277_ (.A1(_11842_[0]),
    .A2(_04052_),
    .B1(_04093_),
    .C1(net4103),
    .D1(_04031_),
    .Y(_04212_));
 sky130_fd_sc_hd__o21ai_0 _13278_ (.A1(net4103),
    .A2(_04211_),
    .B1(_04212_),
    .Y(_04213_));
 sky130_fd_sc_hd__nor2_1 _13279_ (.A(net4066),
    .B(_04213_),
    .Y(_04214_));
 sky130_fd_sc_hd__o21ai_0 _13280_ (.A1(_04208_),
    .A2(_04214_),
    .B1(net3627),
    .Y(_04215_));
 sky130_fd_sc_hd__a21oi_1 _13281_ (.A1(_11833_[0]),
    .A2(_03957_),
    .B1(_04194_),
    .Y(_04216_));
 sky130_fd_sc_hd__o311ai_0 _13282_ (.A1(net4069),
    .A2(_04016_),
    .A3(_04046_),
    .B1(_04083_),
    .C1(_03611_),
    .Y(_04217_));
 sky130_fd_sc_hd__o21ai_0 _13283_ (.A1(_03611_),
    .A2(_04216_),
    .B1(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__nand2_1 _13284_ (.A(_04060_),
    .B(_04122_),
    .Y(_04219_));
 sky130_fd_sc_hd__nand2_1 _13285_ (.A(_03578_),
    .B(_04219_),
    .Y(_04220_));
 sky130_fd_sc_hd__nand3_1 _13286_ (.A(net4108),
    .B(_03945_),
    .C(_03980_),
    .Y(_04221_));
 sky130_fd_sc_hd__nand3_1 _13287_ (.A(net4069),
    .B(_03966_),
    .C(_04197_),
    .Y(_04222_));
 sky130_fd_sc_hd__a21oi_1 _13288_ (.A1(_04221_),
    .A2(_04222_),
    .B1(_03611_),
    .Y(_04223_));
 sky130_fd_sc_hd__a311oi_1 _13289_ (.A1(_03611_),
    .A2(_04034_),
    .A3(_04220_),
    .B1(_04223_),
    .C1(net4066),
    .Y(_04224_));
 sky130_fd_sc_hd__a21oi_1 _13290_ (.A1(net4066),
    .A2(_04218_),
    .B1(_04224_),
    .Y(_04225_));
 sky130_fd_sc_hd__a21oi_1 _13291_ (.A1(_03767_),
    .A2(_04225_),
    .B1(_03758_),
    .Y(_04226_));
 sky130_fd_sc_hd__a22oi_1 _13292_ (.A1(_03758_),
    .A2(_04204_),
    .B1(_04215_),
    .B2(_04226_),
    .Y(_00003_));
 sky130_fd_sc_hd__nor3_1 _13293_ (.A(net4108),
    .B(_04041_),
    .C(_04046_),
    .Y(_04227_));
 sky130_fd_sc_hd__a31oi_1 _13294_ (.A1(net4108),
    .A2(_04032_),
    .A3(_03942_),
    .B1(_04227_),
    .Y(_04228_));
 sky130_fd_sc_hd__nand3_1 _13295_ (.A(net4108),
    .B(_03610_),
    .C(_04054_),
    .Y(_04229_));
 sky130_fd_sc_hd__o21ai_0 _13296_ (.A1(_11840_[0]),
    .A2(_03610_),
    .B1(_03586_),
    .Y(_04230_));
 sky130_fd_sc_hd__nand2_1 _13297_ (.A(net4101),
    .B(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__o2111ai_1 _13298_ (.A1(_03586_),
    .A2(_03610_),
    .B1(_04032_),
    .C1(_04231_),
    .D1(_03579_),
    .Y(_04232_));
 sky130_fd_sc_hd__o2111ai_1 _13299_ (.A1(_03610_),
    .A2(_04228_),
    .B1(_04229_),
    .C1(_03766_),
    .D1(_04232_),
    .Y(_04233_));
 sky130_fd_sc_hd__nor2_1 _13300_ (.A(_03579_),
    .B(_04147_),
    .Y(_04234_));
 sky130_fd_sc_hd__a311oi_1 _13301_ (.A1(_03579_),
    .A2(_04076_),
    .A3(_03942_),
    .B1(_04234_),
    .C1(_03610_),
    .Y(_04235_));
 sky130_fd_sc_hd__a21boi_0 _13302_ (.A1(_04004_),
    .A2(_04164_),
    .B1_N(_04077_),
    .Y(_04236_));
 sky130_fd_sc_hd__o21ai_0 _13303_ (.A1(_04235_),
    .A2(_04236_),
    .B1(_03767_),
    .Y(_04237_));
 sky130_fd_sc_hd__a21oi_2 _13304_ (.A1(_04233_),
    .A2(_04237_),
    .B1(_03602_),
    .Y(_04238_));
 sky130_fd_sc_hd__nor3_1 _13305_ (.A(_03579_),
    .B(_04038_),
    .C(_03972_),
    .Y(_04239_));
 sky130_fd_sc_hd__o21ai_0 _13306_ (.A1(_04047_),
    .A2(_04239_),
    .B1(_03767_),
    .Y(_04240_));
 sky130_fd_sc_hd__a221o_1 _13307_ (.A1(_11828_[0]),
    .A2(net4108),
    .B1(_03957_),
    .B2(_11829_[0]),
    .C1(_03767_),
    .X(_04241_));
 sky130_fd_sc_hd__a21oi_2 _13308_ (.A1(_04240_),
    .A2(_04241_),
    .B1(_03611_),
    .Y(_04242_));
 sky130_fd_sc_hd__mux2i_2 _13309_ (.A0(_11840_[0]),
    .A1(net4105),
    .S(_03618_),
    .Y(_04243_));
 sky130_fd_sc_hd__o22ai_2 _13310_ (.A1(_11833_[0]),
    .A2(_04082_),
    .B1(_04243_),
    .B2(_03578_),
    .Y(_04244_));
 sky130_fd_sc_hd__nand2_1 _13311_ (.A(_03766_),
    .B(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__a21oi_1 _13312_ (.A1(_11835_[0]),
    .A2(net4108),
    .B1(_03618_),
    .Y(_04246_));
 sky130_fd_sc_hd__o21ai_0 _13313_ (.A1(_03944_),
    .A2(net4108),
    .B1(_04246_),
    .Y(_04247_));
 sky130_fd_sc_hd__o211ai_1 _13314_ (.A1(_11840_[0]),
    .A2(net4102),
    .B1(_03767_),
    .C1(_04247_),
    .Y(_04248_));
 sky130_fd_sc_hd__a21oi_2 _13315_ (.A1(_04245_),
    .A2(_04248_),
    .B1(_03610_),
    .Y(_04249_));
 sky130_fd_sc_hd__nor3_4 _13316_ (.A(net4066),
    .B(_04242_),
    .C(_04249_),
    .Y(_04250_));
 sky130_fd_sc_hd__o21ai_0 _13317_ (.A1(_11830_[0]),
    .A2(_03579_),
    .B1(net4101),
    .Y(_04251_));
 sky130_fd_sc_hd__o21ai_0 _13318_ (.A1(_03579_),
    .A2(_04028_),
    .B1(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__nand2_1 _13319_ (.A(_04004_),
    .B(_04098_),
    .Y(_04253_));
 sky130_fd_sc_hd__a211oi_1 _13320_ (.A1(_03578_),
    .A2(_04253_),
    .B1(_04099_),
    .C1(net4103),
    .Y(_04254_));
 sky130_fd_sc_hd__a21oi_1 _13321_ (.A1(net4103),
    .A2(_04252_),
    .B1(_04254_),
    .Y(_04255_));
 sky130_fd_sc_hd__nor2_2 _13322_ (.A(_03611_),
    .B(_03618_),
    .Y(_04256_));
 sky130_fd_sc_hd__a221oi_1 _13323_ (.A1(net4106),
    .A2(_03942_),
    .B1(_04256_),
    .B2(net4105),
    .C1(_03579_),
    .Y(_04257_));
 sky130_fd_sc_hd__nor2_1 _13324_ (.A(_03610_),
    .B(_03618_),
    .Y(_04258_));
 sky130_fd_sc_hd__a221oi_1 _13325_ (.A1(_03610_),
    .A2(_04129_),
    .B1(_04258_),
    .B2(_11842_[0]),
    .C1(net4107),
    .Y(_04259_));
 sky130_fd_sc_hd__nand2_1 _13326_ (.A(_03579_),
    .B(_03610_),
    .Y(_04260_));
 sky130_fd_sc_hd__o22ai_1 _13327_ (.A1(_03610_),
    .A2(_03617_),
    .B1(_04260_),
    .B2(net4106),
    .Y(_04261_));
 sky130_fd_sc_hd__nand2_1 _13328_ (.A(_03593_),
    .B(_04261_),
    .Y(_04262_));
 sky130_fd_sc_hd__o211ai_1 _13329_ (.A1(_04257_),
    .A2(_04259_),
    .B1(_03767_),
    .C1(_04262_),
    .Y(_04263_));
 sky130_fd_sc_hd__o211ai_1 _13330_ (.A1(_03767_),
    .A2(_04255_),
    .B1(_04263_),
    .C1(net4066),
    .Y(_04264_));
 sky130_fd_sc_hd__nor2_1 _13331_ (.A(_11844_[0]),
    .B(_03579_),
    .Y(_04265_));
 sky130_fd_sc_hd__a21oi_1 _13332_ (.A1(_11828_[0]),
    .A2(_03579_),
    .B1(_04265_),
    .Y(_04266_));
 sky130_fd_sc_hd__a21oi_1 _13333_ (.A1(_03945_),
    .A2(_04079_),
    .B1(_03579_),
    .Y(_04267_));
 sky130_fd_sc_hd__o32ai_1 _13334_ (.A1(net4103),
    .A2(_03618_),
    .A3(_04266_),
    .B1(_04267_),
    .B2(_03982_),
    .Y(_04268_));
 sky130_fd_sc_hd__nand2_1 _13335_ (.A(_11858_[0]),
    .B(_03579_),
    .Y(_04269_));
 sky130_fd_sc_hd__o2111ai_1 _13336_ (.A1(_11842_[0]),
    .A2(_03952_),
    .B1(_04269_),
    .C1(_03610_),
    .D1(_04118_),
    .Y(_04270_));
 sky130_fd_sc_hd__o211ai_1 _13337_ (.A1(net4108),
    .A2(_04046_),
    .B1(_03984_),
    .C1(_03611_),
    .Y(_04271_));
 sky130_fd_sc_hd__nand3_1 _13338_ (.A(_03767_),
    .B(_04270_),
    .C(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hd__o211ai_1 _13339_ (.A1(_03767_),
    .A2(_04268_),
    .B1(_04272_),
    .C1(_03602_),
    .Y(_04273_));
 sky130_fd_sc_hd__nand3_2 _13340_ (.A(_03759_),
    .B(_04264_),
    .C(_04273_),
    .Y(_04274_));
 sky130_fd_sc_hd__o31ai_4 _13341_ (.A1(_03759_),
    .A2(_04238_),
    .A3(_04250_),
    .B1(_04274_),
    .Y(_00004_));
 sky130_fd_sc_hd__a32oi_2 _13342_ (.A1(net4069),
    .A2(_03977_),
    .A3(_03996_),
    .B1(_03955_),
    .B2(_03944_),
    .Y(_04275_));
 sky130_fd_sc_hd__a21oi_1 _13343_ (.A1(_04019_),
    .A2(_04024_),
    .B1(net4107),
    .Y(_04276_));
 sky130_fd_sc_hd__a211o_1 _13344_ (.A1(_11830_[0]),
    .A2(_04142_),
    .B1(_04276_),
    .C1(_03759_),
    .X(_04277_));
 sky130_fd_sc_hd__o21ai_0 _13345_ (.A1(_03758_),
    .A2(_04275_),
    .B1(_04277_),
    .Y(_04278_));
 sky130_fd_sc_hd__nor2_1 _13346_ (.A(_11835_[0]),
    .B(net4100),
    .Y(_04279_));
 sky130_fd_sc_hd__nor2_1 _13347_ (.A(net4067),
    .B(_04279_),
    .Y(_04280_));
 sky130_fd_sc_hd__a21oi_1 _13348_ (.A1(_03967_),
    .A2(_04161_),
    .B1(net4069),
    .Y(_04281_));
 sky130_fd_sc_hd__a211o_1 _13349_ (.A1(_11829_[0]),
    .A2(_03957_),
    .B1(_04281_),
    .C1(_03759_),
    .X(_04282_));
 sky130_fd_sc_hd__o311ai_0 _13350_ (.A1(_03758_),
    .A2(_04114_),
    .A3(_04280_),
    .B1(_04282_),
    .C1(_03611_),
    .Y(_04283_));
 sky130_fd_sc_hd__o21ai_0 _13351_ (.A1(_03611_),
    .A2(_04278_),
    .B1(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__nand2_2 _13352_ (.A(_04060_),
    .B(_04026_),
    .Y(_04285_));
 sky130_fd_sc_hd__nand3_1 _13353_ (.A(net4067),
    .B(_04024_),
    .C(_04122_),
    .Y(_04286_));
 sky130_fd_sc_hd__o21ai_0 _13354_ (.A1(net4067),
    .A2(_04285_),
    .B1(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hd__nand2_1 _13355_ (.A(_11838_[0]),
    .B(net4067),
    .Y(_04288_));
 sky130_fd_sc_hd__o21ai_0 _13356_ (.A1(net4067),
    .A2(_03980_),
    .B1(_04288_),
    .Y(_04289_));
 sky130_fd_sc_hd__nand2_1 _13357_ (.A(_03610_),
    .B(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__o21ai_0 _13358_ (.A1(_03610_),
    .A2(_04287_),
    .B1(_04290_),
    .Y(_04291_));
 sky130_fd_sc_hd__a31oi_2 _13359_ (.A1(net4108),
    .A2(_04028_),
    .A3(_04061_),
    .B1(_03982_),
    .Y(_04292_));
 sky130_fd_sc_hd__a21oi_1 _13360_ (.A1(_11830_[0]),
    .A2(net4100),
    .B1(_04115_),
    .Y(_04293_));
 sky130_fd_sc_hd__o22ai_1 _13361_ (.A1(_11838_[0]),
    .A2(_04090_),
    .B1(_04293_),
    .B2(net4067),
    .Y(_04294_));
 sky130_fd_sc_hd__o21ai_0 _13362_ (.A1(_03610_),
    .A2(_04294_),
    .B1(_03759_),
    .Y(_04295_));
 sky130_fd_sc_hd__o221ai_1 _13363_ (.A1(_03759_),
    .A2(_04291_),
    .B1(_04292_),
    .B2(_04295_),
    .C1(_03766_),
    .Y(_04296_));
 sky130_fd_sc_hd__o21ai_2 _13364_ (.A1(_03766_),
    .A2(_04284_),
    .B1(_04296_),
    .Y(_04297_));
 sky130_fd_sc_hd__nor2_1 _13365_ (.A(_03593_),
    .B(_03611_),
    .Y(_04298_));
 sky130_fd_sc_hd__a31oi_1 _13366_ (.A1(_03611_),
    .A2(_04122_),
    .A3(_03980_),
    .B1(_04298_),
    .Y(_04299_));
 sky130_fd_sc_hd__o21ai_0 _13367_ (.A1(_03586_),
    .A2(_03610_),
    .B1(net4105),
    .Y(_04300_));
 sky130_fd_sc_hd__o211ai_1 _13368_ (.A1(net4105),
    .A2(_04256_),
    .B1(_04300_),
    .C1(net4107),
    .Y(_04301_));
 sky130_fd_sc_hd__o21ai_0 _13369_ (.A1(_04142_),
    .A2(_04298_),
    .B1(_03586_),
    .Y(_04302_));
 sky130_fd_sc_hd__o2111ai_2 _13370_ (.A1(net4107),
    .A2(_04299_),
    .B1(_04301_),
    .C1(_03758_),
    .D1(_04302_),
    .Y(_04303_));
 sky130_fd_sc_hd__nor3_1 _13371_ (.A(_03579_),
    .B(_04045_),
    .C(_04046_),
    .Y(_04304_));
 sky130_fd_sc_hd__a311oi_1 _13372_ (.A1(net4069),
    .A2(_04118_),
    .A3(_04061_),
    .B1(_04304_),
    .C1(_03610_),
    .Y(_04305_));
 sky130_fd_sc_hd__nand3_1 _13373_ (.A(net4108),
    .B(_03942_),
    .C(_03984_),
    .Y(_04306_));
 sky130_fd_sc_hd__nand2_1 _13374_ (.A(_03579_),
    .B(_04147_),
    .Y(_04307_));
 sky130_fd_sc_hd__a21oi_1 _13375_ (.A1(_04306_),
    .A2(_04307_),
    .B1(_03611_),
    .Y(_04308_));
 sky130_fd_sc_hd__o21ai_2 _13376_ (.A1(_04305_),
    .A2(_04308_),
    .B1(_03759_),
    .Y(_04309_));
 sky130_fd_sc_hd__a21oi_2 _13377_ (.A1(_04303_),
    .A2(_04309_),
    .B1(_03766_),
    .Y(_04310_));
 sky130_fd_sc_hd__nand2_1 _13378_ (.A(_03586_),
    .B(_03593_),
    .Y(_04311_));
 sky130_fd_sc_hd__nor2_1 _13379_ (.A(net4106),
    .B(_03758_),
    .Y(_04312_));
 sky130_fd_sc_hd__nor2_1 _13380_ (.A(_11828_[0]),
    .B(_03759_),
    .Y(_04313_));
 sky130_fd_sc_hd__o32ai_1 _13381_ (.A1(net4100),
    .A2(_04312_),
    .A3(_04313_),
    .B1(_03759_),
    .B2(_03966_),
    .Y(_04314_));
 sky130_fd_sc_hd__a21oi_1 _13382_ (.A1(_03586_),
    .A2(_03759_),
    .B1(_03578_),
    .Y(_04315_));
 sky130_fd_sc_hd__o21ai_0 _13383_ (.A1(_03759_),
    .A2(_04118_),
    .B1(_04315_),
    .Y(_04316_));
 sky130_fd_sc_hd__o21ai_0 _13384_ (.A1(net4068),
    .A2(_04314_),
    .B1(_04316_),
    .Y(_04317_));
 sky130_fd_sc_hd__o21ai_0 _13385_ (.A1(_03758_),
    .A2(_04311_),
    .B1(_04317_),
    .Y(_04318_));
 sky130_fd_sc_hd__nor2_1 _13386_ (.A(net4068),
    .B(_04243_),
    .Y(_04319_));
 sky130_fd_sc_hd__a31o_1 _13387_ (.A1(net4068),
    .A2(_03966_),
    .A3(_04024_),
    .B1(_04319_),
    .X(_04320_));
 sky130_fd_sc_hd__a221oi_1 _13388_ (.A1(_04025_),
    .A2(_03957_),
    .B1(_04065_),
    .B2(_03578_),
    .C1(_03759_),
    .Y(_04321_));
 sky130_fd_sc_hd__a211oi_1 _13389_ (.A1(_03759_),
    .A2(_04320_),
    .B1(_04321_),
    .C1(_03610_),
    .Y(_04322_));
 sky130_fd_sc_hd__a21oi_1 _13390_ (.A1(_03610_),
    .A2(_04318_),
    .B1(_04322_),
    .Y(_04323_));
 sky130_fd_sc_hd__o21ai_2 _13391_ (.A1(_03767_),
    .A2(_04323_),
    .B1(_03602_),
    .Y(_04324_));
 sky130_fd_sc_hd__o22ai_4 _13392_ (.A1(_03602_),
    .A2(_04297_),
    .B1(_04310_),
    .B2(_04324_),
    .Y(_00005_));
 sky130_fd_sc_hd__a21oi_1 _13393_ (.A1(_11847_[0]),
    .A2(net4069),
    .B1(_04029_),
    .Y(_04325_));
 sky130_fd_sc_hd__a21oi_1 _13394_ (.A1(_03977_),
    .A2(_03996_),
    .B1(net4108),
    .Y(_04326_));
 sky130_fd_sc_hd__a211o_1 _13395_ (.A1(_11829_[0]),
    .A2(_03955_),
    .B1(_04326_),
    .C1(_03611_),
    .X(_04327_));
 sky130_fd_sc_hd__o21ai_0 _13396_ (.A1(net4103),
    .A2(_04325_),
    .B1(_04327_),
    .Y(_04328_));
 sky130_fd_sc_hd__o221ai_1 _13397_ (.A1(_11830_[0]),
    .A2(_04082_),
    .B1(_04311_),
    .B2(_03578_),
    .C1(_04031_),
    .Y(_04329_));
 sky130_fd_sc_hd__nor2_1 _13398_ (.A(net4103),
    .B(_04329_),
    .Y(_04330_));
 sky130_fd_sc_hd__a21oi_1 _13399_ (.A1(_04118_),
    .A2(_04032_),
    .B1(net4107),
    .Y(_04331_));
 sky130_fd_sc_hd__nor4_2 _13400_ (.A(_03611_),
    .B(_04129_),
    .C(_04137_),
    .D(_04331_),
    .Y(_04332_));
 sky130_fd_sc_hd__nor3_1 _13401_ (.A(net4066),
    .B(_04330_),
    .C(_04332_),
    .Y(_04333_));
 sky130_fd_sc_hd__a21oi_1 _13402_ (.A1(net4066),
    .A2(_04328_),
    .B1(_04333_),
    .Y(_04334_));
 sky130_fd_sc_hd__a21oi_1 _13403_ (.A1(_03996_),
    .A2(_04161_),
    .B1(net4108),
    .Y(_04335_));
 sky130_fd_sc_hd__o221ai_1 _13404_ (.A1(net4105),
    .A2(_03957_),
    .B1(_04071_),
    .B2(net4108),
    .C1(net4103),
    .Y(_04336_));
 sky130_fd_sc_hd__o311ai_0 _13405_ (.A1(net4103),
    .A2(_04175_),
    .A3(_04335_),
    .B1(_04336_),
    .C1(_03602_),
    .Y(_04337_));
 sky130_fd_sc_hd__a21oi_1 _13406_ (.A1(_04028_),
    .A2(_03945_),
    .B1(_03579_),
    .Y(_04338_));
 sky130_fd_sc_hd__o211ai_1 _13407_ (.A1(_11844_[0]),
    .A2(net4101),
    .B1(_04087_),
    .C1(_03579_),
    .Y(_04339_));
 sky130_fd_sc_hd__o311ai_0 _13408_ (.A1(_03579_),
    .A2(_04046_),
    .A3(_03972_),
    .B1(_04339_),
    .C1(net4103),
    .Y(_04340_));
 sky130_fd_sc_hd__o311ai_0 _13409_ (.A1(net4103),
    .A2(_04338_),
    .A3(_04326_),
    .B1(_04340_),
    .C1(net4066),
    .Y(_04341_));
 sky130_fd_sc_hd__a21oi_1 _13410_ (.A1(_04337_),
    .A2(_04341_),
    .B1(net3627),
    .Y(_04342_));
 sky130_fd_sc_hd__a21oi_1 _13411_ (.A1(net3627),
    .A2(_04334_),
    .B1(_04342_),
    .Y(_04343_));
 sky130_fd_sc_hd__nor2_1 _13412_ (.A(_11848_[0]),
    .B(_03578_),
    .Y(_04344_));
 sky130_fd_sc_hd__a31oi_1 _13413_ (.A1(_03578_),
    .A2(net4106),
    .A3(net4100),
    .B1(_03610_),
    .Y(_04345_));
 sky130_fd_sc_hd__o21ai_0 _13414_ (.A1(_03578_),
    .A2(_04285_),
    .B1(_04345_),
    .Y(_04346_));
 sky130_fd_sc_hd__o311ai_1 _13415_ (.A1(_03611_),
    .A2(_04319_),
    .A3(_04344_),
    .B1(_04346_),
    .C1(_03602_),
    .Y(_04347_));
 sky130_fd_sc_hd__a221oi_1 _13416_ (.A1(_11838_[0]),
    .A2(_04142_),
    .B1(_04243_),
    .B2(net4067),
    .C1(_03610_),
    .Y(_04348_));
 sky130_fd_sc_hd__o21ai_1 _13417_ (.A1(_04150_),
    .A2(_04348_),
    .B1(net4066),
    .Y(_04349_));
 sky130_fd_sc_hd__nand3_1 _13418_ (.A(_03578_),
    .B(_04118_),
    .C(_04130_),
    .Y(_04350_));
 sky130_fd_sc_hd__o211ai_1 _13419_ (.A1(_03578_),
    .A2(_04006_),
    .B1(_04350_),
    .C1(net4103),
    .Y(_04351_));
 sky130_fd_sc_hd__a311o_1 _13420_ (.A1(net4069),
    .A2(_04076_),
    .A3(_04098_),
    .B1(_03953_),
    .C1(net4103),
    .X(_04352_));
 sky130_fd_sc_hd__nand3_1 _13421_ (.A(net4069),
    .B(_03966_),
    .C(_03967_),
    .Y(_04353_));
 sky130_fd_sc_hd__o211ai_1 _13422_ (.A1(_11844_[0]),
    .A2(_03618_),
    .B1(_04060_),
    .C1(net4108),
    .Y(_04354_));
 sky130_fd_sc_hd__nor2_1 _13423_ (.A(_11852_[0]),
    .B(_03578_),
    .Y(_04355_));
 sky130_fd_sc_hd__a311oi_1 _13424_ (.A1(_03578_),
    .A2(_03966_),
    .A3(_04024_),
    .B1(_04355_),
    .C1(net4103),
    .Y(_04356_));
 sky130_fd_sc_hd__a311oi_1 _13425_ (.A1(net4103),
    .A2(_04353_),
    .A3(_04354_),
    .B1(_04356_),
    .C1(net4066),
    .Y(_04357_));
 sky130_fd_sc_hd__a311oi_1 _13426_ (.A1(net4066),
    .A2(_04351_),
    .A3(_04352_),
    .B1(_04357_),
    .C1(net3627),
    .Y(_04358_));
 sky130_fd_sc_hd__a31oi_1 _13427_ (.A1(net3627),
    .A2(_04347_),
    .A3(_04349_),
    .B1(_04358_),
    .Y(_04359_));
 sky130_fd_sc_hd__nor2_1 _13428_ (.A(_03759_),
    .B(_04359_),
    .Y(_04360_));
 sky130_fd_sc_hd__a21oi_1 _13429_ (.A1(_03759_),
    .A2(_04343_),
    .B1(_04360_),
    .Y(_00006_));
 sky130_fd_sc_hd__nand2_1 _13430_ (.A(_03602_),
    .B(_04243_),
    .Y(_04361_));
 sky130_fd_sc_hd__o311ai_1 _13431_ (.A1(_11849_[0]),
    .A2(_03602_),
    .A3(_04041_),
    .B1(_04361_),
    .C1(_03579_),
    .Y(_04362_));
 sky130_fd_sc_hd__a21oi_1 _13432_ (.A1(net4066),
    .A2(_04046_),
    .B1(_03972_),
    .Y(_04363_));
 sky130_fd_sc_hd__nand2_1 _13433_ (.A(net4108),
    .B(_04363_),
    .Y(_04364_));
 sky130_fd_sc_hd__a21oi_1 _13434_ (.A1(_04362_),
    .A2(_04364_),
    .B1(_03611_),
    .Y(_04365_));
 sky130_fd_sc_hd__nand2_1 _13435_ (.A(net4108),
    .B(_03969_),
    .Y(_04366_));
 sky130_fd_sc_hd__o221ai_1 _13436_ (.A1(_11830_[0]),
    .A2(_04052_),
    .B1(_03958_),
    .B2(_11829_[0]),
    .C1(_04366_),
    .Y(_04367_));
 sky130_fd_sc_hd__nand3_1 _13437_ (.A(_03579_),
    .B(_04004_),
    .C(_04087_),
    .Y(_04368_));
 sky130_fd_sc_hd__o311a_1 _13438_ (.A1(_03579_),
    .A2(_03969_),
    .A3(_04045_),
    .B1(_04368_),
    .C1(_03602_),
    .X(_04369_));
 sky130_fd_sc_hd__a211oi_1 _13439_ (.A1(net4066),
    .A2(_04367_),
    .B1(_04369_),
    .C1(_03610_),
    .Y(_04370_));
 sky130_fd_sc_hd__o21ai_2 _13440_ (.A1(_04365_),
    .A2(_04370_),
    .B1(net3627),
    .Y(_04371_));
 sky130_fd_sc_hd__a221oi_1 _13441_ (.A1(_11835_[0]),
    .A2(net4108),
    .B1(_04032_),
    .B2(_04164_),
    .C1(net4103),
    .Y(_04372_));
 sky130_fd_sc_hd__nor2_1 _13442_ (.A(net4108),
    .B(_03593_),
    .Y(_04373_));
 sky130_fd_sc_hd__o21ai_0 _13443_ (.A1(_04265_),
    .A2(_04373_),
    .B1(net4101),
    .Y(_04374_));
 sky130_fd_sc_hd__a21oi_1 _13444_ (.A1(_04004_),
    .A2(_04374_),
    .B1(_03611_),
    .Y(_04375_));
 sky130_fd_sc_hd__o21ai_0 _13445_ (.A1(_04372_),
    .A2(_04375_),
    .B1(net4066),
    .Y(_04376_));
 sky130_fd_sc_hd__nor3_1 _13446_ (.A(_03579_),
    .B(_04017_),
    .C(_04039_),
    .Y(_04377_));
 sky130_fd_sc_hd__a21oi_1 _13447_ (.A1(_04004_),
    .A2(_04087_),
    .B1(net4069),
    .Y(_04378_));
 sky130_fd_sc_hd__a21oi_1 _13448_ (.A1(net4069),
    .A2(_04219_),
    .B1(_04378_),
    .Y(_04379_));
 sky130_fd_sc_hd__nand2_1 _13449_ (.A(net4103),
    .B(_04379_),
    .Y(_04380_));
 sky130_fd_sc_hd__o311ai_0 _13450_ (.A1(net4103),
    .A2(_04205_),
    .A3(_04377_),
    .B1(_04380_),
    .C1(_03602_),
    .Y(_04381_));
 sky130_fd_sc_hd__a31oi_1 _13451_ (.A1(_03767_),
    .A2(_04376_),
    .A3(_04381_),
    .B1(_03758_),
    .Y(_04382_));
 sky130_fd_sc_hd__nor3_1 _13452_ (.A(net4106),
    .B(_03610_),
    .C(_03617_),
    .Y(_04383_));
 sky130_fd_sc_hd__o21ai_0 _13453_ (.A1(_04091_),
    .A2(_04383_),
    .B1(_03579_),
    .Y(_04384_));
 sky130_fd_sc_hd__o211ai_1 _13454_ (.A1(_04017_),
    .A2(_04129_),
    .B1(net4107),
    .C1(_03610_),
    .Y(_04385_));
 sky130_fd_sc_hd__nand2_1 _13455_ (.A(net4107),
    .B(_03611_),
    .Y(_04386_));
 sky130_fd_sc_hd__o21ai_0 _13456_ (.A1(net4105),
    .A2(_04260_),
    .B1(_04386_),
    .Y(_04387_));
 sky130_fd_sc_hd__a21oi_1 _13457_ (.A1(net4106),
    .A2(_04387_),
    .B1(net4066),
    .Y(_04388_));
 sky130_fd_sc_hd__nand2_1 _13458_ (.A(_03952_),
    .B(_04260_),
    .Y(_04389_));
 sky130_fd_sc_hd__nand2_1 _13459_ (.A(_11829_[0]),
    .B(net4107),
    .Y(_04390_));
 sky130_fd_sc_hd__nand3_1 _13460_ (.A(_11833_[0]),
    .B(_03579_),
    .C(_03611_),
    .Y(_04391_));
 sky130_fd_sc_hd__a21oi_1 _13461_ (.A1(_04390_),
    .A2(_04391_),
    .B1(_03617_),
    .Y(_04392_));
 sky130_fd_sc_hd__a211o_1 _13462_ (.A1(_11828_[0]),
    .A2(_04389_),
    .B1(_04392_),
    .C1(_04256_),
    .X(_04393_));
 sky130_fd_sc_hd__a32oi_1 _13463_ (.A1(_04384_),
    .A2(_04385_),
    .A3(_04388_),
    .B1(_04393_),
    .B2(net4066),
    .Y(_04394_));
 sky130_fd_sc_hd__nand2_1 _13464_ (.A(_11828_[0]),
    .B(_03579_),
    .Y(_04395_));
 sky130_fd_sc_hd__nand2_1 _13465_ (.A(net4107),
    .B(_04161_),
    .Y(_04396_));
 sky130_fd_sc_hd__a21oi_1 _13466_ (.A1(_04076_),
    .A2(_04098_),
    .B1(_03579_),
    .Y(_04397_));
 sky130_fd_sc_hd__nor3_1 _13467_ (.A(_03610_),
    .B(_04099_),
    .C(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__a31oi_1 _13468_ (.A1(_03610_),
    .A2(_04395_),
    .A3(_04396_),
    .B1(_04398_),
    .Y(_04399_));
 sky130_fd_sc_hd__nor2_1 _13469_ (.A(_11858_[0]),
    .B(net4107),
    .Y(_04400_));
 sky130_fd_sc_hd__a311oi_1 _13470_ (.A1(net4107),
    .A2(_03945_),
    .A3(_03996_),
    .B1(_04400_),
    .C1(_03611_),
    .Y(_04401_));
 sky130_fd_sc_hd__a21oi_1 _13471_ (.A1(net4106),
    .A2(net4101),
    .B1(_11854_[0]),
    .Y(_04402_));
 sky130_fd_sc_hd__nor2_1 _13472_ (.A(_03579_),
    .B(_04402_),
    .Y(_04403_));
 sky130_fd_sc_hd__o21a_1 _13473_ (.A1(_04155_),
    .A2(_04403_),
    .B1(_03611_),
    .X(_04404_));
 sky130_fd_sc_hd__o21ai_0 _13474_ (.A1(_04401_),
    .A2(_04404_),
    .B1(net4066),
    .Y(_04405_));
 sky130_fd_sc_hd__o211ai_1 _13475_ (.A1(net4066),
    .A2(_04399_),
    .B1(_04405_),
    .C1(_03767_),
    .Y(_04406_));
 sky130_fd_sc_hd__o21ai_0 _13476_ (.A1(_03767_),
    .A2(_04394_),
    .B1(_04406_),
    .Y(_04407_));
 sky130_fd_sc_hd__a22oi_1 _13477_ (.A1(_04371_),
    .A2(_04382_),
    .B1(_04407_),
    .B2(_03758_),
    .Y(_00007_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1223 ();
 sky130_fd_sc_hd__nor2_4 _13483_ (.A(_03696_),
    .B(_03715_),
    .Y(_04411_));
 sky130_fd_sc_hd__nand2_8 _13484_ (.A(_03696_),
    .B(_03715_),
    .Y(_04412_));
 sky130_fd_sc_hd__nand2b_2 _13485_ (.A_N(_04411_),
    .B(_04412_),
    .Y(_04413_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1222 ();
 sky130_fd_sc_hd__xnor2_1 _13487_ (.A(_03704_),
    .B(net4084),
    .Y(_04415_));
 sky130_fd_sc_hd__nand2_1 _13488_ (.A(net4090),
    .B(_04415_),
    .Y(_04416_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1220 ();
 sky130_fd_sc_hd__o211ai_1 _13491_ (.A1(net4090),
    .A2(_04413_),
    .B1(_04416_),
    .C1(_03735_),
    .Y(_04419_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1217 ();
 sky130_fd_sc_hd__nor2_4 _13495_ (.A(net4088),
    .B(_03715_),
    .Y(_04423_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1214 ();
 sky130_fd_sc_hd__nor2_2 _13499_ (.A(_11863_[0]),
    .B(net4084),
    .Y(_04427_));
 sky130_fd_sc_hd__a21oi_1 _13500_ (.A1(net4061),
    .A2(_04427_),
    .B1(_04411_),
    .Y(_04428_));
 sky130_fd_sc_hd__nor2_1 _13501_ (.A(_03704_),
    .B(_04428_),
    .Y(_04429_));
 sky130_fd_sc_hd__a31oi_1 _13502_ (.A1(_11863_[0]),
    .A2(net4061),
    .A3(_04423_),
    .B1(_04429_),
    .Y(_04430_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1213 ();
 sky130_fd_sc_hd__nor2_4 _13504_ (.A(_03704_),
    .B(_03715_),
    .Y(_04432_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1212 ();
 sky130_fd_sc_hd__nand2_8 _13506_ (.A(_03704_),
    .B(_03715_),
    .Y(_04434_));
 sky130_fd_sc_hd__nor2_4 _13507_ (.A(_11863_[0]),
    .B(_04434_),
    .Y(_04435_));
 sky130_fd_sc_hd__a221oi_1 _13508_ (.A1(_11876_[0]),
    .A2(_04415_),
    .B1(_04432_),
    .B2(_11872_[0]),
    .C1(_04435_),
    .Y(_04436_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1211 ();
 sky130_fd_sc_hd__nor2_1 _13510_ (.A(_11876_[0]),
    .B(net4084),
    .Y(_04438_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1210 ();
 sky130_fd_sc_hd__nor2_4 _13512_ (.A(_11862_[0]),
    .B(_03715_),
    .Y(_04440_));
 sky130_fd_sc_hd__nor3_1 _13513_ (.A(_03704_),
    .B(_04438_),
    .C(_04440_),
    .Y(_04441_));
 sky130_fd_sc_hd__nor2_4 _13514_ (.A(_11872_[0]),
    .B(net4084),
    .Y(_04442_));
 sky130_fd_sc_hd__nand2_4 _13515_ (.A(_11863_[0]),
    .B(net4084),
    .Y(_04443_));
 sky130_fd_sc_hd__nor3b_1 _13516_ (.A(net4086),
    .B(_04442_),
    .C_N(_04443_),
    .Y(_04444_));
 sky130_fd_sc_hd__nor3_1 _13517_ (.A(net4061),
    .B(_04441_),
    .C(_04444_),
    .Y(_04445_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1209 ();
 sky130_fd_sc_hd__a211oi_1 _13519_ (.A1(net4061),
    .A2(_04436_),
    .B1(_04445_),
    .C1(_03725_),
    .Y(_04447_));
 sky130_fd_sc_hd__a31oi_1 _13520_ (.A1(_03725_),
    .A2(_04419_),
    .A3(_04430_),
    .B1(_04447_),
    .Y(_04448_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1208 ();
 sky130_fd_sc_hd__nand2_8 _13522_ (.A(net4086),
    .B(net4084),
    .Y(_04450_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1207 ();
 sky130_fd_sc_hd__nor2_2 _13524_ (.A(_11867_[0]),
    .B(_03715_),
    .Y(_04452_));
 sky130_fd_sc_hd__a21oi_1 _13525_ (.A1(_11878_[0]),
    .A2(_03715_),
    .B1(_04452_),
    .Y(_04453_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1206 ();
 sky130_fd_sc_hd__o221ai_1 _13527_ (.A1(_11872_[0]),
    .A2(_04450_),
    .B1(_04453_),
    .B2(net4086),
    .C1(_03735_),
    .Y(_04455_));
 sky130_fd_sc_hd__a221o_1 _13528_ (.A1(_11888_[0]),
    .A2(_03715_),
    .B1(_04432_),
    .B2(_11863_[0]),
    .C1(_03735_),
    .X(_04456_));
 sky130_fd_sc_hd__nand3_1 _13529_ (.A(_03725_),
    .B(_04455_),
    .C(_04456_),
    .Y(_04457_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1201 ();
 sky130_fd_sc_hd__nand2_1 _13535_ (.A(_11867_[0]),
    .B(_03715_),
    .Y(_04463_));
 sky130_fd_sc_hd__o21ai_2 _13536_ (.A1(_11878_[0]),
    .A2(_03715_),
    .B1(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1200 ();
 sky130_fd_sc_hd__nor2_4 _13538_ (.A(_03704_),
    .B(net4084),
    .Y(_04466_));
 sky130_fd_sc_hd__nand2_1 _13539_ (.A(_11874_[0]),
    .B(_04466_),
    .Y(_04467_));
 sky130_fd_sc_hd__o21ai_0 _13540_ (.A1(net4086),
    .A2(_04464_),
    .B1(_04467_),
    .Y(_04468_));
 sky130_fd_sc_hd__nand2_4 _13541_ (.A(net4090),
    .B(net4084),
    .Y(_04469_));
 sky130_fd_sc_hd__nand2_4 _13542_ (.A(net4063),
    .B(_03715_),
    .Y(_04470_));
 sky130_fd_sc_hd__a21oi_1 _13543_ (.A1(_04469_),
    .A2(_04470_),
    .B1(_03704_),
    .Y(_04471_));
 sky130_fd_sc_hd__nor3_2 _13544_ (.A(net4086),
    .B(_04438_),
    .C(_04452_),
    .Y(_04472_));
 sky130_fd_sc_hd__o21ai_0 _13545_ (.A1(_04471_),
    .A2(_04472_),
    .B1(net4061),
    .Y(_04473_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1198 ();
 sky130_fd_sc_hd__o211ai_1 _13548_ (.A1(net4061),
    .A2(_04468_),
    .B1(_04473_),
    .C1(net4062),
    .Y(_04476_));
 sky130_fd_sc_hd__nand3_1 _13549_ (.A(_03751_),
    .B(_04457_),
    .C(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hd__o21ai_2 _13550_ (.A1(_03751_),
    .A2(_04448_),
    .B1(_04477_),
    .Y(_04478_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1197 ();
 sky130_fd_sc_hd__a211oi_1 _13552_ (.A1(_11864_[0]),
    .A2(_03715_),
    .B1(_04411_),
    .C1(net4086),
    .Y(_04480_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1196 ();
 sky130_fd_sc_hd__nor2_4 _13554_ (.A(net4063),
    .B(net4084),
    .Y(_04482_));
 sky130_fd_sc_hd__nor3_1 _13555_ (.A(_03704_),
    .B(_04482_),
    .C(_04452_),
    .Y(_04483_));
 sky130_fd_sc_hd__nand2_2 _13556_ (.A(_11863_[0]),
    .B(_03715_),
    .Y(_04484_));
 sky130_fd_sc_hd__nand2_2 _13557_ (.A(_11867_[0]),
    .B(net4084),
    .Y(_04485_));
 sky130_fd_sc_hd__nand2b_4 _13558_ (.A_N(_11864_[0]),
    .B(_03715_),
    .Y(_04486_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1195 ();
 sky130_fd_sc_hd__a21oi_1 _13560_ (.A1(_04485_),
    .A2(_04486_),
    .B1(_03704_),
    .Y(_04488_));
 sky130_fd_sc_hd__a311o_1 _13561_ (.A1(_03704_),
    .A2(_04469_),
    .A3(_04484_),
    .B1(_04488_),
    .C1(_03734_),
    .X(_04489_));
 sky130_fd_sc_hd__o311ai_1 _13562_ (.A1(_03735_),
    .A2(_04480_),
    .A3(_04483_),
    .B1(_04489_),
    .C1(_03725_),
    .Y(_04490_));
 sky130_fd_sc_hd__nand2_4 _13563_ (.A(_03696_),
    .B(net4086),
    .Y(_04491_));
 sky130_fd_sc_hd__nand2_1 _13564_ (.A(_11878_[0]),
    .B(_03704_),
    .Y(_04492_));
 sky130_fd_sc_hd__a21oi_1 _13565_ (.A1(_04491_),
    .A2(_04492_),
    .B1(_03715_),
    .Y(_04493_));
 sky130_fd_sc_hd__nor2_1 _13566_ (.A(_03725_),
    .B(_04493_),
    .Y(_04494_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1194 ();
 sky130_fd_sc_hd__nand2_2 _13568_ (.A(_11862_[0]),
    .B(_03704_),
    .Y(_04496_));
 sky130_fd_sc_hd__o211ai_1 _13569_ (.A1(net4090),
    .A2(_03704_),
    .B1(_03715_),
    .C1(_04496_),
    .Y(_04497_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1193 ();
 sky130_fd_sc_hd__inv_2 _13571_ (.A(_11867_[0]),
    .Y(_04499_));
 sky130_fd_sc_hd__nor2_4 _13572_ (.A(_04499_),
    .B(net4084),
    .Y(_04500_));
 sky130_fd_sc_hd__nor2_4 _13573_ (.A(net4090),
    .B(_03715_),
    .Y(_04501_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1192 ();
 sky130_fd_sc_hd__o21ai_0 _13575_ (.A1(_04500_),
    .A2(_04501_),
    .B1(net4086),
    .Y(_04503_));
 sky130_fd_sc_hd__o21ai_2 _13576_ (.A1(_11869_[0]),
    .A2(_04434_),
    .B1(_04503_),
    .Y(_04504_));
 sky130_fd_sc_hd__nor2_4 _13577_ (.A(_03725_),
    .B(_03734_),
    .Y(_04505_));
 sky130_fd_sc_hd__a32oi_1 _13578_ (.A1(_03734_),
    .A2(_04494_),
    .A3(_04497_),
    .B1(_04504_),
    .B2(_04505_),
    .Y(_04506_));
 sky130_fd_sc_hd__nand3_1 _13579_ (.A(_03750_),
    .B(_04490_),
    .C(_04506_),
    .Y(_04507_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1190 ();
 sky130_fd_sc_hd__nor2_4 _13582_ (.A(net4089),
    .B(_03715_),
    .Y(_04510_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1189 ();
 sky130_fd_sc_hd__o21ai_1 _13584_ (.A1(_04482_),
    .A2(_04510_),
    .B1(_03704_),
    .Y(_04512_));
 sky130_fd_sc_hd__nor2_4 _13585_ (.A(_11863_[0]),
    .B(_03715_),
    .Y(_04513_));
 sky130_fd_sc_hd__o21ai_0 _13586_ (.A1(_04442_),
    .A2(_04513_),
    .B1(_03702_),
    .Y(_04514_));
 sky130_fd_sc_hd__nand2_1 _13587_ (.A(_11876_[0]),
    .B(_04432_),
    .Y(_04515_));
 sky130_fd_sc_hd__nor2_1 _13588_ (.A(_11878_[0]),
    .B(_03715_),
    .Y(_04516_));
 sky130_fd_sc_hd__nor2_4 _13589_ (.A(_11869_[0]),
    .B(net4084),
    .Y(_04517_));
 sky130_fd_sc_hd__o21ai_0 _13590_ (.A1(_04516_),
    .A2(_04517_),
    .B1(_03704_),
    .Y(_04518_));
 sky130_fd_sc_hd__a21oi_1 _13591_ (.A1(_04515_),
    .A2(_04518_),
    .B1(net4062),
    .Y(_04519_));
 sky130_fd_sc_hd__a31oi_1 _13592_ (.A1(net4062),
    .A2(_04512_),
    .A3(_04514_),
    .B1(_04519_),
    .Y(_04520_));
 sky130_fd_sc_hd__a21oi_1 _13593_ (.A1(_11874_[0]),
    .A2(_03704_),
    .B1(_03715_),
    .Y(_04521_));
 sky130_fd_sc_hd__or3_1 _13594_ (.A(net4062),
    .B(_04435_),
    .C(_04521_),
    .X(_04522_));
 sky130_fd_sc_hd__nand2_4 _13595_ (.A(_11869_[0]),
    .B(_04432_),
    .Y(_04523_));
 sky130_fd_sc_hd__o2111ai_1 _13596_ (.A1(_03725_),
    .A2(_04497_),
    .B1(_04522_),
    .C1(_04523_),
    .D1(_03734_),
    .Y(_04524_));
 sky130_fd_sc_hd__o211ai_1 _13597_ (.A1(_03734_),
    .A2(_04520_),
    .B1(_04524_),
    .C1(_03751_),
    .Y(_04525_));
 sky130_fd_sc_hd__nand3_1 _13598_ (.A(_03744_),
    .B(_04507_),
    .C(_04525_),
    .Y(_04526_));
 sky130_fd_sc_hd__a21boi_2 _13599_ (.A1(net3711),
    .A2(_04478_),
    .B1_N(_04526_),
    .Y(_00008_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1187 ();
 sky130_fd_sc_hd__nand2_1 _13602_ (.A(_11872_[0]),
    .B(_03702_),
    .Y(_04529_));
 sky130_fd_sc_hd__nor3_1 _13603_ (.A(_11890_[0]),
    .B(net4084),
    .C(_03735_),
    .Y(_04530_));
 sky130_fd_sc_hd__a31oi_1 _13604_ (.A1(net4084),
    .A2(_04496_),
    .A3(_04529_),
    .B1(_04530_),
    .Y(_04531_));
 sky130_fd_sc_hd__nor2_1 _13605_ (.A(_03725_),
    .B(_04531_),
    .Y(_04532_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1186 ();
 sky130_fd_sc_hd__nor2_1 _13607_ (.A(_11867_[0]),
    .B(net4084),
    .Y(_04534_));
 sky130_fd_sc_hd__inv_4 _13608_ (.A(_11876_[0]),
    .Y(_04535_));
 sky130_fd_sc_hd__nand2_8 _13609_ (.A(_04535_),
    .B(net4084),
    .Y(_04536_));
 sky130_fd_sc_hd__nand3b_1 _13610_ (.A_N(_04534_),
    .B(_04536_),
    .C(_03702_),
    .Y(_04537_));
 sky130_fd_sc_hd__nand2_4 _13611_ (.A(net4063),
    .B(net4084),
    .Y(_04538_));
 sky130_fd_sc_hd__nand2_4 _13612_ (.A(_11862_[0]),
    .B(_03715_),
    .Y(_04539_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1185 ();
 sky130_fd_sc_hd__a21o_1 _13614_ (.A1(_04538_),
    .A2(_04539_),
    .B1(net4086),
    .X(_04541_));
 sky130_fd_sc_hd__a21oi_1 _13615_ (.A1(_04537_),
    .A2(_04541_),
    .B1(_03734_),
    .Y(_04542_));
 sky130_fd_sc_hd__nor2_4 _13616_ (.A(net4063),
    .B(_03715_),
    .Y(_04543_));
 sky130_fd_sc_hd__nor3_1 _13617_ (.A(_03702_),
    .B(_04543_),
    .C(_04517_),
    .Y(_04544_));
 sky130_fd_sc_hd__nor2_2 _13618_ (.A(_03704_),
    .B(_04413_),
    .Y(_04545_));
 sky130_fd_sc_hd__nor3_1 _13619_ (.A(_03735_),
    .B(_04544_),
    .C(_04545_),
    .Y(_04546_));
 sky130_fd_sc_hd__nor3_1 _13620_ (.A(net4062),
    .B(_04542_),
    .C(_04546_),
    .Y(_04547_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1184 ();
 sky130_fd_sc_hd__o21ai_0 _13622_ (.A1(_04532_),
    .A2(_04547_),
    .B1(_03750_),
    .Y(_04549_));
 sky130_fd_sc_hd__o21ai_0 _13623_ (.A1(_04411_),
    .A2(_04534_),
    .B1(_03702_),
    .Y(_04550_));
 sky130_fd_sc_hd__nand2_1 _13624_ (.A(net4090),
    .B(_04510_),
    .Y(_04551_));
 sky130_fd_sc_hd__nand2_4 _13625_ (.A(_11869_[0]),
    .B(net4084),
    .Y(_04552_));
 sky130_fd_sc_hd__a21oi_1 _13626_ (.A1(_04484_),
    .A2(_04552_),
    .B1(_03704_),
    .Y(_04553_));
 sky130_fd_sc_hd__a311oi_2 _13627_ (.A1(_03704_),
    .A2(_04485_),
    .A3(_04486_),
    .B1(_04553_),
    .C1(_03735_),
    .Y(_04554_));
 sky130_fd_sc_hd__a31oi_1 _13628_ (.A1(_03735_),
    .A2(_04550_),
    .A3(_04551_),
    .B1(_04554_),
    .Y(_04555_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1183 ();
 sky130_fd_sc_hd__nand2_1 _13630_ (.A(_11881_[0]),
    .B(_03715_),
    .Y(_04557_));
 sky130_fd_sc_hd__nand2_1 _13631_ (.A(_11869_[0]),
    .B(net4087),
    .Y(_04558_));
 sky130_fd_sc_hd__nand2_1 _13632_ (.A(_03696_),
    .B(_03704_),
    .Y(_04559_));
 sky130_fd_sc_hd__nand3_1 _13633_ (.A(net4085),
    .B(_04558_),
    .C(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__a311oi_1 _13634_ (.A1(_03704_),
    .A2(_04484_),
    .A3(_04552_),
    .B1(_04471_),
    .C1(net4061),
    .Y(_04561_));
 sky130_fd_sc_hd__a311o_1 _13635_ (.A1(_03734_),
    .A2(_04557_),
    .A3(_04560_),
    .B1(_04561_),
    .C1(net4062),
    .X(_04562_));
 sky130_fd_sc_hd__o211ai_1 _13636_ (.A1(_03725_),
    .A2(_04555_),
    .B1(_04562_),
    .C1(_03751_),
    .Y(_04563_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1182 ();
 sky130_fd_sc_hd__nand2_4 _13638_ (.A(net4087),
    .B(_03715_),
    .Y(_04565_));
 sky130_fd_sc_hd__a21oi_1 _13639_ (.A1(_11869_[0]),
    .A2(net4084),
    .B1(_04427_),
    .Y(_04566_));
 sky130_fd_sc_hd__o22ai_1 _13640_ (.A1(_11862_[0]),
    .A2(_04565_),
    .B1(_04566_),
    .B2(net4086),
    .Y(_04567_));
 sky130_fd_sc_hd__xnor2_1 _13641_ (.A(_03702_),
    .B(net4084),
    .Y(_04568_));
 sky130_fd_sc_hd__nor2_2 _13642_ (.A(net4090),
    .B(_04568_),
    .Y(_04569_));
 sky130_fd_sc_hd__nor2_1 _13643_ (.A(net4063),
    .B(_04412_),
    .Y(_04570_));
 sky130_fd_sc_hd__a2111oi_0 _13644_ (.A1(_11863_[0]),
    .A2(_04432_),
    .B1(_04569_),
    .C1(_04570_),
    .D1(_03735_),
    .Y(_04571_));
 sky130_fd_sc_hd__a21oi_1 _13645_ (.A1(_03735_),
    .A2(_04567_),
    .B1(_04571_),
    .Y(_04572_));
 sky130_fd_sc_hd__nor3_1 _13646_ (.A(_03704_),
    .B(_04501_),
    .C(_04517_),
    .Y(_04573_));
 sky130_fd_sc_hd__nand2b_4 _13647_ (.A_N(_11863_[0]),
    .B(_03715_),
    .Y(_04574_));
 sky130_fd_sc_hd__a21oi_1 _13648_ (.A1(_04574_),
    .A2(_04536_),
    .B1(_03702_),
    .Y(_04575_));
 sky130_fd_sc_hd__nand2_1 _13649_ (.A(_11864_[0]),
    .B(_04466_),
    .Y(_04576_));
 sky130_fd_sc_hd__nor2_2 _13650_ (.A(_03696_),
    .B(net4084),
    .Y(_04577_));
 sky130_fd_sc_hd__o21ai_0 _13651_ (.A1(_04440_),
    .A2(_04577_),
    .B1(_03704_),
    .Y(_04578_));
 sky130_fd_sc_hd__nand3_1 _13652_ (.A(_03735_),
    .B(_04576_),
    .C(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hd__o311ai_0 _13653_ (.A1(_03735_),
    .A2(_04573_),
    .A3(_04575_),
    .B1(_04579_),
    .C1(_03725_),
    .Y(_04580_));
 sky130_fd_sc_hd__o21ai_1 _13654_ (.A1(_03725_),
    .A2(_04572_),
    .B1(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__nand3_1 _13655_ (.A(_11863_[0]),
    .B(net4086),
    .C(_03715_),
    .Y(_04582_));
 sky130_fd_sc_hd__and2_4 _13656_ (.A(_03725_),
    .B(_04582_),
    .X(_04583_));
 sky130_fd_sc_hd__nand2_2 _13657_ (.A(_04535_),
    .B(_03715_),
    .Y(_04584_));
 sky130_fd_sc_hd__nand2_2 _13658_ (.A(_11878_[0]),
    .B(net4084),
    .Y(_04585_));
 sky130_fd_sc_hd__nand2_1 _13659_ (.A(_04584_),
    .B(_04585_),
    .Y(_04586_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1181 ();
 sky130_fd_sc_hd__a221oi_1 _13661_ (.A1(net4090),
    .A2(_04432_),
    .B1(_04586_),
    .B2(_03704_),
    .C1(_03734_),
    .Y(_04588_));
 sky130_fd_sc_hd__nand2_8 _13662_ (.A(net4089),
    .B(_03715_),
    .Y(_04589_));
 sky130_fd_sc_hd__a21oi_1 _13663_ (.A1(_04536_),
    .A2(_04589_),
    .B1(_03704_),
    .Y(_04590_));
 sky130_fd_sc_hd__o21a_1 _13664_ (.A1(_04544_),
    .A2(_04590_),
    .B1(_03735_),
    .X(_04591_));
 sky130_fd_sc_hd__nand2_4 _13665_ (.A(_11862_[0]),
    .B(net4084),
    .Y(_04592_));
 sky130_fd_sc_hd__a21oi_1 _13666_ (.A1(_04574_),
    .A2(_04592_),
    .B1(_03702_),
    .Y(_04593_));
 sky130_fd_sc_hd__a211oi_1 _13667_ (.A1(net4063),
    .A2(_04432_),
    .B1(_04593_),
    .C1(_03735_),
    .Y(_04594_));
 sky130_fd_sc_hd__o21ai_1 _13668_ (.A1(_11878_[0]),
    .A2(_03715_),
    .B1(_04539_),
    .Y(_04595_));
 sky130_fd_sc_hd__nand2_2 _13669_ (.A(_11864_[0]),
    .B(net4084),
    .Y(_04596_));
 sky130_fd_sc_hd__and3_1 _13670_ (.A(_03704_),
    .B(_04574_),
    .C(_04596_),
    .X(_04597_));
 sky130_fd_sc_hd__a21oi_1 _13671_ (.A1(_03702_),
    .A2(_04595_),
    .B1(_04597_),
    .Y(_04598_));
 sky130_fd_sc_hd__nand2_4 _13672_ (.A(_03725_),
    .B(_03734_),
    .Y(_04599_));
 sky130_fd_sc_hd__o32ai_1 _13673_ (.A1(_03725_),
    .A2(_04591_),
    .A3(_04594_),
    .B1(_04598_),
    .B2(_04599_),
    .Y(_04600_));
 sky130_fd_sc_hd__a211oi_1 _13674_ (.A1(_04583_),
    .A2(_04588_),
    .B1(_03751_),
    .C1(_04600_),
    .Y(_04601_));
 sky130_fd_sc_hd__a211oi_1 _13675_ (.A1(_03751_),
    .A2(_04581_),
    .B1(_04601_),
    .C1(_03743_),
    .Y(_04602_));
 sky130_fd_sc_hd__a31oi_2 _13676_ (.A1(_03743_),
    .A2(_04549_),
    .A3(_04563_),
    .B1(_04602_),
    .Y(_00009_));
 sky130_fd_sc_hd__a21oi_1 _13677_ (.A1(_04484_),
    .A2(_04536_),
    .B1(net4087),
    .Y(_04603_));
 sky130_fd_sc_hd__a211oi_1 _13678_ (.A1(_11869_[0]),
    .A2(_04466_),
    .B1(_04603_),
    .C1(_03734_),
    .Y(_04604_));
 sky130_fd_sc_hd__nor2_2 _13679_ (.A(_04499_),
    .B(_04450_),
    .Y(_04605_));
 sky130_fd_sc_hd__a21oi_1 _13680_ (.A1(_11886_[0]),
    .A2(_03715_),
    .B1(_04605_),
    .Y(_04606_));
 sky130_fd_sc_hd__nor2_1 _13681_ (.A(_03735_),
    .B(_04606_),
    .Y(_04607_));
 sky130_fd_sc_hd__nor3_1 _13682_ (.A(_03725_),
    .B(_04604_),
    .C(_04607_),
    .Y(_04608_));
 sky130_fd_sc_hd__nor2_2 _13683_ (.A(net4063),
    .B(_04434_),
    .Y(_04609_));
 sky130_fd_sc_hd__a221oi_1 _13684_ (.A1(_11862_[0]),
    .A2(_04415_),
    .B1(_04432_),
    .B2(_11872_[0]),
    .C1(_04609_),
    .Y(_04610_));
 sky130_fd_sc_hd__nand2_1 _13685_ (.A(_03735_),
    .B(_04610_),
    .Y(_04611_));
 sky130_fd_sc_hd__o211ai_1 _13686_ (.A1(_11867_[0]),
    .A2(_03704_),
    .B1(_03715_),
    .C1(_04559_),
    .Y(_04612_));
 sky130_fd_sc_hd__o211ai_1 _13687_ (.A1(_11883_[0]),
    .A2(_03715_),
    .B1(_03734_),
    .C1(_04612_),
    .Y(_04613_));
 sky130_fd_sc_hd__a21oi_1 _13688_ (.A1(_04611_),
    .A2(_04613_),
    .B1(net4062),
    .Y(_04614_));
 sky130_fd_sc_hd__nor3_1 _13689_ (.A(_03750_),
    .B(_04608_),
    .C(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hd__a21oi_1 _13690_ (.A1(_04485_),
    .A2(_04539_),
    .B1(_03704_),
    .Y(_04616_));
 sky130_fd_sc_hd__o21ai_0 _13691_ (.A1(_11864_[0]),
    .A2(_04434_),
    .B1(_04505_),
    .Y(_04617_));
 sky130_fd_sc_hd__nand2_1 _13692_ (.A(_11867_[0]),
    .B(_03704_),
    .Y(_04618_));
 sky130_fd_sc_hd__o21ai_0 _13693_ (.A1(_11869_[0]),
    .A2(_03704_),
    .B1(_04618_),
    .Y(_04619_));
 sky130_fd_sc_hd__a21oi_1 _13694_ (.A1(_03715_),
    .A2(_04619_),
    .B1(_03725_),
    .Y(_04620_));
 sky130_fd_sc_hd__nor2_4 _13695_ (.A(net4089),
    .B(net4086),
    .Y(_04621_));
 sky130_fd_sc_hd__nor2_4 _13696_ (.A(_11863_[0]),
    .B(_03704_),
    .Y(_04622_));
 sky130_fd_sc_hd__o21ai_0 _13697_ (.A1(_04621_),
    .A2(_04622_),
    .B1(net4084),
    .Y(_04623_));
 sky130_fd_sc_hd__nand3_1 _13698_ (.A(_03734_),
    .B(_04620_),
    .C(_04623_),
    .Y(_04624_));
 sky130_fd_sc_hd__o21ai_0 _13699_ (.A1(_04616_),
    .A2(_04617_),
    .B1(_04624_),
    .Y(_04625_));
 sky130_fd_sc_hd__nand2_1 _13700_ (.A(_11878_[0]),
    .B(_03715_),
    .Y(_04626_));
 sky130_fd_sc_hd__nand2_2 _13701_ (.A(_03696_),
    .B(net4084),
    .Y(_04627_));
 sky130_fd_sc_hd__nand3_1 _13702_ (.A(net4086),
    .B(_04626_),
    .C(_04627_),
    .Y(_04628_));
 sky130_fd_sc_hd__nand2_8 _13703_ (.A(net4090),
    .B(_03715_),
    .Y(_04629_));
 sky130_fd_sc_hd__nand3_1 _13704_ (.A(_03704_),
    .B(_04443_),
    .C(_04629_),
    .Y(_04630_));
 sky130_fd_sc_hd__a21oi_1 _13705_ (.A1(_04628_),
    .A2(_04630_),
    .B1(net4061),
    .Y(_04631_));
 sky130_fd_sc_hd__nor2_1 _13706_ (.A(_11864_[0]),
    .B(_03715_),
    .Y(_04632_));
 sky130_fd_sc_hd__nor2_1 _13707_ (.A(_04500_),
    .B(_04632_),
    .Y(_04633_));
 sky130_fd_sc_hd__nor2_1 _13708_ (.A(_11869_[0]),
    .B(_03715_),
    .Y(_04634_));
 sky130_fd_sc_hd__nor3_1 _13709_ (.A(net4086),
    .B(_04577_),
    .C(_04634_),
    .Y(_04635_));
 sky130_fd_sc_hd__a211oi_1 _13710_ (.A1(net4086),
    .A2(_04633_),
    .B1(_04635_),
    .C1(_03735_),
    .Y(_04636_));
 sky130_fd_sc_hd__nor3_2 _13711_ (.A(net4062),
    .B(_04631_),
    .C(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__nor3_1 _13712_ (.A(_03751_),
    .B(_04625_),
    .C(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__a211oi_1 _13713_ (.A1(_11867_[0]),
    .A2(_03704_),
    .B1(net4084),
    .C1(_04622_),
    .Y(_04639_));
 sky130_fd_sc_hd__a21oi_1 _13714_ (.A1(_11888_[0]),
    .A2(net4084),
    .B1(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__nand2_1 _13715_ (.A(_11890_[0]),
    .B(net4084),
    .Y(_04641_));
 sky130_fd_sc_hd__nor2_2 _13716_ (.A(_03696_),
    .B(_03704_),
    .Y(_04642_));
 sky130_fd_sc_hd__a211o_1 _13717_ (.A1(net4090),
    .A2(_03696_),
    .B1(net4084),
    .C1(_04642_),
    .X(_04643_));
 sky130_fd_sc_hd__a21oi_1 _13718_ (.A1(_04641_),
    .A2(_04643_),
    .B1(_03735_),
    .Y(_04644_));
 sky130_fd_sc_hd__a21oi_1 _13719_ (.A1(_03735_),
    .A2(_04640_),
    .B1(_04644_),
    .Y(_04645_));
 sky130_fd_sc_hd__nor2_1 _13720_ (.A(_11876_[0]),
    .B(_04450_),
    .Y(_04646_));
 sky130_fd_sc_hd__nor2_1 _13721_ (.A(_03735_),
    .B(_04646_),
    .Y(_04647_));
 sky130_fd_sc_hd__o21ai_0 _13722_ (.A1(_04411_),
    .A2(_04442_),
    .B1(_03704_),
    .Y(_04648_));
 sky130_fd_sc_hd__nor2_1 _13723_ (.A(_11863_[0]),
    .B(_04450_),
    .Y(_04649_));
 sky130_fd_sc_hd__nand2_4 _13724_ (.A(_03725_),
    .B(_03735_),
    .Y(_04650_));
 sky130_fd_sc_hd__a211oi_1 _13725_ (.A1(_11883_[0]),
    .A2(_03715_),
    .B1(_04649_),
    .C1(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__a32oi_1 _13726_ (.A1(_04583_),
    .A2(_04647_),
    .A3(_04648_),
    .B1(_04651_),
    .B2(_04512_),
    .Y(_04652_));
 sky130_fd_sc_hd__o21ai_2 _13727_ (.A1(_03725_),
    .A2(_04645_),
    .B1(_04652_),
    .Y(_04653_));
 sky130_fd_sc_hd__and2_0 _13728_ (.A(_11863_[0]),
    .B(_03715_),
    .X(_04654_));
 sky130_fd_sc_hd__nor2_2 _13729_ (.A(_11874_[0]),
    .B(_03715_),
    .Y(_04655_));
 sky130_fd_sc_hd__nand3_1 _13730_ (.A(_03704_),
    .B(_04574_),
    .C(_04538_),
    .Y(_04656_));
 sky130_fd_sc_hd__o31ai_1 _13731_ (.A1(_03704_),
    .A2(_04654_),
    .A3(_04655_),
    .B1(_04656_),
    .Y(_04657_));
 sky130_fd_sc_hd__nand2_1 _13732_ (.A(_11869_[0]),
    .B(_03715_),
    .Y(_04658_));
 sky130_fd_sc_hd__a21oi_2 _13733_ (.A1(_04658_),
    .A2(_04596_),
    .B1(_03704_),
    .Y(_04659_));
 sky130_fd_sc_hd__o31ai_1 _13734_ (.A1(_03704_),
    .A2(_04577_),
    .A3(_04632_),
    .B1(_03735_),
    .Y(_04660_));
 sky130_fd_sc_hd__nor2_1 _13735_ (.A(_11874_[0]),
    .B(net4084),
    .Y(_04661_));
 sky130_fd_sc_hd__nor3_1 _13736_ (.A(net4086),
    .B(_04501_),
    .C(_04661_),
    .Y(_04662_));
 sky130_fd_sc_hd__o32ai_2 _13737_ (.A1(_03735_),
    .A2(_04609_),
    .A3(_04659_),
    .B1(_04660_),
    .B2(_04662_),
    .Y(_04663_));
 sky130_fd_sc_hd__nor2_1 _13738_ (.A(_03704_),
    .B(_03725_),
    .Y(_04664_));
 sky130_fd_sc_hd__nor3_1 _13739_ (.A(net4087),
    .B(_03725_),
    .C(_04589_),
    .Y(_04665_));
 sky130_fd_sc_hd__a221oi_1 _13740_ (.A1(_11874_[0]),
    .A2(_04423_),
    .B1(_04664_),
    .B2(_11869_[0]),
    .C1(_04665_),
    .Y(_04666_));
 sky130_fd_sc_hd__o22ai_1 _13741_ (.A1(net4062),
    .A2(_04663_),
    .B1(_04666_),
    .B2(_03735_),
    .Y(_04667_));
 sky130_fd_sc_hd__a211oi_1 _13742_ (.A1(_04505_),
    .A2(_04657_),
    .B1(_04667_),
    .C1(_03751_),
    .Y(_04668_));
 sky130_fd_sc_hd__a211o_1 _13743_ (.A1(_03751_),
    .A2(_04653_),
    .B1(_04668_),
    .C1(net3711),
    .X(_04669_));
 sky130_fd_sc_hd__o31ai_2 _13744_ (.A1(_03744_),
    .A2(_04615_),
    .A3(_04638_),
    .B1(_04669_),
    .Y(_00010_));
 sky130_fd_sc_hd__a21boi_0 _13745_ (.A1(_03735_),
    .A2(_04513_),
    .B1_N(_04626_),
    .Y(_04670_));
 sky130_fd_sc_hd__o21ai_0 _13746_ (.A1(net4087),
    .A2(_04670_),
    .B1(_03725_),
    .Y(_04671_));
 sky130_fd_sc_hd__nand2_4 _13747_ (.A(_03704_),
    .B(net4085),
    .Y(_04672_));
 sky130_fd_sc_hd__nor2_1 _13748_ (.A(net4089),
    .B(_04672_),
    .Y(_04673_));
 sky130_fd_sc_hd__nand2b_4 _13749_ (.A_N(_11872_[0]),
    .B(net4084),
    .Y(_04674_));
 sky130_fd_sc_hd__a21oi_1 _13750_ (.A1(_04574_),
    .A2(_04674_),
    .B1(_03704_),
    .Y(_04675_));
 sky130_fd_sc_hd__o21ai_0 _13751_ (.A1(net4090),
    .A2(_03734_),
    .B1(_03704_),
    .Y(_04676_));
 sky130_fd_sc_hd__o31ai_1 _13752_ (.A1(_04482_),
    .A2(_04513_),
    .A3(_04676_),
    .B1(net4062),
    .Y(_04677_));
 sky130_fd_sc_hd__nor2_4 _13753_ (.A(net4063),
    .B(net4087),
    .Y(_04678_));
 sky130_fd_sc_hd__nand2_1 _13754_ (.A(_04538_),
    .B(_04486_),
    .Y(_04679_));
 sky130_fd_sc_hd__o21ai_0 _13755_ (.A1(_04678_),
    .A2(_04679_),
    .B1(_03734_),
    .Y(_04680_));
 sky130_fd_sc_hd__o32ai_1 _13756_ (.A1(_04671_),
    .A2(_04673_),
    .A3(_04675_),
    .B1(_04677_),
    .B2(_04680_),
    .Y(_04681_));
 sky130_fd_sc_hd__a221o_1 _13757_ (.A1(net4090),
    .A2(_04423_),
    .B1(_04568_),
    .B2(_11874_[0]),
    .C1(_04677_),
    .X(_04682_));
 sky130_fd_sc_hd__a21oi_1 _13758_ (.A1(_04671_),
    .A2(_04682_),
    .B1(_03734_),
    .Y(_04683_));
 sky130_fd_sc_hd__nor2_2 _13759_ (.A(net4088),
    .B(net4085),
    .Y(_04684_));
 sky130_fd_sc_hd__a21oi_1 _13760_ (.A1(_04469_),
    .A2(_04589_),
    .B1(_03704_),
    .Y(_04685_));
 sky130_fd_sc_hd__a221oi_1 _13761_ (.A1(_11863_[0]),
    .A2(_04684_),
    .B1(_04510_),
    .B2(net4063),
    .C1(_04685_),
    .Y(_04686_));
 sky130_fd_sc_hd__nor3_1 _13762_ (.A(_03704_),
    .B(_04517_),
    .C(_04510_),
    .Y(_04687_));
 sky130_fd_sc_hd__a311oi_1 _13763_ (.A1(_03704_),
    .A2(_04443_),
    .A3(_04486_),
    .B1(_04687_),
    .C1(_03734_),
    .Y(_04688_));
 sky130_fd_sc_hd__a21oi_1 _13764_ (.A1(_03734_),
    .A2(_04686_),
    .B1(_04688_),
    .Y(_04689_));
 sky130_fd_sc_hd__o32ai_1 _13765_ (.A1(_11883_[0]),
    .A2(_03715_),
    .A3(_04678_),
    .B1(_04565_),
    .B2(_11863_[0]),
    .Y(_04690_));
 sky130_fd_sc_hd__nor3_1 _13766_ (.A(_03704_),
    .B(_04427_),
    .C(_04543_),
    .Y(_04691_));
 sky130_fd_sc_hd__a311o_1 _13767_ (.A1(_03704_),
    .A2(_04584_),
    .A3(_04674_),
    .B1(_04691_),
    .C1(net4061),
    .X(_04692_));
 sky130_fd_sc_hd__o211ai_1 _13768_ (.A1(_03735_),
    .A2(_04690_),
    .B1(_04692_),
    .C1(_03725_),
    .Y(_04693_));
 sky130_fd_sc_hd__o211ai_1 _13769_ (.A1(_03725_),
    .A2(_04689_),
    .B1(_04693_),
    .C1(_03751_),
    .Y(_04694_));
 sky130_fd_sc_hd__o31ai_1 _13770_ (.A1(_03751_),
    .A2(_04681_),
    .A3(_04683_),
    .B1(_04694_),
    .Y(_04695_));
 sky130_fd_sc_hd__o22ai_1 _13771_ (.A1(_03696_),
    .A2(_04450_),
    .B1(_04434_),
    .B2(_11876_[0]),
    .Y(_04696_));
 sky130_fd_sc_hd__a21oi_1 _13772_ (.A1(_03704_),
    .A2(_04627_),
    .B1(net4063),
    .Y(_04697_));
 sky130_fd_sc_hd__nand2_8 _13773_ (.A(_11874_[0]),
    .B(_03715_),
    .Y(_04698_));
 sky130_fd_sc_hd__and3_1 _13774_ (.A(net4086),
    .B(_04674_),
    .C(_04698_),
    .X(_04699_));
 sky130_fd_sc_hd__a21oi_1 _13775_ (.A1(_04629_),
    .A2(_04592_),
    .B1(net4087),
    .Y(_04700_));
 sky130_fd_sc_hd__o21ai_0 _13776_ (.A1(_04699_),
    .A2(_04700_),
    .B1(net4061),
    .Y(_04701_));
 sky130_fd_sc_hd__o311ai_0 _13777_ (.A1(net4061),
    .A2(_04696_),
    .A3(_04697_),
    .B1(_04701_),
    .C1(net4062),
    .Y(_04702_));
 sky130_fd_sc_hd__nand3_1 _13778_ (.A(_03735_),
    .B(_04443_),
    .C(_04698_),
    .Y(_04703_));
 sky130_fd_sc_hd__o21ai_0 _13779_ (.A1(_03735_),
    .A2(_04538_),
    .B1(_04703_),
    .Y(_04704_));
 sky130_fd_sc_hd__a21oi_1 _13780_ (.A1(_03735_),
    .A2(_04482_),
    .B1(_04632_),
    .Y(_04705_));
 sky130_fd_sc_hd__nand2_1 _13781_ (.A(net4087),
    .B(_04705_),
    .Y(_04706_));
 sky130_fd_sc_hd__o21ai_0 _13782_ (.A1(net4087),
    .A2(_04704_),
    .B1(_04706_),
    .Y(_04707_));
 sky130_fd_sc_hd__a21oi_1 _13783_ (.A1(_03725_),
    .A2(_04707_),
    .B1(_03751_),
    .Y(_04708_));
 sky130_fd_sc_hd__o21ai_0 _13784_ (.A1(_11874_[0]),
    .A2(_03715_),
    .B1(_04486_),
    .Y(_04709_));
 sky130_fd_sc_hd__a21oi_1 _13785_ (.A1(_04412_),
    .A2(_04443_),
    .B1(net4087),
    .Y(_04710_));
 sky130_fd_sc_hd__a21oi_1 _13786_ (.A1(net4087),
    .A2(_04709_),
    .B1(_04710_),
    .Y(_04711_));
 sky130_fd_sc_hd__a21oi_1 _13787_ (.A1(_04629_),
    .A2(_04674_),
    .B1(_03704_),
    .Y(_04712_));
 sky130_fd_sc_hd__o22ai_1 _13788_ (.A1(_11863_[0]),
    .A2(_04672_),
    .B1(_04589_),
    .B2(net4090),
    .Y(_04713_));
 sky130_fd_sc_hd__or3_1 _13789_ (.A(_04650_),
    .B(_04712_),
    .C(_04713_),
    .X(_04714_));
 sky130_fd_sc_hd__nand2_1 _13790_ (.A(_11867_[0]),
    .B(_04466_),
    .Y(_04715_));
 sky130_fd_sc_hd__nor2_1 _13791_ (.A(net4090),
    .B(_03696_),
    .Y(_04716_));
 sky130_fd_sc_hd__o21ai_0 _13792_ (.A1(_04678_),
    .A2(_04716_),
    .B1(net4084),
    .Y(_04717_));
 sky130_fd_sc_hd__a21oi_1 _13793_ (.A1(_04715_),
    .A2(_04717_),
    .B1(_03735_),
    .Y(_04718_));
 sky130_fd_sc_hd__o21ai_0 _13794_ (.A1(_04440_),
    .A2(_04442_),
    .B1(_03704_),
    .Y(_04719_));
 sky130_fd_sc_hd__o311a_1 _13795_ (.A1(_03704_),
    .A2(_04500_),
    .A3(_04513_),
    .B1(_04719_),
    .C1(_03735_),
    .X(_04720_));
 sky130_fd_sc_hd__o21ai_0 _13796_ (.A1(_04718_),
    .A2(_04720_),
    .B1(net4062),
    .Y(_04721_));
 sky130_fd_sc_hd__o211ai_1 _13797_ (.A1(_04599_),
    .A2(_04711_),
    .B1(_04714_),
    .C1(_04721_),
    .Y(_04722_));
 sky130_fd_sc_hd__a221oi_1 _13798_ (.A1(_04702_),
    .A2(_04708_),
    .B1(_04722_),
    .B2(_03751_),
    .C1(net3711),
    .Y(_04723_));
 sky130_fd_sc_hd__a21o_4 _13799_ (.A1(net3711),
    .A2(_04695_),
    .B1(_04723_),
    .X(_00011_));
 sky130_fd_sc_hd__o21ai_0 _13800_ (.A1(_04452_),
    .A2(_04577_),
    .B1(_03704_),
    .Y(_04724_));
 sky130_fd_sc_hd__nand3_1 _13801_ (.A(_03743_),
    .B(_04467_),
    .C(_04724_),
    .Y(_04725_));
 sky130_fd_sc_hd__nand3_1 _13802_ (.A(_03702_),
    .B(_03744_),
    .C(_04595_),
    .Y(_04726_));
 sky130_fd_sc_hd__and2_0 _13803_ (.A(_11869_[0]),
    .B(_03704_),
    .X(_04727_));
 sky130_fd_sc_hd__o21ai_0 _13804_ (.A1(_04622_),
    .A2(_04727_),
    .B1(net4084),
    .Y(_04728_));
 sky130_fd_sc_hd__a21oi_1 _13805_ (.A1(_04592_),
    .A2(_04582_),
    .B1(_03744_),
    .Y(_04729_));
 sky130_fd_sc_hd__a311oi_1 _13806_ (.A1(_03744_),
    .A2(_04497_),
    .A3(_04728_),
    .B1(_04729_),
    .C1(_03725_),
    .Y(_04730_));
 sky130_fd_sc_hd__a31oi_1 _13807_ (.A1(_03725_),
    .A2(_04725_),
    .A3(_04726_),
    .B1(_04730_),
    .Y(_04731_));
 sky130_fd_sc_hd__nand2_1 _13808_ (.A(_11892_[0]),
    .B(_03715_),
    .Y(_04732_));
 sky130_fd_sc_hd__nor4b_1 _13809_ (.A(_03743_),
    .B(_04646_),
    .C(_04678_),
    .D_N(_04732_),
    .Y(_04733_));
 sky130_fd_sc_hd__a21oi_1 _13810_ (.A1(_04443_),
    .A2(_04698_),
    .B1(_03704_),
    .Y(_04734_));
 sky130_fd_sc_hd__a211oi_1 _13811_ (.A1(_03704_),
    .A2(_04633_),
    .B1(_04734_),
    .C1(_03744_),
    .Y(_04735_));
 sky130_fd_sc_hd__o21ai_0 _13812_ (.A1(_04733_),
    .A2(_04735_),
    .B1(net4062),
    .Y(_04736_));
 sky130_fd_sc_hd__o2111ai_1 _13813_ (.A1(_03702_),
    .A2(_04516_),
    .B1(_04698_),
    .C1(_03725_),
    .D1(_03744_),
    .Y(_04737_));
 sky130_fd_sc_hd__a21oi_1 _13814_ (.A1(_11874_[0]),
    .A2(_03704_),
    .B1(_03744_),
    .Y(_04738_));
 sky130_fd_sc_hd__nand3_1 _13815_ (.A(_04523_),
    .B(_04583_),
    .C(_04738_),
    .Y(_04739_));
 sky130_fd_sc_hd__nand4_1 _13816_ (.A(_03751_),
    .B(_04736_),
    .C(_04737_),
    .D(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__o21ai_0 _13817_ (.A1(_03751_),
    .A2(_04731_),
    .B1(_04740_),
    .Y(_04741_));
 sky130_fd_sc_hd__nor2_2 _13818_ (.A(net4090),
    .B(_04412_),
    .Y(_04742_));
 sky130_fd_sc_hd__a21oi_1 _13819_ (.A1(_04629_),
    .A2(_04585_),
    .B1(_03702_),
    .Y(_04743_));
 sky130_fd_sc_hd__nor3_1 _13820_ (.A(_04646_),
    .B(_04742_),
    .C(_04743_),
    .Y(_04744_));
 sky130_fd_sc_hd__o221ai_1 _13821_ (.A1(_11864_[0]),
    .A2(_04450_),
    .B1(_04501_),
    .B2(_03702_),
    .C1(_03744_),
    .Y(_04745_));
 sky130_fd_sc_hd__o21ai_0 _13822_ (.A1(_03744_),
    .A2(_04744_),
    .B1(_04745_),
    .Y(_04746_));
 sky130_fd_sc_hd__nand2_1 _13823_ (.A(net4062),
    .B(_04746_),
    .Y(_04747_));
 sky130_fd_sc_hd__a21oi_1 _13824_ (.A1(_04536_),
    .A2(_04658_),
    .B1(_03702_),
    .Y(_04748_));
 sky130_fd_sc_hd__nor2_2 _13825_ (.A(net4090),
    .B(_04411_),
    .Y(_04749_));
 sky130_fd_sc_hd__o21ai_0 _13826_ (.A1(_04543_),
    .A2(_04749_),
    .B1(_03704_),
    .Y(_04750_));
 sky130_fd_sc_hd__o2111ai_1 _13827_ (.A1(_03696_),
    .A2(_04469_),
    .B1(_04467_),
    .C1(_04750_),
    .D1(_03743_),
    .Y(_04751_));
 sky130_fd_sc_hd__o311ai_0 _13828_ (.A1(_03743_),
    .A2(_04545_),
    .A3(_04748_),
    .B1(_04751_),
    .C1(_03725_),
    .Y(_04752_));
 sky130_fd_sc_hd__a21oi_1 _13829_ (.A1(_04747_),
    .A2(_04752_),
    .B1(_03751_),
    .Y(_04753_));
 sky130_fd_sc_hd__o21ai_0 _13830_ (.A1(_04432_),
    .A2(_04678_),
    .B1(net4089),
    .Y(_04754_));
 sky130_fd_sc_hd__o21ai_1 _13831_ (.A1(_04470_),
    .A2(_04642_),
    .B1(_04754_),
    .Y(_04755_));
 sky130_fd_sc_hd__a21oi_1 _13832_ (.A1(_11876_[0]),
    .A2(_04466_),
    .B1(_04621_),
    .Y(_04756_));
 sky130_fd_sc_hd__nor2_1 _13833_ (.A(net4062),
    .B(_04756_),
    .Y(_04757_));
 sky130_fd_sc_hd__a221oi_1 _13834_ (.A1(_04543_),
    .A2(_04491_),
    .B1(_04755_),
    .B2(net4062),
    .C1(_04757_),
    .Y(_04758_));
 sky130_fd_sc_hd__o21ai_1 _13835_ (.A1(_11864_[0]),
    .A2(_03715_),
    .B1(_04412_),
    .Y(_04759_));
 sky130_fd_sc_hd__nand2_1 _13836_ (.A(net4086),
    .B(_04759_),
    .Y(_04760_));
 sky130_fd_sc_hd__o21ai_0 _13837_ (.A1(_04500_),
    .A2(_04634_),
    .B1(_03704_),
    .Y(_04761_));
 sky130_fd_sc_hd__a311oi_1 _13838_ (.A1(net4086),
    .A2(_04552_),
    .A3(_04589_),
    .B1(_03725_),
    .C1(_04472_),
    .Y(_04762_));
 sky130_fd_sc_hd__a311o_1 _13839_ (.A1(_03725_),
    .A2(_04760_),
    .A3(_04761_),
    .B1(_03744_),
    .C1(_04762_),
    .X(_04763_));
 sky130_fd_sc_hd__o21ai_0 _13840_ (.A1(_03743_),
    .A2(_04758_),
    .B1(_04763_),
    .Y(_04764_));
 sky130_fd_sc_hd__o21ai_0 _13841_ (.A1(_03750_),
    .A2(_04764_),
    .B1(_03734_),
    .Y(_04765_));
 sky130_fd_sc_hd__o22a_4 _13842_ (.A1(_03734_),
    .A2(_04741_),
    .B1(_04753_),
    .B2(_04765_),
    .X(_00012_));
 sky130_fd_sc_hd__nand2_1 _13843_ (.A(_11872_[0]),
    .B(_04466_),
    .Y(_04766_));
 sky130_fd_sc_hd__a221oi_1 _13844_ (.A1(net4090),
    .A2(_04411_),
    .B1(_04450_),
    .B2(_03696_),
    .C1(_03725_),
    .Y(_04767_));
 sky130_fd_sc_hd__a41oi_1 _13845_ (.A1(_03725_),
    .A2(_04541_),
    .A3(_04551_),
    .A4(_04766_),
    .B1(_04767_),
    .Y(_04768_));
 sky130_fd_sc_hd__a21oi_1 _13846_ (.A1(_04584_),
    .A2(_04596_),
    .B1(_03704_),
    .Y(_04769_));
 sky130_fd_sc_hd__a21oi_1 _13847_ (.A1(_11878_[0]),
    .A2(_03702_),
    .B1(_04621_),
    .Y(_04770_));
 sky130_fd_sc_hd__o21ai_0 _13848_ (.A1(_03715_),
    .A2(_04770_),
    .B1(_04583_),
    .Y(_04771_));
 sky130_fd_sc_hd__o311ai_0 _13849_ (.A1(_03725_),
    .A2(_04435_),
    .A3(_04769_),
    .B1(_04771_),
    .C1(_03734_),
    .Y(_04772_));
 sky130_fd_sc_hd__o21ai_2 _13850_ (.A1(_03734_),
    .A2(_04768_),
    .B1(_04772_),
    .Y(_04773_));
 sky130_fd_sc_hd__nand2_2 _13851_ (.A(_03751_),
    .B(_04773_),
    .Y(_04774_));
 sky130_fd_sc_hd__o21ai_0 _13852_ (.A1(_11864_[0]),
    .A2(_03704_),
    .B1(_03715_),
    .Y(_04775_));
 sky130_fd_sc_hd__a21oi_1 _13853_ (.A1(_11864_[0]),
    .A2(net4084),
    .B1(_04442_),
    .Y(_04776_));
 sky130_fd_sc_hd__o21ai_0 _13854_ (.A1(_04654_),
    .A2(_04513_),
    .B1(_03704_),
    .Y(_04777_));
 sky130_fd_sc_hd__o21ai_0 _13855_ (.A1(_03704_),
    .A2(_04776_),
    .B1(_04777_),
    .Y(_04778_));
 sky130_fd_sc_hd__nor2_1 _13856_ (.A(_03735_),
    .B(_04778_),
    .Y(_04779_));
 sky130_fd_sc_hd__a31oi_1 _13857_ (.A1(_03735_),
    .A2(_04523_),
    .A3(_04775_),
    .B1(_04779_),
    .Y(_04780_));
 sky130_fd_sc_hd__a21oi_1 _13858_ (.A1(_11872_[0]),
    .A2(_03715_),
    .B1(_03735_),
    .Y(_04781_));
 sky130_fd_sc_hd__o21ai_0 _13859_ (.A1(_03715_),
    .A2(_04496_),
    .B1(_04781_),
    .Y(_04782_));
 sky130_fd_sc_hd__o311ai_0 _13860_ (.A1(_03734_),
    .A2(_04605_),
    .A3(_04700_),
    .B1(_04782_),
    .C1(net4062),
    .Y(_04783_));
 sky130_fd_sc_hd__o211ai_1 _13861_ (.A1(net4062),
    .A2(_04780_),
    .B1(_04783_),
    .C1(_03750_),
    .Y(_04784_));
 sky130_fd_sc_hd__a21oi_1 _13862_ (.A1(net4090),
    .A2(_04423_),
    .B1(_04749_),
    .Y(_04785_));
 sky130_fd_sc_hd__o2111ai_1 _13863_ (.A1(_11862_[0]),
    .A2(_04434_),
    .B1(_04523_),
    .C1(_03734_),
    .D1(_04416_),
    .Y(_04786_));
 sky130_fd_sc_hd__o21ai_0 _13864_ (.A1(_03734_),
    .A2(_04785_),
    .B1(_04786_),
    .Y(_04787_));
 sky130_fd_sc_hd__o221ai_1 _13865_ (.A1(_11862_[0]),
    .A2(_04672_),
    .B1(_04776_),
    .B2(_03704_),
    .C1(_03734_),
    .Y(_04788_));
 sky130_fd_sc_hd__nand3_1 _13866_ (.A(_03704_),
    .B(_04574_),
    .C(_04627_),
    .Y(_04789_));
 sky130_fd_sc_hd__o311ai_1 _13867_ (.A1(_03704_),
    .A2(_04500_),
    .A3(_04655_),
    .B1(_04789_),
    .C1(_03735_),
    .Y(_04790_));
 sky130_fd_sc_hd__nand3_1 _13868_ (.A(_03725_),
    .B(_04788_),
    .C(_04790_),
    .Y(_04791_));
 sky130_fd_sc_hd__o21ai_0 _13869_ (.A1(_03725_),
    .A2(_04787_),
    .B1(_04791_),
    .Y(_04792_));
 sky130_fd_sc_hd__nand2_1 _13870_ (.A(_03750_),
    .B(_04792_),
    .Y(_04793_));
 sky130_fd_sc_hd__nand3_1 _13871_ (.A(_03704_),
    .B(_04443_),
    .C(_04698_),
    .Y(_04794_));
 sky130_fd_sc_hd__nand2_1 _13872_ (.A(net4087),
    .B(_04482_),
    .Y(_04795_));
 sky130_fd_sc_hd__a211oi_1 _13873_ (.A1(_04794_),
    .A2(_04795_),
    .B1(_03725_),
    .C1(_03735_),
    .Y(_04796_));
 sky130_fd_sc_hd__nor3_1 _13874_ (.A(_03704_),
    .B(_04517_),
    .C(_04655_),
    .Y(_04797_));
 sky130_fd_sc_hd__a311oi_1 _13875_ (.A1(_03704_),
    .A2(_04629_),
    .A3(_04485_),
    .B1(_04650_),
    .C1(_04797_),
    .Y(_04798_));
 sky130_fd_sc_hd__o21ai_0 _13876_ (.A1(_03704_),
    .A2(_04500_),
    .B1(_04552_),
    .Y(_04799_));
 sky130_fd_sc_hd__nor2_1 _13877_ (.A(_04599_),
    .B(_04799_),
    .Y(_04800_));
 sky130_fd_sc_hd__nor3_2 _13878_ (.A(_04796_),
    .B(_04798_),
    .C(_04800_),
    .Y(_04801_));
 sky130_fd_sc_hd__a21oi_1 _13879_ (.A1(_11864_[0]),
    .A2(_03702_),
    .B1(_04727_),
    .Y(_04802_));
 sky130_fd_sc_hd__o211ai_1 _13880_ (.A1(net4084),
    .A2(_04802_),
    .B1(_04494_),
    .C1(_03735_),
    .Y(_04803_));
 sky130_fd_sc_hd__a31oi_2 _13881_ (.A1(_03751_),
    .A2(_04801_),
    .A3(_04803_),
    .B1(net3711),
    .Y(_04804_));
 sky130_fd_sc_hd__a32oi_4 _13882_ (.A1(net3711),
    .A2(_04774_),
    .A3(_04784_),
    .B1(_04793_),
    .B2(_04804_),
    .Y(_00013_));
 sky130_fd_sc_hd__a21oi_1 _13883_ (.A1(net4087),
    .A2(_04464_),
    .B1(_04710_),
    .Y(_04805_));
 sky130_fd_sc_hd__nor2_1 _13884_ (.A(_03734_),
    .B(_04805_),
    .Y(_04806_));
 sky130_fd_sc_hd__nor2_1 _13885_ (.A(_11867_[0]),
    .B(_04434_),
    .Y(_04807_));
 sky130_fd_sc_hd__nor4_1 _13886_ (.A(_03735_),
    .B(_04649_),
    .C(_04569_),
    .D(_04807_),
    .Y(_04808_));
 sky130_fd_sc_hd__a21oi_1 _13887_ (.A1(_04412_),
    .A2(_04674_),
    .B1(_03704_),
    .Y(_04809_));
 sky130_fd_sc_hd__nand2_1 _13888_ (.A(_11867_[0]),
    .B(net4088),
    .Y(_04810_));
 sky130_fd_sc_hd__o211ai_1 _13889_ (.A1(_11863_[0]),
    .A2(net4088),
    .B1(net4085),
    .C1(_04810_),
    .Y(_04811_));
 sky130_fd_sc_hd__o211ai_1 _13890_ (.A1(_11886_[0]),
    .A2(net4085),
    .B1(_03735_),
    .C1(_04811_),
    .Y(_04812_));
 sky130_fd_sc_hd__o311ai_0 _13891_ (.A1(_03735_),
    .A2(_04807_),
    .A3(_04809_),
    .B1(_04812_),
    .C1(_03725_),
    .Y(_04813_));
 sky130_fd_sc_hd__o311ai_1 _13892_ (.A1(_03725_),
    .A2(_04806_),
    .A3(_04808_),
    .B1(_03751_),
    .C1(_04813_),
    .Y(_04814_));
 sky130_fd_sc_hd__nor2_1 _13893_ (.A(_11882_[0]),
    .B(net4085),
    .Y(_04815_));
 sky130_fd_sc_hd__nor2_1 _13894_ (.A(_11874_[0]),
    .B(_03704_),
    .Y(_04816_));
 sky130_fd_sc_hd__nor3_1 _13895_ (.A(_03715_),
    .B(_04621_),
    .C(_04816_),
    .Y(_04817_));
 sky130_fd_sc_hd__nor3_1 _13896_ (.A(_03725_),
    .B(_04815_),
    .C(_04817_),
    .Y(_04818_));
 sky130_fd_sc_hd__nor2_1 _13897_ (.A(_03704_),
    .B(_04679_),
    .Y(_04819_));
 sky130_fd_sc_hd__o31ai_1 _13898_ (.A1(net4062),
    .A2(_04435_),
    .A3(_04819_),
    .B1(_03735_),
    .Y(_04820_));
 sky130_fd_sc_hd__nand3_1 _13899_ (.A(net4087),
    .B(_04674_),
    .C(_04698_),
    .Y(_04821_));
 sky130_fd_sc_hd__a21oi_1 _13900_ (.A1(_03696_),
    .A2(_04684_),
    .B1(net4062),
    .Y(_04822_));
 sky130_fd_sc_hd__a21oi_1 _13901_ (.A1(_04821_),
    .A2(_04822_),
    .B1(_04620_),
    .Y(_04823_));
 sky130_fd_sc_hd__o221ai_1 _13902_ (.A1(_04818_),
    .A2(_04820_),
    .B1(_04823_),
    .B2(_03735_),
    .C1(_03750_),
    .Y(_04824_));
 sky130_fd_sc_hd__nand3_2 _13903_ (.A(net3711),
    .B(_04814_),
    .C(_04824_),
    .Y(_04825_));
 sky130_fd_sc_hd__a21oi_1 _13904_ (.A1(_04536_),
    .A2(_04698_),
    .B1(net4087),
    .Y(_04826_));
 sky130_fd_sc_hd__a21oi_1 _13905_ (.A1(_11878_[0]),
    .A2(_04466_),
    .B1(_04826_),
    .Y(_04827_));
 sky130_fd_sc_hd__a2111oi_0 _13906_ (.A1(_11874_[0]),
    .A2(_04684_),
    .B1(_04649_),
    .C1(_04569_),
    .D1(_03735_),
    .Y(_04828_));
 sky130_fd_sc_hd__a21oi_1 _13907_ (.A1(_03735_),
    .A2(_04827_),
    .B1(_04828_),
    .Y(_04829_));
 sky130_fd_sc_hd__nand2_1 _13908_ (.A(_03696_),
    .B(_04565_),
    .Y(_04830_));
 sky130_fd_sc_hd__o211ai_1 _13909_ (.A1(_03696_),
    .A2(_04629_),
    .B1(_04830_),
    .C1(_04505_),
    .Y(_04831_));
 sky130_fd_sc_hd__mux2i_1 _13910_ (.A0(_11864_[0]),
    .A1(_11874_[0]),
    .S(net4088),
    .Y(_04832_));
 sky130_fd_sc_hd__o21ai_0 _13911_ (.A1(_11862_[0]),
    .A2(_03704_),
    .B1(_04492_),
    .Y(_04833_));
 sky130_fd_sc_hd__nand2_1 _13912_ (.A(_03715_),
    .B(_04833_),
    .Y(_04834_));
 sky130_fd_sc_hd__o2111ai_1 _13913_ (.A1(_03715_),
    .A2(_04832_),
    .B1(_04834_),
    .C1(net4062),
    .D1(_03734_),
    .Y(_04835_));
 sky130_fd_sc_hd__nor2_1 _13914_ (.A(net3711),
    .B(_03750_),
    .Y(_04836_));
 sky130_fd_sc_hd__o2111ai_2 _13915_ (.A1(net4062),
    .A2(_04829_),
    .B1(_04831_),
    .C1(_04835_),
    .D1(_04836_),
    .Y(_04837_));
 sky130_fd_sc_hd__o21ai_0 _13916_ (.A1(net4090),
    .A2(net4088),
    .B1(_04810_),
    .Y(_04838_));
 sky130_fd_sc_hd__nand2_1 _13917_ (.A(net4085),
    .B(_04838_),
    .Y(_04839_));
 sky130_fd_sc_hd__o22ai_1 _13918_ (.A1(net4063),
    .A2(_03704_),
    .B1(_04672_),
    .B2(_11864_[0]),
    .Y(_04840_));
 sky130_fd_sc_hd__nor3_2 _13919_ (.A(net4061),
    .B(_04742_),
    .C(_04840_),
    .Y(_04841_));
 sky130_fd_sc_hd__a31oi_1 _13920_ (.A1(_03734_),
    .A2(_04557_),
    .A3(_04839_),
    .B1(_04841_),
    .Y(_04842_));
 sky130_fd_sc_hd__nand2_1 _13921_ (.A(net4087),
    .B(_04470_),
    .Y(_04843_));
 sky130_fd_sc_hd__a2111oi_0 _13922_ (.A1(net4089),
    .A2(_04843_),
    .B1(_04605_),
    .C1(_04609_),
    .D1(_03734_),
    .Y(_04844_));
 sky130_fd_sc_hd__a311oi_1 _13923_ (.A1(_03734_),
    .A2(_04794_),
    .A3(_04843_),
    .B1(_04844_),
    .C1(_03725_),
    .Y(_04845_));
 sky130_fd_sc_hd__a21oi_1 _13924_ (.A1(_03725_),
    .A2(_04842_),
    .B1(_04845_),
    .Y(_04846_));
 sky130_fd_sc_hd__nand3_1 _13925_ (.A(_03744_),
    .B(_03750_),
    .C(_04846_),
    .Y(_04847_));
 sky130_fd_sc_hd__nand3_4 _13926_ (.A(_04825_),
    .B(_04837_),
    .C(_04847_),
    .Y(_00014_));
 sky130_fd_sc_hd__nor3_1 _13927_ (.A(_03704_),
    .B(_04440_),
    .C(_04442_),
    .Y(_04848_));
 sky130_fd_sc_hd__a31oi_1 _13928_ (.A1(_03704_),
    .A2(_04574_),
    .A3(_04536_),
    .B1(_04848_),
    .Y(_04849_));
 sky130_fd_sc_hd__nor2_1 _13929_ (.A(_04535_),
    .B(_03702_),
    .Y(_04850_));
 sky130_fd_sc_hd__a311oi_1 _13930_ (.A1(_03702_),
    .A2(_04412_),
    .A3(_04585_),
    .B1(_04850_),
    .C1(_03735_),
    .Y(_04851_));
 sky130_fd_sc_hd__a21oi_1 _13931_ (.A1(_03735_),
    .A2(_04849_),
    .B1(_04851_),
    .Y(_04852_));
 sky130_fd_sc_hd__nor3b_1 _13932_ (.A(_03704_),
    .B(_04440_),
    .C_N(_04698_),
    .Y(_04853_));
 sky130_fd_sc_hd__a31oi_1 _13933_ (.A1(_03704_),
    .A2(_04470_),
    .A3(_04627_),
    .B1(_04853_),
    .Y(_04854_));
 sky130_fd_sc_hd__o211ai_1 _13934_ (.A1(net4090),
    .A2(_03696_),
    .B1(_03715_),
    .C1(_04491_),
    .Y(_04855_));
 sky130_fd_sc_hd__a31oi_1 _13935_ (.A1(net4061),
    .A2(_04552_),
    .A3(_04855_),
    .B1(net4062),
    .Y(_04856_));
 sky130_fd_sc_hd__o21ai_0 _13936_ (.A1(net4061),
    .A2(_04854_),
    .B1(_04856_),
    .Y(_04857_));
 sky130_fd_sc_hd__o21ai_2 _13937_ (.A1(_03725_),
    .A2(_04852_),
    .B1(_04857_),
    .Y(_04858_));
 sky130_fd_sc_hd__a21oi_1 _13938_ (.A1(_04538_),
    .A2(_04539_),
    .B1(_03704_),
    .Y(_04859_));
 sky130_fd_sc_hd__o21ai_0 _13939_ (.A1(_04472_),
    .A2(_04859_),
    .B1(_03735_),
    .Y(_04860_));
 sky130_fd_sc_hd__o22ai_1 _13940_ (.A1(net4090),
    .A2(_04450_),
    .B1(_04434_),
    .B2(_11864_[0]),
    .Y(_04861_));
 sky130_fd_sc_hd__nor2_1 _13941_ (.A(_11863_[0]),
    .B(_04568_),
    .Y(_04862_));
 sky130_fd_sc_hd__o21ai_0 _13942_ (.A1(_04861_),
    .A2(_04862_),
    .B1(net4061),
    .Y(_04863_));
 sky130_fd_sc_hd__a21oi_1 _13943_ (.A1(_04860_),
    .A2(_04863_),
    .B1(net4062),
    .Y(_04864_));
 sky130_fd_sc_hd__nor2_1 _13944_ (.A(_11874_[0]),
    .B(_04565_),
    .Y(_04865_));
 sky130_fd_sc_hd__a21oi_1 _13945_ (.A1(_03704_),
    .A2(_04759_),
    .B1(_04865_),
    .Y(_04866_));
 sky130_fd_sc_hd__o21ai_0 _13946_ (.A1(_11883_[0]),
    .A2(_04678_),
    .B1(_03715_),
    .Y(_04867_));
 sky130_fd_sc_hd__o2111ai_1 _13947_ (.A1(_03715_),
    .A2(_04832_),
    .B1(_04867_),
    .C1(net4062),
    .D1(_03734_),
    .Y(_04868_));
 sky130_fd_sc_hd__o31ai_1 _13948_ (.A1(_03725_),
    .A2(net4061),
    .A3(_04866_),
    .B1(_04868_),
    .Y(_04869_));
 sky130_fd_sc_hd__o21ai_2 _13949_ (.A1(_04864_),
    .A2(_04869_),
    .B1(_03750_),
    .Y(_04870_));
 sky130_fd_sc_hd__o21ai_4 _13950_ (.A1(_03750_),
    .A2(_04858_),
    .B1(_04870_),
    .Y(_04871_));
 sky130_fd_sc_hd__nor3_1 _13951_ (.A(net4087),
    .B(net4062),
    .C(_04470_),
    .Y(_04872_));
 sky130_fd_sc_hd__a21oi_1 _13952_ (.A1(_04440_),
    .A2(_04664_),
    .B1(_04872_),
    .Y(_04873_));
 sky130_fd_sc_hd__o21ai_0 _13953_ (.A1(_03725_),
    .A2(_04672_),
    .B1(_04565_),
    .Y(_04874_));
 sky130_fd_sc_hd__nand3_1 _13954_ (.A(_03696_),
    .B(_03715_),
    .C(net4062),
    .Y(_04875_));
 sky130_fd_sc_hd__o21ai_0 _13955_ (.A1(_03715_),
    .A2(net4062),
    .B1(_04875_),
    .Y(_04876_));
 sky130_fd_sc_hd__a22oi_1 _13956_ (.A1(net4089),
    .A2(_04874_),
    .B1(_04876_),
    .B2(net4090),
    .Y(_04877_));
 sky130_fd_sc_hd__o21ai_0 _13957_ (.A1(net4084),
    .A2(_03725_),
    .B1(_04450_),
    .Y(_04878_));
 sky130_fd_sc_hd__o21ai_0 _13958_ (.A1(net4062),
    .A2(_04463_),
    .B1(_04443_),
    .Y(_04879_));
 sky130_fd_sc_hd__a221oi_1 _13959_ (.A1(_11862_[0]),
    .A2(_04878_),
    .B1(_04879_),
    .B2(_03704_),
    .C1(_04664_),
    .Y(_04880_));
 sky130_fd_sc_hd__nor2_1 _13960_ (.A(_03735_),
    .B(_04880_),
    .Y(_04881_));
 sky130_fd_sc_hd__a31oi_1 _13961_ (.A1(_03735_),
    .A2(_04873_),
    .A3(_04877_),
    .B1(_04881_),
    .Y(_04882_));
 sky130_fd_sc_hd__a21oi_2 _13962_ (.A1(_11874_[0]),
    .A2(_03704_),
    .B1(_04622_),
    .Y(_04883_));
 sky130_fd_sc_hd__o211ai_1 _13963_ (.A1(_03715_),
    .A2(_04883_),
    .B1(_04732_),
    .C1(_03734_),
    .Y(_04884_));
 sky130_fd_sc_hd__o221ai_1 _13964_ (.A1(_11862_[0]),
    .A2(net4084),
    .B1(_04585_),
    .B2(_03704_),
    .C1(_03735_),
    .Y(_04885_));
 sky130_fd_sc_hd__a21oi_1 _13965_ (.A1(_04884_),
    .A2(_04885_),
    .B1(_03725_),
    .Y(_04886_));
 sky130_fd_sc_hd__a211oi_1 _13966_ (.A1(_11867_[0]),
    .A2(net4084),
    .B1(_04517_),
    .C1(_03702_),
    .Y(_04887_));
 sky130_fd_sc_hd__nor3_1 _13967_ (.A(_04545_),
    .B(_04650_),
    .C(_04887_),
    .Y(_04888_));
 sky130_fd_sc_hd__nor3_1 _13968_ (.A(_03704_),
    .B(_04427_),
    .C(_04501_),
    .Y(_04889_));
 sky130_fd_sc_hd__a2111oi_0 _13969_ (.A1(_11888_[0]),
    .A2(net4084),
    .B1(_04435_),
    .C1(_04599_),
    .D1(_04889_),
    .Y(_04890_));
 sky130_fd_sc_hd__nor4_1 _13970_ (.A(_03750_),
    .B(_04886_),
    .C(_04888_),
    .D(_04890_),
    .Y(_04891_));
 sky130_fd_sc_hd__a211oi_1 _13971_ (.A1(_03750_),
    .A2(_04882_),
    .B1(_04891_),
    .C1(_03744_),
    .Y(_04892_));
 sky130_fd_sc_hd__a21oi_4 _13972_ (.A1(_03744_),
    .A2(_04871_),
    .B1(_04892_),
    .Y(_00015_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1172 ();
 sky130_fd_sc_hd__nor2_4 _13982_ (.A(net4096),
    .B(_03639_),
    .Y(_04899_));
 sky130_fd_sc_hd__a21oi_1 _13983_ (.A1(_11912_[0]),
    .A2(_03639_),
    .B1(_04899_),
    .Y(_04900_));
 sky130_fd_sc_hd__o21a_1 _13984_ (.A1(_03648_),
    .A2(_04900_),
    .B1(_03656_),
    .X(_04901_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1170 ();
 sky130_fd_sc_hd__nand2_2 _13987_ (.A(_03631_),
    .B(_03639_),
    .Y(_04904_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1168 ();
 sky130_fd_sc_hd__nand2_1 _13990_ (.A(_11901_[0]),
    .B(net4093),
    .Y(_04907_));
 sky130_fd_sc_hd__a31oi_1 _13991_ (.A1(net4092),
    .A2(_04904_),
    .A3(_04907_),
    .B1(_03656_),
    .Y(_04908_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1166 ();
 sky130_fd_sc_hd__nor2_1 _13994_ (.A(_11898_[0]),
    .B(net4093),
    .Y(_04911_));
 sky130_fd_sc_hd__a32oi_1 _13995_ (.A1(_11896_[0]),
    .A2(_03639_),
    .A3(_04901_),
    .B1(_04908_),
    .B2(_04911_),
    .Y(_04912_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1165 ();
 sky130_fd_sc_hd__a21oi_1 _13997_ (.A1(net4065),
    .A2(net4093),
    .B1(net4092),
    .Y(_04914_));
 sky130_fd_sc_hd__o21bai_1 _13998_ (.A1(_04901_),
    .A2(_04908_),
    .B1_N(_04914_),
    .Y(_04915_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1164 ();
 sky130_fd_sc_hd__a21oi_1 _14000_ (.A1(_04912_),
    .A2(_04915_),
    .B1(_03667_),
    .Y(_04917_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1159 ();
 sky130_fd_sc_hd__nand2_8 _14006_ (.A(_03639_),
    .B(_03648_),
    .Y(_04923_));
 sky130_fd_sc_hd__nor2_1 _14007_ (.A(_11903_[0]),
    .B(_04923_),
    .Y(_04924_));
 sky130_fd_sc_hd__nand2_8 _14008_ (.A(_11901_[0]),
    .B(net4064),
    .Y(_04925_));
 sky130_fd_sc_hd__nand2_4 _14009_ (.A(_03625_),
    .B(net4092),
    .Y(_04926_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1158 ();
 sky130_fd_sc_hd__a21oi_1 _14011_ (.A1(_04925_),
    .A2(_04926_),
    .B1(_03639_),
    .Y(_04928_));
 sky130_fd_sc_hd__nor3_1 _14012_ (.A(_03658_),
    .B(_04924_),
    .C(_04928_),
    .Y(_04929_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1157 ();
 sky130_fd_sc_hd__nand2b_4 _14014_ (.A_N(_11901_[0]),
    .B(net4092),
    .Y(_04931_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1156 ();
 sky130_fd_sc_hd__nand2_1 _14016_ (.A(_11898_[0]),
    .B(_03648_),
    .Y(_04933_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1155 ();
 sky130_fd_sc_hd__nand2b_4 _14018_ (.A_N(_11897_[0]),
    .B(_03648_),
    .Y(_04935_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1154 ();
 sky130_fd_sc_hd__a21oi_1 _14020_ (.A1(_04926_),
    .A2(_04935_),
    .B1(net4093),
    .Y(_04937_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1153 ();
 sky130_fd_sc_hd__a311oi_1 _14022_ (.A1(net4093),
    .A2(_04931_),
    .A3(_04933_),
    .B1(_04937_),
    .C1(_03656_),
    .Y(_04939_));
 sky130_fd_sc_hd__nor3_1 _14023_ (.A(_03666_),
    .B(_04929_),
    .C(_04939_),
    .Y(_04940_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1152 ();
 sky130_fd_sc_hd__o21ai_0 _14025_ (.A1(_04917_),
    .A2(_04940_),
    .B1(net3628),
    .Y(_04942_));
 sky130_fd_sc_hd__nor2_4 _14026_ (.A(_03639_),
    .B(_03648_),
    .Y(_04943_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1150 ();
 sky130_fd_sc_hd__and2_0 _14029_ (.A(_11908_[0]),
    .B(_03639_),
    .X(_04946_));
 sky130_fd_sc_hd__o22ai_1 _14030_ (.A1(_11897_[0]),
    .A2(_04923_),
    .B1(_04946_),
    .B2(_03648_),
    .Y(_04947_));
 sky130_fd_sc_hd__nand2_1 _14031_ (.A(_11896_[0]),
    .B(_03639_),
    .Y(_04948_));
 sky130_fd_sc_hd__a21oi_2 _14032_ (.A1(_04948_),
    .A2(_04914_),
    .B1(_03658_),
    .Y(_04949_));
 sky130_fd_sc_hd__a21oi_1 _14033_ (.A1(_03658_),
    .A2(_04947_),
    .B1(_04949_),
    .Y(_04950_));
 sky130_fd_sc_hd__a21oi_1 _14034_ (.A1(_11903_[0]),
    .A2(_04943_),
    .B1(_04950_),
    .Y(_04951_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1148 ();
 sky130_fd_sc_hd__nand2b_4 _14037_ (.A_N(_11903_[0]),
    .B(_03648_),
    .Y(_04954_));
 sky130_fd_sc_hd__o21ai_0 _14038_ (.A1(_11912_[0]),
    .A2(_03648_),
    .B1(_04954_),
    .Y(_04955_));
 sky130_fd_sc_hd__a221oi_1 _14039_ (.A1(_11910_[0]),
    .A2(_04943_),
    .B1(_04955_),
    .B2(_03639_),
    .C1(net4091),
    .Y(_04956_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1146 ();
 sky130_fd_sc_hd__nand2b_4 _14042_ (.A_N(_11897_[0]),
    .B(net4092),
    .Y(_04959_));
 sky130_fd_sc_hd__o21ai_0 _14043_ (.A1(_11906_[0]),
    .A2(net4092),
    .B1(_04959_),
    .Y(_04960_));
 sky130_fd_sc_hd__nand2_8 _14044_ (.A(net4097),
    .B(_03648_),
    .Y(_04961_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1145 ();
 sky130_fd_sc_hd__nand2_4 _14046_ (.A(_03631_),
    .B(net4092),
    .Y(_04963_));
 sky130_fd_sc_hd__a21oi_1 _14047_ (.A1(_04961_),
    .A2(_04963_),
    .B1(net4093),
    .Y(_04964_));
 sky130_fd_sc_hd__a21oi_1 _14048_ (.A1(net4093),
    .A2(_04960_),
    .B1(_04964_),
    .Y(_04965_));
 sky130_fd_sc_hd__nor2_1 _14049_ (.A(_03658_),
    .B(_04965_),
    .Y(_04966_));
 sky130_fd_sc_hd__o21ai_0 _14050_ (.A1(_04956_),
    .A2(_04966_),
    .B1(_03667_),
    .Y(_04967_));
 sky130_fd_sc_hd__o211ai_1 _14051_ (.A1(_03667_),
    .A2(_04951_),
    .B1(_04967_),
    .C1(_03685_),
    .Y(_04968_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1144 ();
 sky130_fd_sc_hd__nor2_4 _14053_ (.A(_03639_),
    .B(net4092),
    .Y(_04970_));
 sky130_fd_sc_hd__nand2_4 _14054_ (.A(_11912_[0]),
    .B(net4092),
    .Y(_04971_));
 sky130_fd_sc_hd__o21ai_1 _14055_ (.A1(_11901_[0]),
    .A2(net4092),
    .B1(_04971_),
    .Y(_04972_));
 sky130_fd_sc_hd__a221oi_1 _14056_ (.A1(_11908_[0]),
    .A2(_04970_),
    .B1(_04972_),
    .B2(_03639_),
    .C1(_03666_),
    .Y(_04973_));
 sky130_fd_sc_hd__a21oi_2 _14057_ (.A1(_04961_),
    .A2(_04926_),
    .B1(_03639_),
    .Y(_04974_));
 sky130_fd_sc_hd__nand2b_4 _14058_ (.A_N(_11910_[0]),
    .B(_03648_),
    .Y(_04975_));
 sky130_fd_sc_hd__a21oi_1 _14059_ (.A1(_04975_),
    .A2(_04931_),
    .B1(net4093),
    .Y(_04976_));
 sky130_fd_sc_hd__nor3_1 _14060_ (.A(_03667_),
    .B(_04974_),
    .C(_04976_),
    .Y(_04977_));
 sky130_fd_sc_hd__nor3_1 _14061_ (.A(_03658_),
    .B(_04973_),
    .C(_04977_),
    .Y(_04978_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1143 ();
 sky130_fd_sc_hd__nand2_8 _14063_ (.A(net4093),
    .B(net4092),
    .Y(_04980_));
 sky130_fd_sc_hd__nor2_1 _14064_ (.A(_11906_[0]),
    .B(_04980_),
    .Y(_04981_));
 sky130_fd_sc_hd__nand2_1 _14065_ (.A(_11912_[0]),
    .B(_03648_),
    .Y(_04982_));
 sky130_fd_sc_hd__a21oi_1 _14066_ (.A1(_04931_),
    .A2(_04982_),
    .B1(net4093),
    .Y(_04983_));
 sky130_fd_sc_hd__nor3_1 _14067_ (.A(_03666_),
    .B(_04981_),
    .C(_04983_),
    .Y(_04984_));
 sky130_fd_sc_hd__a221oi_2 _14068_ (.A1(_11922_[0]),
    .A2(_03648_),
    .B1(_04943_),
    .B2(_11897_[0]),
    .C1(_03667_),
    .Y(_04985_));
 sky130_fd_sc_hd__nor3_1 _14069_ (.A(_03656_),
    .B(_04984_),
    .C(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__o21ai_0 _14070_ (.A1(_04978_),
    .A2(_04986_),
    .B1(_03685_),
    .Y(_04987_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1142 ();
 sky130_fd_sc_hd__nor2_2 _14072_ (.A(net4093),
    .B(_03648_),
    .Y(_04989_));
 sky130_fd_sc_hd__nor2_4 _14073_ (.A(_04970_),
    .B(_04989_),
    .Y(_04990_));
 sky130_fd_sc_hd__nor2_2 _14074_ (.A(_03637_),
    .B(net4092),
    .Y(_04991_));
 sky130_fd_sc_hd__nand2_1 _14075_ (.A(_11897_[0]),
    .B(_04991_),
    .Y(_04992_));
 sky130_fd_sc_hd__o221a_1 _14076_ (.A1(_11906_[0]),
    .A2(_04980_),
    .B1(_04990_),
    .B2(_11910_[0]),
    .C1(_04992_),
    .X(_04993_));
 sky130_fd_sc_hd__o211ai_1 _14077_ (.A1(_11896_[0]),
    .A2(_03648_),
    .B1(_04975_),
    .C1(net4093),
    .Y(_04994_));
 sky130_fd_sc_hd__nand2_8 _14078_ (.A(_11897_[0]),
    .B(net4092),
    .Y(_04995_));
 sky130_fd_sc_hd__o211ai_1 _14079_ (.A1(_11906_[0]),
    .A2(net4092),
    .B1(_04995_),
    .C1(_03639_),
    .Y(_04996_));
 sky130_fd_sc_hd__nand3_1 _14080_ (.A(_03667_),
    .B(_04994_),
    .C(_04996_),
    .Y(_04997_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1141 ();
 sky130_fd_sc_hd__o211ai_1 _14082_ (.A1(_03667_),
    .A2(_04993_),
    .B1(_04997_),
    .C1(_03656_),
    .Y(_04999_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1140 ();
 sky130_fd_sc_hd__nand2_8 _14084_ (.A(net4094),
    .B(net4092),
    .Y(_05001_));
 sky130_fd_sc_hd__nand2_8 _14085_ (.A(_03631_),
    .B(_03648_),
    .Y(_05002_));
 sky130_fd_sc_hd__a21oi_1 _14086_ (.A1(_05001_),
    .A2(_05002_),
    .B1(net4098),
    .Y(_05003_));
 sky130_fd_sc_hd__a21oi_1 _14087_ (.A1(net4098),
    .A2(_04990_),
    .B1(_05003_),
    .Y(_05004_));
 sky130_fd_sc_hd__o21ai_0 _14088_ (.A1(_03667_),
    .A2(_04935_),
    .B1(_05001_),
    .Y(_05005_));
 sky130_fd_sc_hd__nor3_1 _14089_ (.A(net4093),
    .B(_03667_),
    .C(_04995_),
    .Y(_05006_));
 sky130_fd_sc_hd__a21oi_1 _14090_ (.A1(net4093),
    .A2(_05005_),
    .B1(_05006_),
    .Y(_05007_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1139 ();
 sky130_fd_sc_hd__o211ai_1 _14092_ (.A1(_03666_),
    .A2(_05004_),
    .B1(_05007_),
    .C1(_03658_),
    .Y(_05009_));
 sky130_fd_sc_hd__nand3_1 _14093_ (.A(_03684_),
    .B(_04999_),
    .C(_05009_),
    .Y(_05010_));
 sky130_fd_sc_hd__a21oi_2 _14094_ (.A1(_04987_),
    .A2(_05010_),
    .B1(_03676_),
    .Y(_05011_));
 sky130_fd_sc_hd__a31o_4 _14095_ (.A1(_03676_),
    .A2(_04942_),
    .A3(_04968_),
    .B1(_05011_),
    .X(_00016_));
 sky130_fd_sc_hd__nor2_1 _14096_ (.A(net4098),
    .B(_04923_),
    .Y(_05012_));
 sky130_fd_sc_hd__nor2_2 _14097_ (.A(_11897_[0]),
    .B(_04980_),
    .Y(_05013_));
 sky130_fd_sc_hd__nand2_2 _14098_ (.A(_03639_),
    .B(net4092),
    .Y(_05014_));
 sky130_fd_sc_hd__nand2_8 _14099_ (.A(net4094),
    .B(_03648_),
    .Y(_05015_));
 sky130_fd_sc_hd__a21oi_1 _14100_ (.A1(_05014_),
    .A2(_05015_),
    .B1(net4065),
    .Y(_05016_));
 sky130_fd_sc_hd__nor4_1 _14101_ (.A(_03667_),
    .B(_05012_),
    .C(_05013_),
    .D(_05016_),
    .Y(_05017_));
 sky130_fd_sc_hd__nand2_4 _14102_ (.A(_03637_),
    .B(net4064),
    .Y(_05018_));
 sky130_fd_sc_hd__nor2_1 _14103_ (.A(_11896_[0]),
    .B(_05018_),
    .Y(_05019_));
 sky130_fd_sc_hd__nand2_4 _14104_ (.A(_11903_[0]),
    .B(net4092),
    .Y(_05020_));
 sky130_fd_sc_hd__a21oi_1 _14105_ (.A1(_04935_),
    .A2(_05020_),
    .B1(net4093),
    .Y(_05021_));
 sky130_fd_sc_hd__nor3_1 _14106_ (.A(_03666_),
    .B(_05019_),
    .C(_05021_),
    .Y(_05022_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1138 ();
 sky130_fd_sc_hd__o21ai_2 _14108_ (.A1(_05017_),
    .A2(_05022_),
    .B1(net4091),
    .Y(_05024_));
 sky130_fd_sc_hd__nand2_4 _14109_ (.A(_11896_[0]),
    .B(net4092),
    .Y(_05025_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1137 ();
 sky130_fd_sc_hd__a32oi_1 _14111_ (.A1(_03639_),
    .A2(_05002_),
    .A3(_05025_),
    .B1(_04970_),
    .B2(_11898_[0]),
    .Y(_05027_));
 sky130_fd_sc_hd__nand3_1 _14112_ (.A(_03658_),
    .B(_03667_),
    .C(_05027_),
    .Y(_05028_));
 sky130_fd_sc_hd__a21oi_1 _14113_ (.A1(_11903_[0]),
    .A2(_04970_),
    .B1(_03667_),
    .Y(_05029_));
 sky130_fd_sc_hd__a21oi_4 _14114_ (.A1(net4099),
    .A2(_04943_),
    .B1(_03656_),
    .Y(_05030_));
 sky130_fd_sc_hd__nor2_2 _14115_ (.A(_11897_[0]),
    .B(net4092),
    .Y(_05031_));
 sky130_fd_sc_hd__nor2_2 _14116_ (.A(_11910_[0]),
    .B(_03648_),
    .Y(_05032_));
 sky130_fd_sc_hd__o21ai_2 _14117_ (.A1(_05031_),
    .A2(_05032_),
    .B1(_03639_),
    .Y(_05033_));
 sky130_fd_sc_hd__a31oi_1 _14118_ (.A1(_05029_),
    .A2(_05030_),
    .A3(_05033_),
    .B1(net3628),
    .Y(_05034_));
 sky130_fd_sc_hd__nand3_1 _14119_ (.A(_05024_),
    .B(_05028_),
    .C(_05034_),
    .Y(_05035_));
 sky130_fd_sc_hd__nand2_1 _14120_ (.A(net4065),
    .B(_04943_),
    .Y(_05036_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1136 ();
 sky130_fd_sc_hd__nand2_1 _14122_ (.A(_04935_),
    .B(_05025_),
    .Y(_05038_));
 sky130_fd_sc_hd__nand2_1 _14123_ (.A(_03639_),
    .B(_05038_),
    .Y(_05039_));
 sky130_fd_sc_hd__nand2b_4 _14124_ (.A_N(_11910_[0]),
    .B(net4092),
    .Y(_05040_));
 sky130_fd_sc_hd__nand2_8 _14125_ (.A(net4098),
    .B(net4092),
    .Y(_05041_));
 sky130_fd_sc_hd__a21oi_1 _14126_ (.A1(_05041_),
    .A2(_04954_),
    .B1(net4093),
    .Y(_05042_));
 sky130_fd_sc_hd__a311oi_1 _14127_ (.A1(net4093),
    .A2(_05040_),
    .A3(_05015_),
    .B1(_05042_),
    .C1(_03666_),
    .Y(_05043_));
 sky130_fd_sc_hd__a31oi_1 _14128_ (.A1(_03666_),
    .A2(_05036_),
    .A3(_05039_),
    .B1(_05043_),
    .Y(_05044_));
 sky130_fd_sc_hd__o21ai_0 _14129_ (.A1(_11896_[0]),
    .A2(net4092),
    .B1(_04971_),
    .Y(_05045_));
 sky130_fd_sc_hd__nand2_4 _14130_ (.A(_11898_[0]),
    .B(net4092),
    .Y(_05046_));
 sky130_fd_sc_hd__a21oi_1 _14131_ (.A1(_04935_),
    .A2(_05046_),
    .B1(net4093),
    .Y(_05047_));
 sky130_fd_sc_hd__a2111oi_0 _14132_ (.A1(net4093),
    .A2(_05045_),
    .B1(_05047_),
    .C1(net4091),
    .D1(_03667_),
    .Y(_05048_));
 sky130_fd_sc_hd__a21oi_1 _14133_ (.A1(net4091),
    .A2(_05044_),
    .B1(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__a21oi_1 _14134_ (.A1(_04971_),
    .A2(_04975_),
    .B1(net4093),
    .Y(_05050_));
 sky130_fd_sc_hd__nand2_1 _14135_ (.A(_11897_[0]),
    .B(_04970_),
    .Y(_05051_));
 sky130_fd_sc_hd__nand4b_1 _14136_ (.A_N(_05050_),
    .B(_05030_),
    .C(_03667_),
    .D(_05051_),
    .Y(_05052_));
 sky130_fd_sc_hd__nand3_1 _14137_ (.A(net3628),
    .B(_05049_),
    .C(_05052_),
    .Y(_05053_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1135 ();
 sky130_fd_sc_hd__a21boi_0 _14139_ (.A1(_11906_[0]),
    .A2(net4093),
    .B1_N(_04948_),
    .Y(_05055_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1134 ();
 sky130_fd_sc_hd__nor3_1 _14141_ (.A(_11924_[0]),
    .B(net4092),
    .C(_03667_),
    .Y(_05057_));
 sky130_fd_sc_hd__a21oi_1 _14142_ (.A1(net4092),
    .A2(_05055_),
    .B1(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__nor2_1 _14143_ (.A(_11901_[0]),
    .B(net4092),
    .Y(_05059_));
 sky130_fd_sc_hd__nor3_1 _14144_ (.A(_03639_),
    .B(_05059_),
    .C(_05032_),
    .Y(_05060_));
 sky130_fd_sc_hd__nand2_2 _14145_ (.A(_11896_[0]),
    .B(_03648_),
    .Y(_05061_));
 sky130_fd_sc_hd__a21oi_1 _14146_ (.A1(_04926_),
    .A2(_05061_),
    .B1(net4093),
    .Y(_05062_));
 sky130_fd_sc_hd__o21ai_0 _14147_ (.A1(_05060_),
    .A2(_05062_),
    .B1(_03667_),
    .Y(_05063_));
 sky130_fd_sc_hd__a21oi_1 _14148_ (.A1(_05001_),
    .A2(_05002_),
    .B1(_03639_),
    .Y(_05064_));
 sky130_fd_sc_hd__o21ai_0 _14149_ (.A1(_05042_),
    .A2(_05064_),
    .B1(_03666_),
    .Y(_05065_));
 sky130_fd_sc_hd__nand3_1 _14150_ (.A(_03658_),
    .B(_05063_),
    .C(_05065_),
    .Y(_05066_));
 sky130_fd_sc_hd__o21ai_0 _14151_ (.A1(_03658_),
    .A2(_05058_),
    .B1(_05066_),
    .Y(_05067_));
 sky130_fd_sc_hd__nor2_1 _14152_ (.A(net4094),
    .B(_03637_),
    .Y(_05068_));
 sky130_fd_sc_hd__and2_4 _14153_ (.A(_11903_[0]),
    .B(_03637_),
    .X(_05069_));
 sky130_fd_sc_hd__nand2_1 _14154_ (.A(_11915_[0]),
    .B(_03648_),
    .Y(_05070_));
 sky130_fd_sc_hd__o31ai_1 _14155_ (.A1(net4064),
    .A2(_05068_),
    .A3(_05069_),
    .B1(_05070_),
    .Y(_05071_));
 sky130_fd_sc_hd__nand2_1 _14156_ (.A(_03666_),
    .B(_05071_),
    .Y(_05072_));
 sky130_fd_sc_hd__nand2_4 _14157_ (.A(_11897_[0]),
    .B(_03648_),
    .Y(_05073_));
 sky130_fd_sc_hd__a21oi_1 _14158_ (.A1(_05073_),
    .A2(_05020_),
    .B1(_03637_),
    .Y(_05074_));
 sky130_fd_sc_hd__or3_4 _14159_ (.A(_03666_),
    .B(_04974_),
    .C(_05074_),
    .X(_05075_));
 sky130_fd_sc_hd__a21oi_1 _14160_ (.A1(_05072_),
    .A2(_05075_),
    .B1(_03656_),
    .Y(_05076_));
 sky130_fd_sc_hd__and2_4 _14161_ (.A(_11901_[0]),
    .B(_03639_),
    .X(_05077_));
 sky130_fd_sc_hd__o21ai_1 _14162_ (.A1(_11903_[0]),
    .A2(_03639_),
    .B1(net4092),
    .Y(_05078_));
 sky130_fd_sc_hd__o21ai_1 _14163_ (.A1(_05077_),
    .A2(_05078_),
    .B1(_03656_),
    .Y(_05079_));
 sky130_fd_sc_hd__nand2_1 _14164_ (.A(_11897_[0]),
    .B(net4093),
    .Y(_05080_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1133 ();
 sky130_fd_sc_hd__nand2_1 _14166_ (.A(_11898_[0]),
    .B(_03639_),
    .Y(_05082_));
 sky130_fd_sc_hd__a21oi_1 _14167_ (.A1(_05080_),
    .A2(_05082_),
    .B1(net4092),
    .Y(_05083_));
 sky130_fd_sc_hd__nor3_1 _14168_ (.A(_03667_),
    .B(_05079_),
    .C(_05083_),
    .Y(_05084_));
 sky130_fd_sc_hd__o211ai_1 _14169_ (.A1(net4094),
    .A2(_05041_),
    .B1(_03667_),
    .C1(_03656_),
    .Y(_05085_));
 sky130_fd_sc_hd__a31oi_1 _14170_ (.A1(_03637_),
    .A2(_04925_),
    .A3(_04963_),
    .B1(_05085_),
    .Y(_05086_));
 sky130_fd_sc_hd__nor4_2 _14171_ (.A(_03684_),
    .B(_05076_),
    .C(_05084_),
    .D(_05086_),
    .Y(_05087_));
 sky130_fd_sc_hd__a211oi_1 _14172_ (.A1(net3628),
    .A2(_05067_),
    .B1(_05087_),
    .C1(_03676_),
    .Y(_05088_));
 sky130_fd_sc_hd__a31oi_1 _14173_ (.A1(_03676_),
    .A2(_05035_),
    .A3(_05053_),
    .B1(_05088_),
    .Y(_00017_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1132 ();
 sky130_fd_sc_hd__nor2_1 _14175_ (.A(net4094),
    .B(_03648_),
    .Y(_05090_));
 sky130_fd_sc_hd__a21oi_1 _14176_ (.A1(_11912_[0]),
    .A2(_03648_),
    .B1(_05090_),
    .Y(_05091_));
 sky130_fd_sc_hd__a21o_1 _14177_ (.A1(_04961_),
    .A2(_04995_),
    .B1(net4093),
    .X(_05092_));
 sky130_fd_sc_hd__o21ai_0 _14178_ (.A1(_03639_),
    .A2(_05091_),
    .B1(_05092_),
    .Y(_05093_));
 sky130_fd_sc_hd__nor2_2 _14179_ (.A(net4098),
    .B(_03648_),
    .Y(_05094_));
 sky130_fd_sc_hd__nor2_1 _14180_ (.A(_11908_[0]),
    .B(net4092),
    .Y(_05095_));
 sky130_fd_sc_hd__nand2b_4 _14181_ (.A_N(_11898_[0]),
    .B(net4092),
    .Y(_05096_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1131 ();
 sky130_fd_sc_hd__nand3_1 _14183_ (.A(net4093),
    .B(_05015_),
    .C(_05096_),
    .Y(_05098_));
 sky130_fd_sc_hd__o311ai_0 _14184_ (.A1(net4093),
    .A2(_05094_),
    .A3(_05095_),
    .B1(_05098_),
    .C1(_03676_),
    .Y(_05099_));
 sky130_fd_sc_hd__o21ai_0 _14185_ (.A1(_03676_),
    .A2(_05093_),
    .B1(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__nor2_4 _14186_ (.A(_11908_[0]),
    .B(net4064),
    .Y(_05101_));
 sky130_fd_sc_hd__nand3b_1 _14187_ (.A_N(_05101_),
    .B(net4093),
    .C(_05073_),
    .Y(_05102_));
 sky130_fd_sc_hd__o311ai_0 _14188_ (.A1(net4093),
    .A2(_05094_),
    .A3(_05031_),
    .B1(_05102_),
    .C1(_03676_),
    .Y(_05103_));
 sky130_fd_sc_hd__nor2_1 _14189_ (.A(_11898_[0]),
    .B(_04923_),
    .Y(_05104_));
 sky130_fd_sc_hd__nand2_1 _14190_ (.A(_11901_[0]),
    .B(net4092),
    .Y(_05105_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1130 ();
 sky130_fd_sc_hd__a21oi_1 _14192_ (.A1(_05105_),
    .A2(_05061_),
    .B1(_03639_),
    .Y(_05107_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1129 ();
 sky130_fd_sc_hd__o21ai_0 _14194_ (.A1(_05104_),
    .A2(_05107_),
    .B1(_03675_),
    .Y(_05109_));
 sky130_fd_sc_hd__nand3_1 _14195_ (.A(net4091),
    .B(_05103_),
    .C(_05109_),
    .Y(_05110_));
 sky130_fd_sc_hd__o21ai_1 _14196_ (.A1(net4091),
    .A2(_05100_),
    .B1(_05110_),
    .Y(_05111_));
 sky130_fd_sc_hd__nor2_1 _14197_ (.A(_11896_[0]),
    .B(_04990_),
    .Y(_05112_));
 sky130_fd_sc_hd__nor4_1 _14198_ (.A(_03676_),
    .B(_04981_),
    .C(_05012_),
    .D(_05112_),
    .Y(_05113_));
 sky130_fd_sc_hd__a2111oi_0 _14199_ (.A1(_11917_[0]),
    .A2(_03648_),
    .B1(_03675_),
    .C1(_04964_),
    .D1(_05013_),
    .Y(_05114_));
 sky130_fd_sc_hd__nor2_1 _14200_ (.A(_11897_[0]),
    .B(_03639_),
    .Y(_05115_));
 sky130_fd_sc_hd__nand2_1 _14201_ (.A(_11922_[0]),
    .B(net4092),
    .Y(_05116_));
 sky130_fd_sc_hd__o311ai_0 _14202_ (.A1(net4092),
    .A2(_05077_),
    .A3(_05115_),
    .B1(_05116_),
    .C1(_03676_),
    .Y(_05117_));
 sky130_fd_sc_hd__nand2_2 _14203_ (.A(_05073_),
    .B(_05040_),
    .Y(_05118_));
 sky130_fd_sc_hd__a221o_1 _14204_ (.A1(_11903_[0]),
    .A2(_04970_),
    .B1(_05118_),
    .B2(_03639_),
    .C1(_03676_),
    .X(_05119_));
 sky130_fd_sc_hd__nand3_1 _14205_ (.A(_03656_),
    .B(_05117_),
    .C(_05119_),
    .Y(_05120_));
 sky130_fd_sc_hd__o311ai_0 _14206_ (.A1(_03656_),
    .A2(_05113_),
    .A3(_05114_),
    .B1(_03685_),
    .C1(_05120_),
    .Y(_05121_));
 sky130_fd_sc_hd__o21ai_2 _14207_ (.A1(_03685_),
    .A2(_05111_),
    .B1(_05121_),
    .Y(_05122_));
 sky130_fd_sc_hd__o211ai_1 _14208_ (.A1(_11901_[0]),
    .A2(_03639_),
    .B1(_03648_),
    .C1(_04904_),
    .Y(_05123_));
 sky130_fd_sc_hd__o211ai_1 _14209_ (.A1(_11917_[0]),
    .A2(_03648_),
    .B1(_03675_),
    .C1(_05123_),
    .Y(_05124_));
 sky130_fd_sc_hd__o211ai_1 _14210_ (.A1(_11906_[0]),
    .A2(net4092),
    .B1(_05001_),
    .C1(_03639_),
    .Y(_05125_));
 sky130_fd_sc_hd__o211ai_1 _14211_ (.A1(_03639_),
    .A2(_05118_),
    .B1(_05125_),
    .C1(_03676_),
    .Y(_05126_));
 sky130_fd_sc_hd__nand2_1 _14212_ (.A(_11924_[0]),
    .B(net4092),
    .Y(_05127_));
 sky130_fd_sc_hd__nand2_1 _14213_ (.A(net4099),
    .B(_03631_),
    .Y(_05128_));
 sky130_fd_sc_hd__o211ai_1 _14214_ (.A1(_03631_),
    .A2(_03639_),
    .B1(_03648_),
    .C1(_05128_),
    .Y(_05129_));
 sky130_fd_sc_hd__a221oi_1 _14215_ (.A1(_11920_[0]),
    .A2(_03648_),
    .B1(_04943_),
    .B2(_11901_[0]),
    .C1(_03676_),
    .Y(_05130_));
 sky130_fd_sc_hd__a311oi_1 _14216_ (.A1(_03676_),
    .A2(_05127_),
    .A3(_05129_),
    .B1(_05130_),
    .C1(_03658_),
    .Y(_05131_));
 sky130_fd_sc_hd__a311oi_1 _14217_ (.A1(_03658_),
    .A2(_05124_),
    .A3(_05126_),
    .B1(net3628),
    .C1(_05131_),
    .Y(_05132_));
 sky130_fd_sc_hd__nand3_1 _14218_ (.A(_03637_),
    .B(_04954_),
    .C(_04959_),
    .Y(_05133_));
 sky130_fd_sc_hd__nand3_1 _14219_ (.A(_03639_),
    .B(_04925_),
    .C(_04963_),
    .Y(_05134_));
 sky130_fd_sc_hd__nor2_1 _14220_ (.A(_03637_),
    .B(_05101_),
    .Y(_05135_));
 sky130_fd_sc_hd__a211oi_1 _14221_ (.A1(_05002_),
    .A2(_05135_),
    .B1(_05069_),
    .C1(_03675_),
    .Y(_05136_));
 sky130_fd_sc_hd__a311o_1 _14222_ (.A1(_03675_),
    .A2(_05133_),
    .A3(_05134_),
    .B1(_05136_),
    .C1(_03658_),
    .X(_05137_));
 sky130_fd_sc_hd__nor2_4 _14223_ (.A(net4098),
    .B(net4092),
    .Y(_05138_));
 sky130_fd_sc_hd__nand3_1 _14224_ (.A(_03637_),
    .B(_04954_),
    .C(_05096_),
    .Y(_05139_));
 sky130_fd_sc_hd__o311ai_0 _14225_ (.A1(_03637_),
    .A2(_05138_),
    .A3(_05101_),
    .B1(_05139_),
    .C1(_03676_),
    .Y(_05140_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1128 ();
 sky130_fd_sc_hd__nand3_1 _14227_ (.A(_03637_),
    .B(_04925_),
    .C(_05096_),
    .Y(_05142_));
 sky130_fd_sc_hd__o211ai_1 _14228_ (.A1(_11903_[0]),
    .A2(_03648_),
    .B1(_05015_),
    .C1(_03639_),
    .Y(_05143_));
 sky130_fd_sc_hd__nand3_1 _14229_ (.A(_03675_),
    .B(_05142_),
    .C(_05143_),
    .Y(_05144_));
 sky130_fd_sc_hd__nand3_1 _14230_ (.A(_03658_),
    .B(_05140_),
    .C(_05144_),
    .Y(_05145_));
 sky130_fd_sc_hd__a21oi_1 _14231_ (.A1(_05137_),
    .A2(_05145_),
    .B1(_03685_),
    .Y(_05146_));
 sky130_fd_sc_hd__o21ai_1 _14232_ (.A1(_05132_),
    .A2(_05146_),
    .B1(_03666_),
    .Y(_05147_));
 sky130_fd_sc_hd__o21ai_4 _14233_ (.A1(_03666_),
    .A2(_05122_),
    .B1(_05147_),
    .Y(_00018_));
 sky130_fd_sc_hd__nand2_8 _14234_ (.A(_11908_[0]),
    .B(net4064),
    .Y(_05148_));
 sky130_fd_sc_hd__nand3_1 _14235_ (.A(_03667_),
    .B(_04995_),
    .C(_05148_),
    .Y(_05149_));
 sky130_fd_sc_hd__o211ai_1 _14236_ (.A1(_03667_),
    .A2(_04926_),
    .B1(_05149_),
    .C1(_03639_),
    .Y(_05150_));
 sky130_fd_sc_hd__o211ai_1 _14237_ (.A1(_03666_),
    .A2(_04961_),
    .B1(_05096_),
    .C1(_03637_),
    .Y(_05151_));
 sky130_fd_sc_hd__a21oi_1 _14238_ (.A1(_05150_),
    .A2(_05151_),
    .B1(_03656_),
    .Y(_05152_));
 sky130_fd_sc_hd__nand2b_4 _14239_ (.A_N(_11906_[0]),
    .B(net4092),
    .Y(_05153_));
 sky130_fd_sc_hd__a21oi_1 _14240_ (.A1(_04961_),
    .A2(_05025_),
    .B1(_03637_),
    .Y(_05154_));
 sky130_fd_sc_hd__a31oi_1 _14241_ (.A1(_03637_),
    .A2(_05153_),
    .A3(_05148_),
    .B1(_05154_),
    .Y(_05155_));
 sky130_fd_sc_hd__nor2_1 _14242_ (.A(_03667_),
    .B(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__o22ai_1 _14243_ (.A1(_03631_),
    .A2(_04980_),
    .B1(_04923_),
    .B2(_11910_[0]),
    .Y(_05157_));
 sky130_fd_sc_hd__a21oi_1 _14244_ (.A1(_03639_),
    .A2(_04963_),
    .B1(_03625_),
    .Y(_05158_));
 sky130_fd_sc_hd__nor3_1 _14245_ (.A(_03666_),
    .B(_05157_),
    .C(_05158_),
    .Y(_05159_));
 sky130_fd_sc_hd__nor3_1 _14246_ (.A(_03658_),
    .B(_05156_),
    .C(_05159_),
    .Y(_05160_));
 sky130_fd_sc_hd__o21ai_2 _14247_ (.A1(_05152_),
    .A2(_05160_),
    .B1(_03684_),
    .Y(_05161_));
 sky130_fd_sc_hd__nor2_2 _14248_ (.A(net4098),
    .B(_05002_),
    .Y(_05162_));
 sky130_fd_sc_hd__a21oi_1 _14249_ (.A1(_11906_[0]),
    .A2(_04943_),
    .B1(_05162_),
    .Y(_05163_));
 sky130_fd_sc_hd__nand3_1 _14250_ (.A(_03667_),
    .B(_05092_),
    .C(_05163_),
    .Y(_05164_));
 sky130_fd_sc_hd__nand3_1 _14251_ (.A(_03639_),
    .B(_04959_),
    .C(_05015_),
    .Y(_05165_));
 sky130_fd_sc_hd__nor2_1 _14252_ (.A(_11898_[0]),
    .B(net4092),
    .Y(_05166_));
 sky130_fd_sc_hd__o21ai_0 _14253_ (.A1(_05101_),
    .A2(_05166_),
    .B1(net4093),
    .Y(_05167_));
 sky130_fd_sc_hd__nand3_1 _14254_ (.A(_03666_),
    .B(_05165_),
    .C(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__a21oi_1 _14255_ (.A1(_05164_),
    .A2(_05168_),
    .B1(_03656_),
    .Y(_05169_));
 sky130_fd_sc_hd__nand2_1 _14256_ (.A(_11901_[0]),
    .B(_04970_),
    .Y(_05170_));
 sky130_fd_sc_hd__nor2_4 _14257_ (.A(net4065),
    .B(net4093),
    .Y(_05171_));
 sky130_fd_sc_hd__nor2_1 _14258_ (.A(net4098),
    .B(_03631_),
    .Y(_05172_));
 sky130_fd_sc_hd__o21ai_0 _14259_ (.A1(_05171_),
    .A2(_05172_),
    .B1(net4092),
    .Y(_05173_));
 sky130_fd_sc_hd__nand3_1 _14260_ (.A(_03637_),
    .B(_04925_),
    .C(_04959_),
    .Y(_05174_));
 sky130_fd_sc_hd__nand2_4 _14261_ (.A(_11906_[0]),
    .B(_03648_),
    .Y(_05175_));
 sky130_fd_sc_hd__nand3_1 _14262_ (.A(_03639_),
    .B(_05025_),
    .C(_05175_),
    .Y(_05176_));
 sky130_fd_sc_hd__a21oi_1 _14263_ (.A1(_05174_),
    .A2(_05176_),
    .B1(_03666_),
    .Y(_05177_));
 sky130_fd_sc_hd__a31oi_1 _14264_ (.A1(_03666_),
    .A2(_05170_),
    .A3(_05173_),
    .B1(_05177_),
    .Y(_05178_));
 sky130_fd_sc_hd__nor2_1 _14265_ (.A(_03658_),
    .B(_05178_),
    .Y(_05179_));
 sky130_fd_sc_hd__o21ai_2 _14266_ (.A1(_05169_),
    .A2(_05179_),
    .B1(_03685_),
    .Y(_05180_));
 sky130_fd_sc_hd__o21ai_0 _14267_ (.A1(_03666_),
    .A2(_04959_),
    .B1(_04982_),
    .Y(_05181_));
 sky130_fd_sc_hd__a21oi_1 _14268_ (.A1(_03639_),
    .A2(_05181_),
    .B1(_03656_),
    .Y(_05182_));
 sky130_fd_sc_hd__a21oi_1 _14269_ (.A1(_04935_),
    .A2(_05153_),
    .B1(_03639_),
    .Y(_05183_));
 sky130_fd_sc_hd__a21oi_1 _14270_ (.A1(_03631_),
    .A2(_04989_),
    .B1(_05183_),
    .Y(_05184_));
 sky130_fd_sc_hd__a21oi_1 _14271_ (.A1(_05182_),
    .A2(_05184_),
    .B1(_03667_),
    .Y(_05185_));
 sky130_fd_sc_hd__o2111ai_1 _14272_ (.A1(net4098),
    .A2(_03666_),
    .B1(_04961_),
    .C1(_04959_),
    .D1(_03639_),
    .Y(_05186_));
 sky130_fd_sc_hd__nand2_1 _14273_ (.A(net4098),
    .B(_04989_),
    .Y(_05187_));
 sky130_fd_sc_hd__nand2_1 _14274_ (.A(_11908_[0]),
    .B(_04990_),
    .Y(_05188_));
 sky130_fd_sc_hd__a41oi_1 _14275_ (.A1(_03656_),
    .A2(_05186_),
    .A3(_05187_),
    .A4(_05188_),
    .B1(_05182_),
    .Y(_05189_));
 sky130_fd_sc_hd__nor3_1 _14276_ (.A(_05094_),
    .B(_05166_),
    .C(_05171_),
    .Y(_05190_));
 sky130_fd_sc_hd__nor2_1 _14277_ (.A(_03667_),
    .B(_05190_),
    .Y(_05191_));
 sky130_fd_sc_hd__a31oi_1 _14278_ (.A1(_03656_),
    .A2(_05186_),
    .A3(_05191_),
    .B1(_03685_),
    .Y(_05192_));
 sky130_fd_sc_hd__o21ai_2 _14279_ (.A1(_05185_),
    .A2(_05189_),
    .B1(_05192_),
    .Y(_05193_));
 sky130_fd_sc_hd__a211oi_1 _14280_ (.A1(_11897_[0]),
    .A2(net4092),
    .B1(_05166_),
    .C1(net4093),
    .Y(_05194_));
 sky130_fd_sc_hd__a31oi_1 _14281_ (.A1(net4093),
    .A2(_04954_),
    .A3(_04963_),
    .B1(_05194_),
    .Y(_05195_));
 sky130_fd_sc_hd__o21ai_0 _14282_ (.A1(net4094),
    .A2(_04926_),
    .B1(_04992_),
    .Y(_05196_));
 sky130_fd_sc_hd__a21oi_1 _14283_ (.A1(_05041_),
    .A2(_05015_),
    .B1(_03639_),
    .Y(_05197_));
 sky130_fd_sc_hd__nor4_1 _14284_ (.A(_03658_),
    .B(_03667_),
    .C(_05196_),
    .D(_05197_),
    .Y(_05198_));
 sky130_fd_sc_hd__a31oi_1 _14285_ (.A1(_03656_),
    .A2(_03667_),
    .A3(_05195_),
    .B1(_05198_),
    .Y(_05199_));
 sky130_fd_sc_hd__o32ai_2 _14286_ (.A1(_11917_[0]),
    .A2(_03648_),
    .A3(_05171_),
    .B1(_05018_),
    .B2(_11897_[0]),
    .Y(_05200_));
 sky130_fd_sc_hd__a21oi_1 _14287_ (.A1(_05041_),
    .A2(_04935_),
    .B1(_03639_),
    .Y(_05201_));
 sky130_fd_sc_hd__a21oi_1 _14288_ (.A1(_04975_),
    .A2(_05153_),
    .B1(net4093),
    .Y(_05202_));
 sky130_fd_sc_hd__o21ai_0 _14289_ (.A1(_05201_),
    .A2(_05202_),
    .B1(_03667_),
    .Y(_05203_));
 sky130_fd_sc_hd__o211ai_1 _14290_ (.A1(_03667_),
    .A2(_05200_),
    .B1(_05203_),
    .C1(_03658_),
    .Y(_05204_));
 sky130_fd_sc_hd__a31oi_1 _14291_ (.A1(_03685_),
    .A2(_05199_),
    .A3(_05204_),
    .B1(_03676_),
    .Y(_05205_));
 sky130_fd_sc_hd__a32oi_4 _14292_ (.A1(_03676_),
    .A2(_05161_),
    .A3(_05180_),
    .B1(_05193_),
    .B2(_05205_),
    .Y(_00019_));
 sky130_fd_sc_hd__o22ai_1 _14293_ (.A1(net4093),
    .A2(_05094_),
    .B1(_04980_),
    .B2(_11898_[0]),
    .Y(_05206_));
 sky130_fd_sc_hd__nor2_1 _14294_ (.A(_03658_),
    .B(_05206_),
    .Y(_05207_));
 sky130_fd_sc_hd__a211oi_1 _14295_ (.A1(_11903_[0]),
    .A2(_03648_),
    .B1(_05032_),
    .C1(net4093),
    .Y(_05208_));
 sky130_fd_sc_hd__nor3_1 _14296_ (.A(net4091),
    .B(_05064_),
    .C(_05208_),
    .Y(_05209_));
 sky130_fd_sc_hd__o21ai_1 _14297_ (.A1(_05207_),
    .A2(_05209_),
    .B1(_03666_),
    .Y(_05210_));
 sky130_fd_sc_hd__a21oi_1 _14298_ (.A1(_11903_[0]),
    .A2(_03639_),
    .B1(_05115_),
    .Y(_05211_));
 sky130_fd_sc_hd__o21ai_1 _14299_ (.A1(_03648_),
    .A2(_05211_),
    .B1(_04949_),
    .Y(_05212_));
 sky130_fd_sc_hd__o311ai_0 _14300_ (.A1(_03639_),
    .A2(net4091),
    .A3(_05045_),
    .B1(_05212_),
    .C1(_03667_),
    .Y(_05213_));
 sky130_fd_sc_hd__nor2_1 _14301_ (.A(_11910_[0]),
    .B(_04980_),
    .Y(_05214_));
 sky130_fd_sc_hd__a21oi_1 _14302_ (.A1(_04971_),
    .A2(_04961_),
    .B1(net4093),
    .Y(_05215_));
 sky130_fd_sc_hd__nor4_1 _14303_ (.A(_03667_),
    .B(_05162_),
    .C(_05214_),
    .D(_05215_),
    .Y(_05216_));
 sky130_fd_sc_hd__a21oi_1 _14304_ (.A1(_05025_),
    .A2(_05051_),
    .B1(_03666_),
    .Y(_05217_));
 sky130_fd_sc_hd__o21ai_0 _14305_ (.A1(_05216_),
    .A2(_05217_),
    .B1(net4091),
    .Y(_05218_));
 sky130_fd_sc_hd__a21oi_1 _14306_ (.A1(_03639_),
    .A2(_05001_),
    .B1(net4099),
    .Y(_05219_));
 sky130_fd_sc_hd__nand2_1 _14307_ (.A(_03666_),
    .B(_04961_),
    .Y(_05220_));
 sky130_fd_sc_hd__a211oi_1 _14308_ (.A1(_04931_),
    .A2(_05015_),
    .B1(net4093),
    .C1(_03666_),
    .Y(_05221_));
 sky130_fd_sc_hd__a21oi_1 _14309_ (.A1(_11908_[0]),
    .A2(_04970_),
    .B1(_05221_),
    .Y(_05222_));
 sky130_fd_sc_hd__o311ai_0 _14310_ (.A1(_04899_),
    .A2(_05219_),
    .A3(_05220_),
    .B1(_05222_),
    .C1(_03658_),
    .Y(_05223_));
 sky130_fd_sc_hd__a21oi_1 _14311_ (.A1(_05218_),
    .A2(_05223_),
    .B1(_03676_),
    .Y(_05224_));
 sky130_fd_sc_hd__a31o_4 _14312_ (.A1(_03676_),
    .A2(_05210_),
    .A3(_05213_),
    .B1(_05224_),
    .X(_05225_));
 sky130_fd_sc_hd__nand2_1 _14313_ (.A(_11926_[0]),
    .B(_03648_),
    .Y(_05226_));
 sky130_fd_sc_hd__nand3_1 _14314_ (.A(_03656_),
    .B(_03676_),
    .C(_05226_),
    .Y(_05227_));
 sky130_fd_sc_hd__nor3_1 _14315_ (.A(_05171_),
    .B(_05214_),
    .C(_05227_),
    .Y(_05228_));
 sky130_fd_sc_hd__nor2_1 _14316_ (.A(_03666_),
    .B(_05228_),
    .Y(_05229_));
 sky130_fd_sc_hd__a21oi_1 _14317_ (.A1(_04995_),
    .A2(_05148_),
    .B1(_03639_),
    .Y(_05230_));
 sky130_fd_sc_hd__a31oi_1 _14318_ (.A1(_03639_),
    .A2(_04925_),
    .A3(_05096_),
    .B1(_05230_),
    .Y(_05231_));
 sky130_fd_sc_hd__nand4_1 _14319_ (.A(_03637_),
    .B(_03675_),
    .C(_05073_),
    .D(_05020_),
    .Y(_05232_));
 sky130_fd_sc_hd__o21ai_0 _14320_ (.A1(net4064),
    .A2(_03675_),
    .B1(_11908_[0]),
    .Y(_05233_));
 sky130_fd_sc_hd__o21ai_0 _14321_ (.A1(_03639_),
    .A2(_03676_),
    .B1(_05233_),
    .Y(_05234_));
 sky130_fd_sc_hd__o21ai_0 _14322_ (.A1(_11912_[0]),
    .A2(net4064),
    .B1(_03639_),
    .Y(_05235_));
 sky130_fd_sc_hd__o21ai_0 _14323_ (.A1(_03675_),
    .A2(_05235_),
    .B1(_03658_),
    .Y(_05236_));
 sky130_fd_sc_hd__a21oi_1 _14324_ (.A1(_05232_),
    .A2(_05234_),
    .B1(_05236_),
    .Y(_05237_));
 sky130_fd_sc_hd__a31oi_1 _14325_ (.A1(_03656_),
    .A2(_03675_),
    .A3(_05231_),
    .B1(_05237_),
    .Y(_05238_));
 sky130_fd_sc_hd__o21ai_0 _14326_ (.A1(_03631_),
    .A2(_03639_),
    .B1(_05138_),
    .Y(_05239_));
 sky130_fd_sc_hd__o21ai_0 _14327_ (.A1(_04943_),
    .A2(_05171_),
    .B1(net4094),
    .Y(_05240_));
 sky130_fd_sc_hd__a211oi_1 _14328_ (.A1(_11910_[0]),
    .A2(_04970_),
    .B1(_05068_),
    .C1(_03656_),
    .Y(_05241_));
 sky130_fd_sc_hd__a31oi_1 _14329_ (.A1(_03656_),
    .A2(_05239_),
    .A3(_05240_),
    .B1(_05241_),
    .Y(_05242_));
 sky130_fd_sc_hd__o21ai_0 _14330_ (.A1(_05041_),
    .A2(_04899_),
    .B1(_03676_),
    .Y(_05243_));
 sky130_fd_sc_hd__o21ai_0 _14331_ (.A1(_11903_[0]),
    .A2(_03648_),
    .B1(_04925_),
    .Y(_05244_));
 sky130_fd_sc_hd__a21oi_1 _14332_ (.A1(_05002_),
    .A2(_05096_),
    .B1(_03639_),
    .Y(_05245_));
 sky130_fd_sc_hd__a21oi_1 _14333_ (.A1(_03639_),
    .A2(_05244_),
    .B1(_05245_),
    .Y(_05246_));
 sky130_fd_sc_hd__o21ai_0 _14334_ (.A1(net4094),
    .A2(_03639_),
    .B1(_03648_),
    .Y(_05247_));
 sky130_fd_sc_hd__a21oi_1 _14335_ (.A1(_11910_[0]),
    .A2(_03639_),
    .B1(_05247_),
    .Y(_05248_));
 sky130_fd_sc_hd__o22ai_1 _14336_ (.A1(_03656_),
    .A2(_05246_),
    .B1(_05248_),
    .B2(_05079_),
    .Y(_05249_));
 sky130_fd_sc_hd__o22ai_1 _14337_ (.A1(_05242_),
    .A2(_05243_),
    .B1(_05249_),
    .B2(_03676_),
    .Y(_05250_));
 sky130_fd_sc_hd__a221oi_1 _14338_ (.A1(_05229_),
    .A2(_05238_),
    .B1(_05250_),
    .B2(_03666_),
    .C1(_03684_),
    .Y(_05251_));
 sky130_fd_sc_hd__a21oi_4 _14339_ (.A1(_03684_),
    .A2(_05225_),
    .B1(_05251_),
    .Y(_00020_));
 sky130_fd_sc_hd__nor3b_1 _14340_ (.A(_05101_),
    .B(_03639_),
    .C_N(_04925_),
    .Y(_05252_));
 sky130_fd_sc_hd__nor3_1 _14341_ (.A(net4093),
    .B(_05031_),
    .C(_05090_),
    .Y(_05253_));
 sky130_fd_sc_hd__o21ai_0 _14342_ (.A1(_05252_),
    .A2(_05253_),
    .B1(_03676_),
    .Y(_05254_));
 sky130_fd_sc_hd__o221ai_1 _14343_ (.A1(_11898_[0]),
    .A2(_05018_),
    .B1(_05069_),
    .B2(net4064),
    .C1(_03675_),
    .Y(_05255_));
 sky130_fd_sc_hd__nand2_1 _14344_ (.A(_03625_),
    .B(_05001_),
    .Y(_05256_));
 sky130_fd_sc_hd__a211oi_1 _14345_ (.A1(_11901_[0]),
    .A2(_04943_),
    .B1(_05154_),
    .C1(_03676_),
    .Y(_05257_));
 sky130_fd_sc_hd__a311oi_1 _14346_ (.A1(_03676_),
    .A2(_05187_),
    .A3(_05256_),
    .B1(_05257_),
    .C1(_03658_),
    .Y(_05258_));
 sky130_fd_sc_hd__a31oi_1 _14347_ (.A1(_03658_),
    .A2(_05254_),
    .A3(_05255_),
    .B1(_05258_),
    .Y(_05259_));
 sky130_fd_sc_hd__nor2_1 _14348_ (.A(_03685_),
    .B(_05259_),
    .Y(_05260_));
 sky130_fd_sc_hd__nand3b_1 _14349_ (.A_N(_05101_),
    .B(_03637_),
    .C(_04954_),
    .Y(_05261_));
 sky130_fd_sc_hd__nand3_1 _14350_ (.A(_03639_),
    .B(_04961_),
    .C(_05105_),
    .Y(_05262_));
 sky130_fd_sc_hd__nand3_1 _14351_ (.A(_03658_),
    .B(_05261_),
    .C(_05262_),
    .Y(_05263_));
 sky130_fd_sc_hd__nand2_1 _14352_ (.A(_11898_[0]),
    .B(net4093),
    .Y(_05264_));
 sky130_fd_sc_hd__a21boi_0 _14353_ (.A1(_11903_[0]),
    .A2(_03639_),
    .B1_N(_05264_),
    .Y(_05265_));
 sky130_fd_sc_hd__o21ai_0 _14354_ (.A1(net4092),
    .A2(_05265_),
    .B1(_04901_),
    .Y(_05266_));
 sky130_fd_sc_hd__nor2_1 _14355_ (.A(net4092),
    .B(_03658_),
    .Y(_05267_));
 sky130_fd_sc_hd__nor2_1 _14356_ (.A(_03656_),
    .B(_05041_),
    .Y(_05268_));
 sky130_fd_sc_hd__o21ai_0 _14357_ (.A1(_05267_),
    .A2(_05268_),
    .B1(net4096),
    .Y(_05269_));
 sky130_fd_sc_hd__o21ai_0 _14358_ (.A1(_03631_),
    .A2(_03658_),
    .B1(_04980_),
    .Y(_05270_));
 sky130_fd_sc_hd__nor2_1 _14359_ (.A(_03648_),
    .B(_03658_),
    .Y(_05271_));
 sky130_fd_sc_hd__nor2_1 _14360_ (.A(net4092),
    .B(_03656_),
    .Y(_05272_));
 sky130_fd_sc_hd__a222oi_1 _14361_ (.A1(net4065),
    .A2(_05270_),
    .B1(_05271_),
    .B2(_04899_),
    .C1(_05272_),
    .C2(_05055_),
    .Y(_05273_));
 sky130_fd_sc_hd__a21oi_1 _14362_ (.A1(_05269_),
    .A2(_05273_),
    .B1(_03676_),
    .Y(_05274_));
 sky130_fd_sc_hd__a311oi_2 _14363_ (.A1(_03676_),
    .A2(_05263_),
    .A3(_05266_),
    .B1(net3628),
    .C1(_05274_),
    .Y(_05275_));
 sky130_fd_sc_hd__nand3_1 _14364_ (.A(_11896_[0]),
    .B(_03639_),
    .C(net4092),
    .Y(_05276_));
 sky130_fd_sc_hd__nand3_1 _14365_ (.A(_03637_),
    .B(_05096_),
    .C(_05175_),
    .Y(_05277_));
 sky130_fd_sc_hd__a21o_1 _14366_ (.A1(_05073_),
    .A2(_04959_),
    .B1(_03637_),
    .X(_05278_));
 sky130_fd_sc_hd__a21oi_1 _14367_ (.A1(_05277_),
    .A2(_05278_),
    .B1(_03656_),
    .Y(_05279_));
 sky130_fd_sc_hd__a311oi_1 _14368_ (.A1(_03656_),
    .A2(_05175_),
    .A3(_05276_),
    .B1(_05279_),
    .C1(_03676_),
    .Y(_05280_));
 sky130_fd_sc_hd__nor2_1 _14369_ (.A(net4099),
    .B(net4093),
    .Y(_05281_));
 sky130_fd_sc_hd__o21ai_2 _14370_ (.A1(_05078_),
    .A2(_05281_),
    .B1(_04949_),
    .Y(_05282_));
 sky130_fd_sc_hd__o211ai_1 _14371_ (.A1(_11896_[0]),
    .A2(_05014_),
    .B1(_05277_),
    .C1(_03658_),
    .Y(_05283_));
 sky130_fd_sc_hd__a21oi_1 _14372_ (.A1(_05282_),
    .A2(_05283_),
    .B1(_03675_),
    .Y(_05284_));
 sky130_fd_sc_hd__o21ai_0 _14373_ (.A1(_05280_),
    .A2(_05284_),
    .B1(_03684_),
    .Y(_05285_));
 sky130_fd_sc_hd__nand2_1 _14374_ (.A(_03639_),
    .B(_05020_),
    .Y(_05286_));
 sky130_fd_sc_hd__a21oi_1 _14375_ (.A1(_04925_),
    .A2(_05286_),
    .B1(_03675_),
    .Y(_05287_));
 sky130_fd_sc_hd__a21oi_1 _14376_ (.A1(_04971_),
    .A2(_05073_),
    .B1(_03639_),
    .Y(_05288_));
 sky130_fd_sc_hd__a211oi_1 _14377_ (.A1(_03631_),
    .A2(_04989_),
    .B1(_05288_),
    .C1(_03676_),
    .Y(_05289_));
 sky130_fd_sc_hd__a21oi_1 _14378_ (.A1(_04975_),
    .A2(_05046_),
    .B1(_03639_),
    .Y(_05290_));
 sky130_fd_sc_hd__o21ai_0 _14379_ (.A1(_11897_[0]),
    .A2(_04923_),
    .B1(_03675_),
    .Y(_05291_));
 sky130_fd_sc_hd__nor2_1 _14380_ (.A(_03639_),
    .B(_04961_),
    .Y(_05292_));
 sky130_fd_sc_hd__a31oi_1 _14381_ (.A1(_03639_),
    .A2(_04995_),
    .A3(_05148_),
    .B1(_05292_),
    .Y(_05293_));
 sky130_fd_sc_hd__o221ai_1 _14382_ (.A1(_05290_),
    .A2(_05291_),
    .B1(_05293_),
    .B2(_03675_),
    .C1(_03656_),
    .Y(_05294_));
 sky130_fd_sc_hd__o311ai_1 _14383_ (.A1(_03656_),
    .A2(_05287_),
    .A3(_05289_),
    .B1(_03685_),
    .C1(_05294_),
    .Y(_05295_));
 sky130_fd_sc_hd__nand3_1 _14384_ (.A(_03666_),
    .B(_05285_),
    .C(_05295_),
    .Y(_05296_));
 sky130_fd_sc_hd__o31ai_2 _14385_ (.A1(_03666_),
    .A2(_05260_),
    .A3(_05275_),
    .B1(_05296_),
    .Y(_00021_));
 sky130_fd_sc_hd__o21ai_0 _14386_ (.A1(_03639_),
    .A2(_04972_),
    .B1(_05165_),
    .Y(_05297_));
 sky130_fd_sc_hd__nand2_1 _14387_ (.A(_05018_),
    .B(_05014_),
    .Y(_05298_));
 sky130_fd_sc_hd__nor2_1 _14388_ (.A(_11901_[0]),
    .B(_04923_),
    .Y(_05299_));
 sky130_fd_sc_hd__a2111oi_0 _14389_ (.A1(_03625_),
    .A2(_05298_),
    .B1(_05013_),
    .C1(_05299_),
    .D1(_03667_),
    .Y(_05300_));
 sky130_fd_sc_hd__a211oi_1 _14390_ (.A1(_03667_),
    .A2(_05297_),
    .B1(_05300_),
    .C1(_03658_),
    .Y(_05301_));
 sky130_fd_sc_hd__a21oi_1 _14391_ (.A1(_05002_),
    .A2(_05153_),
    .B1(_03639_),
    .Y(_05302_));
 sky130_fd_sc_hd__o211ai_1 _14392_ (.A1(_11897_[0]),
    .A2(net4093),
    .B1(net4092),
    .C1(_04907_),
    .Y(_05303_));
 sky130_fd_sc_hd__o211ai_1 _14393_ (.A1(_11920_[0]),
    .A2(net4092),
    .B1(_03667_),
    .C1(_05303_),
    .Y(_05304_));
 sky130_fd_sc_hd__o311a_1 _14394_ (.A1(_03667_),
    .A2(_05299_),
    .A3(_05302_),
    .B1(_05304_),
    .C1(_03658_),
    .X(_05305_));
 sky130_fd_sc_hd__o21ai_2 _14395_ (.A1(_05301_),
    .A2(_05305_),
    .B1(_03685_),
    .Y(_05306_));
 sky130_fd_sc_hd__nor2_1 _14396_ (.A(_11903_[0]),
    .B(_03639_),
    .Y(_05307_));
 sky130_fd_sc_hd__o21ai_0 _14397_ (.A1(_05077_),
    .A2(_05307_),
    .B1(_03648_),
    .Y(_05308_));
 sky130_fd_sc_hd__o211ai_1 _14398_ (.A1(_11908_[0]),
    .A2(_03639_),
    .B1(net4092),
    .C1(_04904_),
    .Y(_05309_));
 sky130_fd_sc_hd__o211ai_1 _14399_ (.A1(_11916_[0]),
    .A2(net4092),
    .B1(_03667_),
    .C1(_05309_),
    .Y(_05310_));
 sky130_fd_sc_hd__o21ai_0 _14400_ (.A1(_03667_),
    .A2(_05308_),
    .B1(_05310_),
    .Y(_05311_));
 sky130_fd_sc_hd__nand2_1 _14401_ (.A(_03656_),
    .B(_05311_),
    .Y(_05312_));
 sky130_fd_sc_hd__o21ai_0 _14402_ (.A1(_11897_[0]),
    .A2(net4093),
    .B1(_05264_),
    .Y(_05313_));
 sky130_fd_sc_hd__nand2_1 _14403_ (.A(_03648_),
    .B(_05313_),
    .Y(_05314_));
 sky130_fd_sc_hd__a32oi_1 _14404_ (.A1(_03637_),
    .A2(_05153_),
    .A3(_05148_),
    .B1(_04991_),
    .B2(_03631_),
    .Y(_05315_));
 sky130_fd_sc_hd__nor3_1 _14405_ (.A(_03656_),
    .B(_03667_),
    .C(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__a31oi_1 _14406_ (.A1(_03667_),
    .A2(_05030_),
    .A3(_05314_),
    .B1(_05316_),
    .Y(_05317_));
 sky130_fd_sc_hd__nand3_2 _14407_ (.A(_03684_),
    .B(_05312_),
    .C(_05317_),
    .Y(_05318_));
 sky130_fd_sc_hd__o21ai_0 _14408_ (.A1(_11908_[0]),
    .A2(_03648_),
    .B1(_05061_),
    .Y(_05319_));
 sky130_fd_sc_hd__o211ai_1 _14409_ (.A1(_11912_[0]),
    .A2(net4092),
    .B1(_05096_),
    .C1(_03639_),
    .Y(_05320_));
 sky130_fd_sc_hd__o21ai_0 _14410_ (.A1(_03639_),
    .A2(_05319_),
    .B1(_05320_),
    .Y(_05321_));
 sky130_fd_sc_hd__o221ai_1 _14411_ (.A1(net4094),
    .A2(_04970_),
    .B1(_05015_),
    .B2(_03625_),
    .C1(_03667_),
    .Y(_05322_));
 sky130_fd_sc_hd__o21ai_0 _14412_ (.A1(_03667_),
    .A2(_05321_),
    .B1(_05322_),
    .Y(_05323_));
 sky130_fd_sc_hd__nor2_1 _14413_ (.A(_03658_),
    .B(_05323_),
    .Y(_05324_));
 sky130_fd_sc_hd__a221oi_1 _14414_ (.A1(_11908_[0]),
    .A2(_04991_),
    .B1(_05298_),
    .B2(_03625_),
    .C1(_05013_),
    .Y(_05325_));
 sky130_fd_sc_hd__a21oi_1 _14415_ (.A1(_05040_),
    .A2(_05148_),
    .B1(net4093),
    .Y(_05326_));
 sky130_fd_sc_hd__a211oi_1 _14416_ (.A1(_11912_[0]),
    .A2(_04970_),
    .B1(_05326_),
    .C1(_03666_),
    .Y(_05327_));
 sky130_fd_sc_hd__a211oi_1 _14417_ (.A1(_03666_),
    .A2(_05325_),
    .B1(_05327_),
    .C1(_03656_),
    .Y(_05328_));
 sky130_fd_sc_hd__o21ai_2 _14418_ (.A1(_05324_),
    .A2(_05328_),
    .B1(_03685_),
    .Y(_05329_));
 sky130_fd_sc_hd__o21ai_0 _14419_ (.A1(net4098),
    .A2(net4093),
    .B1(_04907_),
    .Y(_05330_));
 sky130_fd_sc_hd__nand2_1 _14420_ (.A(net4092),
    .B(_05330_),
    .Y(_05331_));
 sky130_fd_sc_hd__o22ai_1 _14421_ (.A1(net4065),
    .A2(_03639_),
    .B1(_05014_),
    .B2(_11898_[0]),
    .Y(_05332_));
 sky130_fd_sc_hd__nor3_1 _14422_ (.A(_03666_),
    .B(_05162_),
    .C(_05332_),
    .Y(_05333_));
 sky130_fd_sc_hd__a31oi_1 _14423_ (.A1(_03666_),
    .A2(_05070_),
    .A3(_05331_),
    .B1(_05333_),
    .Y(_05334_));
 sky130_fd_sc_hd__o21ai_0 _14424_ (.A1(_03639_),
    .A2(_05138_),
    .B1(net4094),
    .Y(_05335_));
 sky130_fd_sc_hd__a22oi_1 _14425_ (.A1(_11901_[0]),
    .A2(_04943_),
    .B1(_04991_),
    .B2(net4098),
    .Y(_05336_));
 sky130_fd_sc_hd__o21ai_0 _14426_ (.A1(_03639_),
    .A2(_05138_),
    .B1(_03666_),
    .Y(_05337_));
 sky130_fd_sc_hd__a31oi_1 _14427_ (.A1(_03639_),
    .A2(_04995_),
    .A3(_05148_),
    .B1(_05337_),
    .Y(_05338_));
 sky130_fd_sc_hd__a311oi_1 _14428_ (.A1(_03667_),
    .A2(_05335_),
    .A3(_05336_),
    .B1(_05338_),
    .C1(_03658_),
    .Y(_05339_));
 sky130_fd_sc_hd__a21oi_1 _14429_ (.A1(_03658_),
    .A2(_05334_),
    .B1(_05339_),
    .Y(_05340_));
 sky130_fd_sc_hd__a21oi_2 _14430_ (.A1(_03684_),
    .A2(_05340_),
    .B1(_03675_),
    .Y(_05341_));
 sky130_fd_sc_hd__a32oi_4 _14431_ (.A1(_03675_),
    .A2(_05306_),
    .A3(_05318_),
    .B1(_05329_),
    .B2(_05341_),
    .Y(_00022_));
 sky130_fd_sc_hd__a21oi_1 _14432_ (.A1(_05105_),
    .A2(_04954_),
    .B1(net4093),
    .Y(_05342_));
 sky130_fd_sc_hd__o211ai_1 _14433_ (.A1(_11896_[0]),
    .A2(_03648_),
    .B1(_05148_),
    .C1(net4093),
    .Y(_05343_));
 sky130_fd_sc_hd__o311ai_0 _14434_ (.A1(net4093),
    .A2(_05138_),
    .A3(_05090_),
    .B1(_05343_),
    .C1(_03676_),
    .Y(_05344_));
 sky130_fd_sc_hd__o311ai_0 _14435_ (.A1(_03676_),
    .A2(_05064_),
    .A3(_05342_),
    .B1(_05344_),
    .C1(_03658_),
    .Y(_05345_));
 sky130_fd_sc_hd__o22ai_1 _14436_ (.A1(_11896_[0]),
    .A2(net4092),
    .B1(_04971_),
    .B2(_03639_),
    .Y(_05346_));
 sky130_fd_sc_hd__nand3_1 _14437_ (.A(net4093),
    .B(_05025_),
    .C(_05175_),
    .Y(_05347_));
 sky130_fd_sc_hd__nand3_1 _14438_ (.A(_03676_),
    .B(_05033_),
    .C(_05347_),
    .Y(_05348_));
 sky130_fd_sc_hd__o21ai_0 _14439_ (.A1(_03676_),
    .A2(_05346_),
    .B1(_05348_),
    .Y(_05349_));
 sky130_fd_sc_hd__nand2_1 _14440_ (.A(net4091),
    .B(_05349_),
    .Y(_05350_));
 sky130_fd_sc_hd__nand3_2 _14441_ (.A(_03685_),
    .B(_05345_),
    .C(_05350_),
    .Y(_05351_));
 sky130_fd_sc_hd__a31oi_1 _14442_ (.A1(net4093),
    .A2(_04926_),
    .A3(_05061_),
    .B1(_04976_),
    .Y(_05352_));
 sky130_fd_sc_hd__nor2_1 _14443_ (.A(_03656_),
    .B(_05352_),
    .Y(_05353_));
 sky130_fd_sc_hd__a21oi_1 _14444_ (.A1(_05002_),
    .A2(_05096_),
    .B1(net4093),
    .Y(_05354_));
 sky130_fd_sc_hd__nor2_1 _14445_ (.A(_11908_[0]),
    .B(_05018_),
    .Y(_05355_));
 sky130_fd_sc_hd__nor3_1 _14446_ (.A(_03658_),
    .B(_05354_),
    .C(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__a21oi_1 _14447_ (.A1(_03639_),
    .A2(_05271_),
    .B1(_04970_),
    .Y(_05357_));
 sky130_fd_sc_hd__nor4_1 _14448_ (.A(_11896_[0]),
    .B(_03639_),
    .C(_03648_),
    .D(_03658_),
    .Y(_05358_));
 sky130_fd_sc_hd__a21oi_1 _14449_ (.A1(_05281_),
    .A2(_05272_),
    .B1(_05358_),
    .Y(_05359_));
 sky130_fd_sc_hd__a31oi_1 _14450_ (.A1(net4099),
    .A2(_03631_),
    .A3(_05267_),
    .B1(_05268_),
    .Y(_05360_));
 sky130_fd_sc_hd__o2111ai_2 _14451_ (.A1(_03631_),
    .A2(_05357_),
    .B1(_05359_),
    .C1(_03675_),
    .D1(_05360_),
    .Y(_05361_));
 sky130_fd_sc_hd__o311ai_2 _14452_ (.A1(_03675_),
    .A2(_05353_),
    .A3(_05356_),
    .B1(_05361_),
    .C1(net3628),
    .Y(_05362_));
 sky130_fd_sc_hd__o221ai_1 _14453_ (.A1(_11898_[0]),
    .A2(_04923_),
    .B1(_04990_),
    .B2(_11897_[0]),
    .C1(_05036_),
    .Y(_05363_));
 sky130_fd_sc_hd__a21oi_1 _14454_ (.A1(_04961_),
    .A2(_05046_),
    .B1(net4093),
    .Y(_05364_));
 sky130_fd_sc_hd__a22o_1 _14455_ (.A1(_11917_[0]),
    .A2(_03648_),
    .B1(_04943_),
    .B2(_11908_[0]),
    .X(_05365_));
 sky130_fd_sc_hd__nor3_1 _14456_ (.A(_03658_),
    .B(_05364_),
    .C(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__a211o_1 _14457_ (.A1(_03658_),
    .A2(_05363_),
    .B1(_05366_),
    .C1(_03675_),
    .X(_05367_));
 sky130_fd_sc_hd__nand3_1 _14458_ (.A(_11901_[0]),
    .B(_03648_),
    .C(_03658_),
    .Y(_05368_));
 sky130_fd_sc_hd__nand3_1 _14459_ (.A(_03639_),
    .B(_04995_),
    .C(_05368_),
    .Y(_05369_));
 sky130_fd_sc_hd__o21ai_0 _14460_ (.A1(_03639_),
    .A2(_03656_),
    .B1(_05369_),
    .Y(_05370_));
 sky130_fd_sc_hd__o21ai_0 _14461_ (.A1(_04943_),
    .A2(_05267_),
    .B1(_11896_[0]),
    .Y(_05371_));
 sky130_fd_sc_hd__nand3_1 _14462_ (.A(_03675_),
    .B(_05370_),
    .C(_05371_),
    .Y(_05372_));
 sky130_fd_sc_hd__a21oi_1 _14463_ (.A1(_05367_),
    .A2(_05372_),
    .B1(_03685_),
    .Y(_05373_));
 sky130_fd_sc_hd__xnor2_1 _14464_ (.A(_11897_[0]),
    .B(_03639_),
    .Y(_05374_));
 sky130_fd_sc_hd__o2111ai_1 _14465_ (.A1(net4092),
    .A2(_05374_),
    .B1(_05116_),
    .C1(_05030_),
    .D1(_03675_),
    .Y(_05375_));
 sky130_fd_sc_hd__o21ai_0 _14466_ (.A1(_04946_),
    .A2(_05115_),
    .B1(net4092),
    .Y(_05376_));
 sky130_fd_sc_hd__nand2_1 _14467_ (.A(_05226_),
    .B(_05376_),
    .Y(_05377_));
 sky130_fd_sc_hd__a21oi_1 _14468_ (.A1(_11912_[0]),
    .A2(net4092),
    .B1(_03639_),
    .Y(_05378_));
 sky130_fd_sc_hd__a221oi_1 _14469_ (.A1(_11910_[0]),
    .A2(_03639_),
    .B1(_05002_),
    .B2(_05378_),
    .C1(_03675_),
    .Y(_05379_));
 sky130_fd_sc_hd__a211o_1 _14470_ (.A1(_03675_),
    .A2(_05377_),
    .B1(_05379_),
    .C1(_03658_),
    .X(_05380_));
 sky130_fd_sc_hd__o2111ai_1 _14471_ (.A1(_05172_),
    .A2(_05247_),
    .B1(_03658_),
    .C1(_03676_),
    .D1(_05020_),
    .Y(_05381_));
 sky130_fd_sc_hd__and4_1 _14472_ (.A(_03685_),
    .B(_05375_),
    .C(_05380_),
    .D(_05381_),
    .X(_05382_));
 sky130_fd_sc_hd__nor3_2 _14473_ (.A(_03667_),
    .B(_05373_),
    .C(_05382_),
    .Y(_05383_));
 sky130_fd_sc_hd__a31oi_4 _14474_ (.A1(_03667_),
    .A2(_05351_),
    .A3(_05362_),
    .B1(_05383_),
    .Y(_00023_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1121 ();
 sky130_fd_sc_hd__and2_4 _14482_ (.A(_03817_),
    .B(_03824_),
    .X(_05388_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1117 ();
 sky130_fd_sc_hd__nand2_4 _14487_ (.A(_03773_),
    .B(_03792_),
    .Y(_05393_));
 sky130_fd_sc_hd__nand2_8 _14488_ (.A(net4083),
    .B(net4077),
    .Y(_05394_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1116 ();
 sky130_fd_sc_hd__a21oi_2 _14490_ (.A1(_05393_),
    .A2(_05394_),
    .B1(net4080),
    .Y(_05396_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1115 ();
 sky130_fd_sc_hd__nand2_2 _14492_ (.A(_11944_[0]),
    .B(_03792_),
    .Y(_05398_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1113 ();
 sky130_fd_sc_hd__nand2_2 _14495_ (.A(_11935_[0]),
    .B(net4076),
    .Y(_05401_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1111 ();
 sky130_fd_sc_hd__a21oi_2 _14498_ (.A1(_05398_),
    .A2(_05401_),
    .B1(_03784_),
    .Y(_05404_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1109 ();
 sky130_fd_sc_hd__o21ai_0 _14501_ (.A1(_05396_),
    .A2(_05404_),
    .B1(net4060),
    .Y(_05407_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1108 ();
 sky130_fd_sc_hd__and2_4 _14503_ (.A(_11935_[0]),
    .B(_03792_),
    .X(_05409_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1107 ();
 sky130_fd_sc_hd__nor2_4 _14505_ (.A(_11946_[0]),
    .B(_03792_),
    .Y(_05411_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1106 ();
 sky130_fd_sc_hd__nor2_4 _14507_ (.A(net4078),
    .B(net4074),
    .Y(_05413_));
 sky130_fd_sc_hd__a21oi_1 _14508_ (.A1(_11942_[0]),
    .A2(_05413_),
    .B1(net4060),
    .Y(_05414_));
 sky130_fd_sc_hd__o31ai_1 _14509_ (.A1(_03784_),
    .A2(_05409_),
    .A3(_05411_),
    .B1(_05414_),
    .Y(_05415_));
 sky130_fd_sc_hd__nand3_1 _14510_ (.A(net4073),
    .B(_05407_),
    .C(_05415_),
    .Y(_05416_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1105 ();
 sky130_fd_sc_hd__nand2_4 _14512_ (.A(_03784_),
    .B(net4075),
    .Y(_05418_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1104 ();
 sky130_fd_sc_hd__nor2_1 _14514_ (.A(_11935_[0]),
    .B(_03792_),
    .Y(_05420_));
 sky130_fd_sc_hd__a21oi_1 _14515_ (.A1(_11946_[0]),
    .A2(_03792_),
    .B1(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__o221ai_1 _14516_ (.A1(_11940_[0]),
    .A2(_05418_),
    .B1(_05421_),
    .B2(_03784_),
    .C1(_03810_),
    .Y(_05422_));
 sky130_fd_sc_hd__nor2_4 _14517_ (.A(net4078),
    .B(_03792_),
    .Y(_05423_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1102 ();
 sky130_fd_sc_hd__a221o_1 _14520_ (.A1(_11951_[0]),
    .A2(_03792_),
    .B1(_05423_),
    .B2(net395),
    .C1(_03810_),
    .X(_05426_));
 sky130_fd_sc_hd__nand3_1 _14521_ (.A(_03801_),
    .B(_05422_),
    .C(_05426_),
    .Y(_05427_));
 sky130_fd_sc_hd__nand2_8 _14522_ (.A(_00398_),
    .B(_03824_),
    .Y(_05428_));
 sky130_fd_sc_hd__nor2_4 _14523_ (.A(net4074),
    .B(net4073),
    .Y(_05429_));
 sky130_fd_sc_hd__o21ai_0 _14524_ (.A1(net395),
    .A2(_03784_),
    .B1(_05429_),
    .Y(_05430_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1100 ();
 sky130_fd_sc_hd__nand2_4 _14527_ (.A(net4083),
    .B(_03792_),
    .Y(_05433_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1097 ();
 sky130_fd_sc_hd__nand2_4 _14531_ (.A(_11937_[0]),
    .B(net4077),
    .Y(_05437_));
 sky130_fd_sc_hd__o21ai_0 _14532_ (.A1(_03801_),
    .A2(_05433_),
    .B1(_05437_),
    .Y(_05438_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1095 ();
 sky130_fd_sc_hd__nand2_1 _14535_ (.A(_03792_),
    .B(net4073),
    .Y(_05441_));
 sky130_fd_sc_hd__nand2_2 _14536_ (.A(net4074),
    .B(_03801_),
    .Y(_05442_));
 sky130_fd_sc_hd__clkinv_2 _14537_ (.A(_11942_[0]),
    .Y(_05443_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1094 ();
 sky130_fd_sc_hd__o221ai_1 _14539_ (.A1(_11930_[0]),
    .A2(_05441_),
    .B1(_05442_),
    .B2(_05443_),
    .C1(net4078),
    .Y(_05445_));
 sky130_fd_sc_hd__o21ai_0 _14540_ (.A1(net4080),
    .A2(_05438_),
    .B1(_05445_),
    .Y(_05446_));
 sky130_fd_sc_hd__nand2_8 _14541_ (.A(_03778_),
    .B(net4076),
    .Y(_05447_));
 sky130_fd_sc_hd__nor2_2 _14542_ (.A(_11940_[0]),
    .B(net4074),
    .Y(_05448_));
 sky130_fd_sc_hd__nor2_4 _14543_ (.A(net395),
    .B(_03792_),
    .Y(_05449_));
 sky130_fd_sc_hd__nor3_1 _14544_ (.A(net4080),
    .B(_05448_),
    .C(_05449_),
    .Y(_05450_));
 sky130_fd_sc_hd__a31oi_1 _14545_ (.A1(net4080),
    .A2(_05447_),
    .A3(_05433_),
    .B1(_05450_),
    .Y(_05451_));
 sky130_fd_sc_hd__nor2_4 _14546_ (.A(_11937_[0]),
    .B(net4074),
    .Y(_05452_));
 sky130_fd_sc_hd__o21ai_0 _14547_ (.A1(_05452_),
    .A2(_05411_),
    .B1(net4080),
    .Y(_05453_));
 sky130_fd_sc_hd__a21oi_1 _14548_ (.A1(_11944_[0]),
    .A2(_05423_),
    .B1(net4073),
    .Y(_05454_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1093 ();
 sky130_fd_sc_hd__a221oi_1 _14550_ (.A1(net4073),
    .A2(_05451_),
    .B1(_05453_),
    .B2(_05454_),
    .C1(net4060),
    .Y(_05456_));
 sky130_fd_sc_hd__a31oi_1 _14551_ (.A1(net4060),
    .A2(_05430_),
    .A3(_05446_),
    .B1(_05456_),
    .Y(_05457_));
 sky130_fd_sc_hd__nor2_1 _14552_ (.A(_05428_),
    .B(_05457_),
    .Y(_05458_));
 sky130_fd_sc_hd__xnor2_2 _14553_ (.A(_03784_),
    .B(_03792_),
    .Y(_05459_));
 sky130_fd_sc_hd__nand2_8 _14554_ (.A(net4078),
    .B(_03792_),
    .Y(_05460_));
 sky130_fd_sc_hd__nor2_4 _14555_ (.A(net395),
    .B(_05460_),
    .Y(_05461_));
 sky130_fd_sc_hd__a221oi_1 _14556_ (.A1(_11940_[0]),
    .A2(_05423_),
    .B1(_05459_),
    .B2(_11944_[0]),
    .C1(_05461_),
    .Y(_05462_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1092 ();
 sky130_fd_sc_hd__nand2_4 _14558_ (.A(_03778_),
    .B(_03784_),
    .Y(_05464_));
 sky130_fd_sc_hd__nor2_2 _14559_ (.A(net395),
    .B(net4078),
    .Y(_05465_));
 sky130_fd_sc_hd__a32oi_1 _14560_ (.A1(net395),
    .A2(net4074),
    .A3(_05464_),
    .B1(_05447_),
    .B2(_05465_),
    .Y(_05466_));
 sky130_fd_sc_hd__nand2_1 _14561_ (.A(_03801_),
    .B(_05466_),
    .Y(_05467_));
 sky130_fd_sc_hd__o21ai_0 _14562_ (.A1(_03801_),
    .A2(_05462_),
    .B1(_05467_),
    .Y(_05468_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1091 ();
 sky130_fd_sc_hd__nand2_1 _14564_ (.A(_03809_),
    .B(_03817_),
    .Y(_05470_));
 sky130_fd_sc_hd__nor2_4 _14565_ (.A(_03773_),
    .B(_03784_),
    .Y(_05471_));
 sky130_fd_sc_hd__a21oi_1 _14566_ (.A1(_03773_),
    .A2(_03778_),
    .B1(_05471_),
    .Y(_05472_));
 sky130_fd_sc_hd__xnor2_1 _14567_ (.A(net4076),
    .B(_05472_),
    .Y(_05473_));
 sky130_fd_sc_hd__clkinv_8 _14568_ (.A(_11931_[0]),
    .Y(_05474_));
 sky130_fd_sc_hd__nor2_2 _14569_ (.A(_05474_),
    .B(_03792_),
    .Y(_05475_));
 sky130_fd_sc_hd__o21ai_0 _14570_ (.A1(_05448_),
    .A2(_05475_),
    .B1(net4078),
    .Y(_05476_));
 sky130_fd_sc_hd__nand2_2 _14571_ (.A(_11930_[0]),
    .B(net4076),
    .Y(_05477_));
 sky130_fd_sc_hd__nand3_1 _14572_ (.A(_03784_),
    .B(_05398_),
    .C(_05477_),
    .Y(_05478_));
 sky130_fd_sc_hd__nand3_1 _14573_ (.A(net4073),
    .B(_05476_),
    .C(_05478_),
    .Y(_05479_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1090 ();
 sky130_fd_sc_hd__o2111ai_1 _14575_ (.A1(net4073),
    .A2(_05473_),
    .B1(_05479_),
    .C1(_03810_),
    .D1(_03817_),
    .Y(_05481_));
 sky130_fd_sc_hd__o21ai_1 _14576_ (.A1(_05468_),
    .A2(_05470_),
    .B1(_05481_),
    .Y(_05482_));
 sky130_fd_sc_hd__nand2_4 _14577_ (.A(net4060),
    .B(_00398_),
    .Y(_05483_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1089 ();
 sky130_fd_sc_hd__nand2_4 _14579_ (.A(_03777_),
    .B(_03784_),
    .Y(_05485_));
 sky130_fd_sc_hd__nand2b_2 _14580_ (.A_N(_11946_[0]),
    .B(net4081),
    .Y(_05486_));
 sky130_fd_sc_hd__nor2_1 _14581_ (.A(_11930_[0]),
    .B(_03784_),
    .Y(_05487_));
 sky130_fd_sc_hd__a21oi_1 _14582_ (.A1(_03772_),
    .A2(_03784_),
    .B1(_05487_),
    .Y(_05488_));
 sky130_fd_sc_hd__o21ai_2 _14583_ (.A1(net4075),
    .A2(_05488_),
    .B1(net4073),
    .Y(_05489_));
 sky130_fd_sc_hd__a31oi_2 _14584_ (.A1(net4075),
    .A2(_05485_),
    .A3(_05486_),
    .B1(_05489_),
    .Y(_05490_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1087 ();
 sky130_fd_sc_hd__nand2_2 _14587_ (.A(_11932_[0]),
    .B(_03792_),
    .Y(_05493_));
 sky130_fd_sc_hd__nand2_4 _14588_ (.A(net4082),
    .B(net4074),
    .Y(_05494_));
 sky130_fd_sc_hd__a21oi_2 _14589_ (.A1(_05493_),
    .A2(_05494_),
    .B1(_03784_),
    .Y(_05495_));
 sky130_fd_sc_hd__a311oi_1 _14590_ (.A1(_03784_),
    .A2(_05393_),
    .A3(_05401_),
    .B1(net4073),
    .C1(_05495_),
    .Y(_05496_));
 sky130_fd_sc_hd__nor3_1 _14591_ (.A(_05483_),
    .B(_05490_),
    .C(_05496_),
    .Y(_05497_));
 sky130_fd_sc_hd__nor2_2 _14592_ (.A(_11932_[0]),
    .B(net4077),
    .Y(_05498_));
 sky130_fd_sc_hd__and2_4 _14593_ (.A(_11935_[0]),
    .B(net4074),
    .X(_05499_));
 sky130_fd_sc_hd__nor3_1 _14594_ (.A(net4079),
    .B(_05498_),
    .C(_05499_),
    .Y(_05500_));
 sky130_fd_sc_hd__nand2_4 _14595_ (.A(net395),
    .B(_03792_),
    .Y(_05501_));
 sky130_fd_sc_hd__a21oi_1 _14596_ (.A1(_05394_),
    .A2(_05501_),
    .B1(_03784_),
    .Y(_05502_));
 sky130_fd_sc_hd__nand2_4 _14597_ (.A(_03810_),
    .B(_00398_),
    .Y(_05503_));
 sky130_fd_sc_hd__nor2_4 _14598_ (.A(net4073),
    .B(_05503_),
    .Y(_05504_));
 sky130_fd_sc_hd__o21ai_2 _14599_ (.A1(_05500_),
    .A2(_05502_),
    .B1(_05504_),
    .Y(_05505_));
 sky130_fd_sc_hd__nor2_2 _14600_ (.A(_03801_),
    .B(_05503_),
    .Y(_05506_));
 sky130_fd_sc_hd__nand2b_4 _14601_ (.A_N(_11935_[0]),
    .B(_03792_),
    .Y(_05507_));
 sky130_fd_sc_hd__nand3_1 _14602_ (.A(_03784_),
    .B(_05394_),
    .C(_05507_),
    .Y(_05508_));
 sky130_fd_sc_hd__o211ai_1 _14603_ (.A1(_11937_[0]),
    .A2(_05460_),
    .B1(_05506_),
    .C1(_05508_),
    .Y(_05509_));
 sky130_fd_sc_hd__nand2_1 _14604_ (.A(_05505_),
    .B(_05509_),
    .Y(_05510_));
 sky130_fd_sc_hd__nor4_1 _14605_ (.A(net3626),
    .B(_05482_),
    .C(_05497_),
    .D(_05510_),
    .Y(_05511_));
 sky130_fd_sc_hd__a311oi_2 _14606_ (.A1(_05388_),
    .A2(_05416_),
    .A3(_05427_),
    .B1(_05458_),
    .C1(_05511_),
    .Y(_00024_));
 sky130_fd_sc_hd__a31oi_1 _14607_ (.A1(net4079),
    .A2(_05501_),
    .A3(_05437_),
    .B1(_05396_),
    .Y(_05512_));
 sky130_fd_sc_hd__o21ai_0 _14608_ (.A1(_11954_[0]),
    .A2(net4076),
    .B1(net4060),
    .Y(_05513_));
 sky130_fd_sc_hd__nor2_4 _14609_ (.A(_03778_),
    .B(_03784_),
    .Y(_05514_));
 sky130_fd_sc_hd__nor2_2 _14610_ (.A(_11937_[0]),
    .B(net4079),
    .Y(_05515_));
 sky130_fd_sc_hd__nor3_1 _14611_ (.A(_03792_),
    .B(_05514_),
    .C(_05515_),
    .Y(_05516_));
 sky130_fd_sc_hd__o221ai_1 _14612_ (.A1(_03809_),
    .A2(_05512_),
    .B1(_05513_),
    .B2(_05516_),
    .C1(_03801_),
    .Y(_05517_));
 sky130_fd_sc_hd__nand2_4 _14613_ (.A(net4073),
    .B(_03809_),
    .Y(_05518_));
 sky130_fd_sc_hd__o21ai_0 _14614_ (.A1(_05498_),
    .A2(_05499_),
    .B1(net4079),
    .Y(_05519_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1086 ();
 sky130_fd_sc_hd__nand3_2 _14616_ (.A(_03784_),
    .B(_05501_),
    .C(_05437_),
    .Y(_05521_));
 sky130_fd_sc_hd__nand2_1 _14617_ (.A(_05519_),
    .B(_05521_),
    .Y(_05522_));
 sky130_fd_sc_hd__nor2_1 _14618_ (.A(_03773_),
    .B(_05447_),
    .Y(_05523_));
 sky130_fd_sc_hd__a21oi_1 _14619_ (.A1(_05494_),
    .A2(_05507_),
    .B1(net4080),
    .Y(_05524_));
 sky130_fd_sc_hd__nor2_4 _14620_ (.A(_03801_),
    .B(net4060),
    .Y(_05525_));
 sky130_fd_sc_hd__o21ai_0 _14621_ (.A1(_05523_),
    .A2(_05524_),
    .B1(_05525_),
    .Y(_05526_));
 sky130_fd_sc_hd__o21a_1 _14622_ (.A1(_05518_),
    .A2(_05522_),
    .B1(_05526_),
    .X(_05527_));
 sky130_fd_sc_hd__nor2_4 _14623_ (.A(net4073),
    .B(_03809_),
    .Y(_05528_));
 sky130_fd_sc_hd__o21ai_0 _14624_ (.A1(_11930_[0]),
    .A2(net4076),
    .B1(_05394_),
    .Y(_05529_));
 sky130_fd_sc_hd__o211ai_1 _14625_ (.A1(_11944_[0]),
    .A2(_03792_),
    .B1(_05507_),
    .C1(_03784_),
    .Y(_05530_));
 sky130_fd_sc_hd__o21ai_0 _14626_ (.A1(_03784_),
    .A2(_05529_),
    .B1(_05530_),
    .Y(_05531_));
 sky130_fd_sc_hd__a21oi_1 _14627_ (.A1(_05528_),
    .A2(_05531_),
    .B1(_00398_),
    .Y(_05532_));
 sky130_fd_sc_hd__nand3b_1 _14628_ (.A_N(_05452_),
    .B(net4080),
    .C(_05394_),
    .Y(_05533_));
 sky130_fd_sc_hd__nor2_4 _14629_ (.A(net4073),
    .B(_03810_),
    .Y(_05534_));
 sky130_fd_sc_hd__nand2_4 _14630_ (.A(_03778_),
    .B(_03792_),
    .Y(_05535_));
 sky130_fd_sc_hd__nand3_2 _14631_ (.A(_03784_),
    .B(_05494_),
    .C(_05535_),
    .Y(_05536_));
 sky130_fd_sc_hd__nand3_1 _14632_ (.A(_05533_),
    .B(_05534_),
    .C(_05536_),
    .Y(_05537_));
 sky130_fd_sc_hd__mux2i_1 _14633_ (.A0(_11930_[0]),
    .A1(_11940_[0]),
    .S(_03784_),
    .Y(_05538_));
 sky130_fd_sc_hd__a21oi_1 _14634_ (.A1(net4076),
    .A2(_05538_),
    .B1(_03801_),
    .Y(_05539_));
 sky130_fd_sc_hd__o31ai_1 _14635_ (.A1(_11958_[0]),
    .A2(net4076),
    .A3(_03810_),
    .B1(_05539_),
    .Y(_05540_));
 sky130_fd_sc_hd__nand2b_2 _14636_ (.A_N(_11946_[0]),
    .B(net4077),
    .Y(_05541_));
 sky130_fd_sc_hd__a21oi_1 _14637_ (.A1(_05394_),
    .A2(_05501_),
    .B1(net4080),
    .Y(_05542_));
 sky130_fd_sc_hd__a31oi_1 _14638_ (.A1(net4080),
    .A2(_05398_),
    .A3(_05541_),
    .B1(_05542_),
    .Y(_05543_));
 sky130_fd_sc_hd__nand2_4 _14639_ (.A(_05474_),
    .B(_03792_),
    .Y(_05544_));
 sky130_fd_sc_hd__a21oi_1 _14640_ (.A1(_05477_),
    .A2(_05544_),
    .B1(_03784_),
    .Y(_05545_));
 sky130_fd_sc_hd__a211oi_1 _14641_ (.A1(_03773_),
    .A2(_05423_),
    .B1(_05545_),
    .C1(_03810_),
    .Y(_05546_));
 sky130_fd_sc_hd__nand2_8 _14642_ (.A(_11944_[0]),
    .B(net4074),
    .Y(_05547_));
 sky130_fd_sc_hd__nand3_1 _14643_ (.A(_03784_),
    .B(_05547_),
    .C(_05535_),
    .Y(_05548_));
 sky130_fd_sc_hd__a21oi_1 _14644_ (.A1(_05533_),
    .A2(_05548_),
    .B1(net4060),
    .Y(_05549_));
 sky130_fd_sc_hd__nor3_1 _14645_ (.A(_03801_),
    .B(_05546_),
    .C(_05549_),
    .Y(_05550_));
 sky130_fd_sc_hd__a21oi_1 _14646_ (.A1(_11930_[0]),
    .A2(_03792_),
    .B1(_05411_),
    .Y(_05551_));
 sky130_fd_sc_hd__nand2_4 _14647_ (.A(_11932_[0]),
    .B(net4076),
    .Y(_05552_));
 sky130_fd_sc_hd__a21oi_1 _14648_ (.A1(_05544_),
    .A2(_05552_),
    .B1(_03784_),
    .Y(_05553_));
 sky130_fd_sc_hd__a2111oi_0 _14649_ (.A1(_03784_),
    .A2(_05551_),
    .B1(_05553_),
    .C1(net4073),
    .D1(_03810_),
    .Y(_05554_));
 sky130_fd_sc_hd__a2111oi_1 _14650_ (.A1(_05528_),
    .A2(_05543_),
    .B1(_05550_),
    .C1(_05554_),
    .D1(_03817_),
    .Y(_05555_));
 sky130_fd_sc_hd__a311oi_1 _14651_ (.A1(_05532_),
    .A2(_05537_),
    .A3(_05540_),
    .B1(_05555_),
    .C1(_03824_),
    .Y(_05556_));
 sky130_fd_sc_hd__nand2_1 _14652_ (.A(_03773_),
    .B(_05459_),
    .Y(_05557_));
 sky130_fd_sc_hd__o221ai_2 _14653_ (.A1(_05474_),
    .A2(_05418_),
    .B1(_05535_),
    .B2(_03773_),
    .C1(_05557_),
    .Y(_05558_));
 sky130_fd_sc_hd__a21oi_1 _14654_ (.A1(_05544_),
    .A2(_05437_),
    .B1(_03784_),
    .Y(_05559_));
 sky130_fd_sc_hd__nand2_4 _14655_ (.A(_03784_),
    .B(_03792_),
    .Y(_05560_));
 sky130_fd_sc_hd__o21ai_0 _14656_ (.A1(_11930_[0]),
    .A2(_05560_),
    .B1(_03810_),
    .Y(_05561_));
 sky130_fd_sc_hd__nor2_1 _14657_ (.A(_05559_),
    .B(_05561_),
    .Y(_05562_));
 sky130_fd_sc_hd__a21oi_1 _14658_ (.A1(net4060),
    .A2(_05558_),
    .B1(_05562_),
    .Y(_05563_));
 sky130_fd_sc_hd__nand2_1 _14659_ (.A(_11932_[0]),
    .B(_05413_),
    .Y(_05564_));
 sky130_fd_sc_hd__nor2_1 _14660_ (.A(_11930_[0]),
    .B(_03792_),
    .Y(_05565_));
 sky130_fd_sc_hd__nor2_4 _14661_ (.A(_03778_),
    .B(net4076),
    .Y(_05566_));
 sky130_fd_sc_hd__o21ai_0 _14662_ (.A1(_05565_),
    .A2(_05566_),
    .B1(net4079),
    .Y(_05567_));
 sky130_fd_sc_hd__nor2_1 _14663_ (.A(net4083),
    .B(_03792_),
    .Y(_05568_));
 sky130_fd_sc_hd__nand3_1 _14664_ (.A(net4079),
    .B(_05501_),
    .C(_05547_),
    .Y(_05569_));
 sky130_fd_sc_hd__o311a_1 _14665_ (.A1(net4079),
    .A2(_05568_),
    .A3(_05452_),
    .B1(_05569_),
    .C1(_03809_),
    .X(_05570_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1085 ();
 sky130_fd_sc_hd__a311oi_1 _14667_ (.A1(_03810_),
    .A2(_05564_),
    .A3(_05567_),
    .B1(_05570_),
    .C1(net4073),
    .Y(_05572_));
 sky130_fd_sc_hd__a211oi_1 _14668_ (.A1(net4073),
    .A2(_05563_),
    .B1(_05572_),
    .C1(_05428_),
    .Y(_05573_));
 sky130_fd_sc_hd__a311oi_1 _14669_ (.A1(_05388_),
    .A2(_05517_),
    .A3(_05527_),
    .B1(_05556_),
    .C1(_05573_),
    .Y(_00025_));
 sky130_fd_sc_hd__a21oi_1 _14670_ (.A1(_11930_[0]),
    .A2(_03792_),
    .B1(_05499_),
    .Y(_05574_));
 sky130_fd_sc_hd__o221ai_1 _14671_ (.A1(_11932_[0]),
    .A2(_05460_),
    .B1(_05574_),
    .B2(net4078),
    .C1(_05525_),
    .Y(_05575_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1084 ();
 sky130_fd_sc_hd__mux2i_1 _14673_ (.A0(_05474_),
    .A1(_03776_),
    .S(_03781_),
    .Y(_05577_));
 sky130_fd_sc_hd__nand2_1 _14674_ (.A(net47),
    .B(_11931_[0]),
    .Y(_05578_));
 sky130_fd_sc_hd__o211ai_1 _14675_ (.A1(net46),
    .A2(net47),
    .B1(_05578_),
    .C1(net129),
    .Y(_05579_));
 sky130_fd_sc_hd__o21ai_0 _14676_ (.A1(net129),
    .A2(_05577_),
    .B1(_05579_),
    .Y(_05580_));
 sky130_fd_sc_hd__a21oi_1 _14677_ (.A1(_11946_[0]),
    .A2(_03784_),
    .B1(net4074),
    .Y(_05581_));
 sky130_fd_sc_hd__nand2_4 _14678_ (.A(net4083),
    .B(net4081),
    .Y(_05582_));
 sky130_fd_sc_hd__a22oi_1 _14679_ (.A1(net4074),
    .A2(_05580_),
    .B1(_05581_),
    .B2(_05582_),
    .Y(_05583_));
 sky130_fd_sc_hd__nand2_1 _14680_ (.A(_05528_),
    .B(_05583_),
    .Y(_05584_));
 sky130_fd_sc_hd__o21ai_0 _14681_ (.A1(_05474_),
    .A2(net4078),
    .B1(net4074),
    .Y(_05585_));
 sky130_fd_sc_hd__a21o_1 _14682_ (.A1(_11935_[0]),
    .A2(net4079),
    .B1(_05515_),
    .X(_05586_));
 sky130_fd_sc_hd__a21oi_2 _14683_ (.A1(_03792_),
    .A2(_05586_),
    .B1(_03801_),
    .Y(_05587_));
 sky130_fd_sc_hd__o211ai_1 _14684_ (.A1(_05585_),
    .A2(_05514_),
    .B1(_05587_),
    .C1(_03809_),
    .Y(_05588_));
 sky130_fd_sc_hd__nor2_2 _14685_ (.A(_11937_[0]),
    .B(_03792_),
    .Y(_05589_));
 sky130_fd_sc_hd__nor3_1 _14686_ (.A(_03784_),
    .B(_05566_),
    .C(_05589_),
    .Y(_05590_));
 sky130_fd_sc_hd__a21oi_2 _14687_ (.A1(_05507_),
    .A2(_05552_),
    .B1(net4080),
    .Y(_05591_));
 sky130_fd_sc_hd__o21ai_2 _14688_ (.A1(_05590_),
    .A2(_05591_),
    .B1(_05534_),
    .Y(_05592_));
 sky130_fd_sc_hd__nand4_1 _14689_ (.A(_05575_),
    .B(_05584_),
    .C(_05588_),
    .D(_05592_),
    .Y(_05593_));
 sky130_fd_sc_hd__nand2_4 _14690_ (.A(_11942_[0]),
    .B(net4074),
    .Y(_05594_));
 sky130_fd_sc_hd__a21oi_1 _14691_ (.A1(_05544_),
    .A2(_05594_),
    .B1(net4079),
    .Y(_05595_));
 sky130_fd_sc_hd__o21ai_0 _14692_ (.A1(_05502_),
    .A2(_05595_),
    .B1(_05525_),
    .Y(_05596_));
 sky130_fd_sc_hd__nand2_4 _14693_ (.A(net4082),
    .B(_03792_),
    .Y(_05597_));
 sky130_fd_sc_hd__a311oi_1 _14694_ (.A1(net4079),
    .A2(_05597_),
    .A3(_05594_),
    .B1(_05518_),
    .C1(_05515_),
    .Y(_05598_));
 sky130_fd_sc_hd__nor3_1 _14695_ (.A(_03817_),
    .B(_03824_),
    .C(_05598_),
    .Y(_05599_));
 sky130_fd_sc_hd__nor2_2 _14696_ (.A(_11942_[0]),
    .B(net4074),
    .Y(_05600_));
 sky130_fd_sc_hd__nor3_1 _14697_ (.A(_03784_),
    .B(_05568_),
    .C(net3625),
    .Y(_05601_));
 sky130_fd_sc_hd__nor2_4 _14698_ (.A(_11932_[0]),
    .B(_03792_),
    .Y(_05602_));
 sky130_fd_sc_hd__nor3_1 _14699_ (.A(net4079),
    .B(_05602_),
    .C(_05566_),
    .Y(_05603_));
 sky130_fd_sc_hd__o21ai_0 _14700_ (.A1(_05601_),
    .A2(_05603_),
    .B1(_05528_),
    .Y(_05604_));
 sky130_fd_sc_hd__a21oi_1 _14701_ (.A1(_05433_),
    .A2(_05594_),
    .B1(_03784_),
    .Y(_05605_));
 sky130_fd_sc_hd__nor3_1 _14702_ (.A(net4079),
    .B(_05452_),
    .C(_05602_),
    .Y(_05606_));
 sky130_fd_sc_hd__o21ai_0 _14703_ (.A1(_05605_),
    .A2(_05606_),
    .B1(_05534_),
    .Y(_05607_));
 sky130_fd_sc_hd__nand2_1 _14704_ (.A(net4082),
    .B(net4078),
    .Y(_05608_));
 sky130_fd_sc_hd__o211ai_1 _14705_ (.A1(net4083),
    .A2(net4082),
    .B1(_03792_),
    .C1(_05608_),
    .Y(_05609_));
 sky130_fd_sc_hd__o211ai_1 _14706_ (.A1(_11958_[0]),
    .A2(_03792_),
    .B1(net4073),
    .C1(_05609_),
    .Y(_05610_));
 sky130_fd_sc_hd__o21ai_0 _14707_ (.A1(_11944_[0]),
    .A2(_03792_),
    .B1(_05501_),
    .Y(_05611_));
 sky130_fd_sc_hd__nor2_1 _14708_ (.A(net4078),
    .B(_05611_),
    .Y(_05612_));
 sky130_fd_sc_hd__nor2_2 _14709_ (.A(_03778_),
    .B(_03792_),
    .Y(_05613_));
 sky130_fd_sc_hd__nor3_1 _14710_ (.A(_03784_),
    .B(_05448_),
    .C(_05613_),
    .Y(_05614_));
 sky130_fd_sc_hd__o21ai_0 _14711_ (.A1(_05612_),
    .A2(_05614_),
    .B1(_03801_),
    .Y(_05615_));
 sky130_fd_sc_hd__nand2_2 _14712_ (.A(net4076),
    .B(net4073),
    .Y(_05616_));
 sky130_fd_sc_hd__nand2_1 _14713_ (.A(net4082),
    .B(_05429_),
    .Y(_05617_));
 sky130_fd_sc_hd__o21ai_0 _14714_ (.A1(net4082),
    .A2(net4073),
    .B1(_05507_),
    .Y(_05618_));
 sky130_fd_sc_hd__a211o_1 _14715_ (.A1(net395),
    .A2(net4073),
    .B1(_05449_),
    .C1(net4080),
    .X(_05619_));
 sky130_fd_sc_hd__o21ai_0 _14716_ (.A1(_03784_),
    .A2(_05618_),
    .B1(_05619_),
    .Y(_05620_));
 sky130_fd_sc_hd__nor2_4 _14717_ (.A(net4082),
    .B(net4074),
    .Y(_05621_));
 sky130_fd_sc_hd__o211ai_1 _14718_ (.A1(_05621_),
    .A2(_05514_),
    .B1(_03773_),
    .C1(_03801_),
    .Y(_05622_));
 sky130_fd_sc_hd__o211ai_1 _14719_ (.A1(_11951_[0]),
    .A2(_05616_),
    .B1(_05622_),
    .C1(_03810_),
    .Y(_05623_));
 sky130_fd_sc_hd__a31oi_1 _14720_ (.A1(_05616_),
    .A2(_05617_),
    .A3(_05620_),
    .B1(_05623_),
    .Y(_05624_));
 sky130_fd_sc_hd__a311oi_2 _14721_ (.A1(net4060),
    .A2(_05610_),
    .A3(_05615_),
    .B1(_05428_),
    .C1(_05624_),
    .Y(_05625_));
 sky130_fd_sc_hd__a41oi_2 _14722_ (.A1(_05596_),
    .A2(_05599_),
    .A3(_05604_),
    .A4(_05607_),
    .B1(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__a221oi_1 _14723_ (.A1(_11937_[0]),
    .A2(_05413_),
    .B1(_05611_),
    .B2(net4078),
    .C1(net4060),
    .Y(_05627_));
 sky130_fd_sc_hd__nand2_1 _14724_ (.A(_11949_[0]),
    .B(_03792_),
    .Y(_05628_));
 sky130_fd_sc_hd__nand2_2 _14725_ (.A(_11935_[0]),
    .B(_05423_),
    .Y(_05629_));
 sky130_fd_sc_hd__a21oi_1 _14726_ (.A1(_05628_),
    .A2(_05629_),
    .B1(_03810_),
    .Y(_05630_));
 sky130_fd_sc_hd__nor2_2 _14727_ (.A(_03773_),
    .B(_05460_),
    .Y(_05631_));
 sky130_fd_sc_hd__a221oi_1 _14728_ (.A1(_11940_[0]),
    .A2(_05423_),
    .B1(_05459_),
    .B2(_11930_[0]),
    .C1(_05631_),
    .Y(_05632_));
 sky130_fd_sc_hd__and2_4 _14729_ (.A(_11935_[0]),
    .B(_03784_),
    .X(_05633_));
 sky130_fd_sc_hd__nand2_1 _14730_ (.A(_11956_[0]),
    .B(net4074),
    .Y(_05634_));
 sky130_fd_sc_hd__o311ai_0 _14731_ (.A1(net4074),
    .A2(_05514_),
    .A3(_05633_),
    .B1(_05634_),
    .C1(_03809_),
    .Y(_05635_));
 sky130_fd_sc_hd__o211ai_1 _14732_ (.A1(_03809_),
    .A2(_05632_),
    .B1(_05635_),
    .C1(_03801_),
    .Y(_05636_));
 sky130_fd_sc_hd__o311ai_0 _14733_ (.A1(_03801_),
    .A2(_05627_),
    .A3(_05630_),
    .B1(_05388_),
    .C1(_05636_),
    .Y(_05637_));
 sky130_fd_sc_hd__o311a_4 _14734_ (.A1(_00398_),
    .A2(_03824_),
    .A3(_05593_),
    .B1(_05626_),
    .C1(_05637_),
    .X(_00026_));
 sky130_fd_sc_hd__nor2_1 _14735_ (.A(_11944_[0]),
    .B(net4074),
    .Y(_05638_));
 sky130_fd_sc_hd__nor2_1 _14736_ (.A(_11940_[0]),
    .B(_03792_),
    .Y(_05639_));
 sky130_fd_sc_hd__nand3_1 _14737_ (.A(_03784_),
    .B(_05544_),
    .C(_05394_),
    .Y(_05640_));
 sky130_fd_sc_hd__o311ai_0 _14738_ (.A1(_03784_),
    .A2(_05638_),
    .A3(_05639_),
    .B1(_05640_),
    .C1(_05528_),
    .Y(_05641_));
 sky130_fd_sc_hd__nor2_2 _14739_ (.A(_03784_),
    .B(_03792_),
    .Y(_05642_));
 sky130_fd_sc_hd__nand2_4 _14740_ (.A(_03773_),
    .B(_05642_),
    .Y(_05643_));
 sky130_fd_sc_hd__nor2_1 _14741_ (.A(net4082),
    .B(_03792_),
    .Y(_05644_));
 sky130_fd_sc_hd__nor2_1 _14742_ (.A(net395),
    .B(net4074),
    .Y(_05645_));
 sky130_fd_sc_hd__o21ai_0 _14743_ (.A1(_05644_),
    .A2(_05645_),
    .B1(_03784_),
    .Y(_05646_));
 sky130_fd_sc_hd__a31oi_1 _14744_ (.A1(_05534_),
    .A2(_05643_),
    .A3(_05646_),
    .B1(_00398_),
    .Y(_05647_));
 sky130_fd_sc_hd__nand2_1 _14745_ (.A(_11937_[0]),
    .B(_03784_),
    .Y(_05648_));
 sky130_fd_sc_hd__a21oi_1 _14746_ (.A1(_11932_[0]),
    .A2(net4081),
    .B1(net4074),
    .Y(_05649_));
 sky130_fd_sc_hd__nand2_2 _14747_ (.A(net4073),
    .B(_03810_),
    .Y(_05650_));
 sky130_fd_sc_hd__a21oi_1 _14748_ (.A1(_05648_),
    .A2(_05649_),
    .B1(_05650_),
    .Y(_05651_));
 sky130_fd_sc_hd__o21ai_1 _14749_ (.A1(_03792_),
    .A2(_05580_),
    .B1(_05651_),
    .Y(_05652_));
 sky130_fd_sc_hd__nor2_1 _14750_ (.A(_05474_),
    .B(_05460_),
    .Y(_05653_));
 sky130_fd_sc_hd__nor2_1 _14751_ (.A(net4083),
    .B(_05447_),
    .Y(_05654_));
 sky130_fd_sc_hd__a21oi_1 _14752_ (.A1(_05394_),
    .A2(_05597_),
    .B1(net4079),
    .Y(_05655_));
 sky130_fd_sc_hd__o311ai_0 _14753_ (.A1(_05653_),
    .A2(_05654_),
    .A3(_05655_),
    .B1(_03809_),
    .C1(net4073),
    .Y(_05656_));
 sky130_fd_sc_hd__nand4_1 _14754_ (.A(_05641_),
    .B(_05647_),
    .C(_05652_),
    .D(_05656_),
    .Y(_05657_));
 sky130_fd_sc_hd__nand3_1 _14755_ (.A(_03784_),
    .B(_05493_),
    .C(_05594_),
    .Y(_05658_));
 sky130_fd_sc_hd__o311ai_0 _14756_ (.A1(_03784_),
    .A2(_05449_),
    .A3(_05566_),
    .B1(_05534_),
    .C1(_05658_),
    .Y(_05659_));
 sky130_fd_sc_hd__nand2_1 _14757_ (.A(_11940_[0]),
    .B(_05423_),
    .Y(_05660_));
 sky130_fd_sc_hd__nor2_2 _14758_ (.A(_03773_),
    .B(net4074),
    .Y(_05661_));
 sky130_fd_sc_hd__o21ai_0 _14759_ (.A1(_05475_),
    .A2(_05661_),
    .B1(net4078),
    .Y(_05662_));
 sky130_fd_sc_hd__nand2_2 _14760_ (.A(_03773_),
    .B(_05621_),
    .Y(_05663_));
 sky130_fd_sc_hd__nand4_1 _14761_ (.A(_05660_),
    .B(_05528_),
    .C(_05662_),
    .D(_05663_),
    .Y(_05664_));
 sky130_fd_sc_hd__and2_4 _14762_ (.A(_11930_[0]),
    .B(net4074),
    .X(_05665_));
 sky130_fd_sc_hd__a21oi_1 _14763_ (.A1(_11940_[0]),
    .A2(_03792_),
    .B1(_05665_),
    .Y(_05666_));
 sky130_fd_sc_hd__o21ai_0 _14764_ (.A1(_05449_),
    .A2(_05409_),
    .B1(_03784_),
    .Y(_05667_));
 sky130_fd_sc_hd__o211ai_1 _14765_ (.A1(_03784_),
    .A2(_05666_),
    .B1(_05667_),
    .C1(_05525_),
    .Y(_05668_));
 sky130_fd_sc_hd__a21oi_1 _14766_ (.A1(_11935_[0]),
    .A2(_05413_),
    .B1(_05518_),
    .Y(_05669_));
 sky130_fd_sc_hd__nor2_1 _14767_ (.A(net4083),
    .B(_03778_),
    .Y(_05670_));
 sky130_fd_sc_hd__o21ai_1 _14768_ (.A1(_05471_),
    .A2(_05670_),
    .B1(net4076),
    .Y(_05671_));
 sky130_fd_sc_hd__a21oi_1 _14769_ (.A1(_05669_),
    .A2(_05671_),
    .B1(_03817_),
    .Y(_05672_));
 sky130_fd_sc_hd__nand4_1 _14770_ (.A(_05659_),
    .B(_05664_),
    .C(_05668_),
    .D(_05672_),
    .Y(_05673_));
 sky130_fd_sc_hd__nand2_1 _14771_ (.A(_05657_),
    .B(_05673_),
    .Y(_05674_));
 sky130_fd_sc_hd__nor2_1 _14772_ (.A(_03792_),
    .B(_03810_),
    .Y(_05675_));
 sky130_fd_sc_hd__a22oi_1 _14773_ (.A1(_11946_[0]),
    .A2(_03792_),
    .B1(_05675_),
    .B2(_03778_),
    .Y(_05676_));
 sky130_fd_sc_hd__nor2_2 _14774_ (.A(_03792_),
    .B(_03809_),
    .Y(_05677_));
 sky130_fd_sc_hd__nor3_1 _14775_ (.A(net4081),
    .B(net4074),
    .C(_03810_),
    .Y(_05678_));
 sky130_fd_sc_hd__a21oi_1 _14776_ (.A1(net4081),
    .A2(_05677_),
    .B1(_05678_),
    .Y(_05679_));
 sky130_fd_sc_hd__nor2_1 _14777_ (.A(_11940_[0]),
    .B(net4081),
    .Y(_05680_));
 sky130_fd_sc_hd__a21oi_1 _14778_ (.A1(_05675_),
    .A2(_05680_),
    .B1(net4073),
    .Y(_05681_));
 sky130_fd_sc_hd__o221ai_1 _14779_ (.A1(_03784_),
    .A2(_05676_),
    .B1(_05679_),
    .B2(net396),
    .C1(_05681_),
    .Y(_05682_));
 sky130_fd_sc_hd__a21oi_1 _14780_ (.A1(net4083),
    .A2(_03809_),
    .B1(net4074),
    .Y(_05683_));
 sky130_fd_sc_hd__a21oi_1 _14781_ (.A1(_11932_[0]),
    .A2(_03809_),
    .B1(_05560_),
    .Y(_05684_));
 sky130_fd_sc_hd__a21oi_1 _14782_ (.A1(_03773_),
    .A2(_05675_),
    .B1(_05684_),
    .Y(_05685_));
 sky130_fd_sc_hd__o221ai_1 _14783_ (.A1(_11942_[0]),
    .A2(_03809_),
    .B1(_05683_),
    .B2(_03784_),
    .C1(_05685_),
    .Y(_05686_));
 sky130_fd_sc_hd__a21oi_2 _14784_ (.A1(_03773_),
    .A2(_03784_),
    .B1(_05661_),
    .Y(_05687_));
 sky130_fd_sc_hd__a32oi_1 _14785_ (.A1(net395),
    .A2(_03809_),
    .A3(_05687_),
    .B1(_05677_),
    .B2(_05471_),
    .Y(_05688_));
 sky130_fd_sc_hd__nand3_1 _14786_ (.A(net4073),
    .B(_05686_),
    .C(_05688_),
    .Y(_05689_));
 sky130_fd_sc_hd__o21ai_0 _14787_ (.A1(_03784_),
    .A2(_05644_),
    .B1(net4083),
    .Y(_05690_));
 sky130_fd_sc_hd__o221ai_1 _14788_ (.A1(_11944_[0]),
    .A2(_05460_),
    .B1(_05418_),
    .B2(_03778_),
    .C1(_05690_),
    .Y(_05691_));
 sky130_fd_sc_hd__nor2_4 _14789_ (.A(_05449_),
    .B(_05600_),
    .Y(_05692_));
 sky130_fd_sc_hd__nor2_2 _14790_ (.A(_03784_),
    .B(_05692_),
    .Y(_05693_));
 sky130_fd_sc_hd__a31oi_2 _14791_ (.A1(_03784_),
    .A2(_05393_),
    .A3(_05552_),
    .B1(_05693_),
    .Y(_05694_));
 sky130_fd_sc_hd__o211ai_1 _14792_ (.A1(_11942_[0]),
    .A2(net4081),
    .B1(_03792_),
    .C1(_05582_),
    .Y(_05695_));
 sky130_fd_sc_hd__nand2_1 _14793_ (.A(_11932_[0]),
    .B(_03784_),
    .Y(_05696_));
 sky130_fd_sc_hd__nor2_1 _14794_ (.A(_05471_),
    .B(_05442_),
    .Y(_05697_));
 sky130_fd_sc_hd__a221oi_1 _14795_ (.A1(_05539_),
    .A2(_05695_),
    .B1(_05696_),
    .B2(_05697_),
    .C1(_05483_),
    .Y(_05698_));
 sky130_fd_sc_hd__a221o_4 _14796_ (.A1(_05506_),
    .A2(_05691_),
    .B1(_05694_),
    .B2(_05504_),
    .C1(_05698_),
    .X(_05699_));
 sky130_fd_sc_hd__a311oi_1 _14797_ (.A1(_03817_),
    .A2(_05682_),
    .A3(_05689_),
    .B1(net3626),
    .C1(_05699_),
    .Y(_05700_));
 sky130_fd_sc_hd__a21oi_1 _14798_ (.A1(_03824_),
    .A2(_05674_),
    .B1(_05700_),
    .Y(_00027_));
 sky130_fd_sc_hd__a31oi_2 _14799_ (.A1(net395),
    .A2(_03784_),
    .A3(_03792_),
    .B1(_05665_),
    .Y(_05701_));
 sky130_fd_sc_hd__nand2_2 _14800_ (.A(_03778_),
    .B(net4078),
    .Y(_05702_));
 sky130_fd_sc_hd__nand2_4 _14801_ (.A(net4083),
    .B(_03777_),
    .Y(_05703_));
 sky130_fd_sc_hd__a31oi_1 _14802_ (.A1(net4074),
    .A2(_05702_),
    .A3(_05703_),
    .B1(_05631_),
    .Y(_05704_));
 sky130_fd_sc_hd__o21ai_1 _14803_ (.A1(_11942_[0]),
    .A2(_05687_),
    .B1(_05704_),
    .Y(_05705_));
 sky130_fd_sc_hd__o21ai_0 _14804_ (.A1(_05420_),
    .A2(_05566_),
    .B1(net4080),
    .Y(_05706_));
 sky130_fd_sc_hd__a221oi_1 _14805_ (.A1(net4060),
    .A2(_05705_),
    .B1(_05706_),
    .B2(_05414_),
    .C1(net4073),
    .Y(_05707_));
 sky130_fd_sc_hd__a21oi_1 _14806_ (.A1(_05433_),
    .A2(_05547_),
    .B1(net4080),
    .Y(_05708_));
 sky130_fd_sc_hd__nand2_1 _14807_ (.A(net4078),
    .B(net4076),
    .Y(_05709_));
 sky130_fd_sc_hd__o22ai_1 _14808_ (.A1(_11946_[0]),
    .A2(_05709_),
    .B1(_05597_),
    .B2(net4083),
    .Y(_05710_));
 sky130_fd_sc_hd__nor3_1 _14809_ (.A(_05518_),
    .B(_05708_),
    .C(_05710_),
    .Y(_05711_));
 sky130_fd_sc_hd__a2111oi_0 _14810_ (.A1(_05525_),
    .A2(_05701_),
    .B1(_05707_),
    .C1(net3626),
    .D1(_05711_),
    .Y(_05712_));
 sky130_fd_sc_hd__o211ai_1 _14811_ (.A1(_11935_[0]),
    .A2(_03784_),
    .B1(_05485_),
    .C1(_05429_),
    .Y(_05713_));
 sky130_fd_sc_hd__o21ai_0 _14812_ (.A1(_05621_),
    .A2(_05589_),
    .B1(net4073),
    .Y(_05714_));
 sky130_fd_sc_hd__o21ai_0 _14813_ (.A1(_11932_[0]),
    .A2(_05442_),
    .B1(_05714_),
    .Y(_05715_));
 sky130_fd_sc_hd__and3_1 _14814_ (.A(_03801_),
    .B(_05589_),
    .C(_05696_),
    .X(_05716_));
 sky130_fd_sc_hd__a221oi_1 _14815_ (.A1(net4073),
    .A2(_05404_),
    .B1(_05715_),
    .B2(_03784_),
    .C1(_05716_),
    .Y(_05717_));
 sky130_fd_sc_hd__o211ai_1 _14816_ (.A1(_11942_[0]),
    .A2(_03784_),
    .B1(_05528_),
    .C1(_05521_),
    .Y(_05718_));
 sky130_fd_sc_hd__nand3_1 _14817_ (.A(net4080),
    .B(_05507_),
    .C(_05552_),
    .Y(_05719_));
 sky130_fd_sc_hd__o211ai_1 _14818_ (.A1(net4080),
    .A2(_05692_),
    .B1(_05719_),
    .C1(_05525_),
    .Y(_05720_));
 sky130_fd_sc_hd__a31oi_1 _14819_ (.A1(net3626),
    .A2(_05718_),
    .A3(_05720_),
    .B1(_00398_),
    .Y(_05721_));
 sky130_fd_sc_hd__a41oi_1 _14820_ (.A1(net4060),
    .A2(_03817_),
    .A3(_05713_),
    .A4(_05717_),
    .B1(_05721_),
    .Y(_05722_));
 sky130_fd_sc_hd__a21oi_1 _14821_ (.A1(_11942_[0]),
    .A2(_03792_),
    .B1(net4080),
    .Y(_05723_));
 sky130_fd_sc_hd__o21ai_0 _14822_ (.A1(_05411_),
    .A2(_05723_),
    .B1(_03801_),
    .Y(_05724_));
 sky130_fd_sc_hd__a311oi_1 _14823_ (.A1(_03784_),
    .A2(_05547_),
    .A3(_05597_),
    .B1(_03801_),
    .C1(_05471_),
    .Y(_05725_));
 sky130_fd_sc_hd__nor3b_1 _14824_ (.A(_05503_),
    .B(_05725_),
    .C_N(net3626),
    .Y(_05726_));
 sky130_fd_sc_hd__o21ai_0 _14825_ (.A1(net4080),
    .A2(_05602_),
    .B1(_05643_),
    .Y(_05727_));
 sky130_fd_sc_hd__nand3b_1 _14826_ (.A_N(_05452_),
    .B(_05547_),
    .C(net4080),
    .Y(_05728_));
 sky130_fd_sc_hd__a21oi_2 _14827_ (.A1(_05536_),
    .A2(_05728_),
    .B1(net4073),
    .Y(_05729_));
 sky130_fd_sc_hd__a21oi_1 _14828_ (.A1(net4073),
    .A2(_05727_),
    .B1(_05729_),
    .Y(_05730_));
 sky130_fd_sc_hd__nor3_1 _14829_ (.A(net3626),
    .B(_05483_),
    .C(_05730_),
    .Y(_05731_));
 sky130_fd_sc_hd__a21oi_1 _14830_ (.A1(_05724_),
    .A2(_05726_),
    .B1(_05731_),
    .Y(_05732_));
 sky130_fd_sc_hd__o21ai_0 _14831_ (.A1(_03778_),
    .A2(_05413_),
    .B1(_05663_),
    .Y(_05733_));
 sky130_fd_sc_hd__nand3_1 _14832_ (.A(net4073),
    .B(_05643_),
    .C(_05733_),
    .Y(_05734_));
 sky130_fd_sc_hd__nand3_1 _14833_ (.A(_11944_[0]),
    .B(_03784_),
    .C(_03792_),
    .Y(_05735_));
 sky130_fd_sc_hd__a21oi_1 _14834_ (.A1(_05702_),
    .A2(_05735_),
    .B1(net4073),
    .Y(_05736_));
 sky130_fd_sc_hd__a311oi_1 _14835_ (.A1(_03772_),
    .A2(net4074),
    .A3(_05464_),
    .B1(_05483_),
    .C1(_05736_),
    .Y(_05737_));
 sky130_fd_sc_hd__a21o_1 _14836_ (.A1(_11937_[0]),
    .A2(net4078),
    .B1(_05465_),
    .X(_05738_));
 sky130_fd_sc_hd__a21oi_1 _14837_ (.A1(net4074),
    .A2(_05738_),
    .B1(_05489_),
    .Y(_05739_));
 sky130_fd_sc_hd__nor3_1 _14838_ (.A(net4080),
    .B(net4073),
    .C(_05551_),
    .Y(_05740_));
 sky130_fd_sc_hd__nor4_1 _14839_ (.A(net3626),
    .B(_05503_),
    .C(_05739_),
    .D(_05740_),
    .Y(_05741_));
 sky130_fd_sc_hd__a31oi_1 _14840_ (.A1(net3626),
    .A2(_05734_),
    .A3(_05737_),
    .B1(_05741_),
    .Y(_05742_));
 sky130_fd_sc_hd__o211ai_1 _14841_ (.A1(_05712_),
    .A2(_05722_),
    .B1(_05732_),
    .C1(_05742_),
    .Y(_00028_));
 sky130_fd_sc_hd__a21oi_1 _14842_ (.A1(net4079),
    .A2(_05437_),
    .B1(_05409_),
    .Y(_05743_));
 sky130_fd_sc_hd__nor2_1 _14843_ (.A(_11942_[0]),
    .B(_03792_),
    .Y(_05744_));
 sky130_fd_sc_hd__nand3_1 _14844_ (.A(net4080),
    .B(_05401_),
    .C(_05433_),
    .Y(_05745_));
 sky130_fd_sc_hd__o311ai_0 _14845_ (.A1(net4080),
    .A2(_05452_),
    .A3(_05744_),
    .B1(_05745_),
    .C1(_03810_),
    .Y(_05746_));
 sky130_fd_sc_hd__o211ai_1 _14846_ (.A1(_03810_),
    .A2(_05743_),
    .B1(_05746_),
    .C1(_03801_),
    .Y(_05747_));
 sky130_fd_sc_hd__a211oi_1 _14847_ (.A1(net4083),
    .A2(_05413_),
    .B1(_05518_),
    .C1(_05693_),
    .Y(_05748_));
 sky130_fd_sc_hd__o21ai_0 _14848_ (.A1(_05498_),
    .A2(_05613_),
    .B1(_03784_),
    .Y(_05749_));
 sky130_fd_sc_hd__and3_1 _14849_ (.A(_05453_),
    .B(_05525_),
    .C(_05749_),
    .X(_05750_));
 sky130_fd_sc_hd__nor3_1 _14850_ (.A(_05428_),
    .B(_05748_),
    .C(_05750_),
    .Y(_05751_));
 sky130_fd_sc_hd__o22ai_1 _14851_ (.A1(_03778_),
    .A2(_05441_),
    .B1(_05442_),
    .B2(_05703_),
    .Y(_05752_));
 sky130_fd_sc_hd__nand2_1 _14852_ (.A(_05429_),
    .B(_05538_),
    .Y(_05753_));
 sky130_fd_sc_hd__nor2_1 _14853_ (.A(_03778_),
    .B(_03801_),
    .Y(_05754_));
 sky130_fd_sc_hd__o21ai_0 _14854_ (.A1(_05423_),
    .A2(_05754_),
    .B1(_03773_),
    .Y(_05755_));
 sky130_fd_sc_hd__o211ai_1 _14855_ (.A1(_05464_),
    .A2(_05616_),
    .B1(_05753_),
    .C1(_05755_),
    .Y(_05756_));
 sky130_fd_sc_hd__o21ai_0 _14856_ (.A1(_05752_),
    .A2(_05756_),
    .B1(_03810_),
    .Y(_05757_));
 sky130_fd_sc_hd__nand2_1 _14857_ (.A(_11946_[0]),
    .B(net4074),
    .Y(_05758_));
 sky130_fd_sc_hd__a21oi_1 _14858_ (.A1(_05501_),
    .A2(_05758_),
    .B1(net4078),
    .Y(_05759_));
 sky130_fd_sc_hd__a21oi_1 _14859_ (.A1(_03778_),
    .A2(_05642_),
    .B1(_05759_),
    .Y(_05760_));
 sky130_fd_sc_hd__and2_0 _14860_ (.A(_11932_[0]),
    .B(net4074),
    .X(_05761_));
 sky130_fd_sc_hd__o21ai_0 _14861_ (.A1(_05638_),
    .A2(_05761_),
    .B1(_03784_),
    .Y(_05762_));
 sky130_fd_sc_hd__nor2_1 _14862_ (.A(_03801_),
    .B(_05461_),
    .Y(_05763_));
 sky130_fd_sc_hd__a221o_1 _14863_ (.A1(_03801_),
    .A2(_05760_),
    .B1(_05762_),
    .B2(_05763_),
    .C1(_03810_),
    .X(_05764_));
 sky130_fd_sc_hd__nor2_1 _14864_ (.A(net4074),
    .B(_03810_),
    .Y(_05765_));
 sky130_fd_sc_hd__o21ai_2 _14865_ (.A1(_03809_),
    .A2(_05433_),
    .B1(_05477_),
    .Y(_05766_));
 sky130_fd_sc_hd__a222oi_1 _14866_ (.A1(_11940_[0]),
    .A2(_05765_),
    .B1(_05633_),
    .B2(_05677_),
    .C1(_05766_),
    .C2(net4078),
    .Y(_05767_));
 sky130_fd_sc_hd__o21ai_0 _14867_ (.A1(_05448_),
    .A2(_05761_),
    .B1(_03784_),
    .Y(_05768_));
 sky130_fd_sc_hd__o311ai_0 _14868_ (.A1(_03784_),
    .A2(_05475_),
    .A3(_05645_),
    .B1(_05768_),
    .C1(_03809_),
    .Y(_05769_));
 sky130_fd_sc_hd__o2bb2ai_1 _14869_ (.A1_N(net4074),
    .A2_N(_05648_),
    .B1(_05560_),
    .B2(_11932_[0]),
    .Y(_05770_));
 sky130_fd_sc_hd__a21oi_1 _14870_ (.A1(_03810_),
    .A2(_05770_),
    .B1(net4073),
    .Y(_05771_));
 sky130_fd_sc_hd__a221oi_1 _14871_ (.A1(net4073),
    .A2(_05767_),
    .B1(_05769_),
    .B2(_05771_),
    .C1(_03824_),
    .Y(_05772_));
 sky130_fd_sc_hd__a31oi_1 _14872_ (.A1(net3626),
    .A2(_05757_),
    .A3(_05764_),
    .B1(_05772_),
    .Y(_05773_));
 sky130_fd_sc_hd__nor2_1 _14873_ (.A(_00398_),
    .B(_05773_),
    .Y(_05774_));
 sky130_fd_sc_hd__nor3_1 _14874_ (.A(net4079),
    .B(_05409_),
    .C(_05744_),
    .Y(_05775_));
 sky130_fd_sc_hd__a31oi_1 _14875_ (.A1(net4079),
    .A2(_05447_),
    .A3(_05544_),
    .B1(_05775_),
    .Y(_05776_));
 sky130_fd_sc_hd__nor2_1 _14876_ (.A(net4083),
    .B(_05613_),
    .Y(_05777_));
 sky130_fd_sc_hd__a21oi_1 _14877_ (.A1(net4083),
    .A2(_05642_),
    .B1(_05777_),
    .Y(_05778_));
 sky130_fd_sc_hd__o211ai_1 _14878_ (.A1(_11930_[0]),
    .A2(_05709_),
    .B1(_05534_),
    .C1(_05768_),
    .Y(_05779_));
 sky130_fd_sc_hd__o21ai_0 _14879_ (.A1(_05650_),
    .A2(_05778_),
    .B1(_05779_),
    .Y(_05780_));
 sky130_fd_sc_hd__a21oi_1 _14880_ (.A1(_05582_),
    .A2(_05648_),
    .B1(_03792_),
    .Y(_05781_));
 sky130_fd_sc_hd__nor3_1 _14881_ (.A(_03810_),
    .B(_05489_),
    .C(_05781_),
    .Y(_05782_));
 sky130_fd_sc_hd__a211oi_1 _14882_ (.A1(_05528_),
    .A2(_05776_),
    .B1(_05780_),
    .C1(_05782_),
    .Y(_05783_));
 sky130_fd_sc_hd__nor3_1 _14883_ (.A(_03817_),
    .B(net3626),
    .C(_05783_),
    .Y(_05784_));
 sky130_fd_sc_hd__a211oi_1 _14884_ (.A1(_05747_),
    .A2(_05751_),
    .B1(_05774_),
    .C1(_05784_),
    .Y(_00029_));
 sky130_fd_sc_hd__a21oi_1 _14885_ (.A1(_03784_),
    .A2(_05393_),
    .B1(_03778_),
    .Y(_05785_));
 sky130_fd_sc_hd__nand2_1 _14886_ (.A(_05506_),
    .B(_05629_),
    .Y(_05786_));
 sky130_fd_sc_hd__nor3_1 _14887_ (.A(_05631_),
    .B(_05785_),
    .C(_05786_),
    .Y(_05787_));
 sky130_fd_sc_hd__o21a_1 _14888_ (.A1(_11935_[0]),
    .A2(net4078),
    .B1(_05697_),
    .X(_05788_));
 sky130_fd_sc_hd__a221oi_1 _14889_ (.A1(_03773_),
    .A2(_05413_),
    .B1(_05692_),
    .B2(net4080),
    .C1(_03801_),
    .Y(_05789_));
 sky130_fd_sc_hd__a2111oi_0 _14890_ (.A1(_11954_[0]),
    .A2(_05429_),
    .B1(_05788_),
    .C1(_05789_),
    .D1(_05483_),
    .Y(_05790_));
 sky130_fd_sc_hd__o31ai_1 _14891_ (.A1(_11932_[0]),
    .A2(_03784_),
    .A3(_03792_),
    .B1(_05663_),
    .Y(_05791_));
 sky130_fd_sc_hd__o21ai_0 _14892_ (.A1(_03773_),
    .A2(net4078),
    .B1(_05504_),
    .Y(_05792_));
 sky130_fd_sc_hd__nor2_1 _14893_ (.A(_05791_),
    .B(_05792_),
    .Y(_05793_));
 sky130_fd_sc_hd__nor4_1 _14894_ (.A(net3626),
    .B(_05787_),
    .C(_05790_),
    .D(_05793_),
    .Y(_05794_));
 sky130_fd_sc_hd__a21oi_1 _14895_ (.A1(_05493_),
    .A2(_05394_),
    .B1(net4078),
    .Y(_05795_));
 sky130_fd_sc_hd__o21ai_0 _14896_ (.A1(_05461_),
    .A2(_05795_),
    .B1(_03801_),
    .Y(_05796_));
 sky130_fd_sc_hd__nand2_1 _14897_ (.A(_11942_[0]),
    .B(_03784_),
    .Y(_05797_));
 sky130_fd_sc_hd__nand3_1 _14898_ (.A(net4074),
    .B(_05608_),
    .C(_05797_),
    .Y(_05798_));
 sky130_fd_sc_hd__o211ai_1 _14899_ (.A1(_11950_[0]),
    .A2(net4074),
    .B1(net4073),
    .C1(_05798_),
    .Y(_05799_));
 sky130_fd_sc_hd__a21oi_1 _14900_ (.A1(_11940_[0]),
    .A2(net4074),
    .B1(net3625),
    .Y(_05800_));
 sky130_fd_sc_hd__o221ai_1 _14901_ (.A1(net4082),
    .A2(_05460_),
    .B1(_05800_),
    .B2(net4078),
    .C1(_03801_),
    .Y(_05801_));
 sky130_fd_sc_hd__nor2_1 _14902_ (.A(_03810_),
    .B(_05587_),
    .Y(_05802_));
 sky130_fd_sc_hd__a32oi_1 _14903_ (.A1(_03810_),
    .A2(_05796_),
    .A3(_05799_),
    .B1(_05801_),
    .B2(_05802_),
    .Y(_05803_));
 sky130_fd_sc_hd__nand2_2 _14904_ (.A(_03817_),
    .B(_05803_),
    .Y(_05804_));
 sky130_fd_sc_hd__nand2_1 _14905_ (.A(_03817_),
    .B(net3626),
    .Y(_05805_));
 sky130_fd_sc_hd__nor2_1 _14906_ (.A(_11935_[0]),
    .B(_05460_),
    .Y(_05806_));
 sky130_fd_sc_hd__o21ai_1 _14907_ (.A1(net396),
    .A2(_05418_),
    .B1(_05557_),
    .Y(_05807_));
 sky130_fd_sc_hd__o21ai_0 _14908_ (.A1(_05806_),
    .A2(_05807_),
    .B1(_03809_),
    .Y(_05808_));
 sky130_fd_sc_hd__o21ai_0 _14909_ (.A1(_05409_),
    .A2(_05411_),
    .B1(_03784_),
    .Y(_05809_));
 sky130_fd_sc_hd__o311ai_2 _14910_ (.A1(_03784_),
    .A2(_05449_),
    .A3(_05566_),
    .B1(_05809_),
    .C1(_03810_),
    .Y(_05810_));
 sky130_fd_sc_hd__o21ai_0 _14911_ (.A1(_05621_),
    .A2(_05639_),
    .B1(_03784_),
    .Y(_05811_));
 sky130_fd_sc_hd__nand3b_1 _14912_ (.A_N(_05806_),
    .B(_05811_),
    .C(_03809_),
    .Y(_05812_));
 sky130_fd_sc_hd__o21ai_0 _14913_ (.A1(net395),
    .A2(_03784_),
    .B1(net4074),
    .Y(_05813_));
 sky130_fd_sc_hd__o221ai_1 _14914_ (.A1(_11949_[0]),
    .A2(net4074),
    .B1(_05633_),
    .B2(_05813_),
    .C1(_03810_),
    .Y(_05814_));
 sky130_fd_sc_hd__a21oi_1 _14915_ (.A1(_05812_),
    .A2(_05814_),
    .B1(net4073),
    .Y(_05815_));
 sky130_fd_sc_hd__a31oi_1 _14916_ (.A1(net4073),
    .A2(_05808_),
    .A3(_05810_),
    .B1(_05815_),
    .Y(_05816_));
 sky130_fd_sc_hd__a31oi_1 _14917_ (.A1(_11946_[0]),
    .A2(_03810_),
    .A3(_05413_),
    .B1(net4073),
    .Y(_05817_));
 sky130_fd_sc_hd__nor2_1 _14918_ (.A(_05443_),
    .B(_05460_),
    .Y(_05818_));
 sky130_fd_sc_hd__o21ai_0 _14919_ (.A1(_05807_),
    .A2(_05818_),
    .B1(_03809_),
    .Y(_05819_));
 sky130_fd_sc_hd__nor3_1 _14920_ (.A(_03784_),
    .B(_03809_),
    .C(net3625),
    .Y(_05820_));
 sky130_fd_sc_hd__nand2_1 _14921_ (.A(_05547_),
    .B(_05820_),
    .Y(_05821_));
 sky130_fd_sc_hd__a21boi_0 _14922_ (.A1(_11932_[0]),
    .A2(net4081),
    .B1_N(_05797_),
    .Y(_05822_));
 sky130_fd_sc_hd__o21ai_0 _14923_ (.A1(_03792_),
    .A2(_05822_),
    .B1(net4073),
    .Y(_05823_));
 sky130_fd_sc_hd__nand2_1 _14924_ (.A(_03792_),
    .B(_05486_),
    .Y(_05824_));
 sky130_fd_sc_hd__a21oi_1 _14925_ (.A1(_11930_[0]),
    .A2(_03784_),
    .B1(_05824_),
    .Y(_05825_));
 sky130_fd_sc_hd__nor2_1 _14926_ (.A(_03778_),
    .B(_05661_),
    .Y(_05826_));
 sky130_fd_sc_hd__a21oi_1 _14927_ (.A1(_03778_),
    .A2(_05413_),
    .B1(_05826_),
    .Y(_05827_));
 sky130_fd_sc_hd__o32ai_1 _14928_ (.A1(_03810_),
    .A2(_05823_),
    .A3(_05825_),
    .B1(_05827_),
    .B2(_05650_),
    .Y(_05828_));
 sky130_fd_sc_hd__a31oi_1 _14929_ (.A1(_05817_),
    .A2(_05819_),
    .A3(_05821_),
    .B1(_05828_),
    .Y(_05829_));
 sky130_fd_sc_hd__o22ai_2 _14930_ (.A1(_05805_),
    .A2(_05816_),
    .B1(_05829_),
    .B2(_05428_),
    .Y(_05830_));
 sky130_fd_sc_hd__a21oi_4 _14931_ (.A1(net3569),
    .A2(_05804_),
    .B1(_05830_),
    .Y(_00030_));
 sky130_fd_sc_hd__or3_1 _14932_ (.A(_03784_),
    .B(_05499_),
    .C(_05452_),
    .X(_05831_));
 sky130_fd_sc_hd__a2111oi_0 _14933_ (.A1(_11951_[0]),
    .A2(net4077),
    .B1(_03810_),
    .C1(_05461_),
    .D1(_05542_),
    .Y(_05832_));
 sky130_fd_sc_hd__a31oi_1 _14934_ (.A1(_03810_),
    .A2(_05536_),
    .A3(_05831_),
    .B1(_05832_),
    .Y(_05833_));
 sky130_fd_sc_hd__nor2_1 _14935_ (.A(_11960_[0]),
    .B(net4076),
    .Y(_05834_));
 sky130_fd_sc_hd__a211oi_1 _14936_ (.A1(_11942_[0]),
    .A2(net4078),
    .B1(_03792_),
    .C1(_05465_),
    .Y(_05835_));
 sky130_fd_sc_hd__nand3_1 _14937_ (.A(_11946_[0]),
    .B(_03784_),
    .C(net4076),
    .Y(_05836_));
 sky130_fd_sc_hd__o21ai_0 _14938_ (.A1(_11930_[0]),
    .A2(net4076),
    .B1(_05836_),
    .Y(_05837_));
 sky130_fd_sc_hd__nand2_1 _14939_ (.A(_05525_),
    .B(_05837_),
    .Y(_05838_));
 sky130_fd_sc_hd__o311ai_0 _14940_ (.A1(_05518_),
    .A2(_05834_),
    .A3(_05835_),
    .B1(_05838_),
    .C1(_05388_),
    .Y(_05839_));
 sky130_fd_sc_hd__a21oi_1 _14941_ (.A1(_03801_),
    .A2(_05833_),
    .B1(_05839_),
    .Y(_05840_));
 sky130_fd_sc_hd__nand2_1 _14942_ (.A(_03777_),
    .B(_05459_),
    .Y(_05841_));
 sky130_fd_sc_hd__o221ai_1 _14943_ (.A1(_11930_[0]),
    .A2(_05418_),
    .B1(_05535_),
    .B2(_03773_),
    .C1(_05841_),
    .Y(_05842_));
 sky130_fd_sc_hd__a21oi_1 _14944_ (.A1(_03792_),
    .A2(_05464_),
    .B1(_03772_),
    .Y(_05843_));
 sky130_fd_sc_hd__a21oi_1 _14945_ (.A1(_05485_),
    .A2(_05661_),
    .B1(_05843_),
    .Y(_05844_));
 sky130_fd_sc_hd__a22oi_1 _14946_ (.A1(_05525_),
    .A2(_05842_),
    .B1(_05844_),
    .B2(_05528_),
    .Y(_05845_));
 sky130_fd_sc_hd__nor2_2 _14947_ (.A(_00398_),
    .B(_05845_),
    .Y(_05846_));
 sky130_fd_sc_hd__nand2_1 _14948_ (.A(_05418_),
    .B(_05441_),
    .Y(_05847_));
 sky130_fd_sc_hd__a211oi_1 _14949_ (.A1(_11935_[0]),
    .A2(_05429_),
    .B1(_05475_),
    .C1(_03784_),
    .Y(_05848_));
 sky130_fd_sc_hd__a21oi_1 _14950_ (.A1(_03784_),
    .A2(_03801_),
    .B1(_05848_),
    .Y(_05849_));
 sky130_fd_sc_hd__a211oi_1 _14951_ (.A1(_11930_[0]),
    .A2(_05847_),
    .B1(_05849_),
    .C1(_05470_),
    .Y(_05850_));
 sky130_fd_sc_hd__a21oi_1 _14952_ (.A1(_05582_),
    .A2(_05485_),
    .B1(net4075),
    .Y(_05851_));
 sky130_fd_sc_hd__nor2_1 _14953_ (.A(_05823_),
    .B(_05851_),
    .Y(_05852_));
 sky130_fd_sc_hd__o22ai_1 _14954_ (.A1(_11932_[0]),
    .A2(_05460_),
    .B1(_05418_),
    .B2(net4083),
    .Y(_05853_));
 sky130_fd_sc_hd__a21oi_1 _14955_ (.A1(_05474_),
    .A2(_05459_),
    .B1(_05853_),
    .Y(_05854_));
 sky130_fd_sc_hd__nor2_1 _14956_ (.A(net4073),
    .B(_05854_),
    .Y(_05855_));
 sky130_fd_sc_hd__nor2_1 _14957_ (.A(net4080),
    .B(_05529_),
    .Y(_05856_));
 sky130_fd_sc_hd__o21ai_0 _14958_ (.A1(_05602_),
    .A2(_05621_),
    .B1(net4080),
    .Y(_05857_));
 sky130_fd_sc_hd__o211ai_1 _14959_ (.A1(_11942_[0]),
    .A2(_05560_),
    .B1(_05857_),
    .C1(net4073),
    .Y(_05858_));
 sky130_fd_sc_hd__o31a_1 _14960_ (.A1(net4073),
    .A2(_05404_),
    .A3(_05856_),
    .B1(_05858_),
    .X(_05859_));
 sky130_fd_sc_hd__o32ai_2 _14961_ (.A1(_05483_),
    .A2(_05852_),
    .A3(_05855_),
    .B1(_05503_),
    .B2(_05859_),
    .Y(_05860_));
 sky130_fd_sc_hd__nor4_4 _14962_ (.A(net3626),
    .B(_05846_),
    .C(_05850_),
    .D(_05860_),
    .Y(_05861_));
 sky130_fd_sc_hd__nor3_1 _14963_ (.A(net4079),
    .B(_05665_),
    .C(net3625),
    .Y(_05862_));
 sky130_fd_sc_hd__a311oi_1 _14964_ (.A1(net4079),
    .A2(_05494_),
    .A3(_05433_),
    .B1(_05862_),
    .C1(_03809_),
    .Y(_05863_));
 sky130_fd_sc_hd__a31oi_2 _14965_ (.A1(_03792_),
    .A2(_05702_),
    .A3(_05703_),
    .B1(_05589_),
    .Y(_05864_));
 sky130_fd_sc_hd__nor2_1 _14966_ (.A(_03810_),
    .B(_05864_),
    .Y(_05865_));
 sky130_fd_sc_hd__nor3_1 _14967_ (.A(net4073),
    .B(_05863_),
    .C(_05865_),
    .Y(_05866_));
 sky130_fd_sc_hd__nand2_1 _14968_ (.A(_03784_),
    .B(_05666_),
    .Y(_05867_));
 sky130_fd_sc_hd__nor2_1 _14969_ (.A(_11944_[0]),
    .B(_03784_),
    .Y(_05868_));
 sky130_fd_sc_hd__a311oi_1 _14970_ (.A1(_03784_),
    .A2(_05541_),
    .A3(_05597_),
    .B1(_05868_),
    .C1(_03810_),
    .Y(_05869_));
 sky130_fd_sc_hd__a311oi_1 _14971_ (.A1(_03810_),
    .A2(_05569_),
    .A3(_05867_),
    .B1(_05869_),
    .C1(_03801_),
    .Y(_05870_));
 sky130_fd_sc_hd__nor3_1 _14972_ (.A(_05428_),
    .B(_05866_),
    .C(_05870_),
    .Y(_05871_));
 sky130_fd_sc_hd__nor3_1 _14973_ (.A(_05840_),
    .B(_05861_),
    .C(_05871_),
    .Y(_00031_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1082 ();
 sky130_fd_sc_hd__xnor2_1 _14976_ (.A(net4229),
    .B(\sa00_sr[0] ),
    .Y(_05874_));
 sky130_fd_sc_hd__xor2_1 _14977_ (.A(\sa20_sr[1] ),
    .B(\sa30_sr[1] ),
    .X(_05875_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1081 ();
 sky130_fd_sc_hd__xor3_1 _14979_ (.A(\sa10_sr[7] ),
    .B(net4220),
    .C(\sa10_sr[1] ),
    .X(_05877_));
 sky130_fd_sc_hd__xnor3_1 _14980_ (.A(_05874_),
    .B(net4122),
    .C(_05877_),
    .X(_05878_));
 sky130_fd_sc_hd__clkinv_16 _14981_ (.A(ld_r),
    .Y(_05879_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1079 ();
 sky130_fd_sc_hd__mux2i_2 _14984_ (.A0(\text_in_r[121] ),
    .A1(_05878_),
    .S(net4119),
    .Y(_05882_));
 sky130_fd_sc_hd__xor2_4 _14985_ (.A(net4169),
    .B(_05882_),
    .X(_05883_));
 sky130_fd_sc_hd__clkinv_8 _14986_ (.A(_05883_),
    .Y(_05884_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1078 ();
 sky130_fd_sc_hd__xor2_1 _14988_ (.A(\sa10_sr[0] ),
    .B(\sa20_sr[0] ),
    .X(_05885_));
 sky130_fd_sc_hd__xnor3_1 _14989_ (.A(net4229),
    .B(net4216),
    .C(\sa30_sr[0] ),
    .X(_05886_));
 sky130_fd_sc_hd__xnor2_1 _14990_ (.A(net4110),
    .B(_05886_),
    .Y(_05887_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1077 ();
 sky130_fd_sc_hd__mux2i_2 _14992_ (.A0(\text_in_r[120] ),
    .A1(_05887_),
    .S(net4119),
    .Y(_05889_));
 sky130_fd_sc_hd__xor2_4 _14993_ (.A(net4170),
    .B(_05889_),
    .X(_05890_));
 sky130_fd_sc_hd__inv_16 _14994_ (.A(_05890_),
    .Y(_05891_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1075 ();
 sky130_fd_sc_hd__xnor3_1 _14997_ (.A(\sa00_sr[1] ),
    .B(net4219),
    .C(\sa20_sr[2] ),
    .X(_05893_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1074 ();
 sky130_fd_sc_hd__xor2_1 _14999_ (.A(\sa10_sr[1] ),
    .B(\sa30_sr[2] ),
    .X(_05895_));
 sky130_fd_sc_hd__xnor2_2 _15000_ (.A(_05893_),
    .B(_05895_),
    .Y(_05896_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1073 ();
 sky130_fd_sc_hd__mux2i_2 _15002_ (.A0(\text_in_r[122] ),
    .A1(_05896_),
    .S(net4120),
    .Y(_05898_));
 sky130_fd_sc_hd__xnor2_4 _15003_ (.A(net4168),
    .B(_05898_),
    .Y(_05899_));
 sky130_fd_sc_hd__clkinv_16 _15004_ (.A(_05899_),
    .Y(_05900_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1060 ();
 sky130_fd_sc_hd__xnor3_1 _15018_ (.A(\sa10_sr[4] ),
    .B(\sa20_sr[5] ),
    .C(\sa30_sr[5] ),
    .X(_05911_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1059 ();
 sky130_fd_sc_hd__xnor2_1 _15020_ (.A(\sa00_sr[4] ),
    .B(\sa10_sr[5] ),
    .Y(_05913_));
 sky130_fd_sc_hd__xnor2_1 _15021_ (.A(_05911_),
    .B(_05913_),
    .Y(_05914_));
 sky130_fd_sc_hd__nor2_2 _15022_ (.A(net398),
    .B(_05914_),
    .Y(_05915_));
 sky130_fd_sc_hd__a21oi_4 _15023_ (.A1(net398),
    .A2(\text_in_r[125] ),
    .B1(_05915_),
    .Y(_05916_));
 sky130_fd_sc_hd__xnor2_4 _15024_ (.A(net4165),
    .B(_05916_),
    .Y(_05917_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1056 ();
 sky130_fd_sc_hd__nor2_2 _15028_ (.A(net4057),
    .B(net4054),
    .Y(_05921_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1055 ();
 sky130_fd_sc_hd__nor2b_4 _15030_ (.A(net4230),
    .B_N(net4167),
    .Y(_05923_));
 sky130_fd_sc_hd__nor2_2 _15031_ (.A(net4167),
    .B(net4230),
    .Y(_05924_));
 sky130_fd_sc_hd__xnor2_1 _15032_ (.A(net4216),
    .B(\sa10_sr[3] ),
    .Y(_05925_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1054 ();
 sky130_fd_sc_hd__xnor3_1 _15034_ (.A(net4229),
    .B(\sa00_sr[2] ),
    .C(\sa20_sr[3] ),
    .X(_05927_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1053 ();
 sky130_fd_sc_hd__xnor2_1 _15036_ (.A(net4219),
    .B(\sa30_sr[3] ),
    .Y(_05929_));
 sky130_fd_sc_hd__xnor3_1 _15037_ (.A(_05925_),
    .B(_05927_),
    .C(_05929_),
    .X(_05930_));
 sky130_fd_sc_hd__mux2_8 _15038_ (.A0(_05923_),
    .A1(_05924_),
    .S(_05930_),
    .X(_05931_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1051 ();
 sky130_fd_sc_hd__nand2_2 _15041_ (.A(net4167),
    .B(net398),
    .Y(_05934_));
 sky130_fd_sc_hd__nand3b_1 _15042_ (.A_N(net4167),
    .B(net398),
    .C(\text_in_r[123] ),
    .Y(_05935_));
 sky130_fd_sc_hd__o21ai_4 _15043_ (.A1(\text_in_r[123] ),
    .A2(_05934_),
    .B1(_05935_),
    .Y(_05936_));
 sky130_fd_sc_hd__nor2_4 _15044_ (.A(_05936_),
    .B(_05931_),
    .Y(_05937_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1049 ();
 sky130_fd_sc_hd__o21ai_1 _15047_ (.A1(_11966_[0]),
    .A2(net3709),
    .B1(net4048),
    .Y(_05940_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1048 ();
 sky130_fd_sc_hd__nand2_1 _15049_ (.A(net4056),
    .B(net3709),
    .Y(_05942_));
 sky130_fd_sc_hd__mux2i_4 _15050_ (.A0(_05923_),
    .A1(_05924_),
    .S(_05930_),
    .Y(_05943_));
 sky130_fd_sc_hd__o21a_4 _15051_ (.A1(\text_in_r[123] ),
    .A2(_05934_),
    .B1(_05935_),
    .X(_05944_));
 sky130_fd_sc_hd__nand2_8 _15052_ (.A(_05943_),
    .B(_05944_),
    .Y(_05945_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1047 ();
 sky130_fd_sc_hd__nand3_4 _15054_ (.A(net3710),
    .B(_05891_),
    .C(net4054),
    .Y(_05947_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1046 ();
 sky130_fd_sc_hd__xnor3_1 _15056_ (.A(net4229),
    .B(\sa00_sr[3] ),
    .C(\sa20_sr[4] ),
    .X(_05949_));
 sky130_fd_sc_hd__xnor2_1 _15057_ (.A(net4217),
    .B(net4190),
    .Y(_05950_));
 sky130_fd_sc_hd__xnor3_1 _15058_ (.A(_05949_),
    .B(_05925_),
    .C(_05950_),
    .X(_05951_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1045 ();
 sky130_fd_sc_hd__mux2i_4 _15060_ (.A0(\text_in_r[124] ),
    .A1(_05951_),
    .S(net4120),
    .Y(_05953_));
 sky130_fd_sc_hd__xnor2_4 _15061_ (.A(net4166),
    .B(_05953_),
    .Y(_05954_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1044 ();
 sky130_fd_sc_hd__a31oi_2 _15063_ (.A1(_05942_),
    .A2(_05945_),
    .A3(_05947_),
    .B1(_05954_),
    .Y(_05956_));
 sky130_fd_sc_hd__o21ai_0 _15064_ (.A1(_05921_),
    .A2(_05940_),
    .B1(_05956_),
    .Y(_05957_));
 sky130_fd_sc_hd__xor2_4 _15065_ (.A(net4166),
    .B(_05953_),
    .X(_05958_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1043 ();
 sky130_fd_sc_hd__nand2_4 _15067_ (.A(_05917_),
    .B(_05958_),
    .Y(_05960_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1042 ();
 sky130_fd_sc_hd__nor2_1 _15069_ (.A(net3710),
    .B(net4048),
    .Y(_05962_));
 sky130_fd_sc_hd__nand2_8 _15070_ (.A(net4054),
    .B(_05945_),
    .Y(_05963_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1041 ();
 sky130_fd_sc_hd__o22a_1 _15072_ (.A1(_05942_),
    .A2(_05962_),
    .B1(_05963_),
    .B2(_11969_[0]),
    .X(_05965_));
 sky130_fd_sc_hd__o22ai_1 _15073_ (.A1(_05917_),
    .A2(_05957_),
    .B1(_05960_),
    .B2(_05965_),
    .Y(_05966_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1038 ();
 sky130_fd_sc_hd__xnor2_1 _15077_ (.A(\sa10_sr[7] ),
    .B(\sa20_sr[7] ),
    .Y(_05970_));
 sky130_fd_sc_hd__xor2_1 _15078_ (.A(\sa00_sr[6] ),
    .B(net4109),
    .X(_05971_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1036 ();
 sky130_fd_sc_hd__xnor2_1 _15081_ (.A(\sa10_sr[6] ),
    .B(net4189),
    .Y(_05974_));
 sky130_fd_sc_hd__xnor2_1 _15082_ (.A(_05971_),
    .B(_05974_),
    .Y(_05975_));
 sky130_fd_sc_hd__nand2_2 _15083_ (.A(net4119),
    .B(_05975_),
    .Y(_05976_));
 sky130_fd_sc_hd__o21ai_4 _15084_ (.A1(net4119),
    .A2(\text_in_r[127] ),
    .B1(_05976_),
    .Y(_05977_));
 sky130_fd_sc_hd__xor2_4 _15085_ (.A(\u0.w[0][31] ),
    .B(_05977_),
    .X(_05978_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1033 ();
 sky130_fd_sc_hd__xnor3_1 _15089_ (.A(\sa10_sr[5] ),
    .B(\sa20_sr[6] ),
    .C(\sa30_sr[6] ),
    .X(_05982_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1032 ();
 sky130_fd_sc_hd__xnor2_1 _15091_ (.A(\sa00_sr[5] ),
    .B(\sa10_sr[6] ),
    .Y(_05984_));
 sky130_fd_sc_hd__xnor2_1 _15092_ (.A(_05982_),
    .B(_05984_),
    .Y(_05985_));
 sky130_fd_sc_hd__nor2_1 _15093_ (.A(net398),
    .B(_05985_),
    .Y(_05986_));
 sky130_fd_sc_hd__a21oi_4 _15094_ (.A1(net398),
    .A2(\text_in_r[126] ),
    .B1(_05986_),
    .Y(_05987_));
 sky130_fd_sc_hd__xnor2_4 _15095_ (.A(net4164),
    .B(_05987_),
    .Y(_05988_));
 sky130_fd_sc_hd__nand2_4 _15096_ (.A(_05978_),
    .B(_05988_),
    .Y(_05989_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1031 ();
 sky130_fd_sc_hd__nor2_4 _15098_ (.A(_05900_),
    .B(net4051),
    .Y(_05991_));
 sky130_fd_sc_hd__nand2_8 _15099_ (.A(net4059),
    .B(net4048),
    .Y(_05992_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1030 ();
 sky130_fd_sc_hd__nand2_8 _15101_ (.A(_11978_[0]),
    .B(_05945_),
    .Y(_05994_));
 sky130_fd_sc_hd__a21oi_1 _15102_ (.A1(_05992_),
    .A2(_05994_),
    .B1(net4054),
    .Y(_05995_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1029 ();
 sky130_fd_sc_hd__nor2_4 _15104_ (.A(net4056),
    .B(_05945_),
    .Y(_05997_));
 sky130_fd_sc_hd__a211o_1 _15105_ (.A1(net3636),
    .A2(_05991_),
    .B1(_05995_),
    .C1(_05997_),
    .X(_05998_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1028 ();
 sky130_fd_sc_hd__nand2_4 _15107_ (.A(net3710),
    .B(net4050),
    .Y(_06000_));
 sky130_fd_sc_hd__nand3_1 _15108_ (.A(net4054),
    .B(_05994_),
    .C(_06000_),
    .Y(_06001_));
 sky130_fd_sc_hd__a31oi_1 _15109_ (.A1(net4056),
    .A2(net3709),
    .A3(_05992_),
    .B1(_05917_),
    .Y(_06002_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1027 ();
 sky130_fd_sc_hd__a221oi_2 _15111_ (.A1(_05917_),
    .A2(_05998_),
    .B1(_06001_),
    .B2(_06002_),
    .C1(_05958_),
    .Y(_06004_));
 sky130_fd_sc_hd__or3_4 _15112_ (.A(_05966_),
    .B(_05989_),
    .C(_06004_),
    .X(_06005_));
 sky130_fd_sc_hd__nor2_4 _15113_ (.A(_05917_),
    .B(_05978_),
    .Y(_06006_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1026 ();
 sky130_fd_sc_hd__nor3_2 _15115_ (.A(net4059),
    .B(_05891_),
    .C(_05900_),
    .Y(_06008_));
 sky130_fd_sc_hd__nor2_2 _15116_ (.A(_11969_[0]),
    .B(net4054),
    .Y(_06009_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1025 ();
 sky130_fd_sc_hd__o31ai_4 _15118_ (.A1(net4046),
    .A2(_06008_),
    .A3(_06009_),
    .B1(_05958_),
    .Y(_06011_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1024 ();
 sky130_fd_sc_hd__nor2_1 _15120_ (.A(_11964_[0]),
    .B(_05963_),
    .Y(_06013_));
 sky130_fd_sc_hd__nand2_4 _15121_ (.A(_05891_),
    .B(_05945_),
    .Y(_06014_));
 sky130_fd_sc_hd__nand2_4 _15122_ (.A(_11966_[0]),
    .B(net4049),
    .Y(_06015_));
 sky130_fd_sc_hd__a21oi_1 _15123_ (.A1(_06014_),
    .A2(_06015_),
    .B1(net4054),
    .Y(_06016_));
 sky130_fd_sc_hd__nor3_1 _15124_ (.A(_06011_),
    .B(_06013_),
    .C(_06016_),
    .Y(_06017_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1023 ();
 sky130_fd_sc_hd__nor2_4 _15126_ (.A(net4054),
    .B(_05945_),
    .Y(_06019_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1022 ();
 sky130_fd_sc_hd__a221oi_1 _15128_ (.A1(_11985_[0]),
    .A2(_05945_),
    .B1(_06019_),
    .B2(net3636),
    .C1(net4039),
    .Y(_06021_));
 sky130_fd_sc_hd__nor3_1 _15129_ (.A(_05988_),
    .B(_06017_),
    .C(_06021_),
    .Y(_06022_));
 sky130_fd_sc_hd__nand2_8 _15130_ (.A(net4056),
    .B(net4046),
    .Y(_06023_));
 sky130_fd_sc_hd__nor2_2 _15131_ (.A(_05954_),
    .B(_06023_),
    .Y(_06024_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1021 ();
 sky130_fd_sc_hd__nor2_2 _15133_ (.A(_11969_[0]),
    .B(_05945_),
    .Y(_06026_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1020 ();
 sky130_fd_sc_hd__nand2_4 _15135_ (.A(net3636),
    .B(_05945_),
    .Y(_06028_));
 sky130_fd_sc_hd__nand2_8 _15136_ (.A(_11974_[0]),
    .B(net4052),
    .Y(_06029_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1018 ();
 sky130_fd_sc_hd__a21oi_1 _15139_ (.A1(_06028_),
    .A2(_06029_),
    .B1(net3709),
    .Y(_06032_));
 sky130_fd_sc_hd__nor2_1 _15140_ (.A(_05958_),
    .B(_06032_),
    .Y(_06033_));
 sky130_fd_sc_hd__o32ai_1 _15141_ (.A1(net4054),
    .A2(_06024_),
    .A3(_06026_),
    .B1(_05956_),
    .B2(_06033_),
    .Y(_06034_));
 sky130_fd_sc_hd__xor2_4 _15142_ (.A(net4165),
    .B(_05916_),
    .X(_06035_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1017 ();
 sky130_fd_sc_hd__nand2_4 _15144_ (.A(_06035_),
    .B(_05988_),
    .Y(_06037_));
 sky130_fd_sc_hd__nor2_1 _15145_ (.A(_05978_),
    .B(_06037_),
    .Y(_06038_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1016 ();
 sky130_fd_sc_hd__a21oi_2 _15147_ (.A1(_05943_),
    .A2(_05944_),
    .B1(_11972_[0]),
    .Y(_06040_));
 sky130_fd_sc_hd__nor3_4 _15148_ (.A(_11965_[0]),
    .B(_05931_),
    .C(_05936_),
    .Y(_06041_));
 sky130_fd_sc_hd__nor3_1 _15149_ (.A(net4054),
    .B(_06040_),
    .C(_06041_),
    .Y(_06042_));
 sky130_fd_sc_hd__a31oi_1 _15150_ (.A1(net4054),
    .A2(_05992_),
    .A3(_06014_),
    .B1(_06042_),
    .Y(_06043_));
 sky130_fd_sc_hd__nand2_8 _15151_ (.A(_11969_[0]),
    .B(_05945_),
    .Y(_06044_));
 sky130_fd_sc_hd__nand3_2 _15152_ (.A(net4054),
    .B(_06015_),
    .C(_06044_),
    .Y(_06045_));
 sky130_fd_sc_hd__a21oi_1 _15153_ (.A1(_11964_[0]),
    .A2(_06019_),
    .B1(net4040),
    .Y(_06046_));
 sky130_fd_sc_hd__xor2_4 _15154_ (.A(net4164),
    .B(_05987_),
    .X(_06047_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1015 ();
 sky130_fd_sc_hd__a221oi_1 _15156_ (.A1(net4040),
    .A2(_06043_),
    .B1(_06045_),
    .B2(_06046_),
    .C1(_06047_),
    .Y(_06049_));
 sky130_fd_sc_hd__nand2_1 _15157_ (.A(_11966_[0]),
    .B(_05945_),
    .Y(_06050_));
 sky130_fd_sc_hd__o21ai_0 _15158_ (.A1(net4058),
    .A2(_05891_),
    .B1(net4049),
    .Y(_06051_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1014 ();
 sky130_fd_sc_hd__a21oi_2 _15160_ (.A1(_06050_),
    .A2(_06051_),
    .B1(_05900_),
    .Y(_06053_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1013 ();
 sky130_fd_sc_hd__nand2_1 _15162_ (.A(net4042),
    .B(_06047_),
    .Y(_06055_));
 sky130_fd_sc_hd__nand2_4 _15163_ (.A(_05900_),
    .B(net403),
    .Y(_06056_));
 sky130_fd_sc_hd__nor2_2 _15164_ (.A(_11972_[0]),
    .B(_06056_),
    .Y(_06057_));
 sky130_fd_sc_hd__nor3_1 _15165_ (.A(_06053_),
    .B(_06055_),
    .C(_06057_),
    .Y(_06058_));
 sky130_fd_sc_hd__xnor2_4 _15166_ (.A(\u0.w[0][31] ),
    .B(_05977_),
    .Y(_06059_));
 sky130_fd_sc_hd__nand2_4 _15167_ (.A(_05917_),
    .B(_06059_),
    .Y(_06060_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1012 ();
 sky130_fd_sc_hd__nor2_2 _15169_ (.A(net4057),
    .B(_05891_),
    .Y(_06062_));
 sky130_fd_sc_hd__nor2_4 _15170_ (.A(_05900_),
    .B(_05945_),
    .Y(_06063_));
 sky130_fd_sc_hd__a211oi_1 _15171_ (.A1(_11966_[0]),
    .A2(_06063_),
    .B1(_05988_),
    .C1(net4042),
    .Y(_06064_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1011 ();
 sky130_fd_sc_hd__nor2_4 _15173_ (.A(net4054),
    .B(net4053),
    .Y(_06066_));
 sky130_fd_sc_hd__nand2_1 _15174_ (.A(_11974_[0]),
    .B(_06066_),
    .Y(_06067_));
 sky130_fd_sc_hd__o211a_1 _15175_ (.A1(_05963_),
    .A2(_06062_),
    .B1(_06064_),
    .C1(_06067_),
    .X(_06068_));
 sky130_fd_sc_hd__nor4_2 _15176_ (.A(_06049_),
    .B(_06058_),
    .C(_06060_),
    .D(_06068_),
    .Y(_06069_));
 sky130_fd_sc_hd__a221oi_1 _15177_ (.A1(_06006_),
    .A2(_06022_),
    .B1(_06034_),
    .B2(_06038_),
    .C1(_06069_),
    .Y(_06070_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1010 ();
 sky130_fd_sc_hd__nor2_2 _15179_ (.A(net3708),
    .B(_05988_),
    .Y(_06072_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1009 ();
 sky130_fd_sc_hd__nor2_1 _15181_ (.A(_05884_),
    .B(net4054),
    .Y(_06074_));
 sky130_fd_sc_hd__nand2_4 _15182_ (.A(net3636),
    .B(net4048),
    .Y(_06075_));
 sky130_fd_sc_hd__nor2_2 _15183_ (.A(net3636),
    .B(net4054),
    .Y(_06076_));
 sky130_fd_sc_hd__a2bb2oi_1 _15184_ (.A1_N(_06074_),
    .A2_N(_06075_),
    .B1(_06076_),
    .B2(_05992_),
    .Y(_06077_));
 sky130_fd_sc_hd__xnor2_2 _15185_ (.A(_05900_),
    .B(net403),
    .Y(_06078_));
 sky130_fd_sc_hd__nor2_1 _15186_ (.A(_11964_[0]),
    .B(_06078_),
    .Y(_06079_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1008 ();
 sky130_fd_sc_hd__a2111oi_0 _15188_ (.A1(net3636),
    .A2(_05991_),
    .B1(_06057_),
    .C1(_06079_),
    .D1(net4042),
    .Y(_06081_));
 sky130_fd_sc_hd__a21oi_1 _15189_ (.A1(_05954_),
    .A2(_06077_),
    .B1(net3574),
    .Y(_06082_));
 sky130_fd_sc_hd__inv_6 _15190_ (.A(net3636),
    .Y(_06083_));
 sky130_fd_sc_hd__nand2_2 _15191_ (.A(_06083_),
    .B(net403),
    .Y(_06084_));
 sky130_fd_sc_hd__nand2_4 _15192_ (.A(_11972_[0]),
    .B(net4044),
    .Y(_06085_));
 sky130_fd_sc_hd__nand2_4 _15193_ (.A(net3710),
    .B(_05997_),
    .Y(_06086_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1007 ();
 sky130_fd_sc_hd__a21oi_1 _15195_ (.A1(_11964_[0]),
    .A2(_05945_),
    .B1(net4054),
    .Y(_06088_));
 sky130_fd_sc_hd__a32oi_1 _15196_ (.A1(net4054),
    .A2(_06084_),
    .A3(_06085_),
    .B1(_06086_),
    .B2(_06088_),
    .Y(_06089_));
 sky130_fd_sc_hd__nand2_8 _15197_ (.A(_05891_),
    .B(net4054),
    .Y(_06090_));
 sky130_fd_sc_hd__nand2_4 _15198_ (.A(net4057),
    .B(net4056),
    .Y(_06091_));
 sky130_fd_sc_hd__a21oi_2 _15199_ (.A1(_06090_),
    .A2(_06091_),
    .B1(net4049),
    .Y(_06092_));
 sky130_fd_sc_hd__and3_1 _15200_ (.A(net4049),
    .B(_06090_),
    .C(_06091_),
    .X(_06093_));
 sky130_fd_sc_hd__nor3_1 _15201_ (.A(net4039),
    .B(_06092_),
    .C(_06093_),
    .Y(_06094_));
 sky130_fd_sc_hd__nand2_4 _15202_ (.A(_05978_),
    .B(_06047_),
    .Y(_06095_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1006 ();
 sky130_fd_sc_hd__a2111oi_0 _15204_ (.A1(net4039),
    .A2(_06089_),
    .B1(_06094_),
    .C1(_06095_),
    .D1(net3706),
    .Y(_06097_));
 sky130_fd_sc_hd__a31oi_1 _15205_ (.A1(_05978_),
    .A2(_06072_),
    .A3(_06082_),
    .B1(net3573),
    .Y(_06098_));
 sky130_fd_sc_hd__nand3_2 _15206_ (.A(_06005_),
    .B(_06070_),
    .C(_06098_),
    .Y(_00032_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1003 ();
 sky130_fd_sc_hd__nor2_2 _15210_ (.A(_06083_),
    .B(net4054),
    .Y(_06102_));
 sky130_fd_sc_hd__a21oi_1 _15211_ (.A1(_11978_[0]),
    .A2(net4054),
    .B1(_06102_),
    .Y(_06103_));
 sky130_fd_sc_hd__o21bai_2 _15212_ (.A1(net4050),
    .A2(_06103_),
    .B1_N(_06011_),
    .Y(_06104_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1002 ();
 sky130_fd_sc_hd__o22ai_1 _15214_ (.A1(_11969_[0]),
    .A2(_06056_),
    .B1(_06078_),
    .B2(net4057),
    .Y(_06105_));
 sky130_fd_sc_hd__nand2_1 _15215_ (.A(_05954_),
    .B(_06105_),
    .Y(_06106_));
 sky130_fd_sc_hd__nand2_1 _15216_ (.A(net4054),
    .B(net4041),
    .Y(_06107_));
 sky130_fd_sc_hd__nand2_1 _15217_ (.A(net4056),
    .B(_06066_),
    .Y(_06108_));
 sky130_fd_sc_hd__a21oi_1 _15218_ (.A1(_06107_),
    .A2(_06108_),
    .B1(net4057),
    .Y(_06109_));
 sky130_fd_sc_hd__nor2_4 _15219_ (.A(net4054),
    .B(_05958_),
    .Y(_06110_));
 sky130_fd_sc_hd__nor2_1 _15220_ (.A(_05954_),
    .B(_05945_),
    .Y(_06111_));
 sky130_fd_sc_hd__a22oi_1 _15221_ (.A1(_05945_),
    .A2(_06110_),
    .B1(_06111_),
    .B2(net4057),
    .Y(_06112_));
 sky130_fd_sc_hd__nor2_1 _15222_ (.A(_05891_),
    .B(_06112_),
    .Y(_06113_));
 sky130_fd_sc_hd__nand2_8 _15223_ (.A(_05891_),
    .B(_05900_),
    .Y(_06114_));
 sky130_fd_sc_hd__nand2_2 _15224_ (.A(_05954_),
    .B(net4051),
    .Y(_06115_));
 sky130_fd_sc_hd__o21ai_0 _15225_ (.A1(_06083_),
    .A2(_05958_),
    .B1(_05945_),
    .Y(_06116_));
 sky130_fd_sc_hd__o21a_1 _15226_ (.A1(_11969_[0]),
    .A2(_06115_),
    .B1(_06116_),
    .X(_06117_));
 sky130_fd_sc_hd__o22ai_1 _15227_ (.A1(_06114_),
    .A2(_06115_),
    .B1(_06117_),
    .B2(net3709),
    .Y(_06118_));
 sky130_fd_sc_hd__nor4_1 _15228_ (.A(_06060_),
    .B(_06109_),
    .C(_06113_),
    .D(_06118_),
    .Y(_06119_));
 sky130_fd_sc_hd__a31oi_2 _15229_ (.A1(_06006_),
    .A2(_06104_),
    .A3(_06106_),
    .B1(_06119_),
    .Y(_06120_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1001 ();
 sky130_fd_sc_hd__a21oi_1 _15231_ (.A1(_11972_[0]),
    .A2(_05900_),
    .B1(net4044),
    .Y(_06122_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1000 ();
 sky130_fd_sc_hd__a21oi_1 _15233_ (.A1(_05947_),
    .A2(_06122_),
    .B1(net4042),
    .Y(_06124_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_998 ();
 sky130_fd_sc_hd__nor2_1 _15236_ (.A(_11988_[0]),
    .B(net4049),
    .Y(_06127_));
 sky130_fd_sc_hd__a21oi_1 _15237_ (.A1(_06035_),
    .A2(_06127_),
    .B1(_05988_),
    .Y(_06128_));
 sky130_fd_sc_hd__nand2_8 _15238_ (.A(_05884_),
    .B(_05945_),
    .Y(_06129_));
 sky130_fd_sc_hd__a21oi_1 _15239_ (.A1(_05992_),
    .A2(_06129_),
    .B1(net4054),
    .Y(_06130_));
 sky130_fd_sc_hd__nand2_1 _15240_ (.A(net4056),
    .B(net4049),
    .Y(_06131_));
 sky130_fd_sc_hd__a21oi_1 _15241_ (.A1(_06044_),
    .A2(_06131_),
    .B1(_05900_),
    .Y(_06132_));
 sky130_fd_sc_hd__o21ai_0 _15242_ (.A1(_06130_),
    .A2(_06132_),
    .B1(_06035_),
    .Y(_06133_));
 sky130_fd_sc_hd__nand2_1 _15243_ (.A(net4056),
    .B(net4054),
    .Y(_06134_));
 sky130_fd_sc_hd__nand2_1 _15244_ (.A(_11964_[0]),
    .B(_05900_),
    .Y(_06135_));
 sky130_fd_sc_hd__a21o_1 _15245_ (.A1(_06134_),
    .A2(_06135_),
    .B1(net4044),
    .X(_06136_));
 sky130_fd_sc_hd__nor2_2 _15246_ (.A(net4057),
    .B(net4049),
    .Y(_06137_));
 sky130_fd_sc_hd__a31oi_1 _15247_ (.A1(_06134_),
    .A2(_06137_),
    .A3(_06114_),
    .B1(_06035_),
    .Y(_06138_));
 sky130_fd_sc_hd__a21oi_1 _15248_ (.A1(_06136_),
    .A2(_06138_),
    .B1(_06055_),
    .Y(_06139_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_997 ();
 sky130_fd_sc_hd__a221oi_1 _15250_ (.A1(_06124_),
    .A2(_06128_),
    .B1(_06133_),
    .B2(_06139_),
    .C1(_06059_),
    .Y(_06141_));
 sky130_fd_sc_hd__nand2_1 _15251_ (.A(_06047_),
    .B(_06141_),
    .Y(_06142_));
 sky130_fd_sc_hd__nand2_4 _15252_ (.A(_06059_),
    .B(net3707),
    .Y(_06143_));
 sky130_fd_sc_hd__nor2_4 _15253_ (.A(net4057),
    .B(_05900_),
    .Y(_06144_));
 sky130_fd_sc_hd__a21oi_1 _15254_ (.A1(net3598),
    .A2(_05900_),
    .B1(_06144_),
    .Y(_06145_));
 sky130_fd_sc_hd__nor3_1 _15255_ (.A(net4039),
    .B(net4049),
    .C(_06145_),
    .Y(_06146_));
 sky130_fd_sc_hd__nor2_4 _15256_ (.A(net4058),
    .B(net4056),
    .Y(_06147_));
 sky130_fd_sc_hd__o21ai_0 _15257_ (.A1(_11969_[0]),
    .A2(net4043),
    .B1(_06063_),
    .Y(_06148_));
 sky130_fd_sc_hd__o21ai_0 _15258_ (.A1(_06147_),
    .A2(_06148_),
    .B1(net3708),
    .Y(_06149_));
 sky130_fd_sc_hd__o21ai_4 _15259_ (.A1(net4057),
    .A2(net4056),
    .B1(net4047),
    .Y(_06150_));
 sky130_fd_sc_hd__nand2_8 _15260_ (.A(_06083_),
    .B(_05945_),
    .Y(_06151_));
 sky130_fd_sc_hd__nand2_2 _15261_ (.A(_11969_[0]),
    .B(net4050),
    .Y(_06152_));
 sky130_fd_sc_hd__and3_1 _15262_ (.A(net4054),
    .B(_06151_),
    .C(_06152_),
    .X(_06153_));
 sky130_fd_sc_hd__a211oi_1 _15263_ (.A1(_05900_),
    .A2(_06150_),
    .B1(_06153_),
    .C1(net4043),
    .Y(_06154_));
 sky130_fd_sc_hd__nor3_1 _15264_ (.A(_06146_),
    .B(_06149_),
    .C(_06154_),
    .Y(_06155_));
 sky130_fd_sc_hd__nor2_4 _15265_ (.A(net4056),
    .B(net4050),
    .Y(_06156_));
 sky130_fd_sc_hd__nor2_1 _15266_ (.A(_05891_),
    .B(_06078_),
    .Y(_06157_));
 sky130_fd_sc_hd__a221oi_1 _15267_ (.A1(net4057),
    .A2(_06156_),
    .B1(_06019_),
    .B2(net3636),
    .C1(_06157_),
    .Y(_06158_));
 sky130_fd_sc_hd__nand2_4 _15268_ (.A(_05891_),
    .B(net4052),
    .Y(_06159_));
 sky130_fd_sc_hd__nand2_8 _15269_ (.A(_11964_[0]),
    .B(net4050),
    .Y(_06160_));
 sky130_fd_sc_hd__a21oi_1 _15270_ (.A1(_06028_),
    .A2(_06160_),
    .B1(_05900_),
    .Y(_06161_));
 sky130_fd_sc_hd__a311oi_1 _15271_ (.A1(_05900_),
    .A2(_06159_),
    .A3(_06044_),
    .B1(_06161_),
    .C1(net4041),
    .Y(_06162_));
 sky130_fd_sc_hd__a211oi_1 _15272_ (.A1(net4041),
    .A2(_06158_),
    .B1(_06162_),
    .C1(_05917_),
    .Y(_06163_));
 sky130_fd_sc_hd__or3_4 _15273_ (.A(_06143_),
    .B(_06155_),
    .C(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__nor2_2 _15274_ (.A(net3636),
    .B(net4051),
    .Y(_06165_));
 sky130_fd_sc_hd__nand2_4 _15275_ (.A(_11978_[0]),
    .B(net4051),
    .Y(_06166_));
 sky130_fd_sc_hd__nand2_2 _15276_ (.A(net4054),
    .B(_06166_),
    .Y(_06167_));
 sky130_fd_sc_hd__o211ai_1 _15277_ (.A1(_06165_),
    .A2(_06167_),
    .B1(net3705),
    .C1(net4043),
    .Y(_06168_));
 sky130_fd_sc_hd__a31oi_1 _15278_ (.A1(_05900_),
    .A2(_06015_),
    .A3(_06150_),
    .B1(_06168_),
    .Y(_06169_));
 sky130_fd_sc_hd__a21oi_1 _15279_ (.A1(_06086_),
    .A2(_06151_),
    .B1(_05900_),
    .Y(_06170_));
 sky130_fd_sc_hd__a21oi_1 _15280_ (.A1(net4056),
    .A2(_06019_),
    .B1(_05917_),
    .Y(_06171_));
 sky130_fd_sc_hd__nor3b_1 _15281_ (.A(net4043),
    .B(_06170_),
    .C_N(_06171_),
    .Y(_06172_));
 sky130_fd_sc_hd__o21ai_0 _15282_ (.A1(_11964_[0]),
    .A2(_05945_),
    .B1(_06129_),
    .Y(_06173_));
 sky130_fd_sc_hd__a21oi_1 _15283_ (.A1(_05900_),
    .A2(_06173_),
    .B1(_06132_),
    .Y(_06174_));
 sky130_fd_sc_hd__nand2_4 _15284_ (.A(net3708),
    .B(net4042),
    .Y(_06175_));
 sky130_fd_sc_hd__nand2_2 _15285_ (.A(_06159_),
    .B(_06028_),
    .Y(_06176_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_996 ();
 sky130_fd_sc_hd__nor2_1 _15287_ (.A(_11966_[0]),
    .B(net4044),
    .Y(_06178_));
 sky130_fd_sc_hd__a211oi_1 _15288_ (.A1(_11964_[0]),
    .A2(_05945_),
    .B1(_06178_),
    .C1(_05900_),
    .Y(_06179_));
 sky130_fd_sc_hd__a21oi_1 _15289_ (.A1(_05900_),
    .A2(_06176_),
    .B1(_06179_),
    .Y(_06180_));
 sky130_fd_sc_hd__o22ai_1 _15290_ (.A1(_05960_),
    .A2(_06174_),
    .B1(_06175_),
    .B2(_06180_),
    .Y(_06181_));
 sky130_fd_sc_hd__o31ai_1 _15291_ (.A1(_06169_),
    .A2(_06172_),
    .A3(_06181_),
    .B1(_06141_),
    .Y(_06182_));
 sky130_fd_sc_hd__o2111ai_2 _15292_ (.A1(net3707),
    .A2(_06120_),
    .B1(_06142_),
    .C1(_06164_),
    .D1(_06182_),
    .Y(_00033_));
 sky130_fd_sc_hd__or3_4 _15293_ (.A(_11978_[0]),
    .B(_05931_),
    .C(_05936_),
    .X(_06183_));
 sky130_fd_sc_hd__nor2_4 _15294_ (.A(_11974_[0]),
    .B(net4049),
    .Y(_06184_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_995 ();
 sky130_fd_sc_hd__nor3b_1 _15296_ (.A(_06184_),
    .B(_05900_),
    .C_N(_06131_),
    .Y(_06186_));
 sky130_fd_sc_hd__a31oi_1 _15297_ (.A1(_05900_),
    .A2(_06129_),
    .A3(_06183_),
    .B1(_06186_),
    .Y(_06187_));
 sky130_fd_sc_hd__nor2_4 _15298_ (.A(net4057),
    .B(net4044),
    .Y(_06188_));
 sky130_fd_sc_hd__nor2_1 _15299_ (.A(_11966_[0]),
    .B(net4049),
    .Y(_06189_));
 sky130_fd_sc_hd__nor3_1 _15300_ (.A(net4054),
    .B(_06188_),
    .C(_06189_),
    .Y(_06190_));
 sky130_fd_sc_hd__a21oi_2 _15301_ (.A1(_06014_),
    .A2(_06075_),
    .B1(_05900_),
    .Y(_06191_));
 sky130_fd_sc_hd__nor3_1 _15302_ (.A(_05988_),
    .B(_06190_),
    .C(_06191_),
    .Y(_06192_));
 sky130_fd_sc_hd__a21oi_1 _15303_ (.A1(_05988_),
    .A2(_06187_),
    .B1(_06192_),
    .Y(_06193_));
 sky130_fd_sc_hd__o21ai_0 _15304_ (.A1(_06008_),
    .A2(_06009_),
    .B1(net4046),
    .Y(_06194_));
 sky130_fd_sc_hd__nand2_1 _15305_ (.A(_05958_),
    .B(_06194_),
    .Y(_06195_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_994 ();
 sky130_fd_sc_hd__nor3_1 _15307_ (.A(net4046),
    .B(_06102_),
    .C(_06144_),
    .Y(_06197_));
 sky130_fd_sc_hd__a21oi_2 _15308_ (.A1(_06137_),
    .A2(_06114_),
    .B1(net4039),
    .Y(_06198_));
 sky130_fd_sc_hd__nand2_1 _15309_ (.A(_11969_[0]),
    .B(net4054),
    .Y(_06199_));
 sky130_fd_sc_hd__a21oi_1 _15310_ (.A1(net3598),
    .A2(_05900_),
    .B1(net4044),
    .Y(_06200_));
 sky130_fd_sc_hd__nand2_1 _15311_ (.A(_06199_),
    .B(_06200_),
    .Y(_06201_));
 sky130_fd_sc_hd__nand2_1 _15312_ (.A(_06198_),
    .B(_06201_),
    .Y(_06202_));
 sky130_fd_sc_hd__o211ai_1 _15313_ (.A1(_06195_),
    .A2(_06197_),
    .B1(_06072_),
    .C1(_06202_),
    .Y(_06203_));
 sky130_fd_sc_hd__o21ai_0 _15314_ (.A1(_06175_),
    .A2(_06193_),
    .B1(_06203_),
    .Y(_06204_));
 sky130_fd_sc_hd__nor2_1 _15315_ (.A(_05900_),
    .B(_06176_),
    .Y(_06205_));
 sky130_fd_sc_hd__a311oi_1 _15316_ (.A1(_05900_),
    .A2(_06029_),
    .A3(_06151_),
    .B1(_06205_),
    .C1(_06047_),
    .Y(_06206_));
 sky130_fd_sc_hd__o21ai_0 _15317_ (.A1(net3598),
    .A2(_05963_),
    .B1(_06047_),
    .Y(_06207_));
 sky130_fd_sc_hd__a31oi_1 _15318_ (.A1(_05921_),
    .A2(_06159_),
    .A3(_06023_),
    .B1(_06207_),
    .Y(_06208_));
 sky130_fd_sc_hd__nor2_1 _15319_ (.A(_11969_[0]),
    .B(net4048),
    .Y(_06209_));
 sky130_fd_sc_hd__nor2_4 _15320_ (.A(net3598),
    .B(net4044),
    .Y(_06210_));
 sky130_fd_sc_hd__o211ai_1 _15321_ (.A1(_11974_[0]),
    .A2(net4046),
    .B1(_06023_),
    .C1(net4054),
    .Y(_06211_));
 sky130_fd_sc_hd__o31ai_1 _15322_ (.A1(net4054),
    .A2(_06209_),
    .A3(_06210_),
    .B1(_06211_),
    .Y(_06212_));
 sky130_fd_sc_hd__a311oi_1 _15323_ (.A1(net4054),
    .A2(_06029_),
    .A3(_06129_),
    .B1(_05954_),
    .C1(_06009_),
    .Y(_06213_));
 sky130_fd_sc_hd__a211o_1 _15324_ (.A1(_05954_),
    .A2(_06212_),
    .B1(_06213_),
    .C1(_06037_),
    .X(_06214_));
 sky130_fd_sc_hd__o311ai_0 _15325_ (.A1(_05960_),
    .A2(_06206_),
    .A3(_06208_),
    .B1(_06214_),
    .C1(_05978_),
    .Y(_06215_));
 sky130_fd_sc_hd__nand3_1 _15326_ (.A(net4054),
    .B(_05992_),
    .C(_06085_),
    .Y(_06216_));
 sky130_fd_sc_hd__nand3_1 _15327_ (.A(_05900_),
    .B(_06160_),
    .C(_06151_),
    .Y(_06217_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_993 ();
 sky130_fd_sc_hd__a21oi_1 _15329_ (.A1(_06216_),
    .A2(_06217_),
    .B1(net4039),
    .Y(_06219_));
 sky130_fd_sc_hd__nand2_1 _15330_ (.A(net4039),
    .B(net4044),
    .Y(_06220_));
 sky130_fd_sc_hd__nor2_1 _15331_ (.A(_06220_),
    .B(_06144_),
    .Y(_06221_));
 sky130_fd_sc_hd__a21oi_1 _15332_ (.A1(_06091_),
    .A2(_06221_),
    .B1(_06037_),
    .Y(_06222_));
 sky130_fd_sc_hd__o31ai_1 _15333_ (.A1(_11988_[0]),
    .A2(net4042),
    .A3(net4044),
    .B1(_06222_),
    .Y(_06223_));
 sky130_fd_sc_hd__o21ai_0 _15334_ (.A1(_06188_),
    .A2(_06074_),
    .B1(net3636),
    .Y(_06224_));
 sky130_fd_sc_hd__a22oi_1 _15335_ (.A1(_05962_),
    .A2(_06090_),
    .B1(_06014_),
    .B2(_06144_),
    .Y(_06225_));
 sky130_fd_sc_hd__a21oi_1 _15336_ (.A1(_06224_),
    .A2(_06225_),
    .B1(net4039),
    .Y(_06226_));
 sky130_fd_sc_hd__nor3_1 _15337_ (.A(net4048),
    .B(_06008_),
    .C(_06076_),
    .Y(_06227_));
 sky130_fd_sc_hd__a211oi_1 _15338_ (.A1(_11985_[0]),
    .A2(net4048),
    .B1(_06227_),
    .C1(net4042),
    .Y(_06228_));
 sky130_fd_sc_hd__nor2_1 _15339_ (.A(_06035_),
    .B(_06047_),
    .Y(_06229_));
 sky130_fd_sc_hd__o21ai_1 _15340_ (.A1(_06226_),
    .A2(_06228_),
    .B1(_06229_),
    .Y(_06230_));
 sky130_fd_sc_hd__o211ai_1 _15341_ (.A1(_06219_),
    .A2(_06223_),
    .B1(_06230_),
    .C1(_06059_),
    .Y(_06231_));
 sky130_fd_sc_hd__a32oi_1 _15342_ (.A1(net4054),
    .A2(_06160_),
    .A3(_06151_),
    .B1(_06066_),
    .B2(_11969_[0]),
    .Y(_06232_));
 sky130_fd_sc_hd__nor2_1 _15343_ (.A(_11983_[0]),
    .B(net4049),
    .Y(_06233_));
 sky130_fd_sc_hd__a21oi_1 _15344_ (.A1(_05900_),
    .A2(_06062_),
    .B1(net4045),
    .Y(_06234_));
 sky130_fd_sc_hd__o21ai_0 _15345_ (.A1(_06233_),
    .A2(_06234_),
    .B1(net3706),
    .Y(_06235_));
 sky130_fd_sc_hd__o21ai_0 _15346_ (.A1(net3706),
    .A2(_06232_),
    .B1(_06235_),
    .Y(_06236_));
 sky130_fd_sc_hd__nor2_1 _15347_ (.A(net4045),
    .B(_06147_),
    .Y(_06237_));
 sky130_fd_sc_hd__nor2_4 _15348_ (.A(_11966_[0]),
    .B(_11969_[0]),
    .Y(_06238_));
 sky130_fd_sc_hd__nor2_4 _15349_ (.A(net4049),
    .B(_06238_),
    .Y(_06239_));
 sky130_fd_sc_hd__nor3_1 _15350_ (.A(_05900_),
    .B(_06237_),
    .C(_06239_),
    .Y(_06240_));
 sky130_fd_sc_hd__o21ai_0 _15351_ (.A1(_11972_[0]),
    .A2(_05945_),
    .B1(_06150_),
    .Y(_06241_));
 sky130_fd_sc_hd__nor2_1 _15352_ (.A(net4054),
    .B(_06241_),
    .Y(_06242_));
 sky130_fd_sc_hd__o211ai_1 _15353_ (.A1(_11992_[0]),
    .A2(net4044),
    .B1(_06198_),
    .C1(_06035_),
    .Y(_06243_));
 sky130_fd_sc_hd__o311ai_0 _15354_ (.A1(_06175_),
    .A2(_06240_),
    .A3(_06242_),
    .B1(_06243_),
    .C1(_06047_),
    .Y(_06244_));
 sky130_fd_sc_hd__a21oi_1 _15355_ (.A1(net4039),
    .A2(_06236_),
    .B1(_06244_),
    .Y(_06245_));
 sky130_fd_sc_hd__o22ai_1 _15356_ (.A1(_06204_),
    .A2(_06215_),
    .B1(_06231_),
    .B2(_06245_),
    .Y(_00034_));
 sky130_fd_sc_hd__nand2_2 _15357_ (.A(net3709),
    .B(_05958_),
    .Y(_06246_));
 sky130_fd_sc_hd__nor2_1 _15358_ (.A(net3709),
    .B(_05954_),
    .Y(_06247_));
 sky130_fd_sc_hd__nor2_1 _15359_ (.A(_06110_),
    .B(_06247_),
    .Y(_06248_));
 sky130_fd_sc_hd__o221ai_1 _15360_ (.A1(net3710),
    .A2(_06246_),
    .B1(_06248_),
    .B2(net3636),
    .C1(_05945_),
    .Y(_06249_));
 sky130_fd_sc_hd__a21oi_1 _15361_ (.A1(net4056),
    .A2(_05958_),
    .B1(net4054),
    .Y(_06250_));
 sky130_fd_sc_hd__nand2_1 _15362_ (.A(net4057),
    .B(_05954_),
    .Y(_06251_));
 sky130_fd_sc_hd__o2111ai_1 _15363_ (.A1(net4057),
    .A2(_06250_),
    .B1(_06251_),
    .C1(net4050),
    .D1(_06090_),
    .Y(_06252_));
 sky130_fd_sc_hd__o2111ai_1 _15364_ (.A1(_05958_),
    .A2(_06090_),
    .B1(_06006_),
    .C1(_06249_),
    .D1(_06252_),
    .Y(_06253_));
 sky130_fd_sc_hd__nor2_1 _15365_ (.A(_11964_[0]),
    .B(net403),
    .Y(_06254_));
 sky130_fd_sc_hd__nor2_1 _15366_ (.A(_11972_[0]),
    .B(_05945_),
    .Y(_06255_));
 sky130_fd_sc_hd__nor3_1 _15367_ (.A(_05900_),
    .B(_06254_),
    .C(_06255_),
    .Y(_06256_));
 sky130_fd_sc_hd__a311oi_1 _15368_ (.A1(_05900_),
    .A2(_06159_),
    .A3(_06151_),
    .B1(_06256_),
    .C1(net4041),
    .Y(_06257_));
 sky130_fd_sc_hd__a21oi_1 _15369_ (.A1(_05994_),
    .A2(_06084_),
    .B1(_06107_),
    .Y(_06258_));
 sky130_fd_sc_hd__a21oi_1 _15370_ (.A1(_06000_),
    .A2(_06044_),
    .B1(_06246_),
    .Y(_06259_));
 sky130_fd_sc_hd__or4_1 _15371_ (.A(_06060_),
    .B(_06257_),
    .C(_06258_),
    .D(_06259_),
    .X(_06260_));
 sky130_fd_sc_hd__a21oi_1 _15372_ (.A1(_06253_),
    .A2(_06260_),
    .B1(net3707),
    .Y(_06261_));
 sky130_fd_sc_hd__o21ai_2 _15373_ (.A1(net3624),
    .A2(_06184_),
    .B1(net4055),
    .Y(_06262_));
 sky130_fd_sc_hd__o21ai_0 _15374_ (.A1(_06156_),
    .A2(_06210_),
    .B1(_05900_),
    .Y(_06263_));
 sky130_fd_sc_hd__nand2_1 _15375_ (.A(_06262_),
    .B(_06263_),
    .Y(_06264_));
 sky130_fd_sc_hd__a21oi_1 _15376_ (.A1(net4054),
    .A2(_05992_),
    .B1(net4056),
    .Y(_06265_));
 sky130_fd_sc_hd__a211oi_2 _15377_ (.A1(net3710),
    .A2(_06019_),
    .B1(_06013_),
    .C1(_06265_),
    .Y(_06266_));
 sky130_fd_sc_hd__o22ai_1 _15378_ (.A1(_06175_),
    .A2(_06264_),
    .B1(_06266_),
    .B2(_05960_),
    .Y(_06267_));
 sky130_fd_sc_hd__a21oi_1 _15379_ (.A1(net4054),
    .A2(_06238_),
    .B1(net4049),
    .Y(_06268_));
 sky130_fd_sc_hd__o21ai_0 _15380_ (.A1(_11974_[0]),
    .A2(net4054),
    .B1(_06268_),
    .Y(_06269_));
 sky130_fd_sc_hd__nor2_4 _15381_ (.A(net4056),
    .B(net3709),
    .Y(_06270_));
 sky130_fd_sc_hd__a211oi_2 _15382_ (.A1(_11978_[0]),
    .A2(net3709),
    .B1(_06270_),
    .C1(_06115_),
    .Y(_06271_));
 sky130_fd_sc_hd__a211oi_1 _15383_ (.A1(_06124_),
    .A2(_06269_),
    .B1(_06271_),
    .C1(net3708),
    .Y(_06272_));
 sky130_fd_sc_hd__nor3_1 _15384_ (.A(_05989_),
    .B(_06267_),
    .C(_06272_),
    .Y(_06273_));
 sky130_fd_sc_hd__nor2_2 _15385_ (.A(net3709),
    .B(_05958_),
    .Y(_06274_));
 sky130_fd_sc_hd__o21ai_0 _15386_ (.A1(_06035_),
    .A2(_06084_),
    .B1(_06050_),
    .Y(_06275_));
 sky130_fd_sc_hd__nand2_2 _15387_ (.A(net4051),
    .B(_06270_),
    .Y(_06276_));
 sky130_fd_sc_hd__nand2_1 _15388_ (.A(_11974_[0]),
    .B(_06078_),
    .Y(_06277_));
 sky130_fd_sc_hd__a211oi_1 _15389_ (.A1(net4044),
    .A2(_06238_),
    .B1(_06041_),
    .C1(_05900_),
    .Y(_06278_));
 sky130_fd_sc_hd__a21oi_1 _15390_ (.A1(_05994_),
    .A2(_06159_),
    .B1(net4054),
    .Y(_06279_));
 sky130_fd_sc_hd__nor3_1 _15391_ (.A(net3708),
    .B(_06278_),
    .C(_06279_),
    .Y(_06280_));
 sky130_fd_sc_hd__a311oi_1 _15392_ (.A1(net3708),
    .A2(_06276_),
    .A3(_06277_),
    .B1(net4043),
    .C1(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__nand2_1 _15393_ (.A(net4058),
    .B(_06063_),
    .Y(_06282_));
 sky130_fd_sc_hd__o21ai_0 _15394_ (.A1(_06165_),
    .A2(_06255_),
    .B1(_05900_),
    .Y(_06283_));
 sky130_fd_sc_hd__a211oi_1 _15395_ (.A1(_06282_),
    .A2(_06283_),
    .B1(net3708),
    .C1(net4041),
    .Y(_06284_));
 sky130_fd_sc_hd__a2111oi_0 _15396_ (.A1(_06274_),
    .A2(_06275_),
    .B1(_06281_),
    .C1(_06284_),
    .D1(_06095_),
    .Y(_06285_));
 sky130_fd_sc_hd__nor3_1 _15397_ (.A(_05900_),
    .B(net3624),
    .C(_06137_),
    .Y(_06286_));
 sky130_fd_sc_hd__a31oi_1 _15398_ (.A1(_05900_),
    .A2(_05994_),
    .A3(_06029_),
    .B1(_06286_),
    .Y(_06287_));
 sky130_fd_sc_hd__a31oi_1 _15399_ (.A1(_05963_),
    .A2(_06091_),
    .A3(_06114_),
    .B1(net4042),
    .Y(_06288_));
 sky130_fd_sc_hd__a21o_1 _15400_ (.A1(net4042),
    .A2(_06287_),
    .B1(_06288_),
    .X(_06289_));
 sky130_fd_sc_hd__nor2_1 _15401_ (.A(net3636),
    .B(_06056_),
    .Y(_06290_));
 sky130_fd_sc_hd__a21oi_1 _15402_ (.A1(_06108_),
    .A2(_06276_),
    .B1(net4058),
    .Y(_06291_));
 sky130_fd_sc_hd__a2111oi_0 _15403_ (.A1(_11972_[0]),
    .A2(_05991_),
    .B1(_05960_),
    .C1(_06290_),
    .D1(_06291_),
    .Y(_06292_));
 sky130_fd_sc_hd__a21oi_1 _15404_ (.A1(net4044),
    .A2(_06091_),
    .B1(_06122_),
    .Y(_06293_));
 sky130_fd_sc_hd__nor3_1 _15405_ (.A(_06175_),
    .B(_06191_),
    .C(_06293_),
    .Y(_06294_));
 sky130_fd_sc_hd__a2111oi_0 _15406_ (.A1(net3706),
    .A2(_06289_),
    .B1(_06292_),
    .C1(_06294_),
    .D1(_06143_),
    .Y(_06295_));
 sky130_fd_sc_hd__nor4_1 _15407_ (.A(_06261_),
    .B(_06273_),
    .C(_06285_),
    .D(_06295_),
    .Y(_00035_));
 sky130_fd_sc_hd__a21oi_2 _15408_ (.A1(_11964_[0]),
    .A2(net3709),
    .B1(_05940_),
    .Y(_06296_));
 sky130_fd_sc_hd__nand3_1 _15409_ (.A(net4042),
    .B(_06067_),
    .C(_06086_),
    .Y(_06297_));
 sky130_fd_sc_hd__a21oi_1 _15410_ (.A1(_05992_),
    .A2(_06023_),
    .B1(_05900_),
    .Y(_06298_));
 sky130_fd_sc_hd__o32a_1 _15411_ (.A1(net4042),
    .A2(_06092_),
    .A3(_06296_),
    .B1(_06297_),
    .B2(_06298_),
    .X(_06299_));
 sky130_fd_sc_hd__nor3_4 _15412_ (.A(net4057),
    .B(_05891_),
    .C(net4049),
    .Y(_06300_));
 sky130_fd_sc_hd__nor3_1 _15413_ (.A(net3709),
    .B(_06026_),
    .C(_06300_),
    .Y(_06301_));
 sky130_fd_sc_hd__a21oi_1 _15414_ (.A1(_06129_),
    .A2(_06166_),
    .B1(net4054),
    .Y(_06302_));
 sky130_fd_sc_hd__nor2_1 _15415_ (.A(_11964_[0]),
    .B(net3709),
    .Y(_06303_));
 sky130_fd_sc_hd__o21a_1 _15416_ (.A1(_05921_),
    .A2(_06303_),
    .B1(net4047),
    .X(_06304_));
 sky130_fd_sc_hd__o32ai_1 _15417_ (.A1(_05958_),
    .A2(_06301_),
    .A3(_06302_),
    .B1(_06304_),
    .B2(_06011_),
    .Y(_06305_));
 sky130_fd_sc_hd__nand2_1 _15418_ (.A(_06059_),
    .B(_06305_),
    .Y(_06306_));
 sky130_fd_sc_hd__o21ai_0 _15419_ (.A1(_06059_),
    .A2(_06299_),
    .B1(_06306_),
    .Y(_06307_));
 sky130_fd_sc_hd__or3_4 _15420_ (.A(_11966_[0]),
    .B(_05931_),
    .C(_05936_),
    .X(_06308_));
 sky130_fd_sc_hd__nand2_1 _15421_ (.A(_11974_[0]),
    .B(net4047),
    .Y(_06309_));
 sky130_fd_sc_hd__nand2_1 _15422_ (.A(net3709),
    .B(_06309_),
    .Y(_06310_));
 sky130_fd_sc_hd__a21oi_1 _15423_ (.A1(_06308_),
    .A2(_06310_),
    .B1(net4040),
    .Y(_06311_));
 sky130_fd_sc_hd__a311oi_1 _15424_ (.A1(net3709),
    .A2(_06160_),
    .A3(_06129_),
    .B1(net4043),
    .C1(_06270_),
    .Y(_06312_));
 sky130_fd_sc_hd__nor3_1 _15425_ (.A(_06035_),
    .B(_06311_),
    .C(_06312_),
    .Y(_06313_));
 sky130_fd_sc_hd__a22oi_1 _15426_ (.A1(_11964_[0]),
    .A2(_06110_),
    .B1(_06247_),
    .B2(net3710),
    .Y(_06314_));
 sky130_fd_sc_hd__a21oi_1 _15427_ (.A1(net4056),
    .A2(_06246_),
    .B1(net4057),
    .Y(_06315_));
 sky130_fd_sc_hd__o21ai_0 _15428_ (.A1(_06270_),
    .A2(_06315_),
    .B1(net4050),
    .Y(_06316_));
 sky130_fd_sc_hd__o21ai_0 _15429_ (.A1(_06024_),
    .A2(_06274_),
    .B1(net4057),
    .Y(_06317_));
 sky130_fd_sc_hd__o2111a_4 _15430_ (.A1(net4050),
    .A2(_06314_),
    .B1(_06316_),
    .C1(_06317_),
    .D1(net3705),
    .X(_06318_));
 sky130_fd_sc_hd__nand3b_1 _15431_ (.A_N(_06209_),
    .B(_06160_),
    .C(net4054),
    .Y(_06319_));
 sky130_fd_sc_hd__or3b_1 _15432_ (.A(net4039),
    .B(_06130_),
    .C_N(_06319_),
    .X(_06320_));
 sky130_fd_sc_hd__nand2_2 _15433_ (.A(net4054),
    .B(net4049),
    .Y(_06321_));
 sky130_fd_sc_hd__o221ai_1 _15434_ (.A1(_05891_),
    .A2(_06321_),
    .B1(_06210_),
    .B2(net4054),
    .C1(net4039),
    .Y(_06322_));
 sky130_fd_sc_hd__a21oi_1 _15435_ (.A1(_11969_[0]),
    .A2(net4054),
    .B1(_06076_),
    .Y(_06323_));
 sky130_fd_sc_hd__o21ai_1 _15436_ (.A1(_05945_),
    .A2(_06323_),
    .B1(_05956_),
    .Y(_06324_));
 sky130_fd_sc_hd__a31oi_1 _15437_ (.A1(_06015_),
    .A2(_06150_),
    .A3(_06110_),
    .B1(_06035_),
    .Y(_06325_));
 sky130_fd_sc_hd__a32o_1 _15438_ (.A1(_06035_),
    .A2(_06320_),
    .A3(_06322_),
    .B1(_06324_),
    .B2(_06325_),
    .X(_06326_));
 sky130_fd_sc_hd__o32ai_1 _15439_ (.A1(_06143_),
    .A2(_06313_),
    .A3(_06318_),
    .B1(_06326_),
    .B2(_05989_),
    .Y(_06327_));
 sky130_fd_sc_hd__nand3_1 _15440_ (.A(net3709),
    .B(_06028_),
    .C(_06152_),
    .Y(_06328_));
 sky130_fd_sc_hd__o211ai_1 _15441_ (.A1(_11974_[0]),
    .A2(net3709),
    .B1(_06059_),
    .C1(_06328_),
    .Y(_06329_));
 sky130_fd_sc_hd__nand2_1 _15442_ (.A(net4057),
    .B(_05991_),
    .Y(_06330_));
 sky130_fd_sc_hd__nand3_4 _15443_ (.A(net3710),
    .B(net4056),
    .C(net4050),
    .Y(_06331_));
 sky130_fd_sc_hd__nand4_1 _15444_ (.A(_05978_),
    .B(_06310_),
    .C(_06330_),
    .D(_06331_),
    .Y(_06332_));
 sky130_fd_sc_hd__nor3_1 _15445_ (.A(_05900_),
    .B(_06210_),
    .C(_06300_),
    .Y(_06333_));
 sky130_fd_sc_hd__nor3_1 _15446_ (.A(net4054),
    .B(net3624),
    .C(_06184_),
    .Y(_06334_));
 sky130_fd_sc_hd__o21ai_1 _15447_ (.A1(_06333_),
    .A2(_06334_),
    .B1(_06059_),
    .Y(_06335_));
 sky130_fd_sc_hd__nor3_1 _15448_ (.A(_06083_),
    .B(net4054),
    .C(net4050),
    .Y(_06336_));
 sky130_fd_sc_hd__a21oi_1 _15449_ (.A1(_11976_[0]),
    .A2(net4050),
    .B1(_06336_),
    .Y(_06337_));
 sky130_fd_sc_hd__a21oi_1 _15450_ (.A1(_05978_),
    .A2(_06337_),
    .B1(net4043),
    .Y(_06338_));
 sky130_fd_sc_hd__a32oi_1 _15451_ (.A1(net4043),
    .A2(_06329_),
    .A3(_06332_),
    .B1(_06335_),
    .B2(_06338_),
    .Y(_06339_));
 sky130_fd_sc_hd__nor3_1 _15452_ (.A(_06035_),
    .B(net3707),
    .C(_06339_),
    .Y(_06340_));
 sky130_fd_sc_hd__a211oi_1 _15453_ (.A1(_06072_),
    .A2(_06307_),
    .B1(_06327_),
    .C1(_06340_),
    .Y(_00036_));
 sky130_fd_sc_hd__o21ai_0 _15454_ (.A1(_11964_[0]),
    .A2(net4052),
    .B1(_06166_),
    .Y(_06341_));
 sky130_fd_sc_hd__nor2_2 _15455_ (.A(net3636),
    .B(_05963_),
    .Y(_06342_));
 sky130_fd_sc_hd__a21oi_1 _15456_ (.A1(_05900_),
    .A2(_06341_),
    .B1(_06342_),
    .Y(_06343_));
 sky130_fd_sc_hd__nand2_1 _15457_ (.A(net4041),
    .B(_06343_),
    .Y(_06344_));
 sky130_fd_sc_hd__nand2_1 _15458_ (.A(_06015_),
    .B(_06028_),
    .Y(_06345_));
 sky130_fd_sc_hd__nand2_1 _15459_ (.A(_05900_),
    .B(_06345_),
    .Y(_06346_));
 sky130_fd_sc_hd__a31oi_1 _15460_ (.A1(net4042),
    .A2(_06282_),
    .A3(_06346_),
    .B1(net3708),
    .Y(_06347_));
 sky130_fd_sc_hd__a211oi_1 _15461_ (.A1(_05954_),
    .A2(_05991_),
    .B1(_06111_),
    .C1(net4057),
    .Y(_06348_));
 sky130_fd_sc_hd__a21oi_1 _15462_ (.A1(net4057),
    .A2(_06115_),
    .B1(_06348_),
    .Y(_06349_));
 sky130_fd_sc_hd__a221oi_1 _15463_ (.A1(net4056),
    .A2(_06063_),
    .B1(_06066_),
    .B2(_11972_[0]),
    .C1(net4041),
    .Y(_06350_));
 sky130_fd_sc_hd__a21oi_1 _15464_ (.A1(net4058),
    .A2(_06056_),
    .B1(net4043),
    .Y(_06351_));
 sky130_fd_sc_hd__o21ai_0 _15465_ (.A1(_06350_),
    .A2(_06351_),
    .B1(_05917_),
    .Y(_06352_));
 sky130_fd_sc_hd__a21oi_2 _15466_ (.A1(_05891_),
    .A2(_06349_),
    .B1(_06352_),
    .Y(_06353_));
 sky130_fd_sc_hd__a21oi_2 _15467_ (.A1(_06344_),
    .A2(_06347_),
    .B1(_06353_),
    .Y(_06354_));
 sky130_fd_sc_hd__o21ai_0 _15468_ (.A1(net4045),
    .A2(_05947_),
    .B1(_06085_),
    .Y(_06355_));
 sky130_fd_sc_hd__a32oi_1 _15469_ (.A1(_06188_),
    .A2(_06134_),
    .A3(_06114_),
    .B1(_06238_),
    .B2(_05991_),
    .Y(_06356_));
 sky130_fd_sc_hd__nor2_1 _15470_ (.A(net3706),
    .B(_06356_),
    .Y(_06357_));
 sky130_fd_sc_hd__a21oi_1 _15471_ (.A1(net3706),
    .A2(_06355_),
    .B1(_06357_),
    .Y(_06358_));
 sky130_fd_sc_hd__nand3_1 _15472_ (.A(_05900_),
    .B(_06085_),
    .C(_06183_),
    .Y(_06359_));
 sky130_fd_sc_hd__nand3_1 _15473_ (.A(net4054),
    .B(_06075_),
    .C(_06151_),
    .Y(_06360_));
 sky130_fd_sc_hd__nand3_1 _15474_ (.A(_06035_),
    .B(_06359_),
    .C(_06360_),
    .Y(_06361_));
 sky130_fd_sc_hd__o21ai_0 _15475_ (.A1(net3598),
    .A2(net4054),
    .B1(net4045),
    .Y(_06362_));
 sky130_fd_sc_hd__nand2_1 _15476_ (.A(_11969_[0]),
    .B(_06019_),
    .Y(_06363_));
 sky130_fd_sc_hd__a31oi_1 _15477_ (.A1(net3708),
    .A2(_06362_),
    .A3(_06363_),
    .B1(net4039),
    .Y(_06364_));
 sky130_fd_sc_hd__a221oi_1 _15478_ (.A1(net4039),
    .A2(_06358_),
    .B1(_06361_),
    .B2(_06364_),
    .C1(_06095_),
    .Y(_06365_));
 sky130_fd_sc_hd__o21ai_0 _15479_ (.A1(_11974_[0]),
    .A2(net4045),
    .B1(_05900_),
    .Y(_06366_));
 sky130_fd_sc_hd__a31oi_1 _15480_ (.A1(net4054),
    .A2(_05992_),
    .A3(_06151_),
    .B1(net3706),
    .Y(_06367_));
 sky130_fd_sc_hd__o21ai_0 _15481_ (.A1(_06300_),
    .A2(_06366_),
    .B1(_06367_),
    .Y(_06368_));
 sky130_fd_sc_hd__o211ai_1 _15482_ (.A1(_06147_),
    .A2(_06321_),
    .B1(_06359_),
    .C1(_06035_),
    .Y(_06369_));
 sky130_fd_sc_hd__and3_4 _15483_ (.A(net4042),
    .B(_06368_),
    .C(_06369_),
    .X(_06370_));
 sky130_fd_sc_hd__nand2_1 _15484_ (.A(_05991_),
    .B(_06147_),
    .Y(_06371_));
 sky130_fd_sc_hd__o221ai_1 _15485_ (.A1(_11969_[0]),
    .A2(_06056_),
    .B1(_06078_),
    .B2(_05891_),
    .C1(_06371_),
    .Y(_06372_));
 sky130_fd_sc_hd__o21ai_0 _15486_ (.A1(net4056),
    .A2(_06063_),
    .B1(_06331_),
    .Y(_06373_));
 sky130_fd_sc_hd__o21ai_0 _15487_ (.A1(net3706),
    .A2(_06373_),
    .B1(net4040),
    .Y(_06374_));
 sky130_fd_sc_hd__a21oi_1 _15488_ (.A1(net3706),
    .A2(_06372_),
    .B1(_06374_),
    .Y(_06375_));
 sky130_fd_sc_hd__a221oi_1 _15489_ (.A1(_11969_[0]),
    .A2(_05945_),
    .B1(_06019_),
    .B2(_11974_[0]),
    .C1(_06053_),
    .Y(_06376_));
 sky130_fd_sc_hd__nor2_1 _15490_ (.A(_05978_),
    .B(_06047_),
    .Y(_06377_));
 sky130_fd_sc_hd__o21ai_0 _15491_ (.A1(_06175_),
    .A2(_06376_),
    .B1(_06377_),
    .Y(_06378_));
 sky130_fd_sc_hd__nand2_1 _15492_ (.A(_05900_),
    .B(_06156_),
    .Y(_06379_));
 sky130_fd_sc_hd__a211oi_1 _15493_ (.A1(net4054),
    .A2(_06152_),
    .B1(_06300_),
    .C1(net4040),
    .Y(_06380_));
 sky130_fd_sc_hd__a31oi_1 _15494_ (.A1(net4040),
    .A2(_06262_),
    .A3(_06379_),
    .B1(_06380_),
    .Y(_06381_));
 sky130_fd_sc_hd__a31oi_1 _15495_ (.A1(_05900_),
    .A2(_05992_),
    .A3(_05994_),
    .B1(net4042),
    .Y(_06382_));
 sky130_fd_sc_hd__a21oi_1 _15496_ (.A1(_06045_),
    .A2(_06382_),
    .B1(net3706),
    .Y(_06383_));
 sky130_fd_sc_hd__a21oi_1 _15497_ (.A1(net3706),
    .A2(_06381_),
    .B1(_06383_),
    .Y(_06384_));
 sky130_fd_sc_hd__o32ai_1 _15498_ (.A1(_05989_),
    .A2(_06370_),
    .A3(_06375_),
    .B1(_06378_),
    .B2(_06384_),
    .Y(_06385_));
 sky130_fd_sc_hd__a311oi_1 _15499_ (.A1(_06059_),
    .A2(_06047_),
    .A3(_06354_),
    .B1(_06365_),
    .C1(_06385_),
    .Y(_00037_));
 sky130_fd_sc_hd__nor2_1 _15500_ (.A(_06178_),
    .B(_06300_),
    .Y(_06386_));
 sky130_fd_sc_hd__nor2_1 _15501_ (.A(net4054),
    .B(_06386_),
    .Y(_06387_));
 sky130_fd_sc_hd__o21ai_0 _15502_ (.A1(net3636),
    .A2(_05900_),
    .B1(net4049),
    .Y(_06388_));
 sky130_fd_sc_hd__a21oi_1 _15503_ (.A1(_05900_),
    .A2(_06062_),
    .B1(_06388_),
    .Y(_06389_));
 sky130_fd_sc_hd__o21ai_0 _15504_ (.A1(_06233_),
    .A2(_06389_),
    .B1(net4042),
    .Y(_06390_));
 sky130_fd_sc_hd__o311ai_0 _15505_ (.A1(net4042),
    .A2(_06286_),
    .A3(_06387_),
    .B1(_06390_),
    .C1(net3708),
    .Y(_06391_));
 sky130_fd_sc_hd__a21oi_1 _15506_ (.A1(_06084_),
    .A2(_06023_),
    .B1(net4054),
    .Y(_06392_));
 sky130_fd_sc_hd__nor3_1 _15507_ (.A(_05900_),
    .B(net4044),
    .C(_06238_),
    .Y(_06393_));
 sky130_fd_sc_hd__nor4_1 _15508_ (.A(net4042),
    .B(_06092_),
    .C(_06392_),
    .D(_06393_),
    .Y(_06394_));
 sky130_fd_sc_hd__a21oi_1 _15509_ (.A1(net3710),
    .A2(_06090_),
    .B1(net4049),
    .Y(_06395_));
 sky130_fd_sc_hd__nor3_1 _15510_ (.A(net4039),
    .B(_06057_),
    .C(_06395_),
    .Y(_06396_));
 sky130_fd_sc_hd__o21ai_1 _15511_ (.A1(_06394_),
    .A2(_06396_),
    .B1(net3706),
    .Y(_06397_));
 sky130_fd_sc_hd__a21oi_2 _15512_ (.A1(_06391_),
    .A2(_06397_),
    .B1(_05988_),
    .Y(_06398_));
 sky130_fd_sc_hd__a21oi_1 _15513_ (.A1(_11966_[0]),
    .A2(_05945_),
    .B1(_06167_),
    .Y(_06399_));
 sky130_fd_sc_hd__a311oi_1 _15514_ (.A1(net3709),
    .A2(_06029_),
    .A3(_06150_),
    .B1(_06399_),
    .C1(net4043),
    .Y(_06400_));
 sky130_fd_sc_hd__nor3_1 _15515_ (.A(net4055),
    .B(net3624),
    .C(_06239_),
    .Y(_06401_));
 sky130_fd_sc_hd__a311oi_1 _15516_ (.A1(net4055),
    .A2(_06131_),
    .A3(_06309_),
    .B1(_06401_),
    .C1(net4040),
    .Y(_06402_));
 sky130_fd_sc_hd__o21ai_0 _15517_ (.A1(_11964_[0]),
    .A2(net4047),
    .B1(_06309_),
    .Y(_06403_));
 sky130_fd_sc_hd__a22oi_1 _15518_ (.A1(_11966_[0]),
    .A2(_06066_),
    .B1(_06403_),
    .B2(net4055),
    .Y(_06404_));
 sky130_fd_sc_hd__a21oi_1 _15519_ (.A1(net4057),
    .A2(net4054),
    .B1(_06150_),
    .Y(_06405_));
 sky130_fd_sc_hd__o31ai_1 _15520_ (.A1(_11981_[0]),
    .A2(_11990_[0]),
    .A3(net4047),
    .B1(net4040),
    .Y(_06406_));
 sky130_fd_sc_hd__o221ai_1 _15521_ (.A1(net4040),
    .A2(_06404_),
    .B1(_06405_),
    .B2(_06406_),
    .C1(_06229_),
    .Y(_06407_));
 sky130_fd_sc_hd__o311ai_0 _15522_ (.A1(_06037_),
    .A2(_06400_),
    .A3(_06402_),
    .B1(_06407_),
    .C1(_06059_),
    .Y(_06408_));
 sky130_fd_sc_hd__nand2_1 _15523_ (.A(net3636),
    .B(_06111_),
    .Y(_06409_));
 sky130_fd_sc_hd__o21ai_0 _15524_ (.A1(_11974_[0]),
    .A2(_05954_),
    .B1(_05945_),
    .Y(_06410_));
 sky130_fd_sc_hd__nor3b_1 _15525_ (.A(net4054),
    .B(_06024_),
    .C_N(_06251_),
    .Y(_06411_));
 sky130_fd_sc_hd__a31oi_1 _15526_ (.A1(net4054),
    .A2(_06409_),
    .A3(_06410_),
    .B1(_06411_),
    .Y(_06412_));
 sky130_fd_sc_hd__o21ai_0 _15527_ (.A1(net4040),
    .A2(_06159_),
    .B1(net3707),
    .Y(_06413_));
 sky130_fd_sc_hd__a21oi_1 _15528_ (.A1(_11972_[0]),
    .A2(net4049),
    .B1(_06184_),
    .Y(_06414_));
 sky130_fd_sc_hd__o211ai_1 _15529_ (.A1(net4055),
    .A2(_06414_),
    .B1(_06330_),
    .C1(_05954_),
    .Y(_06415_));
 sky130_fd_sc_hd__a311oi_1 _15530_ (.A1(_06047_),
    .A2(_06195_),
    .A3(_06415_),
    .B1(_06059_),
    .C1(net3708),
    .Y(_06416_));
 sky130_fd_sc_hd__o21ai_0 _15531_ (.A1(_06412_),
    .A2(_06413_),
    .B1(_06416_),
    .Y(_06417_));
 sky130_fd_sc_hd__o21ai_0 _15532_ (.A1(net4039),
    .A2(_06210_),
    .B1(net4054),
    .Y(_06418_));
 sky130_fd_sc_hd__o21ai_0 _15533_ (.A1(_05891_),
    .A2(net4042),
    .B1(_06418_),
    .Y(_06419_));
 sky130_fd_sc_hd__a31oi_1 _15534_ (.A1(net4057),
    .A2(net4056),
    .A3(net4055),
    .B1(_05997_),
    .Y(_06420_));
 sky130_fd_sc_hd__o221ai_1 _15535_ (.A1(net3710),
    .A2(_06023_),
    .B1(_06420_),
    .B2(net3598),
    .C1(_06114_),
    .Y(_06421_));
 sky130_fd_sc_hd__nor2_1 _15536_ (.A(_06090_),
    .B(_06220_),
    .Y(_06422_));
 sky130_fd_sc_hd__a221oi_1 _15537_ (.A1(net3710),
    .A2(_06419_),
    .B1(_06421_),
    .B2(net4042),
    .C1(_06422_),
    .Y(_06423_));
 sky130_fd_sc_hd__a211oi_1 _15538_ (.A1(_11974_[0]),
    .A2(_05900_),
    .B1(_05945_),
    .C1(_06144_),
    .Y(_06424_));
 sky130_fd_sc_hd__nand2_1 _15539_ (.A(_11982_[0]),
    .B(net4047),
    .Y(_06425_));
 sky130_fd_sc_hd__nand2_1 _15540_ (.A(net4040),
    .B(_06425_),
    .Y(_06426_));
 sky130_fd_sc_hd__o21ai_2 _15541_ (.A1(_06342_),
    .A2(_06279_),
    .B1(net4043),
    .Y(_06427_));
 sky130_fd_sc_hd__o211ai_1 _15542_ (.A1(_06424_),
    .A2(_06426_),
    .B1(_06427_),
    .C1(_06047_),
    .Y(_06428_));
 sky130_fd_sc_hd__o2111ai_1 _15543_ (.A1(_06047_),
    .A2(_06423_),
    .B1(_06428_),
    .C1(net3708),
    .D1(_05978_),
    .Y(_06429_));
 sky130_fd_sc_hd__o211ai_1 _15544_ (.A1(_06398_),
    .A2(_06408_),
    .B1(_06417_),
    .C1(_06429_),
    .Y(_00038_));
 sky130_fd_sc_hd__nand2_1 _15545_ (.A(_06147_),
    .B(_06066_),
    .Y(_06430_));
 sky130_fd_sc_hd__a221oi_1 _15546_ (.A1(_11964_[0]),
    .A2(_05991_),
    .B1(_06019_),
    .B2(net4056),
    .C1(net3705),
    .Y(_06431_));
 sky130_fd_sc_hd__nand3_1 _15547_ (.A(_06331_),
    .B(_06430_),
    .C(_06431_),
    .Y(_06432_));
 sky130_fd_sc_hd__o221ai_1 _15548_ (.A1(_11978_[0]),
    .A2(_05963_),
    .B1(_06078_),
    .B2(net3636),
    .C1(_06171_),
    .Y(_06433_));
 sky130_fd_sc_hd__nand3_1 _15549_ (.A(net4043),
    .B(_06432_),
    .C(_06433_),
    .Y(_06434_));
 sky130_fd_sc_hd__nor3_1 _15550_ (.A(_11974_[0]),
    .B(net4054),
    .C(net4050),
    .Y(_06435_));
 sky130_fd_sc_hd__a31oi_1 _15551_ (.A1(net4054),
    .A2(_06129_),
    .A3(_06166_),
    .B1(_06435_),
    .Y(_06436_));
 sky130_fd_sc_hd__nor2_1 _15552_ (.A(_06035_),
    .B(_06436_),
    .Y(_06437_));
 sky130_fd_sc_hd__nand4_1 _15553_ (.A(net3709),
    .B(net3705),
    .C(_06029_),
    .D(_06129_),
    .Y(_06438_));
 sky130_fd_sc_hd__o31ai_1 _15554_ (.A1(_05917_),
    .A2(_06156_),
    .A3(_06167_),
    .B1(_06438_),
    .Y(_06439_));
 sky130_fd_sc_hd__o21ai_0 _15555_ (.A1(_06437_),
    .A2(_06439_),
    .B1(_05958_),
    .Y(_06440_));
 sky130_fd_sc_hd__a21oi_1 _15556_ (.A1(_06434_),
    .A2(_06440_),
    .B1(_06047_),
    .Y(_06441_));
 sky130_fd_sc_hd__nand3_1 _15557_ (.A(_06035_),
    .B(_05978_),
    .C(_06246_),
    .Y(_06442_));
 sky130_fd_sc_hd__nor2_2 _15558_ (.A(_05900_),
    .B(_06075_),
    .Y(_06443_));
 sky130_fd_sc_hd__o21ai_0 _15559_ (.A1(net4056),
    .A2(_05954_),
    .B1(_05945_),
    .Y(_06444_));
 sky130_fd_sc_hd__a21oi_1 _15560_ (.A1(net4056),
    .A2(_06274_),
    .B1(_06444_),
    .Y(_06445_));
 sky130_fd_sc_hd__a211oi_1 _15561_ (.A1(net4051),
    .A2(_06114_),
    .B1(_06445_),
    .C1(net4058),
    .Y(_06446_));
 sky130_fd_sc_hd__o21ai_0 _15562_ (.A1(_06156_),
    .A2(_06019_),
    .B1(net4057),
    .Y(_06447_));
 sky130_fd_sc_hd__a21oi_1 _15563_ (.A1(_06331_),
    .A2(_06447_),
    .B1(_05954_),
    .Y(_06448_));
 sky130_fd_sc_hd__a21oi_1 _15564_ (.A1(net4056),
    .A2(_05991_),
    .B1(_05997_),
    .Y(_06449_));
 sky130_fd_sc_hd__a21oi_1 _15565_ (.A1(net4050),
    .A2(_06270_),
    .B1(_06066_),
    .Y(_06450_));
 sky130_fd_sc_hd__o22ai_1 _15566_ (.A1(net4041),
    .A2(_06449_),
    .B1(_06450_),
    .B2(net4058),
    .Y(_06451_));
 sky130_fd_sc_hd__o21ai_0 _15567_ (.A1(_06448_),
    .A2(_06451_),
    .B1(_05917_),
    .Y(_06452_));
 sky130_fd_sc_hd__o311a_1 _15568_ (.A1(_06442_),
    .A2(_06443_),
    .A3(_06446_),
    .B1(_06452_),
    .C1(_06047_),
    .X(_06453_));
 sky130_fd_sc_hd__nand3_1 _15569_ (.A(_05900_),
    .B(_06085_),
    .C(_06086_),
    .Y(_06454_));
 sky130_fd_sc_hd__nand3_1 _15570_ (.A(net4054),
    .B(_06028_),
    .C(_06160_),
    .Y(_06455_));
 sky130_fd_sc_hd__o21ai_0 _15571_ (.A1(_11976_[0]),
    .A2(net4050),
    .B1(_06047_),
    .Y(_06456_));
 sky130_fd_sc_hd__a31oi_1 _15572_ (.A1(_11966_[0]),
    .A2(net3709),
    .A3(net4050),
    .B1(_06456_),
    .Y(_06457_));
 sky130_fd_sc_hd__a311oi_1 _15573_ (.A1(net3707),
    .A2(_06454_),
    .A3(_06455_),
    .B1(_06457_),
    .C1(net4043),
    .Y(_06458_));
 sky130_fd_sc_hd__nor3_1 _15574_ (.A(_06270_),
    .B(net3707),
    .C(_06000_),
    .Y(_06459_));
 sky130_fd_sc_hd__nor3_1 _15575_ (.A(net4055),
    .B(_05997_),
    .C(_06184_),
    .Y(_06460_));
 sky130_fd_sc_hd__nand2_1 _15576_ (.A(_05988_),
    .B(_05992_),
    .Y(_06461_));
 sky130_fd_sc_hd__a211oi_1 _15577_ (.A1(net4055),
    .A2(_06239_),
    .B1(_06460_),
    .C1(_06461_),
    .Y(_06462_));
 sky130_fd_sc_hd__nand3_1 _15578_ (.A(net4044),
    .B(_06047_),
    .C(_06199_),
    .Y(_06463_));
 sky130_fd_sc_hd__nor2_1 _15579_ (.A(_05921_),
    .B(_06463_),
    .Y(_06464_));
 sky130_fd_sc_hd__nor4_1 _15580_ (.A(net4040),
    .B(_06459_),
    .C(_06462_),
    .D(_06464_),
    .Y(_06465_));
 sky130_fd_sc_hd__o21bai_1 _15581_ (.A1(_06458_),
    .A2(_06465_),
    .B1_N(_06060_),
    .Y(_06466_));
 sky130_fd_sc_hd__nor2_1 _15582_ (.A(net4054),
    .B(_06176_),
    .Y(_06467_));
 sky130_fd_sc_hd__a311oi_1 _15583_ (.A1(net4054),
    .A2(_06000_),
    .A3(_06151_),
    .B1(_06467_),
    .C1(_05988_),
    .Y(_06468_));
 sky130_fd_sc_hd__nor3_1 _15584_ (.A(_06047_),
    .B(_06026_),
    .C(_06405_),
    .Y(_06469_));
 sky130_fd_sc_hd__a31oi_1 _15585_ (.A1(net3709),
    .A2(_06308_),
    .A3(_06129_),
    .B1(_06303_),
    .Y(_06470_));
 sky130_fd_sc_hd__a211oi_1 _15586_ (.A1(_11974_[0]),
    .A2(net4054),
    .B1(_05945_),
    .C1(_06076_),
    .Y(_06471_));
 sky130_fd_sc_hd__o21ai_0 _15587_ (.A1(_11990_[0]),
    .A2(net4048),
    .B1(_06047_),
    .Y(_06472_));
 sky130_fd_sc_hd__o221ai_1 _15588_ (.A1(_06047_),
    .A2(_06470_),
    .B1(_06471_),
    .B2(_06472_),
    .C1(_05958_),
    .Y(_06473_));
 sky130_fd_sc_hd__o311ai_0 _15589_ (.A1(_05958_),
    .A2(_06468_),
    .A3(_06469_),
    .B1(_06006_),
    .C1(_06473_),
    .Y(_06474_));
 sky130_fd_sc_hd__o311ai_0 _15590_ (.A1(_06059_),
    .A2(_06441_),
    .A3(_06453_),
    .B1(_06466_),
    .C1(_06474_),
    .Y(_00039_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_991 ();
 sky130_fd_sc_hd__xnor2_1 _15593_ (.A(\sa01_sr[7] ),
    .B(\sa01_sr[0] ),
    .Y(_06477_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_990 ();
 sky130_fd_sc_hd__xnor2_1 _15595_ (.A(\sa21_sr[1] ),
    .B(\sa30_sub[1] ),
    .Y(_06479_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_989 ();
 sky130_fd_sc_hd__xnor3_1 _15597_ (.A(\sa11_sr[7] ),
    .B(net4215),
    .C(\sa11_sr[1] ),
    .X(_06481_));
 sky130_fd_sc_hd__xnor3_1 _15598_ (.A(_06477_),
    .B(_06479_),
    .C(_06481_),
    .X(_06482_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_987 ();
 sky130_fd_sc_hd__mux2i_4 _15601_ (.A0(\text_in_r[89] ),
    .A1(_06482_),
    .S(net4117),
    .Y(_06485_));
 sky130_fd_sc_hd__xor2_4 _15602_ (.A(net4150),
    .B(_06485_),
    .X(_06486_));
 sky130_fd_sc_hd__clkinvlp_4 _15603_ (.A(_06486_),
    .Y(_06487_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_985 ();
 sky130_fd_sc_hd__xor2_2 _15606_ (.A(\sa11_sr[0] ),
    .B(\sa21_sr[0] ),
    .X(_06489_));
 sky130_fd_sc_hd__xnor3_1 _15607_ (.A(\sa01_sr[7] ),
    .B(\sa11_sr[7] ),
    .C(\sa30_sub[0] ),
    .X(_06490_));
 sky130_fd_sc_hd__xnor2_1 _15608_ (.A(_06489_),
    .B(_06490_),
    .Y(_06491_));
 sky130_fd_sc_hd__mux2i_2 _15609_ (.A0(\text_in_r[88] ),
    .A1(_06491_),
    .S(net4117),
    .Y(_06492_));
 sky130_fd_sc_hd__xor2_4 _15610_ (.A(net4151),
    .B(_06492_),
    .X(_06493_));
 sky130_fd_sc_hd__clkinv_16 _15611_ (.A(_06493_),
    .Y(_06494_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_984 ();
 sky130_fd_sc_hd__xnor3_1 _15613_ (.A(net4227),
    .B(\sa11_sr[2] ),
    .C(net4205),
    .X(_06495_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_983 ();
 sky130_fd_sc_hd__xnor2_1 _15615_ (.A(\sa11_sr[1] ),
    .B(\sa30_sub[2] ),
    .Y(_06497_));
 sky130_fd_sc_hd__xor2_1 _15616_ (.A(_06495_),
    .B(_06497_),
    .X(_06498_));
 sky130_fd_sc_hd__nand2b_1 _15617_ (.A_N(\text_in_r[90] ),
    .B(net4230),
    .Y(_06499_));
 sky130_fd_sc_hd__o211ai_1 _15618_ (.A1(net398),
    .A2(_06498_),
    .B1(_06499_),
    .C1(net4149),
    .Y(_06500_));
 sky130_fd_sc_hd__and2_0 _15619_ (.A(net4230),
    .B(\text_in_r[90] ),
    .X(_06501_));
 sky130_fd_sc_hd__a211o_1 _15620_ (.A1(net4117),
    .A2(_06498_),
    .B1(_06501_),
    .C1(net4149),
    .X(_06502_));
 sky130_fd_sc_hd__and2_4 _15621_ (.A(_06500_),
    .B(_06502_),
    .X(_06503_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_982 ();
 sky130_fd_sc_hd__clkinv_16 _15623_ (.A(_06503_),
    .Y(_06505_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_973 ();
 sky130_fd_sc_hd__xnor3_1 _15633_ (.A(\sa01_sr[7] ),
    .B(\sa01_sr[3] ),
    .C(\sa21_sr[4] ),
    .X(_06512_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_972 ();
 sky130_fd_sc_hd__xnor2_1 _15635_ (.A(net4214),
    .B(\sa30_sub[4] ),
    .Y(_06514_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_970 ();
 sky130_fd_sc_hd__xnor2_1 _15638_ (.A(\sa11_sr[3] ),
    .B(\sa11_sr[4] ),
    .Y(_06517_));
 sky130_fd_sc_hd__xnor3_1 _15639_ (.A(_06512_),
    .B(_06514_),
    .C(_06517_),
    .X(_06518_));
 sky130_fd_sc_hd__mux2i_4 _15640_ (.A0(\text_in_r[92] ),
    .A1(_06518_),
    .S(net4120),
    .Y(_06519_));
 sky130_fd_sc_hd__xor2_1 _15641_ (.A(\u0.w[1][28] ),
    .B(_06519_),
    .X(_06520_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_964 ();
 sky130_fd_sc_hd__xnor3_1 _15648_ (.A(\sa01_sr[7] ),
    .B(\sa01_sr[2] ),
    .C(\sa21_sr[3] ),
    .X(_06527_));
 sky130_fd_sc_hd__xnor2_1 _15649_ (.A(\sa11_sr[7] ),
    .B(\sa11_sr[2] ),
    .Y(_06528_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_963 ();
 sky130_fd_sc_hd__xnor2_1 _15651_ (.A(\sa11_sr[3] ),
    .B(net4188),
    .Y(_06530_));
 sky130_fd_sc_hd__xnor3_1 _15652_ (.A(_06527_),
    .B(_06528_),
    .C(_06530_),
    .X(_06531_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_962 ();
 sky130_fd_sc_hd__and2_4 _15654_ (.A(net4230),
    .B(\text_in_r[91] ),
    .X(_06533_));
 sky130_fd_sc_hd__a211oi_4 _15655_ (.A1(net4120),
    .A2(_06531_),
    .B1(_06533_),
    .C1(net4148),
    .Y(_06534_));
 sky130_fd_sc_hd__nor2b_1 _15656_ (.A(net4230),
    .B_N(\u0.w[1][27] ),
    .Y(_06535_));
 sky130_fd_sc_hd__a22o_4 _15657_ (.A1(net4148),
    .A2(_06533_),
    .B1(_06535_),
    .B2(_06531_),
    .X(_06536_));
 sky130_fd_sc_hd__or2_4 _15658_ (.A(_06536_),
    .B(_06534_),
    .X(_06537_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_960 ();
 sky130_fd_sc_hd__nor2_2 _15661_ (.A(_06505_),
    .B(_06537_),
    .Y(_06540_));
 sky130_fd_sc_hd__nor2_4 _15662_ (.A(_06534_),
    .B(_06536_),
    .Y(_06541_));
 sky130_fd_sc_hd__nor2_1 _15663_ (.A(net4035),
    .B(_06541_),
    .Y(_06542_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_955 ();
 sky130_fd_sc_hd__mux2i_1 _15669_ (.A0(_12010_[0]),
    .A1(net4037),
    .S(net4031),
    .Y(_06548_));
 sky130_fd_sc_hd__nor2_1 _15670_ (.A(net4033),
    .B(_06548_),
    .Y(_06549_));
 sky130_fd_sc_hd__a211oi_1 _15671_ (.A1(net3635),
    .A2(net3623),
    .B1(net3699),
    .C1(_06549_),
    .Y(_06550_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_953 ();
 sky130_fd_sc_hd__nand2_8 _15674_ (.A(net4033),
    .B(_06541_),
    .Y(_06553_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_951 ();
 sky130_fd_sc_hd__nand2_2 _15677_ (.A(net4035),
    .B(net3700),
    .Y(_06556_));
 sky130_fd_sc_hd__nor2_4 _15678_ (.A(net3704),
    .B(net4027),
    .Y(_06557_));
 sky130_fd_sc_hd__o221ai_1 _15679_ (.A1(_12001_[0]),
    .A2(_06553_),
    .B1(_06556_),
    .B2(_06557_),
    .C1(net4032),
    .Y(_06558_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_950 ();
 sky130_fd_sc_hd__xnor3_1 _15681_ (.A(\sa01_sr[4] ),
    .B(\sa11_sr[5] ),
    .C(\sa21_sr[5] ),
    .X(_06560_));
 sky130_fd_sc_hd__xor2_1 _15682_ (.A(\sa11_sr[4] ),
    .B(\sa30_sub[5] ),
    .X(_06561_));
 sky130_fd_sc_hd__xnor2_1 _15683_ (.A(_06560_),
    .B(_06561_),
    .Y(_06562_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_949 ();
 sky130_fd_sc_hd__mux2i_4 _15685_ (.A0(\text_in_r[93] ),
    .A1(_06562_),
    .S(net4120),
    .Y(_06564_));
 sky130_fd_sc_hd__xnor2_4 _15686_ (.A(net4146),
    .B(_06564_),
    .Y(_06565_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_947 ();
 sky130_fd_sc_hd__o211ai_1 _15689_ (.A1(net4032),
    .A2(_06550_),
    .B1(_06558_),
    .C1(net4020),
    .Y(_06568_));
 sky130_fd_sc_hd__xnor2_4 _15690_ (.A(net4147),
    .B(_06519_),
    .Y(_06569_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_943 ();
 sky130_fd_sc_hd__nor2_4 _15695_ (.A(net4033),
    .B(net4023),
    .Y(_06573_));
 sky130_fd_sc_hd__a21oi_1 _15696_ (.A1(_06494_),
    .A2(net3623),
    .B1(_06573_),
    .Y(_06574_));
 sky130_fd_sc_hd__nand2_8 _15697_ (.A(net4033),
    .B(net399),
    .Y(_06575_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_940 ();
 sky130_fd_sc_hd__nor2_4 _15701_ (.A(net4033),
    .B(net4026),
    .Y(_06579_));
 sky130_fd_sc_hd__nand2_1 _15702_ (.A(net4035),
    .B(_06579_),
    .Y(_06580_));
 sky130_fd_sc_hd__o221ai_1 _15703_ (.A1(net4037),
    .A2(_06574_),
    .B1(_06575_),
    .B2(_11998_[0]),
    .C1(_06580_),
    .Y(_06581_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_939 ();
 sky130_fd_sc_hd__nor2_4 _15705_ (.A(net3704),
    .B(net4022),
    .Y(_06583_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_937 ();
 sky130_fd_sc_hd__nand2_2 _15708_ (.A(net3704),
    .B(net4026),
    .Y(_06586_));
 sky130_fd_sc_hd__nand2_8 _15709_ (.A(_12010_[0]),
    .B(net4022),
    .Y(_06587_));
 sky130_fd_sc_hd__nand3_1 _15710_ (.A(net4033),
    .B(_06586_),
    .C(_06587_),
    .Y(_06588_));
 sky130_fd_sc_hd__o211ai_1 _15711_ (.A1(_06556_),
    .A2(_06583_),
    .B1(_06588_),
    .C1(net4017),
    .Y(_06589_));
 sky130_fd_sc_hd__xor2_4 _15712_ (.A(net4146),
    .B(_06564_),
    .X(_06590_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_934 ();
 sky130_fd_sc_hd__o211ai_1 _15716_ (.A1(net4017),
    .A2(_06581_),
    .B1(_06589_),
    .C1(_06590_),
    .Y(_06594_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_933 ();
 sky130_fd_sc_hd__xnor3_1 _15718_ (.A(\sa11_sr[5] ),
    .B(\sa21_sr[6] ),
    .C(\sa30_sub[6] ),
    .X(_06596_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_931 ();
 sky130_fd_sc_hd__xnor2_1 _15721_ (.A(\sa01_sr[5] ),
    .B(\sa11_sr[6] ),
    .Y(_06599_));
 sky130_fd_sc_hd__xnor2_1 _15722_ (.A(_06596_),
    .B(_06599_),
    .Y(_06600_));
 sky130_fd_sc_hd__nor2_2 _15723_ (.A(net398),
    .B(_06600_),
    .Y(_06601_));
 sky130_fd_sc_hd__a21oi_4 _15724_ (.A1(net398),
    .A2(\text_in_r[94] ),
    .B1(_06601_),
    .Y(_06602_));
 sky130_fd_sc_hd__xnor2_4 _15725_ (.A(net4145),
    .B(_06602_),
    .Y(_06603_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_930 ();
 sky130_fd_sc_hd__xnor3_1 _15727_ (.A(net4214),
    .B(\sa01_sr[6] ),
    .C(\sa21_sr[7] ),
    .X(_06605_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_929 ();
 sky130_fd_sc_hd__xnor2_1 _15729_ (.A(\sa11_sr[6] ),
    .B(net4186),
    .Y(_06607_));
 sky130_fd_sc_hd__xnor2_1 _15730_ (.A(_06605_),
    .B(_06607_),
    .Y(_06608_));
 sky130_fd_sc_hd__nor2_2 _15731_ (.A(net398),
    .B(_06608_),
    .Y(_06609_));
 sky130_fd_sc_hd__a21oi_4 _15732_ (.A1(net398),
    .A2(\text_in_r[95] ),
    .B1(_06609_),
    .Y(_06610_));
 sky130_fd_sc_hd__xor2_4 _15733_ (.A(\u0.w[1][31] ),
    .B(_06610_),
    .X(_06611_));
 sky130_fd_sc_hd__nand2_8 _15734_ (.A(_06603_),
    .B(_06611_),
    .Y(_06612_));
 sky130_fd_sc_hd__a21oi_1 _15735_ (.A1(_06568_),
    .A2(_06594_),
    .B1(_06612_),
    .Y(_06613_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_928 ();
 sky130_fd_sc_hd__nand2_8 _15737_ (.A(_06565_),
    .B(net4032),
    .Y(_06615_));
 sky130_fd_sc_hd__nand2b_4 _15738_ (.A_N(_11998_[0]),
    .B(net4027),
    .Y(_06616_));
 sky130_fd_sc_hd__nand3_4 _15739_ (.A(net3704),
    .B(net4035),
    .C(net4022),
    .Y(_06617_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_927 ();
 sky130_fd_sc_hd__a32oi_1 _15741_ (.A1(net4033),
    .A2(_06616_),
    .A3(_06617_),
    .B1(_06579_),
    .B2(_12006_[0]),
    .Y(_06619_));
 sky130_fd_sc_hd__nand2_4 _15742_ (.A(_11998_[0]),
    .B(net4021),
    .Y(_06620_));
 sky130_fd_sc_hd__o21ai_0 _15743_ (.A1(net4037),
    .A2(_06494_),
    .B1(_06537_),
    .Y(_06621_));
 sky130_fd_sc_hd__a21oi_2 _15744_ (.A1(_06620_),
    .A2(_06621_),
    .B1(net3702),
    .Y(_06622_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_925 ();
 sky130_fd_sc_hd__nor3_2 _15747_ (.A(_12004_[0]),
    .B(net4033),
    .C(net4021),
    .Y(_06625_));
 sky130_fd_sc_hd__nand2_8 _15748_ (.A(_06565_),
    .B(_06569_),
    .Y(_06626_));
 sky130_fd_sc_hd__o21bai_1 _15749_ (.A1(_06622_),
    .A2(_06625_),
    .B1_N(_06626_),
    .Y(_06627_));
 sky130_fd_sc_hd__o21ai_0 _15750_ (.A1(_06615_),
    .A2(_06619_),
    .B1(_06627_),
    .Y(_06628_));
 sky130_fd_sc_hd__xor2_4 _15751_ (.A(net4145),
    .B(_06602_),
    .X(_06629_));
 sky130_fd_sc_hd__xnor2_4 _15752_ (.A(\u0.w[1][31] ),
    .B(_06610_),
    .Y(_06630_));
 sky130_fd_sc_hd__nand2_4 _15753_ (.A(_06629_),
    .B(_06630_),
    .Y(_06631_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_923 ();
 sky130_fd_sc_hd__nand2_1 _15756_ (.A(_12017_[0]),
    .B(net4021),
    .Y(_06634_));
 sky130_fd_sc_hd__and2_4 _15757_ (.A(net3635),
    .B(net3702),
    .X(_06635_));
 sky130_fd_sc_hd__nand2_1 _15758_ (.A(net4027),
    .B(_06635_),
    .Y(_06636_));
 sky130_fd_sc_hd__xnor2_2 _15759_ (.A(_06505_),
    .B(net4029),
    .Y(_06637_));
 sky130_fd_sc_hd__nor2_1 _15760_ (.A(net4036),
    .B(_06637_),
    .Y(_06638_));
 sky130_fd_sc_hd__nand2_8 _15761_ (.A(net4038),
    .B(net4029),
    .Y(_06639_));
 sky130_fd_sc_hd__or3_4 _15762_ (.A(_11996_[0]),
    .B(_06534_),
    .C(_06536_),
    .X(_06640_));
 sky130_fd_sc_hd__a21oi_1 _15763_ (.A1(_06639_),
    .A2(_06640_),
    .B1(net3702),
    .Y(_06641_));
 sky130_fd_sc_hd__nand2_8 _15764_ (.A(_06505_),
    .B(net4031),
    .Y(_06642_));
 sky130_fd_sc_hd__nor2_1 _15765_ (.A(_11998_[0]),
    .B(_12001_[0]),
    .Y(_06643_));
 sky130_fd_sc_hd__o21ai_0 _15766_ (.A1(_06642_),
    .A2(net3589),
    .B1(net4032),
    .Y(_06644_));
 sky130_fd_sc_hd__nor3_1 _15767_ (.A(_06638_),
    .B(_06641_),
    .C(_06644_),
    .Y(_06645_));
 sky130_fd_sc_hd__a311oi_1 _15768_ (.A1(net4017),
    .A2(_06634_),
    .A3(_06636_),
    .B1(_06645_),
    .C1(net4020),
    .Y(_06646_));
 sky130_fd_sc_hd__nand2_2 _15769_ (.A(_06494_),
    .B(net4023),
    .Y(_06647_));
 sky130_fd_sc_hd__nand2_4 _15770_ (.A(_12004_[0]),
    .B(net4023),
    .Y(_06648_));
 sky130_fd_sc_hd__nand2_4 _15771_ (.A(net3635),
    .B(net399),
    .Y(_06649_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_922 ();
 sky130_fd_sc_hd__a21oi_1 _15773_ (.A1(_06648_),
    .A2(_06649_),
    .B1(net4033),
    .Y(_06651_));
 sky130_fd_sc_hd__a311o_1 _15774_ (.A1(net4033),
    .A2(_06639_),
    .A3(_06647_),
    .B1(_06651_),
    .C1(_06615_),
    .X(_06652_));
 sky130_fd_sc_hd__a21oi_2 _15775_ (.A1(net3704),
    .A2(_06494_),
    .B1(net399),
    .Y(_06653_));
 sky130_fd_sc_hd__nand2_4 _15776_ (.A(_12001_[0]),
    .B(net399),
    .Y(_06654_));
 sky130_fd_sc_hd__nand3_1 _15777_ (.A(net3701),
    .B(_06647_),
    .C(_06654_),
    .Y(_06655_));
 sky130_fd_sc_hd__nor2_4 _15778_ (.A(net4019),
    .B(_06569_),
    .Y(_06656_));
 sky130_fd_sc_hd__o211ai_1 _15779_ (.A1(net3701),
    .A2(_06653_),
    .B1(_06655_),
    .C1(_06656_),
    .Y(_06657_));
 sky130_fd_sc_hd__nor2_4 _15780_ (.A(net3635),
    .B(net399),
    .Y(_06658_));
 sky130_fd_sc_hd__nor2_2 _15781_ (.A(_12006_[0]),
    .B(net4021),
    .Y(_06659_));
 sky130_fd_sc_hd__o21ai_0 _15782_ (.A1(_06658_),
    .A2(_06659_),
    .B1(net4033),
    .Y(_06660_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_920 ();
 sky130_fd_sc_hd__nor2_4 _15785_ (.A(net4019),
    .B(net4032),
    .Y(_06663_));
 sky130_fd_sc_hd__o211ai_1 _15786_ (.A1(_12001_[0]),
    .A2(_06642_),
    .B1(_06660_),
    .C1(_06663_),
    .Y(_06664_));
 sky130_fd_sc_hd__nor2_4 _15787_ (.A(_11998_[0]),
    .B(net4021),
    .Y(_06665_));
 sky130_fd_sc_hd__nor2_1 _15788_ (.A(_12001_[0]),
    .B(net4027),
    .Y(_06666_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_919 ();
 sky130_fd_sc_hd__o21ai_0 _15790_ (.A1(_06665_),
    .A2(_06666_),
    .B1(net4033),
    .Y(_06668_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_918 ();
 sky130_fd_sc_hd__a21oi_1 _15792_ (.A1(_11996_[0]),
    .A2(_06573_),
    .B1(_06626_),
    .Y(_06670_));
 sky130_fd_sc_hd__nand2_8 _15793_ (.A(_06603_),
    .B(_06630_),
    .Y(_06671_));
 sky130_fd_sc_hd__a21oi_1 _15794_ (.A1(_06668_),
    .A2(_06670_),
    .B1(_06671_),
    .Y(_06672_));
 sky130_fd_sc_hd__nand4_1 _15795_ (.A(_06652_),
    .B(_06657_),
    .C(_06664_),
    .D(_06672_),
    .Y(_06673_));
 sky130_fd_sc_hd__o31ai_1 _15796_ (.A1(_06628_),
    .A2(_06631_),
    .A3(_06646_),
    .B1(_06673_),
    .Y(_06674_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_917 ();
 sky130_fd_sc_hd__nand2_1 _15798_ (.A(net4020),
    .B(net4026),
    .Y(_06676_));
 sky130_fd_sc_hd__nand2_1 _15799_ (.A(_06590_),
    .B(_06541_),
    .Y(_06677_));
 sky130_fd_sc_hd__nand2_1 _15800_ (.A(_06676_),
    .B(_06677_),
    .Y(_06678_));
 sky130_fd_sc_hd__nor3_1 _15801_ (.A(_12004_[0]),
    .B(_06590_),
    .C(net4026),
    .Y(_06679_));
 sky130_fd_sc_hd__a21oi_1 _15802_ (.A1(net3635),
    .A2(_06678_),
    .B1(_06679_),
    .Y(_06680_));
 sky130_fd_sc_hd__nand2_1 _15803_ (.A(_12004_[0]),
    .B(net4016),
    .Y(_06681_));
 sky130_fd_sc_hd__nor2_4 _15804_ (.A(net4038),
    .B(net4036),
    .Y(_06682_));
 sky130_fd_sc_hd__nand2_1 _15805_ (.A(net4020),
    .B(_06682_),
    .Y(_06683_));
 sky130_fd_sc_hd__nand2_2 _15806_ (.A(_06505_),
    .B(net4021),
    .Y(_06684_));
 sky130_fd_sc_hd__o211ai_1 _15807_ (.A1(net3635),
    .A2(net4016),
    .B1(net4027),
    .C1(net4033),
    .Y(_06685_));
 sky130_fd_sc_hd__a21oi_1 _15808_ (.A1(_06684_),
    .A2(_06685_),
    .B1(_11996_[0]),
    .Y(_06686_));
 sky130_fd_sc_hd__a31oi_1 _15809_ (.A1(_06573_),
    .A2(_06681_),
    .A3(_06683_),
    .B1(_06686_),
    .Y(_06687_));
 sky130_fd_sc_hd__o21ai_0 _15810_ (.A1(net3700),
    .A2(_06680_),
    .B1(_06687_),
    .Y(_06688_));
 sky130_fd_sc_hd__nand2_4 _15811_ (.A(_06505_),
    .B(_06565_),
    .Y(_06689_));
 sky130_fd_sc_hd__nor2_1 _15812_ (.A(net4035),
    .B(_06689_),
    .Y(_06690_));
 sky130_fd_sc_hd__a31oi_1 _15813_ (.A1(net3635),
    .A2(net4033),
    .A3(_06590_),
    .B1(_06690_),
    .Y(_06691_));
 sky130_fd_sc_hd__nor2_1 _15814_ (.A(_06494_),
    .B(_06590_),
    .Y(_06692_));
 sky130_fd_sc_hd__o21ai_0 _15815_ (.A1(net3700),
    .A2(_06692_),
    .B1(net3704),
    .Y(_06693_));
 sky130_fd_sc_hd__nor2_4 _15816_ (.A(net3635),
    .B(net4033),
    .Y(_06694_));
 sky130_fd_sc_hd__nand2_1 _15817_ (.A(net4037),
    .B(net4035),
    .Y(_06695_));
 sky130_fd_sc_hd__nand2_4 _15818_ (.A(_06494_),
    .B(net4033),
    .Y(_06696_));
 sky130_fd_sc_hd__a21oi_1 _15819_ (.A1(_06695_),
    .A2(_06696_),
    .B1(net4016),
    .Y(_06697_));
 sky130_fd_sc_hd__a211oi_1 _15820_ (.A1(net4016),
    .A2(_06694_),
    .B1(_06697_),
    .C1(net4027),
    .Y(_06698_));
 sky130_fd_sc_hd__a311oi_1 _15821_ (.A1(net4026),
    .A2(_06691_),
    .A3(_06693_),
    .B1(_06698_),
    .C1(net4032),
    .Y(_06699_));
 sky130_fd_sc_hd__nand2_4 _15822_ (.A(_06629_),
    .B(_06611_),
    .Y(_06700_));
 sky130_fd_sc_hd__a211oi_1 _15823_ (.A1(net4032),
    .A2(_06688_),
    .B1(_06699_),
    .C1(_06700_),
    .Y(_06701_));
 sky130_fd_sc_hd__nor3_2 _15824_ (.A(_06613_),
    .B(_06674_),
    .C(_06701_),
    .Y(_00040_));
 sky130_fd_sc_hd__nor2_4 _15825_ (.A(_06603_),
    .B(_06630_),
    .Y(_06702_));
 sky130_fd_sc_hd__nor3_1 _15826_ (.A(net3701),
    .B(net3699),
    .C(_06666_),
    .Y(_06703_));
 sky130_fd_sc_hd__nor2_2 _15827_ (.A(net4037),
    .B(net4021),
    .Y(_06704_));
 sky130_fd_sc_hd__nor3_1 _15828_ (.A(net4033),
    .B(_06704_),
    .C(_06557_),
    .Y(_06705_));
 sky130_fd_sc_hd__o21ai_0 _15829_ (.A1(_12020_[0]),
    .A2(net4031),
    .B1(net4032),
    .Y(_06706_));
 sky130_fd_sc_hd__o311ai_0 _15830_ (.A1(net4032),
    .A2(_06703_),
    .A3(_06705_),
    .B1(_06706_),
    .C1(net4016),
    .Y(_06707_));
 sky130_fd_sc_hd__nand2_1 _15831_ (.A(net4033),
    .B(_06682_),
    .Y(_06708_));
 sky130_fd_sc_hd__a21oi_1 _15832_ (.A1(_12004_[0]),
    .A2(_06505_),
    .B1(net4025),
    .Y(_06709_));
 sky130_fd_sc_hd__nand2_1 _15833_ (.A(net4036),
    .B(net4033),
    .Y(_06710_));
 sky130_fd_sc_hd__nand2_1 _15834_ (.A(_11996_[0]),
    .B(net3702),
    .Y(_06711_));
 sky130_fd_sc_hd__a21oi_1 _15835_ (.A1(_06710_),
    .A2(_06711_),
    .B1(net4025),
    .Y(_06712_));
 sky130_fd_sc_hd__nand2_8 _15836_ (.A(net3704),
    .B(net4023),
    .Y(_06713_));
 sky130_fd_sc_hd__nor2_2 _15837_ (.A(_06494_),
    .B(_06505_),
    .Y(_06714_));
 sky130_fd_sc_hd__nor2_1 _15838_ (.A(net4035),
    .B(net4033),
    .Y(_06715_));
 sky130_fd_sc_hd__nor3_2 _15839_ (.A(_06713_),
    .B(_06714_),
    .C(_06715_),
    .Y(_06716_));
 sky130_fd_sc_hd__nor3_1 _15840_ (.A(_06626_),
    .B(_06712_),
    .C(_06716_),
    .Y(_06717_));
 sky130_fd_sc_hd__a31oi_2 _15841_ (.A1(net4032),
    .A2(_06708_),
    .A3(_06709_),
    .B1(_06717_),
    .Y(_06718_));
 sky130_fd_sc_hd__nor2_4 _15842_ (.A(_06494_),
    .B(net4021),
    .Y(_06719_));
 sky130_fd_sc_hd__nand2_4 _15843_ (.A(net3635),
    .B(net4023),
    .Y(_06720_));
 sky130_fd_sc_hd__nand2_8 _15844_ (.A(_11996_[0]),
    .B(net399),
    .Y(_06721_));
 sky130_fd_sc_hd__nand3_1 _15845_ (.A(net4033),
    .B(_06720_),
    .C(_06721_),
    .Y(_06722_));
 sky130_fd_sc_hd__o311ai_0 _15846_ (.A1(net4033),
    .A2(_06666_),
    .A3(_06719_),
    .B1(_06722_),
    .C1(net4017),
    .Y(_06723_));
 sky130_fd_sc_hd__nand2_1 _15847_ (.A(net4036),
    .B(_06540_),
    .Y(_06724_));
 sky130_fd_sc_hd__nor2_4 _15848_ (.A(_06505_),
    .B(net4021),
    .Y(_06725_));
 sky130_fd_sc_hd__nor2_1 _15849_ (.A(net4037),
    .B(_06537_),
    .Y(_06726_));
 sky130_fd_sc_hd__o21ai_0 _15850_ (.A1(_06725_),
    .A2(_06726_),
    .B1(_06494_),
    .Y(_06727_));
 sky130_fd_sc_hd__o2111ai_1 _15851_ (.A1(net3635),
    .A2(_06642_),
    .B1(_06724_),
    .C1(_06727_),
    .D1(net4032),
    .Y(_06728_));
 sky130_fd_sc_hd__a211oi_1 _15852_ (.A1(_06723_),
    .A2(_06728_),
    .B1(net4019),
    .C1(_06671_),
    .Y(_06729_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_916 ();
 sky130_fd_sc_hd__or3_4 _15854_ (.A(_11997_[0]),
    .B(_06534_),
    .C(_06536_),
    .X(_06731_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_915 ();
 sky130_fd_sc_hd__nor2_1 _15856_ (.A(net4033),
    .B(_06653_),
    .Y(_06733_));
 sky130_fd_sc_hd__a311oi_1 _15857_ (.A1(net4033),
    .A2(_06654_),
    .A3(_06731_),
    .B1(_06733_),
    .C1(net4017),
    .Y(_06734_));
 sky130_fd_sc_hd__nor2_1 _15858_ (.A(net3704),
    .B(_06553_),
    .Y(_06735_));
 sky130_fd_sc_hd__nand2_8 _15859_ (.A(_06494_),
    .B(net4029),
    .Y(_06736_));
 sky130_fd_sc_hd__nor2_4 _15860_ (.A(net4037),
    .B(_06736_),
    .Y(_06737_));
 sky130_fd_sc_hd__a2111oi_0 _15861_ (.A1(_06505_),
    .A2(_06587_),
    .B1(_06735_),
    .C1(_06737_),
    .D1(net4032),
    .Y(_06738_));
 sky130_fd_sc_hd__nor4_1 _15862_ (.A(net4016),
    .B(_06671_),
    .C(_06734_),
    .D(_06738_),
    .Y(_06739_));
 sky130_fd_sc_hd__a311o_1 _15863_ (.A1(_06702_),
    .A2(_06707_),
    .A3(_06718_),
    .B1(_06729_),
    .C1(_06739_),
    .X(_06740_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_912 ();
 sky130_fd_sc_hd__a21oi_1 _15867_ (.A1(_11996_[0]),
    .A2(net4021),
    .B1(_06665_),
    .Y(_06744_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_911 ();
 sky130_fd_sc_hd__o21ai_1 _15869_ (.A1(_06658_),
    .A2(_06719_),
    .B1(_06505_),
    .Y(_06746_));
 sky130_fd_sc_hd__o21ai_0 _15870_ (.A1(_06505_),
    .A2(_06744_),
    .B1(_06746_),
    .Y(_06747_));
 sky130_fd_sc_hd__o21ai_0 _15871_ (.A1(_11996_[0]),
    .A2(net4021),
    .B1(_06713_),
    .Y(_06748_));
 sky130_fd_sc_hd__or3_4 _15872_ (.A(_12001_[0]),
    .B(_06534_),
    .C(_06536_),
    .X(_06749_));
 sky130_fd_sc_hd__nand3_1 _15873_ (.A(net4033),
    .B(_06736_),
    .C(_06749_),
    .Y(_06750_));
 sky130_fd_sc_hd__a21boi_0 _15874_ (.A1(net3701),
    .A2(_06748_),
    .B1_N(_06750_),
    .Y(_06751_));
 sky130_fd_sc_hd__o22ai_1 _15875_ (.A1(_06626_),
    .A2(_06747_),
    .B1(_06751_),
    .B2(_06615_),
    .Y(_06752_));
 sky130_fd_sc_hd__o21ai_0 _15876_ (.A1(_06658_),
    .A2(_06737_),
    .B1(net4033),
    .Y(_06753_));
 sky130_fd_sc_hd__nand2_2 _15877_ (.A(net4036),
    .B(_06573_),
    .Y(_06754_));
 sky130_fd_sc_hd__nor3_4 _15878_ (.A(net4037),
    .B(net4035),
    .C(net4026),
    .Y(_06755_));
 sky130_fd_sc_hd__o21ai_0 _15879_ (.A1(_06665_),
    .A2(_06755_),
    .B1(net3701),
    .Y(_06756_));
 sky130_fd_sc_hd__nand2_4 _15880_ (.A(_12010_[0]),
    .B(net4031),
    .Y(_06757_));
 sky130_fd_sc_hd__nand2_4 _15881_ (.A(_06590_),
    .B(_06569_),
    .Y(_06758_));
 sky130_fd_sc_hd__a31oi_1 _15882_ (.A1(net4033),
    .A2(_06731_),
    .A3(_06757_),
    .B1(_06758_),
    .Y(_06759_));
 sky130_fd_sc_hd__a32o_1 _15883_ (.A1(_06656_),
    .A2(_06753_),
    .A3(_06754_),
    .B1(_06756_),
    .B2(_06759_),
    .X(_06760_));
 sky130_fd_sc_hd__nor3_1 _15884_ (.A(_06612_),
    .B(_06752_),
    .C(_06760_),
    .Y(_06761_));
 sky130_fd_sc_hd__nand2_8 _15885_ (.A(net4035),
    .B(net4024),
    .Y(_06762_));
 sky130_fd_sc_hd__a21oi_1 _15886_ (.A1(net3702),
    .A2(_06762_),
    .B1(net4037),
    .Y(_06763_));
 sky130_fd_sc_hd__a2111oi_0 _15887_ (.A1(net4037),
    .A2(_06719_),
    .B1(_06763_),
    .C1(net3622),
    .D1(_06615_),
    .Y(_06764_));
 sky130_fd_sc_hd__a21oi_1 _15888_ (.A1(_12010_[0]),
    .A2(net4033),
    .B1(_06635_),
    .Y(_06765_));
 sky130_fd_sc_hd__nor2_2 _15889_ (.A(_12001_[0]),
    .B(net4033),
    .Y(_06766_));
 sky130_fd_sc_hd__nor3_2 _15890_ (.A(net4037),
    .B(_06494_),
    .C(_06505_),
    .Y(_06767_));
 sky130_fd_sc_hd__o31ai_2 _15891_ (.A1(net4021),
    .A2(_06766_),
    .A3(net3621),
    .B1(net4032),
    .Y(_06768_));
 sky130_fd_sc_hd__o21bai_2 _15892_ (.A1(net4027),
    .A2(_06765_),
    .B1_N(_06768_),
    .Y(_06769_));
 sky130_fd_sc_hd__o22ai_1 _15893_ (.A1(_12001_[0]),
    .A2(_06642_),
    .B1(_06637_),
    .B2(net4038),
    .Y(_06770_));
 sky130_fd_sc_hd__a21oi_1 _15894_ (.A1(_06569_),
    .A2(_06770_),
    .B1(_06565_),
    .Y(_06771_));
 sky130_fd_sc_hd__a21oi_1 _15895_ (.A1(_06654_),
    .A2(_06720_),
    .B1(net3701),
    .Y(_06772_));
 sky130_fd_sc_hd__a31oi_1 _15896_ (.A1(net3701),
    .A2(_06736_),
    .A3(_06762_),
    .B1(_06772_),
    .Y(_06773_));
 sky130_fd_sc_hd__o2bb2ai_1 _15897_ (.A1_N(_06769_),
    .A2_N(_06771_),
    .B1(_06773_),
    .B2(_06626_),
    .Y(_06774_));
 sky130_fd_sc_hd__nor3_1 _15898_ (.A(_06631_),
    .B(_06764_),
    .C(_06774_),
    .Y(_06775_));
 sky130_fd_sc_hd__nor3_1 _15899_ (.A(_06740_),
    .B(_06761_),
    .C(_06775_),
    .Y(_00041_));
 sky130_fd_sc_hd__nor2_4 _15900_ (.A(_06494_),
    .B(net399),
    .Y(_06776_));
 sky130_fd_sc_hd__nand2_2 _15901_ (.A(net3704),
    .B(net3700),
    .Y(_06777_));
 sky130_fd_sc_hd__o32ai_1 _15902_ (.A1(net3699),
    .A2(_06776_),
    .A3(_06777_),
    .B1(_06553_),
    .B2(_12010_[0]),
    .Y(_06778_));
 sky130_fd_sc_hd__nand2_1 _15903_ (.A(_06639_),
    .B(_06620_),
    .Y(_06779_));
 sky130_fd_sc_hd__nor2_2 _15904_ (.A(net3635),
    .B(net4021),
    .Y(_06780_));
 sky130_fd_sc_hd__nor3_1 _15905_ (.A(_06505_),
    .B(_06776_),
    .C(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_910 ();
 sky130_fd_sc_hd__a211oi_2 _15907_ (.A1(_06505_),
    .A2(_06779_),
    .B1(_06781_),
    .C1(net4032),
    .Y(_06783_));
 sky130_fd_sc_hd__a21oi_1 _15908_ (.A1(net4032),
    .A2(_06778_),
    .B1(_06783_),
    .Y(_06784_));
 sky130_fd_sc_hd__nor2_4 _15909_ (.A(_12010_[0]),
    .B(net4023),
    .Y(_06785_));
 sky130_fd_sc_hd__nor2_1 _15910_ (.A(_06776_),
    .B(_06785_),
    .Y(_06786_));
 sky130_fd_sc_hd__a221oi_1 _15911_ (.A1(_12001_[0]),
    .A2(_06725_),
    .B1(_06786_),
    .B2(net3701),
    .C1(_06557_),
    .Y(_06787_));
 sky130_fd_sc_hd__nor2_2 _15912_ (.A(net4037),
    .B(_06505_),
    .Y(_06788_));
 sky130_fd_sc_hd__o21ai_2 _15913_ (.A1(_06766_),
    .A2(net3621),
    .B1(net4021),
    .Y(_06789_));
 sky130_fd_sc_hd__o311ai_0 _15914_ (.A1(net4021),
    .A2(_06635_),
    .A3(_06788_),
    .B1(_06789_),
    .C1(net4032),
    .Y(_06790_));
 sky130_fd_sc_hd__o211ai_1 _15915_ (.A1(net4032),
    .A2(_06787_),
    .B1(_06790_),
    .C1(net4016),
    .Y(_06791_));
 sky130_fd_sc_hd__o21ai_1 _15916_ (.A1(net4016),
    .A2(_06784_),
    .B1(_06791_),
    .Y(_06792_));
 sky130_fd_sc_hd__nand2_4 _15917_ (.A(_12006_[0]),
    .B(net4027),
    .Y(_06793_));
 sky130_fd_sc_hd__nand3_1 _15918_ (.A(net3701),
    .B(_06731_),
    .C(_06793_),
    .Y(_06794_));
 sky130_fd_sc_hd__o21ai_0 _15919_ (.A1(_06658_),
    .A2(_06719_),
    .B1(net4033),
    .Y(_06795_));
 sky130_fd_sc_hd__nand3_1 _15920_ (.A(net4032),
    .B(_06794_),
    .C(_06795_),
    .Y(_06796_));
 sky130_fd_sc_hd__nor2_1 _15921_ (.A(net4037),
    .B(net4033),
    .Y(_06797_));
 sky130_fd_sc_hd__nor2_2 _15922_ (.A(_12006_[0]),
    .B(net3701),
    .Y(_06798_));
 sky130_fd_sc_hd__o21ai_0 _15923_ (.A1(_06797_),
    .A2(_06798_),
    .B1(net4021),
    .Y(_06799_));
 sky130_fd_sc_hd__nand2_1 _15924_ (.A(_12010_[0]),
    .B(net3702),
    .Y(_06800_));
 sky130_fd_sc_hd__a21oi_2 _15925_ (.A1(_06494_),
    .A2(net4033),
    .B1(net4021),
    .Y(_06801_));
 sky130_fd_sc_hd__nand2_1 _15926_ (.A(_06800_),
    .B(_06801_),
    .Y(_06802_));
 sky130_fd_sc_hd__nand3_1 _15927_ (.A(net4017),
    .B(_06799_),
    .C(_06802_),
    .Y(_06803_));
 sky130_fd_sc_hd__nand3_2 _15928_ (.A(net4019),
    .B(_06796_),
    .C(_06803_),
    .Y(_06804_));
 sky130_fd_sc_hd__nand2b_1 _15929_ (.A_N(_12010_[0]),
    .B(net399),
    .Y(_06805_));
 sky130_fd_sc_hd__nor3_1 _15930_ (.A(net3700),
    .B(_06776_),
    .C(_06659_),
    .Y(_06806_));
 sky130_fd_sc_hd__a31oi_1 _15931_ (.A1(net3700),
    .A2(_06749_),
    .A3(_06805_),
    .B1(_06806_),
    .Y(_06807_));
 sky130_fd_sc_hd__a311o_1 _15932_ (.A1(net4033),
    .A2(_06793_),
    .A3(_06713_),
    .B1(net4017),
    .C1(_06766_),
    .X(_06808_));
 sky130_fd_sc_hd__o211ai_1 _15933_ (.A1(net4032),
    .A2(_06807_),
    .B1(_06808_),
    .C1(net4016),
    .Y(_06809_));
 sky130_fd_sc_hd__a21oi_2 _15934_ (.A1(_06804_),
    .A2(_06809_),
    .B1(_06612_),
    .Y(_06810_));
 sky130_fd_sc_hd__o21ai_0 _15935_ (.A1(_06590_),
    .A2(_06575_),
    .B1(_06677_),
    .Y(_06811_));
 sky130_fd_sc_hd__a2111oi_0 _15936_ (.A1(_06541_),
    .A2(_06643_),
    .B1(_06542_),
    .C1(_06505_),
    .D1(_06590_),
    .Y(_06812_));
 sky130_fd_sc_hd__nand3_4 _15937_ (.A(_06494_),
    .B(_06505_),
    .C(_06541_),
    .Y(_06813_));
 sky130_fd_sc_hd__nand2_1 _15938_ (.A(_12024_[0]),
    .B(net4028),
    .Y(_06814_));
 sky130_fd_sc_hd__a21oi_1 _15939_ (.A1(_06813_),
    .A2(_06814_),
    .B1(_06565_),
    .Y(_06815_));
 sky130_fd_sc_hd__nand2_1 _15940_ (.A(_12004_[0]),
    .B(_06537_),
    .Y(_06816_));
 sky130_fd_sc_hd__nor3b_1 _15941_ (.A(_06689_),
    .B(_06755_),
    .C_N(_06816_),
    .Y(_06817_));
 sky130_fd_sc_hd__a2111oi_0 _15942_ (.A1(net4037),
    .A2(_06811_),
    .B1(_06812_),
    .C1(_06815_),
    .D1(_06817_),
    .Y(_06818_));
 sky130_fd_sc_hd__nor3_1 _15943_ (.A(_06603_),
    .B(net4032),
    .C(_06818_),
    .Y(_06819_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_909 ();
 sky130_fd_sc_hd__nor3_1 _15945_ (.A(net4027),
    .B(_06694_),
    .C(_06767_),
    .Y(_06821_));
 sky130_fd_sc_hd__a211oi_1 _15946_ (.A1(_12017_[0]),
    .A2(net4027),
    .B1(_06821_),
    .C1(net4016),
    .Y(_06822_));
 sky130_fd_sc_hd__nand2_1 _15947_ (.A(net3704),
    .B(net4033),
    .Y(_06823_));
 sky130_fd_sc_hd__nor2_1 _15948_ (.A(_12020_[0]),
    .B(net4021),
    .Y(_06824_));
 sky130_fd_sc_hd__a311oi_1 _15949_ (.A1(net4021),
    .A2(_06823_),
    .A3(_06695_),
    .B1(_06824_),
    .C1(net4020),
    .Y(_06825_));
 sky130_fd_sc_hd__nor4_1 _15950_ (.A(_06629_),
    .B(net4017),
    .C(_06822_),
    .D(_06825_),
    .Y(_06826_));
 sky130_fd_sc_hd__o32ai_1 _15951_ (.A1(net3704),
    .A2(net3700),
    .A3(_06776_),
    .B1(_06713_),
    .B2(_06714_),
    .Y(_06827_));
 sky130_fd_sc_hd__a21oi_1 _15952_ (.A1(_06639_),
    .A2(_06777_),
    .B1(net3635),
    .Y(_06828_));
 sky130_fd_sc_hd__nor2_1 _15953_ (.A(_06629_),
    .B(net4032),
    .Y(_06829_));
 sky130_fd_sc_hd__nand3_1 _15954_ (.A(net4033),
    .B(_06639_),
    .C(_06648_),
    .Y(_06830_));
 sky130_fd_sc_hd__nand3_1 _15955_ (.A(net3700),
    .B(_06731_),
    .C(_06721_),
    .Y(_06831_));
 sky130_fd_sc_hd__nand3_1 _15956_ (.A(_06590_),
    .B(_06830_),
    .C(_06831_),
    .Y(_06832_));
 sky130_fd_sc_hd__o311a_1 _15957_ (.A1(_06590_),
    .A2(_06827_),
    .A3(_06828_),
    .B1(_06829_),
    .C1(_06832_),
    .X(_06833_));
 sky130_fd_sc_hd__a32oi_1 _15958_ (.A1(net4033),
    .A2(_06731_),
    .A3(_06721_),
    .B1(_06579_),
    .B2(_12001_[0]),
    .Y(_06834_));
 sky130_fd_sc_hd__nand2_2 _15959_ (.A(net3703),
    .B(net4036),
    .Y(_06835_));
 sky130_fd_sc_hd__nand2_1 _15960_ (.A(_12015_[0]),
    .B(net4021),
    .Y(_06836_));
 sky130_fd_sc_hd__o311ai_0 _15961_ (.A1(net4033),
    .A2(net4021),
    .A3(_06835_),
    .B1(_06836_),
    .C1(net4016),
    .Y(_06837_));
 sky130_fd_sc_hd__o21ai_0 _15962_ (.A1(net4016),
    .A2(_06834_),
    .B1(_06837_),
    .Y(_06838_));
 sky130_fd_sc_hd__a31oi_1 _15963_ (.A1(_06629_),
    .A2(net4032),
    .A3(_06838_),
    .B1(_06611_),
    .Y(_06839_));
 sky130_fd_sc_hd__nor4b_1 _15964_ (.A(_06819_),
    .B(_06826_),
    .C(_06833_),
    .D_N(_06839_),
    .Y(_06840_));
 sky130_fd_sc_hd__a211oi_1 _15965_ (.A1(_06702_),
    .A2(_06792_),
    .B1(_06810_),
    .C1(_06840_),
    .Y(_00042_));
 sky130_fd_sc_hd__nand2_1 _15966_ (.A(net4036),
    .B(_06537_),
    .Y(_06841_));
 sky130_fd_sc_hd__a222oi_1 _15967_ (.A1(net3635),
    .A2(_06540_),
    .B1(_06841_),
    .B2(_06797_),
    .C1(_06801_),
    .C2(net4037),
    .Y(_06842_));
 sky130_fd_sc_hd__nand2_1 _15968_ (.A(net4036),
    .B(_06725_),
    .Y(_06843_));
 sky130_fd_sc_hd__o21ai_0 _15969_ (.A1(_06583_),
    .A2(_06658_),
    .B1(_06505_),
    .Y(_06844_));
 sky130_fd_sc_hd__a21oi_1 _15970_ (.A1(_06843_),
    .A2(_06844_),
    .B1(net4032),
    .Y(_06845_));
 sky130_fd_sc_hd__a21oi_1 _15971_ (.A1(net4032),
    .A2(_06842_),
    .B1(_06845_),
    .Y(_06846_));
 sky130_fd_sc_hd__nor2_2 _15972_ (.A(_12004_[0]),
    .B(net4025),
    .Y(_06847_));
 sky130_fd_sc_hd__nor3b_1 _15973_ (.A(_06847_),
    .B(net3702),
    .C_N(_06640_),
    .Y(_06848_));
 sky130_fd_sc_hd__a311oi_1 _15974_ (.A1(net3702),
    .A2(_06736_),
    .A3(_06731_),
    .B1(_06848_),
    .C1(_06626_),
    .Y(_06849_));
 sky130_fd_sc_hd__nand2b_4 _15975_ (.A_N(net3635),
    .B(net4030),
    .Y(_06850_));
 sky130_fd_sc_hd__a21oi_1 _15976_ (.A1(_06639_),
    .A2(_06749_),
    .B1(net4034),
    .Y(_06851_));
 sky130_fd_sc_hd__a311oi_1 _15977_ (.A1(net4034),
    .A2(_06587_),
    .A3(_06850_),
    .B1(_06851_),
    .C1(_06615_),
    .Y(_06852_));
 sky130_fd_sc_hd__a2111oi_0 _15978_ (.A1(net4016),
    .A2(_06846_),
    .B1(_06849_),
    .C1(_06852_),
    .D1(_06631_),
    .Y(_06853_));
 sky130_fd_sc_hd__nand3_1 _15979_ (.A(_06505_),
    .B(_06617_),
    .C(_06850_),
    .Y(_06854_));
 sky130_fd_sc_hd__nand2_2 _15980_ (.A(net4032),
    .B(net4025),
    .Y(_06855_));
 sky130_fd_sc_hd__a21oi_1 _15981_ (.A1(_06682_),
    .A2(_06855_),
    .B1(_12004_[0]),
    .Y(_06856_));
 sky130_fd_sc_hd__nand2_1 _15982_ (.A(net4032),
    .B(net4028),
    .Y(_06857_));
 sky130_fd_sc_hd__nor2_1 _15983_ (.A(_06682_),
    .B(_06857_),
    .Y(_06858_));
 sky130_fd_sc_hd__o21ai_0 _15984_ (.A1(_06856_),
    .A2(_06858_),
    .B1(net4033),
    .Y(_06859_));
 sky130_fd_sc_hd__a21oi_1 _15985_ (.A1(_06854_),
    .A2(_06859_),
    .B1(_06615_),
    .Y(_06860_));
 sky130_fd_sc_hd__nor3_2 _15986_ (.A(_06505_),
    .B(_06780_),
    .C(_06726_),
    .Y(_06861_));
 sky130_fd_sc_hd__a311oi_1 _15987_ (.A1(_06505_),
    .A2(_06587_),
    .A3(_06793_),
    .B1(_06758_),
    .C1(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__nor2_1 _15988_ (.A(net4036),
    .B(net4027),
    .Y(_06863_));
 sky130_fd_sc_hd__o21ai_0 _15989_ (.A1(_06863_),
    .A2(_06847_),
    .B1(_06505_),
    .Y(_06864_));
 sky130_fd_sc_hd__o211a_1 _15990_ (.A1(net3635),
    .A2(_06575_),
    .B1(_06617_),
    .C1(_06864_),
    .X(_06865_));
 sky130_fd_sc_hd__a21o_1 _15991_ (.A1(_06835_),
    .A2(_06696_),
    .B1(net3622),
    .X(_06866_));
 sky130_fd_sc_hd__a21oi_1 _15992_ (.A1(_06656_),
    .A2(_06866_),
    .B1(_06671_),
    .Y(_06867_));
 sky130_fd_sc_hd__o21ai_0 _15993_ (.A1(_06626_),
    .A2(_06865_),
    .B1(_06867_),
    .Y(_06868_));
 sky130_fd_sc_hd__nand2_4 _15994_ (.A(_12006_[0]),
    .B(net4021),
    .Y(_06869_));
 sky130_fd_sc_hd__a21oi_2 _15995_ (.A1(_06649_),
    .A2(_06869_),
    .B1(net3701),
    .Y(_06870_));
 sky130_fd_sc_hd__a21oi_1 _15996_ (.A1(_06762_),
    .A2(_06757_),
    .B1(net4033),
    .Y(_06871_));
 sky130_fd_sc_hd__o32ai_2 _15997_ (.A1(_06626_),
    .A2(_06870_),
    .A3(_06871_),
    .B1(_06758_),
    .B2(_06802_),
    .Y(_06872_));
 sky130_fd_sc_hd__a21oi_1 _15998_ (.A1(net4034),
    .A2(_06639_),
    .B1(net4036),
    .Y(_06873_));
 sky130_fd_sc_hd__o22ai_1 _15999_ (.A1(_11996_[0]),
    .A2(_06553_),
    .B1(_06642_),
    .B2(net4038),
    .Y(_06874_));
 sky130_fd_sc_hd__nor3_1 _16000_ (.A(_06615_),
    .B(_06873_),
    .C(_06874_),
    .Y(_06875_));
 sky130_fd_sc_hd__nor2_1 _16001_ (.A(_12006_[0]),
    .B(net4034),
    .Y(_06876_));
 sky130_fd_sc_hd__a211oi_1 _16002_ (.A1(net4034),
    .A2(net3589),
    .B1(_06876_),
    .C1(net4030),
    .Y(_06877_));
 sky130_fd_sc_hd__a2111oi_0 _16003_ (.A1(_06708_),
    .A2(_06709_),
    .B1(_06877_),
    .C1(_06569_),
    .D1(_06565_),
    .Y(_06878_));
 sky130_fd_sc_hd__nor3_1 _16004_ (.A(_06872_),
    .B(_06875_),
    .C(_06878_),
    .Y(_06879_));
 sky130_fd_sc_hd__o32ai_1 _16005_ (.A1(_06860_),
    .A2(_06862_),
    .A3(_06868_),
    .B1(_06879_),
    .B2(_06612_),
    .Y(_06880_));
 sky130_fd_sc_hd__a22oi_1 _16006_ (.A1(_06494_),
    .A2(_06725_),
    .B1(_06637_),
    .B2(_12006_[0]),
    .Y(_06881_));
 sky130_fd_sc_hd__nor2_1 _16007_ (.A(_06505_),
    .B(net4032),
    .Y(_06882_));
 sky130_fd_sc_hd__nand2_1 _16008_ (.A(_06620_),
    .B(_06850_),
    .Y(_06883_));
 sky130_fd_sc_hd__a21oi_1 _16009_ (.A1(_06882_),
    .A2(_06883_),
    .B1(net4016),
    .Y(_06884_));
 sky130_fd_sc_hd__o21ai_0 _16010_ (.A1(net4018),
    .A2(_06881_),
    .B1(_06884_),
    .Y(_06885_));
 sky130_fd_sc_hd__or3_1 _16011_ (.A(net4034),
    .B(_06658_),
    .C(_06847_),
    .X(_06886_));
 sky130_fd_sc_hd__o21ai_0 _16012_ (.A1(_06505_),
    .A2(_06779_),
    .B1(_06886_),
    .Y(_06887_));
 sky130_fd_sc_hd__a21oi_1 _16013_ (.A1(net4021),
    .A2(net3589),
    .B1(_06780_),
    .Y(_06888_));
 sky130_fd_sc_hd__a21oi_1 _16014_ (.A1(_06736_),
    .A2(_06587_),
    .B1(net4034),
    .Y(_06889_));
 sky130_fd_sc_hd__a21oi_1 _16015_ (.A1(net4034),
    .A2(_06888_),
    .B1(_06889_),
    .Y(_06890_));
 sky130_fd_sc_hd__a22oi_1 _16016_ (.A1(_06663_),
    .A2(_06887_),
    .B1(_06890_),
    .B2(_06656_),
    .Y(_06891_));
 sky130_fd_sc_hd__a21oi_2 _16017_ (.A1(_06885_),
    .A2(_06891_),
    .B1(_06700_),
    .Y(_06892_));
 sky130_fd_sc_hd__nor3_1 _16018_ (.A(_06853_),
    .B(_06880_),
    .C(_06892_),
    .Y(_00043_));
 sky130_fd_sc_hd__a31oi_1 _16019_ (.A1(net3701),
    .A2(_06654_),
    .A3(_06720_),
    .B1(_06798_),
    .Y(_06893_));
 sky130_fd_sc_hd__nor2_1 _16020_ (.A(net4032),
    .B(_06893_),
    .Y(_06894_));
 sky130_fd_sc_hd__nand2_1 _16021_ (.A(_06649_),
    .B(_06869_),
    .Y(_06895_));
 sky130_fd_sc_hd__nor3_2 _16022_ (.A(net4037),
    .B(_06494_),
    .C(net399),
    .Y(_06896_));
 sky130_fd_sc_hd__nor3_1 _16023_ (.A(net3700),
    .B(_06896_),
    .C(_06785_),
    .Y(_06897_));
 sky130_fd_sc_hd__a211oi_1 _16024_ (.A1(net3700),
    .A2(_06895_),
    .B1(_06897_),
    .C1(net4017),
    .Y(_06898_));
 sky130_fd_sc_hd__o21ai_0 _16025_ (.A1(_11996_[0]),
    .A2(net3700),
    .B1(_06777_),
    .Y(_06899_));
 sky130_fd_sc_hd__a21oi_1 _16026_ (.A1(net4024),
    .A2(_06899_),
    .B1(_06768_),
    .Y(_06900_));
 sky130_fd_sc_hd__nor2_4 _16027_ (.A(_12001_[0]),
    .B(net4023),
    .Y(_06901_));
 sky130_fd_sc_hd__nor3_1 _16028_ (.A(net3700),
    .B(_06896_),
    .C(_06901_),
    .Y(_06902_));
 sky130_fd_sc_hd__o31ai_1 _16029_ (.A1(net4033),
    .A2(_06557_),
    .A3(_06785_),
    .B1(net4017),
    .Y(_06903_));
 sky130_fd_sc_hd__o21ai_0 _16030_ (.A1(_06902_),
    .A2(_06903_),
    .B1(_06590_),
    .Y(_06904_));
 sky130_fd_sc_hd__o32ai_1 _16031_ (.A1(_06590_),
    .A2(_06894_),
    .A3(_06898_),
    .B1(_06900_),
    .B2(_06904_),
    .Y(_06905_));
 sky130_fd_sc_hd__o21ai_2 _16032_ (.A1(_11998_[0]),
    .A2(_06575_),
    .B1(_06617_),
    .Y(_06906_));
 sky130_fd_sc_hd__a21oi_1 _16033_ (.A1(_06647_),
    .A2(_06721_),
    .B1(net4033),
    .Y(_06907_));
 sky130_fd_sc_hd__o21a_1 _16034_ (.A1(_06906_),
    .A2(_06907_),
    .B1(net4032),
    .X(_06908_));
 sky130_fd_sc_hd__a21oi_1 _16035_ (.A1(_06639_),
    .A2(_06762_),
    .B1(net3700),
    .Y(_06909_));
 sky130_fd_sc_hd__a2111oi_0 _16036_ (.A1(_12006_[0]),
    .A2(_06579_),
    .B1(_06737_),
    .C1(_06909_),
    .D1(net4032),
    .Y(_06910_));
 sky130_fd_sc_hd__nand2_2 _16037_ (.A(net3703),
    .B(_06719_),
    .Y(_06911_));
 sky130_fd_sc_hd__a221oi_1 _16038_ (.A1(net4037),
    .A2(_06540_),
    .B1(_06869_),
    .B2(_06505_),
    .C1(_06626_),
    .Y(_06912_));
 sky130_fd_sc_hd__mux2i_1 _16039_ (.A0(_12008_[0]),
    .A1(_06635_),
    .S(net4021),
    .Y(_06913_));
 sky130_fd_sc_hd__nor2_2 _16040_ (.A(net4016),
    .B(net4018),
    .Y(_06914_));
 sky130_fd_sc_hd__a22oi_2 _16041_ (.A1(_06911_),
    .A2(_06912_),
    .B1(_06913_),
    .B2(_06914_),
    .Y(_06915_));
 sky130_fd_sc_hd__o311ai_0 _16042_ (.A1(net4020),
    .A2(_06908_),
    .A3(_06910_),
    .B1(_06915_),
    .C1(_06611_),
    .Y(_06916_));
 sky130_fd_sc_hd__o21ai_0 _16043_ (.A1(_06611_),
    .A2(_06905_),
    .B1(_06916_),
    .Y(_06917_));
 sky130_fd_sc_hd__a311oi_1 _16044_ (.A1(net4033),
    .A2(_06749_),
    .A3(_06721_),
    .B1(_06705_),
    .C1(net4020),
    .Y(_06918_));
 sky130_fd_sc_hd__nor2_1 _16045_ (.A(_06665_),
    .B(_06755_),
    .Y(_06919_));
 sky130_fd_sc_hd__o21ai_0 _16046_ (.A1(_06689_),
    .A2(_06919_),
    .B1(net4017),
    .Y(_06920_));
 sky130_fd_sc_hd__nor2_1 _16047_ (.A(_06918_),
    .B(_06920_),
    .Y(_06921_));
 sky130_fd_sc_hd__nor3_1 _16048_ (.A(net3701),
    .B(_06901_),
    .C(_06755_),
    .Y(_06922_));
 sky130_fd_sc_hd__a31oi_1 _16049_ (.A1(net3701),
    .A2(_06762_),
    .A3(_06649_),
    .B1(_06922_),
    .Y(_06923_));
 sky130_fd_sc_hd__o22ai_1 _16050_ (.A1(_06494_),
    .A2(_06575_),
    .B1(_06785_),
    .B2(net4033),
    .Y(_06924_));
 sky130_fd_sc_hd__a21oi_1 _16051_ (.A1(_06656_),
    .A2(_06924_),
    .B1(_06612_),
    .Y(_06925_));
 sky130_fd_sc_hd__o21ai_1 _16052_ (.A1(_06615_),
    .A2(_06923_),
    .B1(_06925_),
    .Y(_06926_));
 sky130_fd_sc_hd__a21oi_1 _16053_ (.A1(_06505_),
    .A2(_06869_),
    .B1(_06665_),
    .Y(_06927_));
 sky130_fd_sc_hd__nor2_1 _16054_ (.A(net4032),
    .B(_06927_),
    .Y(_06928_));
 sky130_fd_sc_hd__nand2_1 _16055_ (.A(net4032),
    .B(_06696_),
    .Y(_06929_));
 sky130_fd_sc_hd__a31oi_1 _16056_ (.A1(_06505_),
    .A2(_06721_),
    .A3(_06713_),
    .B1(_06929_),
    .Y(_06930_));
 sky130_fd_sc_hd__a21oi_1 _16057_ (.A1(net4032),
    .A2(_06776_),
    .B1(_06882_),
    .Y(_06931_));
 sky130_fd_sc_hd__o21ai_0 _16058_ (.A1(net3703),
    .A2(_06931_),
    .B1(net4016),
    .Y(_06932_));
 sky130_fd_sc_hd__nand2_1 _16059_ (.A(net4032),
    .B(_06788_),
    .Y(_06933_));
 sky130_fd_sc_hd__nand3_1 _16060_ (.A(_11996_[0]),
    .B(_06505_),
    .C(net4017),
    .Y(_06934_));
 sky130_fd_sc_hd__nor2_1 _16061_ (.A(net4033),
    .B(net4017),
    .Y(_06935_));
 sky130_fd_sc_hd__o21ai_0 _16062_ (.A1(_06494_),
    .A2(_06935_),
    .B1(net3703),
    .Y(_06936_));
 sky130_fd_sc_hd__a32oi_1 _16063_ (.A1(net4021),
    .A2(_06933_),
    .A3(_06934_),
    .B1(_06801_),
    .B2(_06936_),
    .Y(_06937_));
 sky130_fd_sc_hd__o32ai_2 _16064_ (.A1(net4016),
    .A2(_06928_),
    .A3(_06930_),
    .B1(_06932_),
    .B2(_06937_),
    .Y(_06938_));
 sky130_fd_sc_hd__o22ai_2 _16065_ (.A1(_06921_),
    .A2(_06926_),
    .B1(_06938_),
    .B2(_06671_),
    .Y(_06939_));
 sky130_fd_sc_hd__a21oi_1 _16066_ (.A1(_06629_),
    .A2(_06917_),
    .B1(_06939_),
    .Y(_00044_));
 sky130_fd_sc_hd__nor2_4 _16067_ (.A(_06629_),
    .B(_06630_),
    .Y(_06940_));
 sky130_fd_sc_hd__nand3_1 _16068_ (.A(net4033),
    .B(_06639_),
    .C(_06731_),
    .Y(_06941_));
 sky130_fd_sc_hd__o311ai_0 _16069_ (.A1(net4033),
    .A2(_06896_),
    .A3(_06659_),
    .B1(_06941_),
    .C1(net4020),
    .Y(_06942_));
 sky130_fd_sc_hd__nand3_1 _16070_ (.A(net3700),
    .B(_06648_),
    .C(_06805_),
    .Y(_06943_));
 sky130_fd_sc_hd__o311ai_0 _16071_ (.A1(net3700),
    .A2(net4024),
    .A3(_06682_),
    .B1(_06943_),
    .C1(_06590_),
    .Y(_06944_));
 sky130_fd_sc_hd__nand3_1 _16072_ (.A(net4017),
    .B(_06942_),
    .C(_06944_),
    .Y(_06945_));
 sky130_fd_sc_hd__a21oi_1 _16073_ (.A1(_06590_),
    .A2(_06901_),
    .B1(_06776_),
    .Y(_06946_));
 sky130_fd_sc_hd__o21ai_0 _16074_ (.A1(net4020),
    .A2(_06713_),
    .B1(_06676_),
    .Y(_06947_));
 sky130_fd_sc_hd__o21ai_0 _16075_ (.A1(net4020),
    .A2(net4024),
    .B1(net4035),
    .Y(_06948_));
 sky130_fd_sc_hd__o211ai_1 _16076_ (.A1(net4035),
    .A2(_06947_),
    .B1(_06948_),
    .C1(net4033),
    .Y(_06949_));
 sky130_fd_sc_hd__a21oi_1 _16077_ (.A1(_06586_),
    .A2(_06692_),
    .B1(net4017),
    .Y(_06950_));
 sky130_fd_sc_hd__o211ai_1 _16078_ (.A1(net4033),
    .A2(_06946_),
    .B1(_06949_),
    .C1(_06950_),
    .Y(_06951_));
 sky130_fd_sc_hd__nand3_1 _16079_ (.A(_06940_),
    .B(_06945_),
    .C(_06951_),
    .Y(_06952_));
 sky130_fd_sc_hd__a221o_1 _16080_ (.A1(_12001_[0]),
    .A2(net4023),
    .B1(_06573_),
    .B2(_12006_[0]),
    .C1(net4016),
    .X(_06953_));
 sky130_fd_sc_hd__a21oi_1 _16081_ (.A1(net4033),
    .A2(_06654_),
    .B1(_06896_),
    .Y(_06954_));
 sky130_fd_sc_hd__o22ai_1 _16082_ (.A1(_06622_),
    .A2(_06953_),
    .B1(_06954_),
    .B2(net4020),
    .Y(_06955_));
 sky130_fd_sc_hd__o211ai_1 _16083_ (.A1(net3701),
    .A2(_06895_),
    .B1(_06813_),
    .C1(_06656_),
    .Y(_06956_));
 sky130_fd_sc_hd__nand2_1 _16084_ (.A(net3702),
    .B(_06548_),
    .Y(_06957_));
 sky130_fd_sc_hd__nand3_1 _16085_ (.A(_06914_),
    .B(_06668_),
    .C(_06957_),
    .Y(_06958_));
 sky130_fd_sc_hd__o211a_1 _16086_ (.A1(net4032),
    .A2(_06955_),
    .B1(_06956_),
    .C1(_06958_),
    .X(_06959_));
 sky130_fd_sc_hd__a21oi_1 _16087_ (.A1(_06640_),
    .A2(_06757_),
    .B1(net4033),
    .Y(_06960_));
 sky130_fd_sc_hd__o21ai_0 _16088_ (.A1(net3635),
    .A2(_06553_),
    .B1(net4032),
    .Y(_06961_));
 sky130_fd_sc_hd__a21boi_0 _16089_ (.A1(_11998_[0]),
    .A2(net4028),
    .B1_N(_06720_),
    .Y(_06962_));
 sky130_fd_sc_hd__o221ai_1 _16090_ (.A1(net3703),
    .A2(_06575_),
    .B1(_06962_),
    .B2(net4033),
    .C1(_06569_),
    .Y(_06963_));
 sky130_fd_sc_hd__o2111ai_2 _16091_ (.A1(_06960_),
    .A2(_06961_),
    .B1(_06963_),
    .C1(net4016),
    .D1(_06629_),
    .Y(_06964_));
 sky130_fd_sc_hd__o21ai_0 _16092_ (.A1(net4032),
    .A2(_06553_),
    .B1(_06857_),
    .Y(_06965_));
 sky130_fd_sc_hd__a22oi_1 _16093_ (.A1(_06569_),
    .A2(_06583_),
    .B1(_06965_),
    .B2(net3703),
    .Y(_06966_));
 sky130_fd_sc_hd__a22oi_1 _16094_ (.A1(_12004_[0]),
    .A2(_06579_),
    .B1(_06725_),
    .B2(net4036),
    .Y(_06967_));
 sky130_fd_sc_hd__nand2_1 _16095_ (.A(_06569_),
    .B(net4021),
    .Y(_06968_));
 sky130_fd_sc_hd__a311oi_1 _16096_ (.A1(net4038),
    .A2(_06642_),
    .A3(_06968_),
    .B1(_06603_),
    .C1(net4016),
    .Y(_06969_));
 sky130_fd_sc_hd__o221ai_2 _16097_ (.A1(net4036),
    .A2(_06966_),
    .B1(_06967_),
    .B2(net4032),
    .C1(_06969_),
    .Y(_06970_));
 sky130_fd_sc_hd__o2111ai_1 _16098_ (.A1(_06629_),
    .A2(_06959_),
    .B1(_06964_),
    .C1(_06970_),
    .D1(_06630_),
    .Y(_06971_));
 sky130_fd_sc_hd__nand2_1 _16099_ (.A(_06725_),
    .B(_06682_),
    .Y(_06972_));
 sky130_fd_sc_hd__a31oi_1 _16100_ (.A1(_06648_),
    .A2(_06656_),
    .A3(_06972_),
    .B1(_06700_),
    .Y(_06973_));
 sky130_fd_sc_hd__a21oi_1 _16101_ (.A1(net3623),
    .A2(net3589),
    .B1(_06615_),
    .Y(_06974_));
 sky130_fd_sc_hd__o31ai_1 _16102_ (.A1(_06586_),
    .A2(_06714_),
    .A3(_06715_),
    .B1(_06974_),
    .Y(_06975_));
 sky130_fd_sc_hd__nand3_1 _16103_ (.A(net4033),
    .B(_06649_),
    .C(_06731_),
    .Y(_06976_));
 sky130_fd_sc_hd__nand3_1 _16104_ (.A(_06590_),
    .B(_06943_),
    .C(_06976_),
    .Y(_06977_));
 sky130_fd_sc_hd__nand2_1 _16105_ (.A(_12001_[0]),
    .B(_06573_),
    .Y(_06978_));
 sky130_fd_sc_hd__o21ai_0 _16106_ (.A1(_12010_[0]),
    .A2(net4033),
    .B1(net4024),
    .Y(_06979_));
 sky130_fd_sc_hd__a31oi_1 _16107_ (.A1(net4020),
    .A2(_06978_),
    .A3(_06979_),
    .B1(net4032),
    .Y(_06980_));
 sky130_fd_sc_hd__nand2_1 _16108_ (.A(_06977_),
    .B(_06980_),
    .Y(_06981_));
 sky130_fd_sc_hd__nand3_1 _16109_ (.A(_06973_),
    .B(_06975_),
    .C(_06981_),
    .Y(_06982_));
 sky130_fd_sc_hd__and3_1 _16110_ (.A(_06952_),
    .B(_06971_),
    .C(_06982_),
    .X(_00045_));
 sky130_fd_sc_hd__o21ai_0 _16111_ (.A1(_12006_[0]),
    .A2(net4026),
    .B1(_06816_),
    .Y(_06983_));
 sky130_fd_sc_hd__a211oi_1 _16112_ (.A1(net3700),
    .A2(_06983_),
    .B1(_06735_),
    .C1(net4032),
    .Y(_06984_));
 sky130_fd_sc_hd__a21oi_1 _16113_ (.A1(net4032),
    .A2(_06789_),
    .B1(_06984_),
    .Y(_06985_));
 sky130_fd_sc_hd__a211oi_1 _16114_ (.A1(_12006_[0]),
    .A2(_06505_),
    .B1(net4021),
    .C1(_06788_),
    .Y(_06986_));
 sky130_fd_sc_hd__a21oi_1 _16115_ (.A1(_12014_[0]),
    .A2(net4021),
    .B1(_06986_),
    .Y(_06987_));
 sky130_fd_sc_hd__o21ai_0 _16116_ (.A1(net3635),
    .A2(_06553_),
    .B1(net4018),
    .Y(_06988_));
 sky130_fd_sc_hd__o221ai_1 _16117_ (.A1(net4018),
    .A2(_06987_),
    .B1(_06988_),
    .B2(_06889_),
    .C1(net4019),
    .Y(_06989_));
 sky130_fd_sc_hd__o21ai_0 _16118_ (.A1(net4019),
    .A2(_06985_),
    .B1(_06989_),
    .Y(_06990_));
 sky130_fd_sc_hd__nand2_1 _16119_ (.A(net4032),
    .B(_06580_),
    .Y(_06991_));
 sky130_fd_sc_hd__nand2_1 _16120_ (.A(net4037),
    .B(net3701),
    .Y(_06992_));
 sky130_fd_sc_hd__nand3_1 _16121_ (.A(_06553_),
    .B(_06736_),
    .C(_06992_),
    .Y(_06993_));
 sky130_fd_sc_hd__o22ai_1 _16122_ (.A1(_06870_),
    .A2(_06991_),
    .B1(_06993_),
    .B2(net4032),
    .Y(_06994_));
 sky130_fd_sc_hd__a21oi_1 _16123_ (.A1(_06616_),
    .A2(_06617_),
    .B1(net4033),
    .Y(_06995_));
 sky130_fd_sc_hd__nor3_1 _16124_ (.A(net4017),
    .B(_06861_),
    .C(_06995_),
    .Y(_06996_));
 sky130_fd_sc_hd__o211ai_1 _16125_ (.A1(net3635),
    .A2(net3702),
    .B1(_06569_),
    .C1(net4028),
    .Y(_06997_));
 sky130_fd_sc_hd__nor2_1 _16126_ (.A(net4033),
    .B(_06835_),
    .Y(_06998_));
 sky130_fd_sc_hd__o221ai_1 _16127_ (.A1(_12015_[0]),
    .A2(_06968_),
    .B1(_06997_),
    .B2(_06998_),
    .C1(_06565_),
    .Y(_06999_));
 sky130_fd_sc_hd__nand2_1 _16128_ (.A(net4030),
    .B(net3589),
    .Y(_07000_));
 sky130_fd_sc_hd__nand3_1 _16129_ (.A(net4033),
    .B(_06617_),
    .C(_07000_),
    .Y(_07001_));
 sky130_fd_sc_hd__o21ai_0 _16130_ (.A1(_06776_),
    .A2(_06780_),
    .B1(_06505_),
    .Y(_07002_));
 sky130_fd_sc_hd__o21ai_0 _16131_ (.A1(net4036),
    .A2(net3702),
    .B1(net3703),
    .Y(_07003_));
 sky130_fd_sc_hd__a211oi_1 _16132_ (.A1(net4021),
    .A2(_07003_),
    .B1(_06758_),
    .C1(_06625_),
    .Y(_07004_));
 sky130_fd_sc_hd__a311oi_1 _16133_ (.A1(_06656_),
    .A2(_07001_),
    .A3(_07002_),
    .B1(_07004_),
    .C1(_06631_),
    .Y(_07005_));
 sky130_fd_sc_hd__o21ai_0 _16134_ (.A1(_06996_),
    .A2(_06999_),
    .B1(_07005_),
    .Y(_07006_));
 sky130_fd_sc_hd__a21oi_1 _16135_ (.A1(net4037),
    .A2(_06714_),
    .B1(net3699),
    .Y(_07007_));
 sky130_fd_sc_hd__o22ai_1 _16136_ (.A1(net4035),
    .A2(net4033),
    .B1(_07007_),
    .B2(_12010_[0]),
    .Y(_07008_));
 sky130_fd_sc_hd__nand2_1 _16137_ (.A(net3703),
    .B(net4032),
    .Y(_07009_));
 sky130_fd_sc_hd__o21ai_0 _16138_ (.A1(net3703),
    .A2(_06968_),
    .B1(_07009_),
    .Y(_07010_));
 sky130_fd_sc_hd__o21ai_1 _16139_ (.A1(net4032),
    .A2(_06785_),
    .B1(_06788_),
    .Y(_07011_));
 sky130_fd_sc_hd__o2111ai_1 _16140_ (.A1(_06696_),
    .A2(_06855_),
    .B1(_07011_),
    .C1(net4019),
    .D1(_06940_),
    .Y(_07012_));
 sky130_fd_sc_hd__a221o_1 _16141_ (.A1(_06569_),
    .A2(_07008_),
    .B1(_07010_),
    .B2(net4036),
    .C1(_07012_),
    .X(_07013_));
 sky130_fd_sc_hd__o311ai_0 _16142_ (.A1(_06612_),
    .A2(net4019),
    .A3(_06994_),
    .B1(_07006_),
    .C1(_07013_),
    .Y(_07014_));
 sky130_fd_sc_hd__o21ai_0 _16143_ (.A1(_06659_),
    .A2(_06755_),
    .B1(net3701),
    .Y(_07015_));
 sky130_fd_sc_hd__nand3_1 _16144_ (.A(net4033),
    .B(_06620_),
    .C(_06757_),
    .Y(_07016_));
 sky130_fd_sc_hd__nand3_1 _16145_ (.A(_06656_),
    .B(_07015_),
    .C(_07016_),
    .Y(_07017_));
 sky130_fd_sc_hd__a21oi_2 _16146_ (.A1(_12006_[0]),
    .A2(net4021),
    .B1(_06719_),
    .Y(_07018_));
 sky130_fd_sc_hd__nor2_1 _16147_ (.A(net399),
    .B(net3589),
    .Y(_07019_));
 sky130_fd_sc_hd__nor3_1 _16148_ (.A(net4034),
    .B(_06780_),
    .C(_07019_),
    .Y(_07020_));
 sky130_fd_sc_hd__a21oi_2 _16149_ (.A1(net4034),
    .A2(_07018_),
    .B1(_07020_),
    .Y(_07021_));
 sky130_fd_sc_hd__o21ai_0 _16150_ (.A1(_11996_[0]),
    .A2(net4021),
    .B1(_06869_),
    .Y(_07022_));
 sky130_fd_sc_hd__a221o_1 _16151_ (.A1(_11998_[0]),
    .A2(_06579_),
    .B1(_07022_),
    .B2(net4033),
    .C1(net4016),
    .X(_07023_));
 sky130_fd_sc_hd__o211ai_1 _16152_ (.A1(net4019),
    .A2(_07021_),
    .B1(_07023_),
    .C1(net4017),
    .Y(_07024_));
 sky130_fd_sc_hd__o21ai_2 _16153_ (.A1(net3704),
    .A2(net3701),
    .B1(_06653_),
    .Y(_07025_));
 sky130_fd_sc_hd__o311ai_1 _16154_ (.A1(_12013_[0]),
    .A2(_12022_[0]),
    .A3(net4021),
    .B1(_06914_),
    .C1(_07025_),
    .Y(_07026_));
 sky130_fd_sc_hd__a31oi_1 _16155_ (.A1(_07017_),
    .A2(_07024_),
    .A3(_07026_),
    .B1(_06671_),
    .Y(_07027_));
 sky130_fd_sc_hd__a211o_1 _16156_ (.A1(_06702_),
    .A2(_06990_),
    .B1(_07014_),
    .C1(_07027_),
    .X(_00046_));
 sky130_fd_sc_hd__o221ai_1 _16157_ (.A1(_12010_[0]),
    .A2(_06553_),
    .B1(_06637_),
    .B2(net3635),
    .C1(_06754_),
    .Y(_07028_));
 sky130_fd_sc_hd__a21oi_1 _16158_ (.A1(_06793_),
    .A2(_06713_),
    .B1(net4033),
    .Y(_07029_));
 sky130_fd_sc_hd__a211oi_1 _16159_ (.A1(net4033),
    .A2(_06786_),
    .B1(_07029_),
    .C1(net4017),
    .Y(_07030_));
 sky130_fd_sc_hd__a21o_1 _16160_ (.A1(net4017),
    .A2(_07028_),
    .B1(_07030_),
    .X(_07031_));
 sky130_fd_sc_hd__a21oi_1 _16161_ (.A1(_06841_),
    .A2(_06813_),
    .B1(net4037),
    .Y(_07032_));
 sky130_fd_sc_hd__a221oi_1 _16162_ (.A1(_11996_[0]),
    .A2(_06540_),
    .B1(_06573_),
    .B2(net4036),
    .C1(_07032_),
    .Y(_07033_));
 sky130_fd_sc_hd__o21ai_0 _16163_ (.A1(_12006_[0]),
    .A2(_06684_),
    .B1(net4032),
    .Y(_07034_));
 sky130_fd_sc_hd__a31oi_1 _16164_ (.A1(net4034),
    .A2(_06713_),
    .A3(_06757_),
    .B1(_07034_),
    .Y(_07035_));
 sky130_fd_sc_hd__a2111oi_0 _16165_ (.A1(net4018),
    .A2(_07033_),
    .B1(_07035_),
    .C1(net4016),
    .D1(_06612_),
    .Y(_07036_));
 sky130_fd_sc_hd__a31oi_1 _16166_ (.A1(_06940_),
    .A2(net4016),
    .A3(_07031_),
    .B1(net3572),
    .Y(_07037_));
 sky130_fd_sc_hd__nand2_1 _16167_ (.A(_11998_[0]),
    .B(_06573_),
    .Y(_07038_));
 sky130_fd_sc_hd__o21ai_0 _16168_ (.A1(_12008_[0]),
    .A2(net4031),
    .B1(_07038_),
    .Y(_07039_));
 sky130_fd_sc_hd__a21oi_1 _16169_ (.A1(_06914_),
    .A2(_07039_),
    .B1(_06631_),
    .Y(_07040_));
 sky130_fd_sc_hd__o311ai_0 _16170_ (.A1(_06505_),
    .A2(_06704_),
    .A3(_06658_),
    .B1(_06663_),
    .C1(_06746_),
    .Y(_07041_));
 sky130_fd_sc_hd__a21oi_1 _16171_ (.A1(_12006_[0]),
    .A2(net4033),
    .B1(_06694_),
    .Y(_07042_));
 sky130_fd_sc_hd__nor2_1 _16172_ (.A(_12022_[0]),
    .B(net4031),
    .Y(_07043_));
 sky130_fd_sc_hd__a21oi_1 _16173_ (.A1(net4031),
    .A2(_07042_),
    .B1(_07043_),
    .Y(_07044_));
 sky130_fd_sc_hd__o21ai_1 _16174_ (.A1(_12001_[0]),
    .A2(net3701),
    .B1(_06992_),
    .Y(_07045_));
 sky130_fd_sc_hd__a221oi_1 _16175_ (.A1(_06704_),
    .A2(_06696_),
    .B1(_07045_),
    .B2(net4021),
    .C1(_06626_),
    .Y(_07046_));
 sky130_fd_sc_hd__a21oi_1 _16176_ (.A1(_06656_),
    .A2(_07044_),
    .B1(_07046_),
    .Y(_07047_));
 sky130_fd_sc_hd__nand3_2 _16177_ (.A(_07040_),
    .B(_07041_),
    .C(_07047_),
    .Y(_07048_));
 sky130_fd_sc_hd__mux2i_1 _16178_ (.A0(net3635),
    .A1(_12004_[0]),
    .S(_06505_),
    .Y(_07049_));
 sky130_fd_sc_hd__o21ai_0 _16179_ (.A1(_06855_),
    .A2(_07049_),
    .B1(net4019),
    .Y(_07050_));
 sky130_fd_sc_hd__nor3_1 _16180_ (.A(net4038),
    .B(net4036),
    .C(net4033),
    .Y(_07051_));
 sky130_fd_sc_hd__a21oi_1 _16181_ (.A1(_11996_[0]),
    .A2(net4033),
    .B1(_07051_),
    .Y(_07052_));
 sky130_fd_sc_hd__nor2_1 _16182_ (.A(net4032),
    .B(_06583_),
    .Y(_07053_));
 sky130_fd_sc_hd__o221ai_1 _16183_ (.A1(_06553_),
    .A2(net3589),
    .B1(_07018_),
    .B2(net4034),
    .C1(_07053_),
    .Y(_07054_));
 sky130_fd_sc_hd__o21ai_0 _16184_ (.A1(_06857_),
    .A2(_07052_),
    .B1(_07054_),
    .Y(_07055_));
 sky130_fd_sc_hd__nor2_1 _16185_ (.A(net4032),
    .B(_06901_),
    .Y(_07056_));
 sky130_fd_sc_hd__nand3_1 _16186_ (.A(net3702),
    .B(_06616_),
    .C(_06713_),
    .Y(_07057_));
 sky130_fd_sc_hd__o21ai_0 _16187_ (.A1(_11996_[0]),
    .A2(net3702),
    .B1(_07057_),
    .Y(_07058_));
 sky130_fd_sc_hd__a22oi_1 _16188_ (.A1(_07025_),
    .A2(_07056_),
    .B1(_07058_),
    .B2(net4032),
    .Y(_07059_));
 sky130_fd_sc_hd__inv_1 _16189_ (.A(_06671_),
    .Y(_07060_));
 sky130_fd_sc_hd__o221ai_1 _16190_ (.A1(_07050_),
    .A2(_07055_),
    .B1(_07059_),
    .B2(net4019),
    .C1(_07060_),
    .Y(_07061_));
 sky130_fd_sc_hd__o21ai_0 _16191_ (.A1(net4036),
    .A2(_06575_),
    .B1(_06684_),
    .Y(_07062_));
 sky130_fd_sc_hd__a21oi_1 _16192_ (.A1(_06736_),
    .A2(_06724_),
    .B1(net4032),
    .Y(_07063_));
 sky130_fd_sc_hd__o21ai_0 _16193_ (.A1(_06573_),
    .A2(_06863_),
    .B1(net4037),
    .Y(_07064_));
 sky130_fd_sc_hd__a21oi_1 _16194_ (.A1(_06911_),
    .A2(_07064_),
    .B1(net4018),
    .Y(_07065_));
 sky130_fd_sc_hd__a211oi_1 _16195_ (.A1(net3703),
    .A2(_07062_),
    .B1(_07063_),
    .C1(_07065_),
    .Y(_07066_));
 sky130_fd_sc_hd__a21oi_1 _16196_ (.A1(_06642_),
    .A2(_06855_),
    .B1(net4036),
    .Y(_07067_));
 sky130_fd_sc_hd__a31oi_1 _16197_ (.A1(net4036),
    .A2(net4018),
    .A3(net3622),
    .B1(_07067_),
    .Y(_07068_));
 sky130_fd_sc_hd__a211oi_1 _16198_ (.A1(net3635),
    .A2(_06725_),
    .B1(_06935_),
    .C1(net4019),
    .Y(_07069_));
 sky130_fd_sc_hd__o21ai_0 _16199_ (.A1(net4037),
    .A2(_07068_),
    .B1(_07069_),
    .Y(_07070_));
 sky130_fd_sc_hd__o211ai_1 _16200_ (.A1(net4016),
    .A2(_07066_),
    .B1(_07070_),
    .C1(_06702_),
    .Y(_07071_));
 sky130_fd_sc_hd__and4_4 _16201_ (.A(_07037_),
    .B(_07048_),
    .C(_07061_),
    .D(_07071_),
    .X(_00047_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_907 ();
 sky130_fd_sc_hd__xnor2_1 _16204_ (.A(\sa02_sr[7] ),
    .B(\sa02_sr[0] ),
    .Y(_07074_));
 sky130_fd_sc_hd__xor2_1 _16205_ (.A(\sa20_sub[1] ),
    .B(\sa31_sub[1] ),
    .X(_07075_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_905 ();
 sky130_fd_sc_hd__xor3_1 _16208_ (.A(\sa12_sr[7] ),
    .B(\sa12_sr[0] ),
    .C(\sa12_sr[1] ),
    .X(_07078_));
 sky130_fd_sc_hd__xnor3_1 _16209_ (.A(_07074_),
    .B(_07075_),
    .C(_07078_),
    .X(_07079_));
 sky130_fd_sc_hd__mux2i_2 _16210_ (.A0(\text_in_r[57] ),
    .A1(_07079_),
    .S(net4111),
    .Y(_07080_));
 sky130_fd_sc_hd__xor2_4 _16211_ (.A(net4137),
    .B(_07080_),
    .X(_07081_));
 sky130_fd_sc_hd__inv_16 _16212_ (.A(net406),
    .Y(_07082_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_903 ();
 sky130_fd_sc_hd__xor2_2 _16215_ (.A(net4223),
    .B(net4212),
    .X(_07084_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_902 ();
 sky130_fd_sc_hd__xnor3_1 _16217_ (.A(\sa12_sr[0] ),
    .B(net4201),
    .C(\sa31_sub[0] ),
    .X(_07086_));
 sky130_fd_sc_hd__xnor2_1 _16218_ (.A(_07084_),
    .B(_07086_),
    .Y(_07087_));
 sky130_fd_sc_hd__mux2i_1 _16219_ (.A0(\text_in_r[56] ),
    .A1(_07087_),
    .S(net4111),
    .Y(_07088_));
 sky130_fd_sc_hd__xor2_1 _16220_ (.A(\u0.w[2][24] ),
    .B(_07088_),
    .X(_07089_));
 sky130_fd_sc_hd__clkinv_16 _16221_ (.A(net4012),
    .Y(_07090_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_898 ();
 sky130_fd_sc_hd__xnor3_1 _16226_ (.A(\sa02_sr[1] ),
    .B(net4213),
    .C(net4200),
    .X(_07094_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_897 ();
 sky130_fd_sc_hd__xnor2_1 _16228_ (.A(\sa12_sr[1] ),
    .B(net4184),
    .Y(_07096_));
 sky130_fd_sc_hd__xor2_1 _16229_ (.A(_07094_),
    .B(_07096_),
    .X(_07097_));
 sky130_fd_sc_hd__mux2i_2 _16230_ (.A0(\text_in_r[58] ),
    .A1(_07097_),
    .S(net4114),
    .Y(_07098_));
 sky130_fd_sc_hd__xnor2_4 _16231_ (.A(\u0.w[2][26] ),
    .B(_07098_),
    .Y(_07099_));
 sky130_fd_sc_hd__clkinv_16 _16232_ (.A(_07099_),
    .Y(_07100_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_887 ();
 sky130_fd_sc_hd__xor2_2 _16243_ (.A(\sa12_sr[7] ),
    .B(net4196),
    .X(_07108_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_886 ();
 sky130_fd_sc_hd__xnor2_1 _16245_ (.A(\sa02_sr[6] ),
    .B(\sa31_sub[7] ),
    .Y(_07110_));
 sky130_fd_sc_hd__xnor2_1 _16246_ (.A(_07108_),
    .B(_07110_),
    .Y(_07111_));
 sky130_fd_sc_hd__xnor2_1 _16247_ (.A(\sa12_sr[6] ),
    .B(_07111_),
    .Y(_07112_));
 sky130_fd_sc_hd__nand2_1 _16248_ (.A(net4231),
    .B(\text_in_r[63] ),
    .Y(_07113_));
 sky130_fd_sc_hd__o21a_4 _16249_ (.A1(net4231),
    .A2(_07112_),
    .B1(_07113_),
    .X(_07114_));
 sky130_fd_sc_hd__xor2_4 _16250_ (.A(\u0.w[2][31] ),
    .B(_07114_),
    .X(_07115_));
 sky130_fd_sc_hd__xnor3_1 _16251_ (.A(\sa02_sr[5] ),
    .B(\sa12_sr[6] ),
    .C(\sa20_sub[6] ),
    .X(_07116_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_885 ();
 sky130_fd_sc_hd__xnor2_1 _16253_ (.A(\sa12_sr[5] ),
    .B(\sa31_sub[6] ),
    .Y(_07118_));
 sky130_fd_sc_hd__xnor2_1 _16254_ (.A(_07116_),
    .B(_07118_),
    .Y(_07119_));
 sky130_fd_sc_hd__nor2_2 _16255_ (.A(net4231),
    .B(_07119_),
    .Y(_07120_));
 sky130_fd_sc_hd__a21oi_4 _16256_ (.A1(net4231),
    .A2(\text_in_r[62] ),
    .B1(_07120_),
    .Y(_07121_));
 sky130_fd_sc_hd__xor2_4 _16257_ (.A(\u0.w[2][30] ),
    .B(_07121_),
    .X(_07122_));
 sky130_fd_sc_hd__nand2_2 _16258_ (.A(_07115_),
    .B(_07122_),
    .Y(_07123_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_883 ();
 sky130_fd_sc_hd__xnor3_1 _16261_ (.A(\sa12_sr[4] ),
    .B(\sa20_sub[5] ),
    .C(\sa31_sub[5] ),
    .X(_07126_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_882 ();
 sky130_fd_sc_hd__xor2_1 _16263_ (.A(\sa02_sr[4] ),
    .B(\sa12_sr[5] ),
    .X(_07128_));
 sky130_fd_sc_hd__xnor2_1 _16264_ (.A(_07126_),
    .B(_07128_),
    .Y(_07129_));
 sky130_fd_sc_hd__mux2i_4 _16265_ (.A0(\text_in_r[61] ),
    .A1(_07129_),
    .S(net4111),
    .Y(_07130_));
 sky130_fd_sc_hd__xnor2_2 _16266_ (.A(\u0.w[2][29] ),
    .B(_07130_),
    .Y(_07131_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_879 ();
 sky130_fd_sc_hd__xnor3_1 _16270_ (.A(net4223),
    .B(\sa02_sr[3] ),
    .C(\sa20_sub[4] ),
    .X(_07135_));
 sky130_fd_sc_hd__xnor2_1 _16271_ (.A(\sa12_sr[3] ),
    .B(\sa31_sub[4] ),
    .Y(_07136_));
 sky130_fd_sc_hd__xnor2_1 _16272_ (.A(net4212),
    .B(\sa12_sr[4] ),
    .Y(_07137_));
 sky130_fd_sc_hd__xnor3_1 _16273_ (.A(_07135_),
    .B(_07136_),
    .C(_07137_),
    .X(_07138_));
 sky130_fd_sc_hd__mux2i_4 _16274_ (.A0(\text_in_r[60] ),
    .A1(_07138_),
    .S(net4111),
    .Y(_07139_));
 sky130_fd_sc_hd__xor2_4 _16275_ (.A(\u0.w[2][28] ),
    .B(_07139_),
    .X(_07140_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_875 ();
 sky130_fd_sc_hd__xnor3_1 _16280_ (.A(\sa02_sr[7] ),
    .B(\sa02_sr[2] ),
    .C(net4199),
    .X(_07145_));
 sky130_fd_sc_hd__nor2b_1 _16281_ (.A(net4230),
    .B_N(\u0.w[2][27] ),
    .Y(_07146_));
 sky130_fd_sc_hd__nand2_1 _16282_ (.A(_07145_),
    .B(_07146_),
    .Y(_07147_));
 sky130_fd_sc_hd__xor3_1 _16283_ (.A(\sa02_sr[7] ),
    .B(\sa02_sr[2] ),
    .C(\sa20_sub[3] ),
    .X(_07148_));
 sky130_fd_sc_hd__nor2_1 _16284_ (.A(\u0.w[2][27] ),
    .B(net4230),
    .Y(_07149_));
 sky130_fd_sc_hd__nand2_1 _16285_ (.A(_07148_),
    .B(_07149_),
    .Y(_07150_));
 sky130_fd_sc_hd__xnor2_1 _16286_ (.A(net4212),
    .B(net4213),
    .Y(_07151_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_874 ();
 sky130_fd_sc_hd__xnor2_1 _16288_ (.A(\sa12_sr[3] ),
    .B(net4183),
    .Y(_07153_));
 sky130_fd_sc_hd__xnor2_1 _16289_ (.A(_07151_),
    .B(_07153_),
    .Y(_07154_));
 sky130_fd_sc_hd__a21oi_2 _16290_ (.A1(_07147_),
    .A2(_07150_),
    .B1(_07154_),
    .Y(_07155_));
 sky130_fd_sc_hd__nand2_1 _16291_ (.A(_07145_),
    .B(_07149_),
    .Y(_07156_));
 sky130_fd_sc_hd__nand2_1 _16292_ (.A(_07148_),
    .B(_07146_),
    .Y(_07157_));
 sky130_fd_sc_hd__a21boi_2 _16293_ (.A1(_07156_),
    .A2(_07157_),
    .B1_N(_07154_),
    .Y(_07158_));
 sky130_fd_sc_hd__nand2b_1 _16294_ (.A_N(\u0.w[2][27] ),
    .B(net4230),
    .Y(_07159_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_873 ();
 sky130_fd_sc_hd__nand3_1 _16296_ (.A(\u0.w[2][27] ),
    .B(net4230),
    .C(\text_in_r[59] ),
    .Y(_07161_));
 sky130_fd_sc_hd__o21ai_2 _16297_ (.A1(\text_in_r[59] ),
    .A2(_07159_),
    .B1(_07161_),
    .Y(_07162_));
 sky130_fd_sc_hd__nor3_4 _16298_ (.A(_07155_),
    .B(_07158_),
    .C(_07162_),
    .Y(_07163_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_871 ();
 sky130_fd_sc_hd__nor2_2 _16301_ (.A(_07082_),
    .B(_07090_),
    .Y(_07166_));
 sky130_fd_sc_hd__nor2_4 _16302_ (.A(net4013),
    .B(_07100_),
    .Y(_07167_));
 sky130_fd_sc_hd__nor2_1 _16303_ (.A(_07166_),
    .B(_07167_),
    .Y(_07168_));
 sky130_fd_sc_hd__xnor2_1 _16304_ (.A(net4005),
    .B(_07168_),
    .Y(_07169_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_868 ();
 sky130_fd_sc_hd__a21oi_4 _16308_ (.A1(_07082_),
    .A2(_07090_),
    .B1(net4005),
    .Y(_07173_));
 sky130_fd_sc_hd__or3_4 _16309_ (.A(_07155_),
    .B(_07158_),
    .C(_07162_),
    .X(_07174_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_865 ();
 sky130_fd_sc_hd__nor2_1 _16313_ (.A(_12028_[0]),
    .B(_07174_),
    .Y(_07178_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_862 ();
 sky130_fd_sc_hd__nor2_2 _16317_ (.A(_12036_[0]),
    .B(net4004),
    .Y(_07182_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_859 ();
 sky130_fd_sc_hd__nand2_8 _16321_ (.A(_12029_[0]),
    .B(net4004),
    .Y(_07186_));
 sky130_fd_sc_hd__nand3b_1 _16322_ (.A_N(_07182_),
    .B(net4011),
    .C(_07186_),
    .Y(_07187_));
 sky130_fd_sc_hd__o311ai_0 _16323_ (.A1(net4011),
    .A2(_07173_),
    .A3(_07178_),
    .B1(net4007),
    .C1(_07187_),
    .Y(_07188_));
 sky130_fd_sc_hd__o21ai_2 _16324_ (.A1(net4007),
    .A2(_07169_),
    .B1(_07188_),
    .Y(_07189_));
 sky130_fd_sc_hd__xnor2_1 _16325_ (.A(\u0.w[2][28] ),
    .B(_07139_),
    .Y(_07190_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_857 ();
 sky130_fd_sc_hd__nor2_2 _16328_ (.A(_07082_),
    .B(net4011),
    .Y(_07193_));
 sky130_fd_sc_hd__nor2_4 _16329_ (.A(_12029_[0]),
    .B(_07099_),
    .Y(_07194_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_856 ();
 sky130_fd_sc_hd__nand2_8 _16331_ (.A(net4015),
    .B(_07174_),
    .Y(_07196_));
 sky130_fd_sc_hd__a2bb2oi_1 _16332_ (.A1_N(_07193_),
    .A2_N(_07186_),
    .B1(_07194_),
    .B2(_07196_),
    .Y(_07197_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_855 ();
 sky130_fd_sc_hd__nor2_4 _16334_ (.A(_07100_),
    .B(_07174_),
    .Y(_07199_));
 sky130_fd_sc_hd__nand2_8 _16335_ (.A(_07100_),
    .B(_07174_),
    .Y(_07200_));
 sky130_fd_sc_hd__nor2_4 _16336_ (.A(_12036_[0]),
    .B(_07200_),
    .Y(_07201_));
 sky130_fd_sc_hd__xnor2_2 _16337_ (.A(_07100_),
    .B(_07174_),
    .Y(_07202_));
 sky130_fd_sc_hd__nor2_1 _16338_ (.A(_12028_[0]),
    .B(_07202_),
    .Y(_07203_));
 sky130_fd_sc_hd__a2111oi_0 _16339_ (.A1(_12029_[0]),
    .A2(_07199_),
    .B1(_07201_),
    .C1(_07203_),
    .D1(net4001),
    .Y(_07204_));
 sky130_fd_sc_hd__a211oi_1 _16340_ (.A1(net4001),
    .A2(_07197_),
    .B1(_07204_),
    .C1(net4009),
    .Y(_07205_));
 sky130_fd_sc_hd__a21oi_1 _16341_ (.A1(net4009),
    .A2(_07189_),
    .B1(_07205_),
    .Y(_07206_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_852 ();
 sky130_fd_sc_hd__nor2_4 _16345_ (.A(_12033_[0]),
    .B(_07174_),
    .Y(_07210_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_851 ();
 sky130_fd_sc_hd__nor2_4 _16347_ (.A(_12030_[0]),
    .B(net4005),
    .Y(_07212_));
 sky130_fd_sc_hd__o21ai_2 _16348_ (.A1(_07210_),
    .A2(_07212_),
    .B1(net4010),
    .Y(_07213_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_850 ();
 sky130_fd_sc_hd__nor2_4 _16350_ (.A(net4011),
    .B(net4005),
    .Y(_07215_));
 sky130_fd_sc_hd__nand2_1 _16351_ (.A(_12028_[0]),
    .B(_07215_),
    .Y(_07216_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_849 ();
 sky130_fd_sc_hd__nand2_8 _16353_ (.A(_07090_),
    .B(net4005),
    .Y(_07218_));
 sky130_fd_sc_hd__nor2_4 _16354_ (.A(_12029_[0]),
    .B(net4005),
    .Y(_07219_));
 sky130_fd_sc_hd__nor3_2 _16355_ (.A(net4011),
    .B(_07182_),
    .C(_07219_),
    .Y(_07220_));
 sky130_fd_sc_hd__a311oi_1 _16356_ (.A1(net4011),
    .A2(_07196_),
    .A3(_07218_),
    .B1(_07220_),
    .C1(net4001),
    .Y(_07221_));
 sky130_fd_sc_hd__a311oi_1 _16357_ (.A1(net4001),
    .A2(_07213_),
    .A3(_07216_),
    .B1(_07221_),
    .C1(net3697),
    .Y(_07222_));
 sky130_fd_sc_hd__nand2_4 _16358_ (.A(net4013),
    .B(_07174_),
    .Y(_07223_));
 sky130_fd_sc_hd__nor2_4 _16359_ (.A(net4015),
    .B(_07223_),
    .Y(_07224_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_848 ();
 sky130_fd_sc_hd__nor2_2 _16361_ (.A(_12030_[0]),
    .B(_07174_),
    .Y(_07226_));
 sky130_fd_sc_hd__nor3_1 _16362_ (.A(_07100_),
    .B(_07224_),
    .C(_07226_),
    .Y(_07227_));
 sky130_fd_sc_hd__nand2_1 _16363_ (.A(_07122_),
    .B(net4001),
    .Y(_07228_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_847 ();
 sky130_fd_sc_hd__nand3_4 _16365_ (.A(_07082_),
    .B(net4013),
    .C(net4005),
    .Y(_07230_));
 sky130_fd_sc_hd__o21ai_2 _16366_ (.A1(_12030_[0]),
    .A2(net4005),
    .B1(_07230_),
    .Y(_07231_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_845 ();
 sky130_fd_sc_hd__nor2_4 _16369_ (.A(_07099_),
    .B(_07174_),
    .Y(_07234_));
 sky130_fd_sc_hd__nand2_1 _16370_ (.A(_12038_[0]),
    .B(_07234_),
    .Y(_07235_));
 sky130_fd_sc_hd__o2111ai_1 _16371_ (.A1(_07100_),
    .A2(_07231_),
    .B1(_07235_),
    .C1(_07122_),
    .D1(_07140_),
    .Y(_07236_));
 sky130_fd_sc_hd__xor2_4 _16372_ (.A(\u0.w[2][29] ),
    .B(_07130_),
    .X(_07237_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_844 ();
 sky130_fd_sc_hd__nor2_1 _16374_ (.A(_07115_),
    .B(net4000),
    .Y(_07239_));
 sky130_fd_sc_hd__o311ai_1 _16375_ (.A1(_07201_),
    .A2(_07227_),
    .A3(_07228_),
    .B1(_07236_),
    .C1(_07239_),
    .Y(_07240_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_841 ();
 sky130_fd_sc_hd__a221oi_1 _16379_ (.A1(_12049_[0]),
    .A2(net4005),
    .B1(_07215_),
    .B2(net3634),
    .C1(_07228_),
    .Y(_07244_));
 sky130_fd_sc_hd__nor3_2 _16380_ (.A(net4015),
    .B(_07090_),
    .C(_07100_),
    .Y(_07245_));
 sky130_fd_sc_hd__o21ai_0 _16381_ (.A1(_12033_[0]),
    .A2(net4011),
    .B1(_07174_),
    .Y(_07246_));
 sky130_fd_sc_hd__o21ai_2 _16382_ (.A1(_07245_),
    .A2(_07246_),
    .B1(_07140_),
    .Y(_07247_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_840 ();
 sky130_fd_sc_hd__nand2_1 _16384_ (.A(_12030_[0]),
    .B(_07174_),
    .Y(_07249_));
 sky130_fd_sc_hd__a21oi_1 _16385_ (.A1(_07218_),
    .A2(_07249_),
    .B1(net4011),
    .Y(_07250_));
 sky130_fd_sc_hd__nand2_8 _16386_ (.A(net4010),
    .B(net4005),
    .Y(_07251_));
 sky130_fd_sc_hd__o21ai_0 _16387_ (.A1(_12028_[0]),
    .A2(_07251_),
    .B1(_07122_),
    .Y(_07252_));
 sky130_fd_sc_hd__nor3_1 _16388_ (.A(_07247_),
    .B(_07250_),
    .C(_07252_),
    .Y(_07253_));
 sky130_fd_sc_hd__nor4_1 _16389_ (.A(_07115_),
    .B(net4009),
    .C(_07244_),
    .D(_07253_),
    .Y(_07254_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_839 ();
 sky130_fd_sc_hd__a21oi_4 _16391_ (.A1(_07082_),
    .A2(_07090_),
    .B1(net4004),
    .Y(_07256_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_837 ();
 sky130_fd_sc_hd__nand2_1 _16394_ (.A(net4013),
    .B(_07234_),
    .Y(_07259_));
 sky130_fd_sc_hd__o221ai_1 _16395_ (.A1(_12033_[0]),
    .A2(net4005),
    .B1(_07256_),
    .B2(_07100_),
    .C1(_07259_),
    .Y(_07260_));
 sky130_fd_sc_hd__nor2_4 _16396_ (.A(_12029_[0]),
    .B(_07174_),
    .Y(_07261_));
 sky130_fd_sc_hd__nor2_4 _16397_ (.A(_12038_[0]),
    .B(net4005),
    .Y(_07262_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_836 ();
 sky130_fd_sc_hd__o21ai_0 _16399_ (.A1(_07261_),
    .A2(_07262_),
    .B1(net4011),
    .Y(_07264_));
 sky130_fd_sc_hd__o211ai_1 _16400_ (.A1(_12033_[0]),
    .A2(_07200_),
    .B1(_07264_),
    .C1(net4001),
    .Y(_07265_));
 sky130_fd_sc_hd__xnor2_4 _16401_ (.A(\u0.w[2][30] ),
    .B(_07121_),
    .Y(_07266_));
 sky130_fd_sc_hd__o211ai_1 _16402_ (.A1(net4001),
    .A2(_07260_),
    .B1(_07265_),
    .C1(_07266_),
    .Y(_07267_));
 sky130_fd_sc_hd__a2bb2oi_1 _16403_ (.A1_N(_07222_),
    .A2_N(_07240_),
    .B1(_07254_),
    .B2(_07267_),
    .Y(_07268_));
 sky130_fd_sc_hd__xnor2_4 _16404_ (.A(\u0.w[2][31] ),
    .B(_07114_),
    .Y(_07269_));
 sky130_fd_sc_hd__nor2_2 _16405_ (.A(_07269_),
    .B(net3697),
    .Y(_07270_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_835 ();
 sky130_fd_sc_hd__nand2_8 _16407_ (.A(_12042_[0]),
    .B(net4005),
    .Y(_07272_));
 sky130_fd_sc_hd__nand2_1 _16408_ (.A(_07082_),
    .B(_07174_),
    .Y(_07273_));
 sky130_fd_sc_hd__nor2_1 _16409_ (.A(_07090_),
    .B(net4011),
    .Y(_07274_));
 sky130_fd_sc_hd__a32oi_1 _16410_ (.A1(net4011),
    .A2(_07272_),
    .A3(_07273_),
    .B1(_07274_),
    .B2(_07196_),
    .Y(_07275_));
 sky130_fd_sc_hd__nor2_1 _16411_ (.A(net4009),
    .B(_07275_),
    .Y(_07276_));
 sky130_fd_sc_hd__a21oi_1 _16412_ (.A1(_07196_),
    .A2(_07272_),
    .B1(net4011),
    .Y(_07277_));
 sky130_fd_sc_hd__nor2_4 _16413_ (.A(net4013),
    .B(net4005),
    .Y(_07278_));
 sky130_fd_sc_hd__a2111oi_0 _16414_ (.A1(_12029_[0]),
    .A2(_07199_),
    .B1(_07277_),
    .C1(_07278_),
    .D1(net4000),
    .Y(_07279_));
 sky130_fd_sc_hd__o21ai_0 _16415_ (.A1(_07276_),
    .A2(_07279_),
    .B1(net4001),
    .Y(_07280_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_834 ();
 sky130_fd_sc_hd__a21oi_1 _16417_ (.A1(_07090_),
    .A2(net3620),
    .B1(_07215_),
    .Y(_07281_));
 sky130_fd_sc_hd__nand2_2 _16418_ (.A(net4011),
    .B(_07174_),
    .Y(_07282_));
 sky130_fd_sc_hd__o221ai_1 _16419_ (.A1(net407),
    .A2(_07281_),
    .B1(_07282_),
    .B2(_12030_[0]),
    .C1(_07259_),
    .Y(_07283_));
 sky130_fd_sc_hd__nor2_4 _16420_ (.A(_07082_),
    .B(_07174_),
    .Y(_07284_));
 sky130_fd_sc_hd__o32a_1 _16421_ (.A1(_07090_),
    .A2(net4011),
    .A3(_07284_),
    .B1(_07251_),
    .B2(_12033_[0]),
    .X(_07285_));
 sky130_fd_sc_hd__a21oi_1 _16422_ (.A1(net4009),
    .A2(_07285_),
    .B1(net4001),
    .Y(_07286_));
 sky130_fd_sc_hd__o21ai_0 _16423_ (.A1(net4009),
    .A2(_07283_),
    .B1(_07286_),
    .Y(_07287_));
 sky130_fd_sc_hd__nand3_1 _16424_ (.A(_07270_),
    .B(_07280_),
    .C(_07287_),
    .Y(_07288_));
 sky130_fd_sc_hd__o211ai_1 _16425_ (.A1(_07123_),
    .A2(_07206_),
    .B1(_07268_),
    .C1(_07288_),
    .Y(_00048_));
 sky130_fd_sc_hd__nand2b_4 _16426_ (.A_N(_12029_[0]),
    .B(net4005),
    .Y(_07289_));
 sky130_fd_sc_hd__nand2_4 _16427_ (.A(_07289_),
    .B(_07223_),
    .Y(_07290_));
 sky130_fd_sc_hd__a211o_1 _16428_ (.A1(_12028_[0]),
    .A2(net4005),
    .B1(_07212_),
    .C1(_07100_),
    .X(_07291_));
 sky130_fd_sc_hd__o21ai_0 _16429_ (.A1(net4010),
    .A2(_07290_),
    .B1(_07291_),
    .Y(_07292_));
 sky130_fd_sc_hd__nor3_1 _16430_ (.A(net4014),
    .B(net4013),
    .C(_07174_),
    .Y(_07293_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_833 ();
 sky130_fd_sc_hd__o21ai_0 _16432_ (.A1(_07212_),
    .A2(_07293_),
    .B1(_07100_),
    .Y(_07295_));
 sky130_fd_sc_hd__nand2_4 _16433_ (.A(_12042_[0]),
    .B(net4004),
    .Y(_07296_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_832 ();
 sky130_fd_sc_hd__a31oi_1 _16435_ (.A1(net4010),
    .A2(_07289_),
    .A3(_07296_),
    .B1(net4009),
    .Y(_07298_));
 sky130_fd_sc_hd__a221oi_1 _16436_ (.A1(net4009),
    .A2(_07292_),
    .B1(_07295_),
    .B2(_07298_),
    .C1(net4007),
    .Y(_07299_));
 sky130_fd_sc_hd__nor2_2 _16437_ (.A(net4011),
    .B(_07223_),
    .Y(_07300_));
 sky130_fd_sc_hd__nand3_4 _16438_ (.A(_07082_),
    .B(_07090_),
    .C(net4004),
    .Y(_07301_));
 sky130_fd_sc_hd__a21oi_1 _16439_ (.A1(_07289_),
    .A2(_07301_),
    .B1(_07100_),
    .Y(_07302_));
 sky130_fd_sc_hd__o21ai_2 _16440_ (.A1(_07300_),
    .A2(_07302_),
    .B1(net4000),
    .Y(_07303_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_831 ();
 sky130_fd_sc_hd__nor2_2 _16442_ (.A(_12028_[0]),
    .B(net4005),
    .Y(_07305_));
 sky130_fd_sc_hd__o21ai_2 _16443_ (.A1(net4014),
    .A2(_07174_),
    .B1(_07100_),
    .Y(_07306_));
 sky130_fd_sc_hd__nand3_4 _16444_ (.A(_07090_),
    .B(net4010),
    .C(_07174_),
    .Y(_07307_));
 sky130_fd_sc_hd__o221ai_1 _16445_ (.A1(_12033_[0]),
    .A2(_07251_),
    .B1(_07305_),
    .B2(_07306_),
    .C1(_07307_),
    .Y(_07308_));
 sky130_fd_sc_hd__nand2_1 _16446_ (.A(net4009),
    .B(_07308_),
    .Y(_07309_));
 sky130_fd_sc_hd__a21oi_1 _16447_ (.A1(_07303_),
    .A2(_07309_),
    .B1(net4002),
    .Y(_07310_));
 sky130_fd_sc_hd__nor3_1 _16448_ (.A(net3697),
    .B(_07299_),
    .C(_07310_),
    .Y(_07311_));
 sky130_fd_sc_hd__nand2_1 _16449_ (.A(_12036_[0]),
    .B(_07100_),
    .Y(_07312_));
 sky130_fd_sc_hd__nand2_1 _16450_ (.A(_07082_),
    .B(_07167_),
    .Y(_07313_));
 sky130_fd_sc_hd__a31oi_1 _16451_ (.A1(net4004),
    .A2(_07312_),
    .A3(_07313_),
    .B1(net4001),
    .Y(_07314_));
 sky130_fd_sc_hd__o31a_1 _16452_ (.A1(_12052_[0]),
    .A2(net4009),
    .A3(net4004),
    .B1(_07314_),
    .X(_07315_));
 sky130_fd_sc_hd__o21ai_0 _16453_ (.A1(_07278_),
    .A2(_07210_),
    .B1(net4011),
    .Y(_07316_));
 sky130_fd_sc_hd__nor2_4 _16454_ (.A(net4015),
    .B(net4005),
    .Y(_07317_));
 sky130_fd_sc_hd__o21ai_2 _16455_ (.A1(_07284_),
    .A2(_07317_),
    .B1(_07100_),
    .Y(_07318_));
 sky130_fd_sc_hd__nand2_8 _16456_ (.A(net4001),
    .B(net4000),
    .Y(_07319_));
 sky130_fd_sc_hd__a21oi_2 _16457_ (.A1(_07316_),
    .A2(_07318_),
    .B1(_07319_),
    .Y(_07320_));
 sky130_fd_sc_hd__nor2_2 _16458_ (.A(net4015),
    .B(net4004),
    .Y(_07321_));
 sky130_fd_sc_hd__nor2_1 _16459_ (.A(_07090_),
    .B(net3698),
    .Y(_07322_));
 sky130_fd_sc_hd__nor2_2 _16460_ (.A(net4013),
    .B(net4011),
    .Y(_07323_));
 sky130_fd_sc_hd__nor2_2 _16461_ (.A(_07322_),
    .B(_07323_),
    .Y(_07324_));
 sky130_fd_sc_hd__nand2_4 _16462_ (.A(_07321_),
    .B(_07324_),
    .Y(_07325_));
 sky130_fd_sc_hd__nor2_4 _16463_ (.A(_07100_),
    .B(net4005),
    .Y(_07326_));
 sky130_fd_sc_hd__nand2_4 _16464_ (.A(net4013),
    .B(_07326_),
    .Y(_07327_));
 sky130_fd_sc_hd__nand2_8 _16465_ (.A(net4001),
    .B(net4009),
    .Y(_07328_));
 sky130_fd_sc_hd__a31oi_1 _16466_ (.A1(_07216_),
    .A2(_07325_),
    .A3(_07327_),
    .B1(_07328_),
    .Y(_07329_));
 sky130_fd_sc_hd__o41ai_1 _16467_ (.A1(_07266_),
    .A2(_07315_),
    .A3(_07320_),
    .A4(_07329_),
    .B1(_07115_),
    .Y(_07330_));
 sky130_fd_sc_hd__o22ai_1 _16468_ (.A1(_12033_[0]),
    .A2(_07200_),
    .B1(_07202_),
    .B2(net4015),
    .Y(_07331_));
 sky130_fd_sc_hd__nor2_4 _16469_ (.A(_07131_),
    .B(_07163_),
    .Y(_07332_));
 sky130_fd_sc_hd__o21ai_0 _16470_ (.A1(_12033_[0]),
    .A2(net4011),
    .B1(_07332_),
    .Y(_07333_));
 sky130_fd_sc_hd__mux2i_1 _16471_ (.A0(_12029_[0]),
    .A1(_12042_[0]),
    .S(net4011),
    .Y(_07334_));
 sky130_fd_sc_hd__o21ai_0 _16472_ (.A1(_07174_),
    .A2(_07334_),
    .B1(_07140_),
    .Y(_07335_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_830 ();
 sky130_fd_sc_hd__a2bb2oi_1 _16474_ (.A1_N(_07245_),
    .A2_N(_07333_),
    .B1(_07335_),
    .B2(net4000),
    .Y(_07337_));
 sky130_fd_sc_hd__a211oi_1 _16475_ (.A1(net4003),
    .A2(_07331_),
    .B1(_07337_),
    .C1(_07266_),
    .Y(_07338_));
 sky130_fd_sc_hd__nand2_2 _16476_ (.A(net4001),
    .B(net4004),
    .Y(_07339_));
 sky130_fd_sc_hd__nor3_1 _16477_ (.A(_12033_[0]),
    .B(_07100_),
    .C(_07339_),
    .Y(_07340_));
 sky130_fd_sc_hd__a21oi_1 _16478_ (.A1(_12029_[0]),
    .A2(net4002),
    .B1(_07251_),
    .Y(_07341_));
 sky130_fd_sc_hd__a22oi_1 _16479_ (.A1(net4011),
    .A2(_07140_),
    .B1(_07234_),
    .B2(net4013),
    .Y(_07342_));
 sky130_fd_sc_hd__nor2_4 _16480_ (.A(_07090_),
    .B(_07174_),
    .Y(_07343_));
 sky130_fd_sc_hd__o211ai_1 _16481_ (.A1(_07278_),
    .A2(_07343_),
    .B1(_07100_),
    .C1(net4003),
    .Y(_07344_));
 sky130_fd_sc_hd__a311oi_1 _16482_ (.A1(net4008),
    .A2(net4004),
    .A3(_07166_),
    .B1(net4000),
    .C1(_07266_),
    .Y(_07345_));
 sky130_fd_sc_hd__o211ai_1 _16483_ (.A1(net4015),
    .A2(_07342_),
    .B1(_07344_),
    .C1(_07345_),
    .Y(_07346_));
 sky130_fd_sc_hd__nor3_1 _16484_ (.A(_07340_),
    .B(_07341_),
    .C(_07346_),
    .Y(_07347_));
 sky130_fd_sc_hd__nor3_1 _16485_ (.A(_07115_),
    .B(_07338_),
    .C(_07347_),
    .Y(_07348_));
 sky130_fd_sc_hd__nor2_4 _16486_ (.A(_07090_),
    .B(net4005),
    .Y(_07349_));
 sky130_fd_sc_hd__nor2_2 _16487_ (.A(net4006),
    .B(net4009),
    .Y(_07350_));
 sky130_fd_sc_hd__o21ai_0 _16488_ (.A1(_07261_),
    .A2(_07305_),
    .B1(net4010),
    .Y(_07351_));
 sky130_fd_sc_hd__o311ai_0 _16489_ (.A1(net4010),
    .A2(_07210_),
    .A3(_07349_),
    .B1(_07350_),
    .C1(_07351_),
    .Y(_07352_));
 sky130_fd_sc_hd__nor2_1 _16490_ (.A(net4011),
    .B(_07256_),
    .Y(_07353_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_829 ();
 sky130_fd_sc_hd__nand2_2 _16492_ (.A(net4010),
    .B(_07289_),
    .Y(_07355_));
 sky130_fd_sc_hd__a21oi_1 _16493_ (.A1(_12033_[0]),
    .A2(net4004),
    .B1(_07355_),
    .Y(_07356_));
 sky130_fd_sc_hd__a22oi_1 _16494_ (.A1(net4015),
    .A2(_07199_),
    .B1(_07272_),
    .B2(_07100_),
    .Y(_07357_));
 sky130_fd_sc_hd__nand3_1 _16495_ (.A(net4002),
    .B(_07301_),
    .C(_07357_),
    .Y(_07358_));
 sky130_fd_sc_hd__o311ai_0 _16496_ (.A1(net4002),
    .A2(_07353_),
    .A3(_07356_),
    .B1(_07358_),
    .C1(net4009),
    .Y(_07359_));
 sky130_fd_sc_hd__nand2_1 _16497_ (.A(_12029_[0]),
    .B(_07215_),
    .Y(_07360_));
 sky130_fd_sc_hd__o221ai_1 _16498_ (.A1(_07090_),
    .A2(_07202_),
    .B1(_07218_),
    .B2(_07082_),
    .C1(_07360_),
    .Y(_07361_));
 sky130_fd_sc_hd__nor2_4 _16499_ (.A(net4001),
    .B(net4009),
    .Y(_07362_));
 sky130_fd_sc_hd__a21oi_1 _16500_ (.A1(_07361_),
    .A2(_07362_),
    .B1(net3697),
    .Y(_07363_));
 sky130_fd_sc_hd__nand3_1 _16501_ (.A(_07352_),
    .B(_07359_),
    .C(_07363_),
    .Y(_07364_));
 sky130_fd_sc_hd__a2bb2oi_1 _16502_ (.A1_N(_07311_),
    .A2_N(_07330_),
    .B1(_07348_),
    .B2(_07364_),
    .Y(_00049_));
 sky130_fd_sc_hd__and2_4 _16503_ (.A(_12033_[0]),
    .B(net3698),
    .X(_07365_));
 sky130_fd_sc_hd__a211oi_1 _16504_ (.A1(net3634),
    .A2(net4010),
    .B1(_07237_),
    .C1(_07365_),
    .Y(_07366_));
 sky130_fd_sc_hd__a21oi_1 _16505_ (.A1(_12047_[0]),
    .A2(_07237_),
    .B1(_07366_),
    .Y(_07367_));
 sky130_fd_sc_hd__o21ai_0 _16506_ (.A1(net4015),
    .A2(_07090_),
    .B1(_07237_),
    .Y(_07368_));
 sky130_fd_sc_hd__a221oi_1 _16507_ (.A1(_12028_[0]),
    .A2(net4009),
    .B1(_07368_),
    .B2(net3698),
    .C1(net4005),
    .Y(_07369_));
 sky130_fd_sc_hd__a21oi_1 _16508_ (.A1(net4005),
    .A2(_07367_),
    .B1(_07369_),
    .Y(_07370_));
 sky130_fd_sc_hd__nand2_4 _16509_ (.A(_07269_),
    .B(_07122_),
    .Y(_07371_));
 sky130_fd_sc_hd__nor2_2 _16510_ (.A(net4001),
    .B(_07371_),
    .Y(_07372_));
 sky130_fd_sc_hd__nand3_2 _16511_ (.A(_07269_),
    .B(_07122_),
    .C(net4003),
    .Y(_07373_));
 sky130_fd_sc_hd__nor2_4 _16512_ (.A(_12030_[0]),
    .B(_12033_[0]),
    .Y(_07374_));
 sky130_fd_sc_hd__nor2_2 _16513_ (.A(net4004),
    .B(_07374_),
    .Y(_07375_));
 sky130_fd_sc_hd__nor3_1 _16514_ (.A(_07100_),
    .B(_07173_),
    .C(_07375_),
    .Y(_07376_));
 sky130_fd_sc_hd__nor2_1 _16515_ (.A(_12036_[0]),
    .B(net4005),
    .Y(_07377_));
 sky130_fd_sc_hd__nor3_1 _16516_ (.A(net4010),
    .B(_07256_),
    .C(_07377_),
    .Y(_07378_));
 sky130_fd_sc_hd__nand2_4 _16517_ (.A(_07082_),
    .B(net4005),
    .Y(_07379_));
 sky130_fd_sc_hd__o221ai_1 _16518_ (.A1(_12056_[0]),
    .A2(net4005),
    .B1(_07379_),
    .B2(_07323_),
    .C1(_07237_),
    .Y(_07380_));
 sky130_fd_sc_hd__o31ai_1 _16519_ (.A1(_07237_),
    .A2(_07376_),
    .A3(_07378_),
    .B1(_07380_),
    .Y(_07381_));
 sky130_fd_sc_hd__o2bb2ai_1 _16520_ (.A1_N(_07370_),
    .A2_N(_07372_),
    .B1(_07373_),
    .B2(_07381_),
    .Y(_07382_));
 sky130_fd_sc_hd__nand2_1 _16521_ (.A(_07082_),
    .B(_07100_),
    .Y(_07383_));
 sky130_fd_sc_hd__o32ai_1 _16522_ (.A1(_07278_),
    .A2(_07343_),
    .A3(_07383_),
    .B1(_07251_),
    .B2(_12042_[0]),
    .Y(_07384_));
 sky130_fd_sc_hd__nor3_1 _16523_ (.A(net4011),
    .B(_07219_),
    .C(_07210_),
    .Y(_07385_));
 sky130_fd_sc_hd__a311oi_1 _16524_ (.A1(net4011),
    .A2(_07196_),
    .A3(_07230_),
    .B1(_07385_),
    .C1(net4009),
    .Y(_07386_));
 sky130_fd_sc_hd__a21oi_1 _16525_ (.A1(net4009),
    .A2(_07384_),
    .B1(_07386_),
    .Y(_07387_));
 sky130_fd_sc_hd__nor3_1 _16526_ (.A(_07100_),
    .B(_07219_),
    .C(_07343_),
    .Y(_07388_));
 sky130_fd_sc_hd__nor3_1 _16527_ (.A(net4011),
    .B(_07317_),
    .C(_07226_),
    .Y(_07389_));
 sky130_fd_sc_hd__nor2_1 _16528_ (.A(_07388_),
    .B(_07389_),
    .Y(_07390_));
 sky130_fd_sc_hd__nor2_4 _16529_ (.A(_12042_[0]),
    .B(net4005),
    .Y(_07391_));
 sky130_fd_sc_hd__nor2_2 _16530_ (.A(_07343_),
    .B(_07391_),
    .Y(_07392_));
 sky130_fd_sc_hd__a221oi_1 _16531_ (.A1(_12033_[0]),
    .A2(_07326_),
    .B1(_07392_),
    .B2(_07100_),
    .C1(_07284_),
    .Y(_07393_));
 sky130_fd_sc_hd__nor2_4 _16532_ (.A(_07269_),
    .B(_07266_),
    .Y(_07394_));
 sky130_fd_sc_hd__o221ai_1 _16533_ (.A1(_07328_),
    .A2(_07390_),
    .B1(_07393_),
    .B2(_07319_),
    .C1(_07394_),
    .Y(_07395_));
 sky130_fd_sc_hd__a21oi_1 _16534_ (.A1(_07140_),
    .A2(_07387_),
    .B1(_07395_),
    .Y(_07396_));
 sky130_fd_sc_hd__nand2_4 _16535_ (.A(_07115_),
    .B(_07266_),
    .Y(_07397_));
 sky130_fd_sc_hd__nand2_2 _16536_ (.A(_12038_[0]),
    .B(net4004),
    .Y(_07398_));
 sky130_fd_sc_hd__o21ai_0 _16537_ (.A1(_12033_[0]),
    .A2(net4011),
    .B1(_07362_),
    .Y(_07399_));
 sky130_fd_sc_hd__a31oi_1 _16538_ (.A1(net4011),
    .A2(_07379_),
    .A3(_07398_),
    .B1(_07399_),
    .Y(_07400_));
 sky130_fd_sc_hd__nor2_1 _16539_ (.A(net4011),
    .B(_07261_),
    .Y(_07401_));
 sky130_fd_sc_hd__nand2_2 _16540_ (.A(_07140_),
    .B(net4009),
    .Y(_07402_));
 sky130_fd_sc_hd__a221oi_1 _16541_ (.A1(net4011),
    .A2(_07290_),
    .B1(_07401_),
    .B2(_07398_),
    .C1(_07402_),
    .Y(_07403_));
 sky130_fd_sc_hd__o211ai_1 _16542_ (.A1(_12038_[0]),
    .A2(_07174_),
    .B1(_07223_),
    .C1(net4011),
    .Y(_07404_));
 sky130_fd_sc_hd__nand2b_2 _16543_ (.A_N(_12042_[0]),
    .B(net4004),
    .Y(_07405_));
 sky130_fd_sc_hd__nand3_1 _16544_ (.A(_07100_),
    .B(_07379_),
    .C(_07405_),
    .Y(_07406_));
 sky130_fd_sc_hd__nor3_1 _16545_ (.A(_07100_),
    .B(_07343_),
    .C(_07262_),
    .Y(_07407_));
 sky130_fd_sc_hd__nor3_1 _16546_ (.A(net4011),
    .B(_07210_),
    .C(_07391_),
    .Y(_07408_));
 sky130_fd_sc_hd__nor3_1 _16547_ (.A(net4009),
    .B(_07407_),
    .C(_07408_),
    .Y(_07409_));
 sky130_fd_sc_hd__a311oi_1 _16548_ (.A1(net4009),
    .A2(_07404_),
    .A3(_07406_),
    .B1(_07409_),
    .C1(net4008),
    .Y(_07410_));
 sky130_fd_sc_hd__nor4_1 _16549_ (.A(_07397_),
    .B(_07400_),
    .C(_07403_),
    .D(_07410_),
    .Y(_07411_));
 sky130_fd_sc_hd__a21oi_1 _16550_ (.A1(_12049_[0]),
    .A2(_07174_),
    .B1(net4000),
    .Y(_07412_));
 sky130_fd_sc_hd__o31ai_1 _16551_ (.A1(_07174_),
    .A2(_07194_),
    .A3(_07245_),
    .B1(_07412_),
    .Y(_07413_));
 sky130_fd_sc_hd__nand2_1 _16552_ (.A(_07082_),
    .B(net4010),
    .Y(_07414_));
 sky130_fd_sc_hd__o211ai_1 _16553_ (.A1(_07082_),
    .A2(_07090_),
    .B1(net4005),
    .C1(_07414_),
    .Y(_07415_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_828 ();
 sky130_fd_sc_hd__o211ai_1 _16555_ (.A1(_12052_[0]),
    .A2(net4005),
    .B1(_07415_),
    .C1(_07237_),
    .Y(_07417_));
 sky130_fd_sc_hd__nand2_2 _16556_ (.A(_12036_[0]),
    .B(net4005),
    .Y(_07418_));
 sky130_fd_sc_hd__nand2_1 _16557_ (.A(_12028_[0]),
    .B(net4004),
    .Y(_07419_));
 sky130_fd_sc_hd__a32oi_1 _16558_ (.A1(net4011),
    .A2(_07196_),
    .A3(_07418_),
    .B1(_07419_),
    .B2(_07401_),
    .Y(_07420_));
 sky130_fd_sc_hd__o21ai_0 _16559_ (.A1(_07317_),
    .A2(_07193_),
    .B1(_12029_[0]),
    .Y(_07421_));
 sky130_fd_sc_hd__nand2_4 _16560_ (.A(_07090_),
    .B(net4011),
    .Y(_07422_));
 sky130_fd_sc_hd__a32oi_1 _16561_ (.A1(_07082_),
    .A2(net4011),
    .A3(_07218_),
    .B1(_07422_),
    .B2(_07284_),
    .Y(_07423_));
 sky130_fd_sc_hd__a21oi_1 _16562_ (.A1(_07421_),
    .A2(_07423_),
    .B1(net4000),
    .Y(_07424_));
 sky130_fd_sc_hd__a211oi_1 _16563_ (.A1(net4000),
    .A2(_07420_),
    .B1(_07424_),
    .C1(net4008),
    .Y(_07425_));
 sky130_fd_sc_hd__nand2_4 _16564_ (.A(_07269_),
    .B(_07266_),
    .Y(_07426_));
 sky130_fd_sc_hd__a311oi_1 _16565_ (.A1(net4008),
    .A2(_07413_),
    .A3(_07417_),
    .B1(_07425_),
    .C1(_07426_),
    .Y(_07427_));
 sky130_fd_sc_hd__nor4_1 _16566_ (.A(_07382_),
    .B(_07396_),
    .C(_07411_),
    .D(_07427_),
    .Y(_00050_));
 sky130_fd_sc_hd__nand2_2 _16567_ (.A(_12030_[0]),
    .B(net4005),
    .Y(_07428_));
 sky130_fd_sc_hd__nand2_1 _16568_ (.A(net3634),
    .B(net4009),
    .Y(_07429_));
 sky130_fd_sc_hd__o211ai_1 _16569_ (.A1(net4015),
    .A2(net4009),
    .B1(net4004),
    .C1(_07429_),
    .Y(_07430_));
 sky130_fd_sc_hd__nand2_1 _16570_ (.A(net3634),
    .B(net4005),
    .Y(_07431_));
 sky130_fd_sc_hd__a21oi_1 _16571_ (.A1(_12036_[0]),
    .A2(_07174_),
    .B1(net4009),
    .Y(_07432_));
 sky130_fd_sc_hd__a21oi_1 _16572_ (.A1(_07431_),
    .A2(_07432_),
    .B1(net4011),
    .Y(_07433_));
 sky130_fd_sc_hd__a31oi_1 _16573_ (.A1(net4011),
    .A2(_07428_),
    .A3(_07430_),
    .B1(_07433_),
    .Y(_07434_));
 sky130_fd_sc_hd__nor2_1 _16574_ (.A(_12042_[0]),
    .B(net4004),
    .Y(_07435_));
 sky130_fd_sc_hd__a21oi_1 _16575_ (.A1(net4005),
    .A2(_07374_),
    .B1(_07219_),
    .Y(_07436_));
 sky130_fd_sc_hd__nand2_1 _16576_ (.A(net4010),
    .B(_07436_),
    .Y(_07437_));
 sky130_fd_sc_hd__o311ai_1 _16577_ (.A1(net4010),
    .A2(_07435_),
    .A3(_07349_),
    .B1(_07437_),
    .C1(_07237_),
    .Y(_07438_));
 sky130_fd_sc_hd__nand2_1 _16578_ (.A(_12038_[0]),
    .B(_07202_),
    .Y(_07439_));
 sky130_fd_sc_hd__a31oi_2 _16579_ (.A1(net4009),
    .A2(_07307_),
    .A3(_07439_),
    .B1(net4001),
    .Y(_07440_));
 sky130_fd_sc_hd__a221oi_1 _16580_ (.A1(net4003),
    .A2(_07434_),
    .B1(_07438_),
    .B2(_07440_),
    .C1(_07123_),
    .Y(_07441_));
 sky130_fd_sc_hd__o21ai_0 _16581_ (.A1(_07234_),
    .A2(_07332_),
    .B1(net4013),
    .Y(_07442_));
 sky130_fd_sc_hd__a21oi_1 _16582_ (.A1(_07307_),
    .A2(_07442_),
    .B1(net4015),
    .Y(_07443_));
 sky130_fd_sc_hd__a22oi_1 _16583_ (.A1(_12036_[0]),
    .A2(_07199_),
    .B1(_07194_),
    .B2(_07174_),
    .Y(_07444_));
 sky130_fd_sc_hd__nor2_1 _16584_ (.A(_07237_),
    .B(_07444_),
    .Y(_07445_));
 sky130_fd_sc_hd__a2111oi_2 _16585_ (.A1(_07167_),
    .A2(_07332_),
    .B1(_07443_),
    .C1(_07445_),
    .D1(net4001),
    .Y(_07446_));
 sky130_fd_sc_hd__nor3_1 _16586_ (.A(_07100_),
    .B(_07219_),
    .C(_07321_),
    .Y(_07447_));
 sky130_fd_sc_hd__a311oi_1 _16587_ (.A1(_07100_),
    .A2(_07272_),
    .A3(_07398_),
    .B1(_07447_),
    .C1(_07319_),
    .Y(_07448_));
 sky130_fd_sc_hd__nand2_4 _16588_ (.A(net4013),
    .B(net4005),
    .Y(_07449_));
 sky130_fd_sc_hd__nor2_4 _16589_ (.A(_07082_),
    .B(_07449_),
    .Y(_07450_));
 sky130_fd_sc_hd__a2111oi_0 _16590_ (.A1(_12036_[0]),
    .A2(_07215_),
    .B1(_07328_),
    .C1(_07388_),
    .D1(_07450_),
    .Y(_07451_));
 sky130_fd_sc_hd__nor4_1 _16591_ (.A(_07426_),
    .B(_07446_),
    .C(_07448_),
    .D(_07451_),
    .Y(_07452_));
 sky130_fd_sc_hd__nor2_1 _16592_ (.A(net3698),
    .B(_07374_),
    .Y(_07453_));
 sky130_fd_sc_hd__a21oi_1 _16593_ (.A1(_12038_[0]),
    .A2(net3698),
    .B1(_07453_),
    .Y(_07454_));
 sky130_fd_sc_hd__a211oi_1 _16594_ (.A1(_12042_[0]),
    .A2(net3698),
    .B1(_07167_),
    .C1(_07339_),
    .Y(_07455_));
 sky130_fd_sc_hd__o221ai_1 _16595_ (.A1(net4004),
    .A2(_07454_),
    .B1(_07455_),
    .B2(_07314_),
    .C1(_07237_),
    .Y(_07456_));
 sky130_fd_sc_hd__nor2_4 _16596_ (.A(_07082_),
    .B(net4005),
    .Y(_07457_));
 sky130_fd_sc_hd__o21ai_0 _16597_ (.A1(net3698),
    .A2(_07457_),
    .B1(_07090_),
    .Y(_07458_));
 sky130_fd_sc_hd__a21oi_1 _16598_ (.A1(_07082_),
    .A2(_07215_),
    .B1(_07402_),
    .Y(_07459_));
 sky130_fd_sc_hd__o211ai_1 _16599_ (.A1(_12028_[0]),
    .A2(_07251_),
    .B1(_07458_),
    .C1(_07459_),
    .Y(_07460_));
 sky130_fd_sc_hd__nand2_2 _16600_ (.A(_12038_[0]),
    .B(net4005),
    .Y(_07461_));
 sky130_fd_sc_hd__nand3_1 _16601_ (.A(net4011),
    .B(_07186_),
    .C(_07461_),
    .Y(_07462_));
 sky130_fd_sc_hd__nand3_1 _16602_ (.A(_07100_),
    .B(_07449_),
    .C(_07296_),
    .Y(_07463_));
 sky130_fd_sc_hd__a21o_1 _16603_ (.A1(_07462_),
    .A2(_07463_),
    .B1(_07328_),
    .X(_07464_));
 sky130_fd_sc_hd__a31oi_1 _16604_ (.A1(_07456_),
    .A2(_07460_),
    .A3(_07464_),
    .B1(_07397_),
    .Y(_07465_));
 sky130_fd_sc_hd__nor3_1 _16605_ (.A(_07100_),
    .B(_07178_),
    .C(_07377_),
    .Y(_07466_));
 sky130_fd_sc_hd__o31ai_1 _16606_ (.A1(net4011),
    .A2(_07278_),
    .A3(_07261_),
    .B1(net4009),
    .Y(_07467_));
 sky130_fd_sc_hd__nor2_1 _16607_ (.A(_07457_),
    .B(_07261_),
    .Y(_07468_));
 sky130_fd_sc_hd__o21ai_2 _16608_ (.A1(net4011),
    .A2(_07468_),
    .B1(_07327_),
    .Y(_07469_));
 sky130_fd_sc_hd__o22ai_1 _16609_ (.A1(_07466_),
    .A2(_07467_),
    .B1(_07469_),
    .B2(net4009),
    .Y(_07470_));
 sky130_fd_sc_hd__nand2_4 _16610_ (.A(net3698),
    .B(net4005),
    .Y(_07471_));
 sky130_fd_sc_hd__nand2_1 _16611_ (.A(_07196_),
    .B(_07383_),
    .Y(_07472_));
 sky130_fd_sc_hd__nor2_2 _16612_ (.A(net4015),
    .B(_07090_),
    .Y(_07473_));
 sky130_fd_sc_hd__o21ai_0 _16613_ (.A1(_07167_),
    .A2(_07473_),
    .B1(net4004),
    .Y(_07474_));
 sky130_fd_sc_hd__o221ai_1 _16614_ (.A1(_07082_),
    .A2(_07471_),
    .B1(_07472_),
    .B2(net3634),
    .C1(_07474_),
    .Y(_07475_));
 sky130_fd_sc_hd__and2_4 _16615_ (.A(_12033_[0]),
    .B(net4005),
    .X(_07476_));
 sky130_fd_sc_hd__nand3b_1 _16616_ (.A_N(_07219_),
    .B(net4011),
    .C(_07272_),
    .Y(_07477_));
 sky130_fd_sc_hd__o311ai_0 _16617_ (.A1(net4011),
    .A2(_07317_),
    .A3(_07476_),
    .B1(_07477_),
    .C1(net4009),
    .Y(_07478_));
 sky130_fd_sc_hd__o211ai_1 _16618_ (.A1(net4009),
    .A2(_07475_),
    .B1(_07478_),
    .C1(_07372_),
    .Y(_07479_));
 sky130_fd_sc_hd__o21ai_0 _16619_ (.A1(_07373_),
    .A2(_07470_),
    .B1(_07479_),
    .Y(_07480_));
 sky130_fd_sc_hd__nor4_1 _16620_ (.A(_07441_),
    .B(_07452_),
    .C(_07465_),
    .D(_07480_),
    .Y(_00051_));
 sky130_fd_sc_hd__a21oi_1 _16621_ (.A1(_12038_[0]),
    .A2(net4005),
    .B1(net4010),
    .Y(_07481_));
 sky130_fd_sc_hd__a21oi_1 _16622_ (.A1(_12028_[0]),
    .A2(_07174_),
    .B1(_07306_),
    .Y(_07482_));
 sky130_fd_sc_hd__o21ai_0 _16623_ (.A1(_07167_),
    .A2(_07482_),
    .B1(net4006),
    .Y(_07483_));
 sky130_fd_sc_hd__o31ai_1 _16624_ (.A1(net4006),
    .A2(_07212_),
    .A3(_07481_),
    .B1(_07483_),
    .Y(_07484_));
 sky130_fd_sc_hd__a21oi_1 _16625_ (.A1(_07100_),
    .A2(net4007),
    .B1(_07090_),
    .Y(_07485_));
 sky130_fd_sc_hd__o211ai_1 _16626_ (.A1(net4014),
    .A2(_07485_),
    .B1(_07422_),
    .C1(_07174_),
    .Y(_07486_));
 sky130_fd_sc_hd__nand3_1 _16627_ (.A(_12028_[0]),
    .B(_07100_),
    .C(net4001),
    .Y(_07487_));
 sky130_fd_sc_hd__o311ai_0 _16628_ (.A1(net4014),
    .A2(_07100_),
    .A3(net4001),
    .B1(net4005),
    .C1(_07487_),
    .Y(_07488_));
 sky130_fd_sc_hd__nand2_4 _16629_ (.A(_07140_),
    .B(net4005),
    .Y(_07489_));
 sky130_fd_sc_hd__o22ai_1 _16630_ (.A1(_07100_),
    .A2(net4007),
    .B1(_07489_),
    .B2(_07090_),
    .Y(_07490_));
 sky130_fd_sc_hd__a221oi_1 _16631_ (.A1(_07486_),
    .A2(_07488_),
    .B1(_07490_),
    .B2(net4014),
    .C1(net4009),
    .Y(_07491_));
 sky130_fd_sc_hd__a21oi_1 _16632_ (.A1(net4009),
    .A2(_07484_),
    .B1(_07491_),
    .Y(_07492_));
 sky130_fd_sc_hd__nor2_2 _16633_ (.A(_12033_[0]),
    .B(net4005),
    .Y(_07493_));
 sky130_fd_sc_hd__nor3_1 _16634_ (.A(_07100_),
    .B(_07493_),
    .C(_07293_),
    .Y(_07494_));
 sky130_fd_sc_hd__a31oi_1 _16635_ (.A1(_07100_),
    .A2(_07186_),
    .A3(_07449_),
    .B1(_07494_),
    .Y(_07495_));
 sky130_fd_sc_hd__o221ai_1 _16636_ (.A1(_12042_[0]),
    .A2(_07200_),
    .B1(_07349_),
    .B2(_07100_),
    .C1(net4000),
    .Y(_07496_));
 sky130_fd_sc_hd__o211ai_1 _16637_ (.A1(net4000),
    .A2(_07495_),
    .B1(_07496_),
    .C1(net4008),
    .Y(_07497_));
 sky130_fd_sc_hd__o311ai_0 _16638_ (.A1(_07100_),
    .A2(_07476_),
    .A3(_07305_),
    .B1(_07318_),
    .C1(net4000),
    .Y(_07498_));
 sky130_fd_sc_hd__a21oi_1 _16639_ (.A1(net4009),
    .A2(_07295_),
    .B1(net4007),
    .Y(_07499_));
 sky130_fd_sc_hd__a21oi_1 _16640_ (.A1(_07498_),
    .A2(_07499_),
    .B1(_07397_),
    .Y(_07500_));
 sky130_fd_sc_hd__nor2_1 _16641_ (.A(_07100_),
    .B(_07493_),
    .Y(_07501_));
 sky130_fd_sc_hd__a21oi_1 _16642_ (.A1(_07296_),
    .A2(_07379_),
    .B1(net4011),
    .Y(_07502_));
 sky130_fd_sc_hd__a21oi_1 _16643_ (.A1(_07230_),
    .A2(_07501_),
    .B1(_07502_),
    .Y(_07503_));
 sky130_fd_sc_hd__o21ai_0 _16644_ (.A1(_12028_[0]),
    .A2(_07100_),
    .B1(_07383_),
    .Y(_07504_));
 sky130_fd_sc_hd__a21oi_1 _16645_ (.A1(net4005),
    .A2(_07504_),
    .B1(_07247_),
    .Y(_07505_));
 sky130_fd_sc_hd__a2111oi_0 _16646_ (.A1(net4003),
    .A2(_07503_),
    .B1(_07505_),
    .C1(net4009),
    .D1(_07371_),
    .Y(_07506_));
 sky130_fd_sc_hd__nand2_1 _16647_ (.A(_12033_[0]),
    .B(_07174_),
    .Y(_07507_));
 sky130_fd_sc_hd__a21oi_1 _16648_ (.A1(_07431_),
    .A2(_07507_),
    .B1(net4011),
    .Y(_07508_));
 sky130_fd_sc_hd__a21oi_1 _16649_ (.A1(_12038_[0]),
    .A2(net4011),
    .B1(_07508_),
    .Y(_07509_));
 sky130_fd_sc_hd__a21oi_1 _16650_ (.A1(_07186_),
    .A2(_07461_),
    .B1(net4011),
    .Y(_07510_));
 sky130_fd_sc_hd__a311oi_1 _16651_ (.A1(net4011),
    .A2(_07230_),
    .A3(_07405_),
    .B1(_07510_),
    .C1(net4003),
    .Y(_07511_));
 sky130_fd_sc_hd__a2111oi_0 _16652_ (.A1(net4003),
    .A2(_07509_),
    .B1(_07511_),
    .C1(net4000),
    .D1(_07371_),
    .Y(_07512_));
 sky130_fd_sc_hd__a211oi_1 _16653_ (.A1(_07497_),
    .A2(_07500_),
    .B1(_07506_),
    .C1(_07512_),
    .Y(_07513_));
 sky130_fd_sc_hd__a21oi_1 _16654_ (.A1(_07218_),
    .A2(_07249_),
    .B1(_07100_),
    .Y(_07514_));
 sky130_fd_sc_hd__nor2_1 _16655_ (.A(_12028_[0]),
    .B(_07200_),
    .Y(_07515_));
 sky130_fd_sc_hd__nor4_1 _16656_ (.A(net4009),
    .B(_07450_),
    .C(_07514_),
    .D(_07515_),
    .Y(_07516_));
 sky130_fd_sc_hd__nand3_1 _16657_ (.A(_12029_[0]),
    .B(_07100_),
    .C(net4005),
    .Y(_07517_));
 sky130_fd_sc_hd__nand2_1 _16658_ (.A(_12040_[0]),
    .B(net4004),
    .Y(_07518_));
 sky130_fd_sc_hd__a21oi_1 _16659_ (.A1(_07517_),
    .A2(_07518_),
    .B1(_07237_),
    .Y(_07519_));
 sky130_fd_sc_hd__o21ai_0 _16660_ (.A1(_07516_),
    .A2(_07519_),
    .B1(_07140_),
    .Y(_07520_));
 sky130_fd_sc_hd__a2111oi_0 _16661_ (.A1(net4015),
    .A2(_07199_),
    .B1(_07224_),
    .C1(_07328_),
    .D1(_07481_),
    .Y(_07521_));
 sky130_fd_sc_hd__o21ai_0 _16662_ (.A1(_07457_),
    .A2(_07343_),
    .B1(net4011),
    .Y(_07522_));
 sky130_fd_sc_hd__a31oi_1 _16663_ (.A1(_07235_),
    .A2(_07301_),
    .A3(_07522_),
    .B1(net4009),
    .Y(_07523_));
 sky130_fd_sc_hd__or3_1 _16664_ (.A(_07140_),
    .B(_07521_),
    .C(_07523_),
    .X(_07524_));
 sky130_fd_sc_hd__nand3_1 _16665_ (.A(_07394_),
    .B(_07520_),
    .C(_07524_),
    .Y(_07525_));
 sky130_fd_sc_hd__o211ai_1 _16666_ (.A1(_07426_),
    .A2(_07492_),
    .B1(_07513_),
    .C1(_07525_),
    .Y(_00052_));
 sky130_fd_sc_hd__o22ai_1 _16667_ (.A1(_12042_[0]),
    .A2(_07471_),
    .B1(_07365_),
    .B2(net4005),
    .Y(_07526_));
 sky130_fd_sc_hd__nand3_2 _16668_ (.A(_07100_),
    .B(_07405_),
    .C(_07418_),
    .Y(_07527_));
 sky130_fd_sc_hd__a31oi_1 _16669_ (.A1(net4011),
    .A2(_07186_),
    .A3(_07289_),
    .B1(net4009),
    .Y(_07528_));
 sky130_fd_sc_hd__a221oi_1 _16670_ (.A1(net4009),
    .A2(_07526_),
    .B1(_07527_),
    .B2(_07528_),
    .C1(_07140_),
    .Y(_07529_));
 sky130_fd_sc_hd__a221o_1 _16671_ (.A1(_07317_),
    .A2(_07324_),
    .B1(_07374_),
    .B2(_07199_),
    .C1(_07237_),
    .X(_07530_));
 sky130_fd_sc_hd__o211ai_1 _16672_ (.A1(net3698),
    .A2(_07301_),
    .B1(_07418_),
    .C1(_07237_),
    .Y(_07531_));
 sky130_fd_sc_hd__a21oi_1 _16673_ (.A1(_07530_),
    .A2(_07531_),
    .B1(net4001),
    .Y(_07532_));
 sky130_fd_sc_hd__o21ai_2 _16674_ (.A1(_07529_),
    .A2(_07532_),
    .B1(_07394_),
    .Y(_07533_));
 sky130_fd_sc_hd__a21oi_1 _16675_ (.A1(_07249_),
    .A2(_07431_),
    .B1(net4011),
    .Y(_07534_));
 sky130_fd_sc_hd__o21ai_0 _16676_ (.A1(_07082_),
    .A2(_07282_),
    .B1(_07350_),
    .Y(_07535_));
 sky130_fd_sc_hd__or3_4 _16677_ (.A(_12029_[0]),
    .B(_07100_),
    .C(net4004),
    .X(_07536_));
 sky130_fd_sc_hd__inv_1 _16678_ (.A(_07296_),
    .Y(_07537_));
 sky130_fd_sc_hd__o21ai_0 _16679_ (.A1(_07178_),
    .A2(_07537_),
    .B1(_07100_),
    .Y(_07538_));
 sky130_fd_sc_hd__a31oi_1 _16680_ (.A1(_07536_),
    .A2(_07362_),
    .A3(_07538_),
    .B1(_07371_),
    .Y(_07539_));
 sky130_fd_sc_hd__o211ai_1 _16681_ (.A1(_07082_),
    .A2(_07215_),
    .B1(_07301_),
    .C1(_07140_),
    .Y(_07540_));
 sky130_fd_sc_hd__a21oi_1 _16682_ (.A1(_07082_),
    .A2(net3620),
    .B1(_07457_),
    .Y(_07541_));
 sky130_fd_sc_hd__nand2_1 _16683_ (.A(_12036_[0]),
    .B(_07234_),
    .Y(_07542_));
 sky130_fd_sc_hd__o2111ai_1 _16684_ (.A1(net4013),
    .A2(_07541_),
    .B1(_07542_),
    .C1(_07327_),
    .D1(net4001),
    .Y(_07543_));
 sky130_fd_sc_hd__nand3_1 _16685_ (.A(net4009),
    .B(_07540_),
    .C(_07543_),
    .Y(_07544_));
 sky130_fd_sc_hd__o211ai_1 _16686_ (.A1(_07534_),
    .A2(_07535_),
    .B1(_07539_),
    .C1(_07544_),
    .Y(_07545_));
 sky130_fd_sc_hd__o21ai_2 _16687_ (.A1(net4013),
    .A2(_07471_),
    .B1(_07462_),
    .Y(_07546_));
 sky130_fd_sc_hd__nand3_1 _16688_ (.A(_07100_),
    .B(_07196_),
    .C(_07272_),
    .Y(_07547_));
 sky130_fd_sc_hd__a21oi_1 _16689_ (.A1(_07213_),
    .A2(_07547_),
    .B1(net4000),
    .Y(_07548_));
 sky130_fd_sc_hd__a21oi_1 _16690_ (.A1(net4000),
    .A2(_07546_),
    .B1(_07548_),
    .Y(_07549_));
 sky130_fd_sc_hd__a21oi_1 _16691_ (.A1(_12038_[0]),
    .A2(_07215_),
    .B1(_07476_),
    .Y(_07550_));
 sky130_fd_sc_hd__o311a_1 _16692_ (.A1(_07100_),
    .A2(_07224_),
    .A3(_07226_),
    .B1(_07550_),
    .C1(net4009),
    .X(_07551_));
 sky130_fd_sc_hd__nand2_1 _16693_ (.A(net4011),
    .B(_07507_),
    .Y(_07552_));
 sky130_fd_sc_hd__a21oi_1 _16694_ (.A1(_07230_),
    .A2(_07552_),
    .B1(net4009),
    .Y(_07553_));
 sky130_fd_sc_hd__o21ai_1 _16695_ (.A1(_07551_),
    .A2(_07553_),
    .B1(net4001),
    .Y(_07554_));
 sky130_fd_sc_hd__o2111ai_1 _16696_ (.A1(net4003),
    .A2(_07549_),
    .B1(_07554_),
    .C1(_07269_),
    .D1(_07266_),
    .Y(_07555_));
 sky130_fd_sc_hd__nor2_1 _16697_ (.A(net4011),
    .B(_07262_),
    .Y(_07556_));
 sky130_fd_sc_hd__a221oi_1 _16698_ (.A1(net4011),
    .A2(_07468_),
    .B1(_07556_),
    .B2(_07230_),
    .C1(_07140_),
    .Y(_07557_));
 sky130_fd_sc_hd__a211oi_1 _16699_ (.A1(_07090_),
    .A2(_07282_),
    .B1(_07224_),
    .C1(net4003),
    .Y(_07558_));
 sky130_fd_sc_hd__o21ai_0 _16700_ (.A1(_07557_),
    .A2(_07558_),
    .B1(net4009),
    .Y(_07559_));
 sky130_fd_sc_hd__nand3_1 _16701_ (.A(_07260_),
    .B(_07307_),
    .C(_07362_),
    .Y(_07560_));
 sky130_fd_sc_hd__a21oi_1 _16702_ (.A1(net4011),
    .A2(_07173_),
    .B1(_07319_),
    .Y(_07561_));
 sky130_fd_sc_hd__a21oi_2 _16703_ (.A1(_07527_),
    .A2(_07561_),
    .B1(_07397_),
    .Y(_07562_));
 sky130_fd_sc_hd__nand3_1 _16704_ (.A(_07559_),
    .B(_07560_),
    .C(_07562_),
    .Y(_07563_));
 sky130_fd_sc_hd__nand4_1 _16705_ (.A(_07533_),
    .B(_07545_),
    .C(_07555_),
    .D(_07563_),
    .Y(_00053_));
 sky130_fd_sc_hd__o31ai_1 _16706_ (.A1(net4010),
    .A2(_07435_),
    .A3(_07349_),
    .B1(_07536_),
    .Y(_07564_));
 sky130_fd_sc_hd__a21oi_1 _16707_ (.A1(_12038_[0]),
    .A2(_07100_),
    .B1(net4005),
    .Y(_07565_));
 sky130_fd_sc_hd__a221oi_1 _16708_ (.A1(_12046_[0]),
    .A2(net4005),
    .B1(_07414_),
    .B2(_07565_),
    .C1(net4001),
    .Y(_07566_));
 sky130_fd_sc_hd__a21oi_1 _16709_ (.A1(net4001),
    .A2(_07564_),
    .B1(_07566_),
    .Y(_07567_));
 sky130_fd_sc_hd__nor2_1 _16710_ (.A(_07237_),
    .B(_07567_),
    .Y(_07568_));
 sky130_fd_sc_hd__nand2_1 _16711_ (.A(_12033_[0]),
    .B(net4007),
    .Y(_07569_));
 sky130_fd_sc_hd__nand2_1 _16712_ (.A(_12038_[0]),
    .B(net4001),
    .Y(_07570_));
 sky130_fd_sc_hd__nand3_1 _16713_ (.A(_07234_),
    .B(_07569_),
    .C(_07570_),
    .Y(_07571_));
 sky130_fd_sc_hd__o21ai_0 _16714_ (.A1(_07312_),
    .A2(_07339_),
    .B1(_07571_),
    .Y(_07572_));
 sky130_fd_sc_hd__nand2_1 _16715_ (.A(net4015),
    .B(net4001),
    .Y(_07573_));
 sky130_fd_sc_hd__nand2_1 _16716_ (.A(_07140_),
    .B(_07473_),
    .Y(_07574_));
 sky130_fd_sc_hd__a21oi_1 _16717_ (.A1(_07573_),
    .A2(_07574_),
    .B1(_07251_),
    .Y(_07575_));
 sky130_fd_sc_hd__nor3_1 _16718_ (.A(net4009),
    .B(_07572_),
    .C(_07575_),
    .Y(_07576_));
 sky130_fd_sc_hd__o21ai_0 _16719_ (.A1(_07568_),
    .A2(_07576_),
    .B1(_07394_),
    .Y(_07577_));
 sky130_fd_sc_hd__a21oi_1 _16720_ (.A1(net4011),
    .A2(_07166_),
    .B1(_07278_),
    .Y(_07578_));
 sky130_fd_sc_hd__nor2_1 _16721_ (.A(_12042_[0]),
    .B(_07578_),
    .Y(_07579_));
 sky130_fd_sc_hd__nor3_1 _16722_ (.A(_07323_),
    .B(_07450_),
    .C(_07579_),
    .Y(_07580_));
 sky130_fd_sc_hd__o21ai_0 _16723_ (.A1(_07140_),
    .A2(_07391_),
    .B1(net4011),
    .Y(_07581_));
 sky130_fd_sc_hd__o221ai_1 _16724_ (.A1(_07422_),
    .A2(_07489_),
    .B1(_07581_),
    .B2(net4015),
    .C1(_07574_),
    .Y(_07582_));
 sky130_fd_sc_hd__o21ai_0 _16725_ (.A1(net4001),
    .A2(_07449_),
    .B1(_07573_),
    .Y(_07583_));
 sky130_fd_sc_hd__a21oi_1 _16726_ (.A1(_12029_[0]),
    .A2(_07140_),
    .B1(net4005),
    .Y(_07584_));
 sky130_fd_sc_hd__nor3_1 _16727_ (.A(_12038_[0]),
    .B(net4001),
    .C(net4004),
    .Y(_07585_));
 sky130_fd_sc_hd__o32ai_1 _16728_ (.A1(_07100_),
    .A2(_07584_),
    .A3(_07585_),
    .B1(_07339_),
    .B2(net4013),
    .Y(_07586_));
 sky130_fd_sc_hd__a211oi_1 _16729_ (.A1(_07100_),
    .A2(_07583_),
    .B1(_07586_),
    .C1(net4009),
    .Y(_07587_));
 sky130_fd_sc_hd__a211oi_1 _16730_ (.A1(net4009),
    .A2(_07582_),
    .B1(_07587_),
    .C1(_07397_),
    .Y(_07588_));
 sky130_fd_sc_hd__o21ai_0 _16731_ (.A1(_07328_),
    .A2(_07580_),
    .B1(_07588_),
    .Y(_07589_));
 sky130_fd_sc_hd__nor2_1 _16732_ (.A(_07262_),
    .B(_07293_),
    .Y(_07590_));
 sky130_fd_sc_hd__nor2_1 _16733_ (.A(net4010),
    .B(_07590_),
    .Y(_07591_));
 sky130_fd_sc_hd__a311oi_1 _16734_ (.A1(net4010),
    .A2(_07428_),
    .A3(_07296_),
    .B1(_07591_),
    .C1(net4009),
    .Y(_07592_));
 sky130_fd_sc_hd__o21ai_0 _16735_ (.A1(_07082_),
    .A2(_07100_),
    .B1(_07256_),
    .Y(_07593_));
 sky130_fd_sc_hd__o311ai_0 _16736_ (.A1(_12045_[0]),
    .A2(_12054_[0]),
    .A3(net4005),
    .B1(_07593_),
    .C1(net4009),
    .Y(_07594_));
 sky130_fd_sc_hd__nand2_1 _16737_ (.A(net4007),
    .B(_07594_),
    .Y(_07595_));
 sky130_fd_sc_hd__a21oi_1 _16738_ (.A1(_12038_[0]),
    .A2(net4005),
    .B1(_07349_),
    .Y(_07596_));
 sky130_fd_sc_hd__nor3_1 _16739_ (.A(net4010),
    .B(_07219_),
    .C(_07375_),
    .Y(_07597_));
 sky130_fd_sc_hd__a21oi_1 _16740_ (.A1(net4010),
    .A2(_07596_),
    .B1(_07597_),
    .Y(_07598_));
 sky130_fd_sc_hd__o21ai_0 _16741_ (.A1(_12028_[0]),
    .A2(net4005),
    .B1(_07461_),
    .Y(_07599_));
 sky130_fd_sc_hd__a221oi_1 _16742_ (.A1(_12030_[0]),
    .A2(_07234_),
    .B1(_07599_),
    .B2(net4010),
    .C1(_07328_),
    .Y(_07600_));
 sky130_fd_sc_hd__nor2_1 _16743_ (.A(_07426_),
    .B(_07600_),
    .Y(_07601_));
 sky130_fd_sc_hd__o221ai_1 _16744_ (.A1(_07592_),
    .A2(_07595_),
    .B1(_07598_),
    .B2(_07319_),
    .C1(_07601_),
    .Y(_07602_));
 sky130_fd_sc_hd__a21o_1 _16745_ (.A1(_07100_),
    .A2(_07231_),
    .B1(_07447_),
    .X(_07603_));
 sky130_fd_sc_hd__nand2_1 _16746_ (.A(net4009),
    .B(_07603_),
    .Y(_07604_));
 sky130_fd_sc_hd__a21oi_1 _16747_ (.A1(net4004),
    .A2(_07374_),
    .B1(net3698),
    .Y(_07605_));
 sky130_fd_sc_hd__a32oi_1 _16748_ (.A1(net3698),
    .A2(_07186_),
    .A3(_07218_),
    .B1(_07230_),
    .B2(_07605_),
    .Y(_07606_));
 sky130_fd_sc_hd__nand2_1 _16749_ (.A(_07237_),
    .B(_07606_),
    .Y(_07607_));
 sky130_fd_sc_hd__nor2_1 _16750_ (.A(_12047_[0]),
    .B(net4004),
    .Y(_07608_));
 sky130_fd_sc_hd__o21ai_0 _16751_ (.A1(net3634),
    .A2(net3698),
    .B1(net4004),
    .Y(_07609_));
 sky130_fd_sc_hd__a21oi_1 _16752_ (.A1(net3698),
    .A2(_07473_),
    .B1(_07609_),
    .Y(_07610_));
 sky130_fd_sc_hd__o21ai_0 _16753_ (.A1(_07608_),
    .A2(_07610_),
    .B1(net4009),
    .Y(_07611_));
 sky130_fd_sc_hd__a21oi_1 _16754_ (.A1(_07082_),
    .A2(_07422_),
    .B1(net4004),
    .Y(_07612_));
 sky130_fd_sc_hd__o21ai_0 _16755_ (.A1(_07201_),
    .A2(_07612_),
    .B1(_07237_),
    .Y(_07613_));
 sky130_fd_sc_hd__a21oi_1 _16756_ (.A1(_07611_),
    .A2(_07613_),
    .B1(_07373_),
    .Y(_07614_));
 sky130_fd_sc_hd__a31oi_2 _16757_ (.A1(_07372_),
    .A2(_07604_),
    .A3(_07607_),
    .B1(_07614_),
    .Y(_07615_));
 sky130_fd_sc_hd__nand4_1 _16758_ (.A(_07577_),
    .B(_07589_),
    .C(_07602_),
    .D(_07615_),
    .Y(_00054_));
 sky130_fd_sc_hd__a21oi_1 _16759_ (.A1(_07174_),
    .A2(_07167_),
    .B1(_07234_),
    .Y(_07616_));
 sky130_fd_sc_hd__a21oi_1 _16760_ (.A1(net4013),
    .A2(_07199_),
    .B1(_07278_),
    .Y(_07617_));
 sky130_fd_sc_hd__a21oi_1 _16761_ (.A1(_07200_),
    .A2(_07218_),
    .B1(_07082_),
    .Y(_07618_));
 sky130_fd_sc_hd__o21ai_0 _16762_ (.A1(_07224_),
    .A2(_07618_),
    .B1(_07140_),
    .Y(_07619_));
 sky130_fd_sc_hd__o221ai_1 _16763_ (.A1(net4015),
    .A2(_07616_),
    .B1(_07617_),
    .B2(_07140_),
    .C1(_07619_),
    .Y(_07620_));
 sky130_fd_sc_hd__nor3_1 _16764_ (.A(_07090_),
    .B(_07140_),
    .C(_07251_),
    .Y(_07621_));
 sky130_fd_sc_hd__a21oi_1 _16765_ (.A1(_07200_),
    .A2(_07489_),
    .B1(net4013),
    .Y(_07622_));
 sky130_fd_sc_hd__o21ai_0 _16766_ (.A1(_07621_),
    .A2(_07622_),
    .B1(_07082_),
    .Y(_07623_));
 sky130_fd_sc_hd__a221oi_1 _16767_ (.A1(_07100_),
    .A2(_07140_),
    .B1(_07326_),
    .B2(_12029_[0]),
    .C1(net4009),
    .Y(_07624_));
 sky130_fd_sc_hd__a221oi_1 _16768_ (.A1(net4009),
    .A2(_07620_),
    .B1(_07623_),
    .B2(_07624_),
    .C1(_07269_),
    .Y(_07625_));
 sky130_fd_sc_hd__a211o_1 _16769_ (.A1(_12038_[0]),
    .A2(net4010),
    .B1(net4005),
    .C1(_07194_),
    .X(_07626_));
 sky130_fd_sc_hd__o21ai_0 _16770_ (.A1(_12054_[0]),
    .A2(_07174_),
    .B1(_07626_),
    .Y(_07627_));
 sky130_fd_sc_hd__nor2_1 _16771_ (.A(_12040_[0]),
    .B(_07174_),
    .Y(_07628_));
 sky130_fd_sc_hd__a311oi_1 _16772_ (.A1(_12030_[0]),
    .A2(_07100_),
    .A3(_07174_),
    .B1(_07628_),
    .C1(_07237_),
    .Y(_07629_));
 sky130_fd_sc_hd__a211oi_1 _16773_ (.A1(_07237_),
    .A2(_07627_),
    .B1(_07629_),
    .C1(net4002),
    .Y(_07630_));
 sky130_fd_sc_hd__o21ai_0 _16774_ (.A1(_07317_),
    .A2(_07355_),
    .B1(_07350_),
    .Y(_07631_));
 sky130_fd_sc_hd__a21oi_1 _16775_ (.A1(_07100_),
    .A2(_07290_),
    .B1(_07631_),
    .Y(_07632_));
 sky130_fd_sc_hd__o21bai_1 _16776_ (.A1(_12033_[0]),
    .A2(_07100_),
    .B1_N(_07193_),
    .Y(_07633_));
 sky130_fd_sc_hd__a221oi_1 _16777_ (.A1(_07317_),
    .A2(_07422_),
    .B1(_07633_),
    .B2(net4005),
    .C1(_07328_),
    .Y(_07634_));
 sky130_fd_sc_hd__nor4_1 _16778_ (.A(_07115_),
    .B(_07630_),
    .C(_07632_),
    .D(_07634_),
    .Y(_07635_));
 sky130_fd_sc_hd__o32a_1 _16779_ (.A1(net4010),
    .A2(_07182_),
    .A3(_07173_),
    .B1(_07355_),
    .B2(_07305_),
    .X(_07636_));
 sky130_fd_sc_hd__o221ai_1 _16780_ (.A1(_12028_[0]),
    .A2(_07100_),
    .B1(_07212_),
    .B2(_07306_),
    .C1(_07237_),
    .Y(_07637_));
 sky130_fd_sc_hd__o21ai_0 _16781_ (.A1(_07237_),
    .A2(_07636_),
    .B1(_07637_),
    .Y(_07638_));
 sky130_fd_sc_hd__a21oi_1 _16782_ (.A1(net4010),
    .A2(_07375_),
    .B1(_07457_),
    .Y(_07639_));
 sky130_fd_sc_hd__o21ai_1 _16783_ (.A1(net4010),
    .A2(_07596_),
    .B1(_07639_),
    .Y(_07640_));
 sky130_fd_sc_hd__nor2_1 _16784_ (.A(net4009),
    .B(_07493_),
    .Y(_07641_));
 sky130_fd_sc_hd__a221oi_1 _16785_ (.A1(net4009),
    .A2(_07640_),
    .B1(_07641_),
    .B2(_07593_),
    .C1(net4007),
    .Y(_07642_));
 sky130_fd_sc_hd__a211o_1 _16786_ (.A1(net4007),
    .A2(_07638_),
    .B1(_07642_),
    .C1(_07426_),
    .X(_07643_));
 sky130_fd_sc_hd__nor2_1 _16787_ (.A(_12042_[0]),
    .B(_07251_),
    .Y(_07644_));
 sky130_fd_sc_hd__nor2_2 _16788_ (.A(_12029_[0]),
    .B(_07202_),
    .Y(_07645_));
 sky130_fd_sc_hd__nor4_1 _16789_ (.A(_07300_),
    .B(_07319_),
    .C(_07644_),
    .D(_07645_),
    .Y(_07646_));
 sky130_fd_sc_hd__a21oi_1 _16790_ (.A1(_07090_),
    .A2(_07234_),
    .B1(_07349_),
    .Y(_07647_));
 sky130_fd_sc_hd__nor2_1 _16791_ (.A(net4015),
    .B(_07647_),
    .Y(_07648_));
 sky130_fd_sc_hd__a2111oi_0 _16792_ (.A1(_12028_[0]),
    .A2(_07199_),
    .B1(_07300_),
    .C1(_07328_),
    .D1(_07648_),
    .Y(_07649_));
 sky130_fd_sc_hd__nor2_1 _16793_ (.A(_12038_[0]),
    .B(_07471_),
    .Y(_07650_));
 sky130_fd_sc_hd__a311oi_2 _16794_ (.A1(net4011),
    .A2(_07296_),
    .A3(_07379_),
    .B1(_07402_),
    .C1(_07650_),
    .Y(_07651_));
 sky130_fd_sc_hd__o21ai_0 _16795_ (.A1(_07284_),
    .A2(_07262_),
    .B1(_07100_),
    .Y(_07652_));
 sky130_fd_sc_hd__o211a_4 _16796_ (.A1(_07100_),
    .A2(_07392_),
    .B1(_07652_),
    .C1(_07362_),
    .X(_07653_));
 sky130_fd_sc_hd__o41ai_2 _16797_ (.A1(_07646_),
    .A2(_07649_),
    .A3(_07651_),
    .A4(_07653_),
    .B1(_07270_),
    .Y(_07654_));
 sky130_fd_sc_hd__o311ai_0 _16798_ (.A1(_07266_),
    .A2(_07625_),
    .A3(_07635_),
    .B1(_07643_),
    .C1(_07654_),
    .Y(_00055_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_826 ();
 sky130_fd_sc_hd__xnor2_1 _16801_ (.A(net4221),
    .B(\sa03_sr[0] ),
    .Y(_07657_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_824 ();
 sky130_fd_sc_hd__xnor2_2 _16804_ (.A(\sa21_sub[1] ),
    .B(\sa32_sub[1] ),
    .Y(_07660_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_821 ();
 sky130_fd_sc_hd__xnor3_1 _16808_ (.A(\sa10_sub[7] ),
    .B(net4211),
    .C(net4210),
    .X(_07664_));
 sky130_fd_sc_hd__xnor3_1 _16809_ (.A(_07657_),
    .B(_07660_),
    .C(_07664_),
    .X(_07665_));
 sky130_fd_sc_hd__mux2i_2 _16810_ (.A0(\text_in_r[25] ),
    .A1(_07665_),
    .S(_05879_),
    .Y(_07666_));
 sky130_fd_sc_hd__xor2_4 _16811_ (.A(net4130),
    .B(_07666_),
    .X(_07667_));
 sky130_fd_sc_hd__inv_16 _16812_ (.A(_07667_),
    .Y(_07668_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_819 ();
 sky130_fd_sc_hd__xnor2_2 _16815_ (.A(\sa03_sr[7] ),
    .B(\sa10_sub[7] ),
    .Y(_07670_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_818 ();
 sky130_fd_sc_hd__xnor3_1 _16817_ (.A(net4211),
    .B(net4195),
    .C(\sa32_sub[0] ),
    .X(_07672_));
 sky130_fd_sc_hd__xor2_1 _16818_ (.A(_07670_),
    .B(_07672_),
    .X(_07673_));
 sky130_fd_sc_hd__mux2i_2 _16819_ (.A0(\text_in_r[24] ),
    .A1(_07673_),
    .S(_05879_),
    .Y(_07674_));
 sky130_fd_sc_hd__xor2_4 _16820_ (.A(net4131),
    .B(_07674_),
    .X(_07675_));
 sky130_fd_sc_hd__clkinv_16 _16821_ (.A(_07675_),
    .Y(_07676_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_816 ();
 sky130_fd_sc_hd__xnor3_1 _16824_ (.A(\sa03_sr[1] ),
    .B(\sa10_sub[2] ),
    .C(net4193),
    .X(_07678_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_815 ();
 sky130_fd_sc_hd__xor2_1 _16826_ (.A(net4210),
    .B(\sa32_sub[2] ),
    .X(_07680_));
 sky130_fd_sc_hd__xnor2_1 _16827_ (.A(_07678_),
    .B(_07680_),
    .Y(_07681_));
 sky130_fd_sc_hd__mux2i_2 _16828_ (.A0(\text_in_r[26] ),
    .A1(_07681_),
    .S(net4116),
    .Y(_07682_));
 sky130_fd_sc_hd__xnor2_4 _16829_ (.A(\u0.tmp_w[26] ),
    .B(_07682_),
    .Y(_07683_));
 sky130_fd_sc_hd__clkinv_16 _16830_ (.A(_07683_),
    .Y(_07684_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_805 ();
 sky130_fd_sc_hd__xnor2_2 _16841_ (.A(\sa10_sub[7] ),
    .B(\sa21_sub[7] ),
    .Y(_07692_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_804 ();
 sky130_fd_sc_hd__xnor2_1 _16843_ (.A(\sa03_sr[6] ),
    .B(net4179),
    .Y(_07694_));
 sky130_fd_sc_hd__xnor2_1 _16844_ (.A(_07692_),
    .B(_07694_),
    .Y(_07695_));
 sky130_fd_sc_hd__xnor2_1 _16845_ (.A(\sa10_sub[6] ),
    .B(_07695_),
    .Y(_07696_));
 sky130_fd_sc_hd__mux2i_4 _16846_ (.A0(\text_in_r[31] ),
    .A1(_07696_),
    .S(net4116),
    .Y(_07697_));
 sky130_fd_sc_hd__xor2_4 _16847_ (.A(\u0.tmp_w[31] ),
    .B(_07697_),
    .X(_07698_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_803 ();
 sky130_fd_sc_hd__xnor2_2 _16849_ (.A(\sa10_sub[5] ),
    .B(\sa21_sub[5] ),
    .Y(_07700_));
 sky130_fd_sc_hd__xor2_1 _16850_ (.A(\sa10_sub[4] ),
    .B(\sa03_sr[4] ),
    .X(_07701_));
 sky130_fd_sc_hd__xnor3_1 _16851_ (.A(\sa32_sub[5] ),
    .B(_07700_),
    .C(_07701_),
    .X(_07702_));
 sky130_fd_sc_hd__mux2i_4 _16852_ (.A0(\text_in_r[29] ),
    .A1(_07702_),
    .S(net4116),
    .Y(_07703_));
 sky130_fd_sc_hd__xnor2_4 _16853_ (.A(net4128),
    .B(_07703_),
    .Y(_07704_));
 sky130_fd_sc_hd__xnor3_1 _16854_ (.A(\sa03_sr[5] ),
    .B(\sa10_sub[6] ),
    .C(\sa21_sub[6] ),
    .X(_07705_));
 sky130_fd_sc_hd__xor2_1 _16855_ (.A(\sa10_sub[5] ),
    .B(\sa32_sub[6] ),
    .X(_07706_));
 sky130_fd_sc_hd__xnor2_1 _16856_ (.A(_07705_),
    .B(_07706_),
    .Y(_07707_));
 sky130_fd_sc_hd__mux2i_4 _16857_ (.A0(\text_in_r[30] ),
    .A1(_07707_),
    .S(net4116),
    .Y(_07708_));
 sky130_fd_sc_hd__xor2_4 _16858_ (.A(\u0.tmp_w[30] ),
    .B(_07708_),
    .X(_07709_));
 sky130_fd_sc_hd__nand2_2 _16859_ (.A(net3994),
    .B(_07709_),
    .Y(_07710_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_802 ();
 sky130_fd_sc_hd__xnor3_1 _16861_ (.A(\sa03_sr[7] ),
    .B(\sa03_sr[3] ),
    .C(\sa21_sub[4] ),
    .X(_07712_));
 sky130_fd_sc_hd__xnor2_1 _16862_ (.A(\sa10_sub[7] ),
    .B(\sa10_sub[3] ),
    .Y(_07713_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_801 ();
 sky130_fd_sc_hd__xnor2_1 _16864_ (.A(\sa10_sub[4] ),
    .B(\sa32_sub[4] ),
    .Y(_07715_));
 sky130_fd_sc_hd__xnor3_1 _16865_ (.A(_07712_),
    .B(_07713_),
    .C(_07715_),
    .X(_07716_));
 sky130_fd_sc_hd__mux2i_4 _16866_ (.A0(\text_in_r[28] ),
    .A1(_07716_),
    .S(net4116),
    .Y(_07717_));
 sky130_fd_sc_hd__xnor2_4 _16867_ (.A(\u0.tmp_w[28] ),
    .B(_07717_),
    .Y(_07718_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_797 ();
 sky130_fd_sc_hd__xnor3_1 _16872_ (.A(\sa03_sr[7] ),
    .B(\sa03_sr[2] ),
    .C(\sa21_sub[3] ),
    .X(_07723_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_796 ();
 sky130_fd_sc_hd__xnor2_1 _16874_ (.A(net4209),
    .B(net4180),
    .Y(_07725_));
 sky130_fd_sc_hd__xnor3_1 _16875_ (.A(_07713_),
    .B(_07723_),
    .C(_07725_),
    .X(_07726_));
 sky130_fd_sc_hd__mux2i_2 _16876_ (.A0(\text_in_r[27] ),
    .A1(_07726_),
    .S(net4116),
    .Y(_07727_));
 sky130_fd_sc_hd__xor2_1 _16877_ (.A(\u0.tmp_w[27] ),
    .B(_07727_),
    .X(_07728_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_793 ();
 sky130_fd_sc_hd__nand2_8 _16881_ (.A(_07676_),
    .B(net3995),
    .Y(_07732_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_792 ();
 sky130_fd_sc_hd__nand2_1 _16883_ (.A(net3999),
    .B(net3998),
    .Y(_07734_));
 sky130_fd_sc_hd__nand2_1 _16884_ (.A(_07732_),
    .B(_07734_),
    .Y(_07735_));
 sky130_fd_sc_hd__xnor2_1 _16885_ (.A(net3989),
    .B(_07735_),
    .Y(_07736_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_789 ();
 sky130_fd_sc_hd__xnor2_1 _16889_ (.A(\u0.tmp_w[27] ),
    .B(_07727_),
    .Y(_07740_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_787 ();
 sky130_fd_sc_hd__nand2_1 _16892_ (.A(_12060_[0]),
    .B(net3986),
    .Y(_07743_));
 sky130_fd_sc_hd__nor2_4 _16893_ (.A(net3997),
    .B(net3986),
    .Y(_07744_));
 sky130_fd_sc_hd__nand2_2 _16894_ (.A(_07668_),
    .B(_07744_),
    .Y(_07745_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_784 ();
 sky130_fd_sc_hd__nor2_4 _16898_ (.A(_12061_[0]),
    .B(net3986),
    .Y(_07749_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_783 ();
 sky130_fd_sc_hd__a211oi_1 _16900_ (.A1(_12068_[0]),
    .A2(net3986),
    .B1(_07749_),
    .C1(net3694),
    .Y(_07751_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_781 ();
 sky130_fd_sc_hd__a311oi_1 _16903_ (.A1(net3694),
    .A2(_07743_),
    .A3(_07745_),
    .B1(_07751_),
    .C1(net3993),
    .Y(_07754_));
 sky130_fd_sc_hd__a21oi_1 _16904_ (.A1(net3993),
    .A2(_07736_),
    .B1(_07754_),
    .Y(_07755_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_779 ();
 sky130_fd_sc_hd__xnor2_4 _16907_ (.A(\u0.tmp_w[30] ),
    .B(_07708_),
    .Y(_07758_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_777 ();
 sky130_fd_sc_hd__nand2_8 _16910_ (.A(net3695),
    .B(net3988),
    .Y(_07761_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_775 ();
 sky130_fd_sc_hd__nand3_2 _16913_ (.A(_12061_[0]),
    .B(net3996),
    .C(net3986),
    .Y(_07764_));
 sky130_fd_sc_hd__nand2_1 _16914_ (.A(_07761_),
    .B(_07764_),
    .Y(_07765_));
 sky130_fd_sc_hd__nand2_8 _16915_ (.A(net3999),
    .B(net3987),
    .Y(_07766_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_774 ();
 sky130_fd_sc_hd__nand2_4 _16917_ (.A(_12074_[0]),
    .B(net3986),
    .Y(_07768_));
 sky130_fd_sc_hd__a21oi_1 _16918_ (.A1(_07766_),
    .A2(_07768_),
    .B1(net3996),
    .Y(_07769_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_773 ();
 sky130_fd_sc_hd__o21ai_0 _16920_ (.A1(_07765_),
    .A2(_07769_),
    .B1(net3993),
    .Y(_07771_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_772 ();
 sky130_fd_sc_hd__nand2_8 _16922_ (.A(net3996),
    .B(net3986),
    .Y(_07773_));
 sky130_fd_sc_hd__nand2_2 _16923_ (.A(net3998),
    .B(net3691),
    .Y(_07774_));
 sky130_fd_sc_hd__nor2_4 _16924_ (.A(_07668_),
    .B(net3990),
    .Y(_07775_));
 sky130_fd_sc_hd__xor2_4 _16925_ (.A(net4129),
    .B(_07717_),
    .X(_07776_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_770 ();
 sky130_fd_sc_hd__o221ai_1 _16928_ (.A1(_12065_[0]),
    .A2(_07773_),
    .B1(_07774_),
    .B2(_07775_),
    .C1(_07776_),
    .Y(_07779_));
 sky130_fd_sc_hd__nand4_1 _16929_ (.A(_07704_),
    .B(_07758_),
    .C(_07771_),
    .D(_07779_),
    .Y(_07780_));
 sky130_fd_sc_hd__nand2_8 _16930_ (.A(net3693),
    .B(net3989),
    .Y(_07781_));
 sky130_fd_sc_hd__nor2_4 _16931_ (.A(_07683_),
    .B(net3987),
    .Y(_07782_));
 sky130_fd_sc_hd__nor2_4 _16932_ (.A(_07684_),
    .B(net3986),
    .Y(_07783_));
 sky130_fd_sc_hd__nor2_4 _16933_ (.A(_07782_),
    .B(_07783_),
    .Y(_07784_));
 sky130_fd_sc_hd__o221a_1 _16934_ (.A1(_12068_[0]),
    .A2(_07781_),
    .B1(_07784_),
    .B2(_12060_[0]),
    .C1(_07764_),
    .X(_07785_));
 sky130_fd_sc_hd__nor2_2 _16935_ (.A(_12061_[0]),
    .B(net3995),
    .Y(_07786_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_769 ();
 sky130_fd_sc_hd__nor2_4 _16937_ (.A(net3696),
    .B(net3995),
    .Y(_07788_));
 sky130_fd_sc_hd__nand2_4 _16938_ (.A(_12061_[0]),
    .B(net3988),
    .Y(_07789_));
 sky130_fd_sc_hd__o2bb2ai_1 _16939_ (.A1_N(_07766_),
    .A2_N(_07786_),
    .B1(_07788_),
    .B2(_07789_),
    .Y(_07790_));
 sky130_fd_sc_hd__xor2_4 _16940_ (.A(net4128),
    .B(_07703_),
    .X(_07791_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_767 ();
 sky130_fd_sc_hd__nand2_4 _16943_ (.A(net3983),
    .B(_07709_),
    .Y(_07794_));
 sky130_fd_sc_hd__a21oi_1 _16944_ (.A1(net3993),
    .A2(_07790_),
    .B1(_07794_),
    .Y(_07795_));
 sky130_fd_sc_hd__o21ai_0 _16945_ (.A1(net3993),
    .A2(_07785_),
    .B1(_07795_),
    .Y(_07796_));
 sky130_fd_sc_hd__o211ai_1 _16946_ (.A1(_07710_),
    .A2(_07755_),
    .B1(_07780_),
    .C1(_07796_),
    .Y(_07797_));
 sky130_fd_sc_hd__nand2_8 _16947_ (.A(_07758_),
    .B(_07698_),
    .Y(_07798_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_765 ();
 sky130_fd_sc_hd__o21ai_0 _16950_ (.A1(net3990),
    .A2(_07732_),
    .B1(_07781_),
    .Y(_07801_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_764 ();
 sky130_fd_sc_hd__nand2_4 _16952_ (.A(net3996),
    .B(net3990),
    .Y(_07803_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_763 ();
 sky130_fd_sc_hd__o21ai_0 _16954_ (.A1(_12062_[0]),
    .A2(_07803_),
    .B1(_07776_),
    .Y(_07805_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_762 ();
 sky130_fd_sc_hd__nor3_4 _16956_ (.A(_07676_),
    .B(net3995),
    .C(net3989),
    .Y(_07807_));
 sky130_fd_sc_hd__a211oi_1 _16957_ (.A1(_07668_),
    .A2(_07801_),
    .B1(_07805_),
    .C1(_07807_),
    .Y(_07808_));
 sky130_fd_sc_hd__nand2_4 _16958_ (.A(_07668_),
    .B(net3987),
    .Y(_07809_));
 sky130_fd_sc_hd__nor2_2 _16959_ (.A(_07668_),
    .B(net3986),
    .Y(_07810_));
 sky130_fd_sc_hd__o21ai_0 _16960_ (.A1(_07774_),
    .A2(_07810_),
    .B1(net3993),
    .Y(_07811_));
 sky130_fd_sc_hd__a31oi_1 _16961_ (.A1(net3996),
    .A2(_07768_),
    .A3(_07809_),
    .B1(_07811_),
    .Y(_07812_));
 sky130_fd_sc_hd__nor4_1 _16962_ (.A(_07704_),
    .B(_07798_),
    .C(_07808_),
    .D(_07812_),
    .Y(_07813_));
 sky130_fd_sc_hd__nand2_4 _16963_ (.A(_12061_[0]),
    .B(net3693),
    .Y(_07814_));
 sky130_fd_sc_hd__nand2_2 _16964_ (.A(net3989),
    .B(_07814_),
    .Y(_07815_));
 sky130_fd_sc_hd__o21ai_2 _16965_ (.A1(_12081_[0]),
    .A2(net3989),
    .B1(_07815_),
    .Y(_07816_));
 sky130_fd_sc_hd__nor2_2 _16966_ (.A(_12065_[0]),
    .B(net3996),
    .Y(_07817_));
 sky130_fd_sc_hd__nor3_2 _16967_ (.A(net3999),
    .B(_07676_),
    .C(net3693),
    .Y(_07818_));
 sky130_fd_sc_hd__nor2_2 _16968_ (.A(_07817_),
    .B(_07818_),
    .Y(_07819_));
 sky130_fd_sc_hd__a21oi_2 _16969_ (.A1(net3989),
    .A2(_07819_),
    .B1(net3993),
    .Y(_07820_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_761 ();
 sky130_fd_sc_hd__nor2_1 _16971_ (.A(_12060_[0]),
    .B(_07684_),
    .Y(_07822_));
 sky130_fd_sc_hd__nand2_8 _16972_ (.A(_07676_),
    .B(net3986),
    .Y(_07823_));
 sky130_fd_sc_hd__nand2_2 _16973_ (.A(_12062_[0]),
    .B(net3988),
    .Y(_07824_));
 sky130_fd_sc_hd__nand2_2 _16974_ (.A(_07823_),
    .B(_07824_),
    .Y(_07825_));
 sky130_fd_sc_hd__a22oi_1 _16975_ (.A1(net3986),
    .A2(_07822_),
    .B1(_07825_),
    .B2(net3694),
    .Y(_07826_));
 sky130_fd_sc_hd__a221oi_1 _16976_ (.A1(net3993),
    .A2(_07816_),
    .B1(_07820_),
    .B2(_07826_),
    .C1(_07794_),
    .Y(_07827_));
 sky130_fd_sc_hd__nand2_1 _16977_ (.A(_07704_),
    .B(_07758_),
    .Y(_07828_));
 sky130_fd_sc_hd__nor2_2 _16978_ (.A(_12065_[0]),
    .B(net3987),
    .Y(_07829_));
 sky130_fd_sc_hd__o21ai_2 _16979_ (.A1(_12062_[0]),
    .A2(net3986),
    .B1(net3996),
    .Y(_07830_));
 sky130_fd_sc_hd__nor2_1 _16980_ (.A(_07829_),
    .B(_07830_),
    .Y(_07831_));
 sky130_fd_sc_hd__a21oi_2 _16981_ (.A1(_12060_[0]),
    .A2(net3990),
    .B1(_07683_),
    .Y(_07832_));
 sky130_fd_sc_hd__nor2_2 _16982_ (.A(_07684_),
    .B(_07718_),
    .Y(_07833_));
 sky130_fd_sc_hd__nand3_2 _16983_ (.A(_07823_),
    .B(_07766_),
    .C(_07833_),
    .Y(_07834_));
 sky130_fd_sc_hd__nand2_2 _16984_ (.A(net3692),
    .B(_07776_),
    .Y(_07835_));
 sky130_fd_sc_hd__nor2_4 _16985_ (.A(_12068_[0]),
    .B(net3989),
    .Y(_07836_));
 sky130_fd_sc_hd__or3_4 _16986_ (.A(_07835_),
    .B(_07836_),
    .C(_07749_),
    .X(_07837_));
 sky130_fd_sc_hd__o311ai_0 _16987_ (.A1(_07776_),
    .A2(_07831_),
    .A3(_07832_),
    .B1(_07834_),
    .C1(_07837_),
    .Y(_07838_));
 sky130_fd_sc_hd__nand2_2 _16988_ (.A(net3990),
    .B(_07817_),
    .Y(_07839_));
 sky130_fd_sc_hd__nor2_4 _16989_ (.A(_07704_),
    .B(_07776_),
    .Y(_07840_));
 sky130_fd_sc_hd__nor2_4 _16990_ (.A(_12061_[0]),
    .B(net3989),
    .Y(_07841_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_760 ();
 sky130_fd_sc_hd__nor2_1 _16992_ (.A(_12070_[0]),
    .B(net3986),
    .Y(_07843_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_759 ();
 sky130_fd_sc_hd__o21ai_0 _16994_ (.A1(_07841_),
    .A2(_07843_),
    .B1(net3995),
    .Y(_07845_));
 sky130_fd_sc_hd__a41oi_1 _16995_ (.A1(_07758_),
    .A2(_07839_),
    .A3(_07840_),
    .A4(_07845_),
    .B1(_07698_),
    .Y(_07846_));
 sky130_fd_sc_hd__nor2_4 _16996_ (.A(net3999),
    .B(net3997),
    .Y(_07847_));
 sky130_fd_sc_hd__nor2_1 _16997_ (.A(net3990),
    .B(_07847_),
    .Y(_07848_));
 sky130_fd_sc_hd__nor2_4 _16998_ (.A(_12065_[0]),
    .B(net3986),
    .Y(_07849_));
 sky130_fd_sc_hd__nand3_1 _16999_ (.A(_07791_),
    .B(_07758_),
    .C(_07776_),
    .Y(_07850_));
 sky130_fd_sc_hd__nor3_1 _17000_ (.A(_07849_),
    .B(_07850_),
    .C(_07807_),
    .Y(_07851_));
 sky130_fd_sc_hd__o21ai_0 _17001_ (.A1(net3691),
    .A2(_07848_),
    .B1(_07851_),
    .Y(_07852_));
 sky130_fd_sc_hd__o211ai_1 _17002_ (.A1(_07828_),
    .A2(_07838_),
    .B1(_07846_),
    .C1(_07852_),
    .Y(_07853_));
 sky130_fd_sc_hd__o21ai_0 _17003_ (.A1(_12068_[0]),
    .A2(_07781_),
    .B1(net3993),
    .Y(_07854_));
 sky130_fd_sc_hd__nand2_4 _17004_ (.A(_12062_[0]),
    .B(net3986),
    .Y(_07855_));
 sky130_fd_sc_hd__nor2_4 _17005_ (.A(net3999),
    .B(_07676_),
    .Y(_07856_));
 sky130_fd_sc_hd__o22ai_2 _17006_ (.A1(_07684_),
    .A2(_07855_),
    .B1(_07803_),
    .B2(_07856_),
    .Y(_07857_));
 sky130_fd_sc_hd__nor2_1 _17007_ (.A(_07854_),
    .B(_07857_),
    .Y(_07858_));
 sky130_fd_sc_hd__nor2_2 _17008_ (.A(_12062_[0]),
    .B(net3986),
    .Y(_07859_));
 sky130_fd_sc_hd__nor3_4 _17009_ (.A(net3999),
    .B(_07676_),
    .C(net3987),
    .Y(_07860_));
 sky130_fd_sc_hd__nor3_1 _17010_ (.A(net3691),
    .B(_07859_),
    .C(_07860_),
    .Y(_07861_));
 sky130_fd_sc_hd__a211oi_1 _17011_ (.A1(_12070_[0]),
    .A2(_07782_),
    .B1(_07861_),
    .C1(net3993),
    .Y(_07862_));
 sky130_fd_sc_hd__nor3_1 _17012_ (.A(_07858_),
    .B(_07862_),
    .C(_07710_),
    .Y(_07863_));
 sky130_fd_sc_hd__nor3_1 _17013_ (.A(_07827_),
    .B(_07853_),
    .C(_07863_),
    .Y(_07864_));
 sky130_fd_sc_hd__a211oi_2 _17014_ (.A1(_07698_),
    .A2(_07797_),
    .B1(_07813_),
    .C1(_07864_),
    .Y(_00056_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_758 ();
 sky130_fd_sc_hd__nand2_1 _17016_ (.A(_12074_[0]),
    .B(net3996),
    .Y(_07866_));
 sky130_fd_sc_hd__nand2_1 _17017_ (.A(_07814_),
    .B(_07866_),
    .Y(_07867_));
 sky130_fd_sc_hd__nand2_1 _17018_ (.A(net3986),
    .B(_07867_),
    .Y(_07868_));
 sky130_fd_sc_hd__nand2_1 _17019_ (.A(_07820_),
    .B(_07868_),
    .Y(_07869_));
 sky130_fd_sc_hd__xnor2_4 _17020_ (.A(\u0.tmp_w[31] ),
    .B(_07697_),
    .Y(_07870_));
 sky130_fd_sc_hd__nand2_8 _17021_ (.A(_07709_),
    .B(_07870_),
    .Y(_07871_));
 sky130_fd_sc_hd__nor2_2 _17022_ (.A(net3994),
    .B(_07871_),
    .Y(_07872_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_756 ();
 sky130_fd_sc_hd__o21ai_0 _17025_ (.A1(_07667_),
    .A2(_07784_),
    .B1(_07839_),
    .Y(_07874_));
 sky130_fd_sc_hd__nand2_1 _17026_ (.A(_07718_),
    .B(_07874_),
    .Y(_07875_));
 sky130_fd_sc_hd__nand2b_4 _17027_ (.A_N(_12061_[0]),
    .B(net3986),
    .Y(_07876_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_755 ();
 sky130_fd_sc_hd__nand2_2 _17029_ (.A(_12065_[0]),
    .B(net3987),
    .Y(_07878_));
 sky130_fd_sc_hd__nand3_1 _17030_ (.A(net3996),
    .B(_07876_),
    .C(_07878_),
    .Y(_07879_));
 sky130_fd_sc_hd__o21ai_0 _17031_ (.A1(_07683_),
    .A2(_07848_),
    .B1(_07879_),
    .Y(_07880_));
 sky130_fd_sc_hd__nand2_8 _17032_ (.A(_07758_),
    .B(_07870_),
    .Y(_07881_));
 sky130_fd_sc_hd__o22ai_1 _17033_ (.A1(net3695),
    .A2(_07773_),
    .B1(_07781_),
    .B2(_12061_[0]),
    .Y(_07882_));
 sky130_fd_sc_hd__nand2_4 _17034_ (.A(_07668_),
    .B(net3986),
    .Y(_07883_));
 sky130_fd_sc_hd__a21oi_1 _17035_ (.A1(_07803_),
    .A2(_07883_),
    .B1(net3998),
    .Y(_07884_));
 sky130_fd_sc_hd__nor3_1 _17036_ (.A(_07704_),
    .B(_07882_),
    .C(_07884_),
    .Y(_07885_));
 sky130_fd_sc_hd__a2111oi_0 _17037_ (.A1(_07704_),
    .A2(_07880_),
    .B1(_07881_),
    .C1(net3993),
    .D1(_07885_),
    .Y(_07886_));
 sky130_fd_sc_hd__nand2_2 _17038_ (.A(net3997),
    .B(net3995),
    .Y(_07887_));
 sky130_fd_sc_hd__nor2_4 _17039_ (.A(net3999),
    .B(net3988),
    .Y(_07888_));
 sky130_fd_sc_hd__nand2_4 _17040_ (.A(net3695),
    .B(_07684_),
    .Y(_07889_));
 sky130_fd_sc_hd__nand2_1 _17041_ (.A(_12060_[0]),
    .B(net3692),
    .Y(_07890_));
 sky130_fd_sc_hd__a21oi_1 _17042_ (.A1(_07887_),
    .A2(_07890_),
    .B1(net3986),
    .Y(_07891_));
 sky130_fd_sc_hd__a311o_1 _17043_ (.A1(_07887_),
    .A2(_07888_),
    .A3(_07889_),
    .B1(_07891_),
    .C1(net3985),
    .X(_07892_));
 sky130_fd_sc_hd__nor2_4 _17044_ (.A(net3997),
    .B(_07684_),
    .Y(_07893_));
 sky130_fd_sc_hd__a221oi_2 _17045_ (.A1(_12068_[0]),
    .A2(net3693),
    .B1(_07893_),
    .B2(_07668_),
    .C1(net3986),
    .Y(_07894_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_754 ();
 sky130_fd_sc_hd__a21oi_1 _17047_ (.A1(_07776_),
    .A2(_07894_),
    .B1(net3983),
    .Y(_07896_));
 sky130_fd_sc_hd__o21ai_0 _17048_ (.A1(_12084_[0]),
    .A2(net3989),
    .B1(_07776_),
    .Y(_07897_));
 sky130_fd_sc_hd__nand2_8 _17049_ (.A(_07709_),
    .B(_07698_),
    .Y(_07898_));
 sky130_fd_sc_hd__o21bai_1 _17050_ (.A1(_07894_),
    .A2(_07897_),
    .B1_N(_07898_),
    .Y(_07899_));
 sky130_fd_sc_hd__nor2_4 _17051_ (.A(net3999),
    .B(net3986),
    .Y(_07900_));
 sky130_fd_sc_hd__o21ai_2 _17052_ (.A1(_07900_),
    .A2(_07775_),
    .B1(net3694),
    .Y(_07901_));
 sky130_fd_sc_hd__o21ai_0 _17053_ (.A1(_07829_),
    .A2(_07744_),
    .B1(net3995),
    .Y(_07902_));
 sky130_fd_sc_hd__a21boi_0 _17054_ (.A1(_07901_),
    .A2(_07902_),
    .B1_N(_07840_),
    .Y(_07903_));
 sky130_fd_sc_hd__a211oi_1 _17055_ (.A1(_07892_),
    .A2(_07896_),
    .B1(_07899_),
    .C1(_07903_),
    .Y(_07904_));
 sky130_fd_sc_hd__a311oi_1 _17056_ (.A1(_07869_),
    .A2(_07872_),
    .A3(_07875_),
    .B1(_07886_),
    .C1(_07904_),
    .Y(_07905_));
 sky130_fd_sc_hd__nor2_1 _17057_ (.A(_07709_),
    .B(_07870_),
    .Y(_07906_));
 sky130_fd_sc_hd__a21oi_1 _17058_ (.A1(_07876_),
    .A2(_07745_),
    .B1(net3693),
    .Y(_07907_));
 sky130_fd_sc_hd__nor2_4 _17059_ (.A(net3995),
    .B(net3986),
    .Y(_07908_));
 sky130_fd_sc_hd__nand2_2 _17060_ (.A(net3998),
    .B(_07908_),
    .Y(_07909_));
 sky130_fd_sc_hd__nand2_1 _17061_ (.A(net3983),
    .B(_07909_),
    .Y(_07910_));
 sky130_fd_sc_hd__nor2_1 _17062_ (.A(_12060_[0]),
    .B(net3986),
    .Y(_07911_));
 sky130_fd_sc_hd__o311ai_0 _17063_ (.A1(net3995),
    .A2(_07888_),
    .A3(_07911_),
    .B1(_07902_),
    .C1(net3994),
    .Y(_07912_));
 sky130_fd_sc_hd__o21ai_0 _17064_ (.A1(_07907_),
    .A2(_07910_),
    .B1(_07912_),
    .Y(_07913_));
 sky130_fd_sc_hd__nand3_1 _17065_ (.A(net3985),
    .B(_07906_),
    .C(_07913_),
    .Y(_07914_));
 sky130_fd_sc_hd__a21oi_1 _17066_ (.A1(_12060_[0]),
    .A2(net3986),
    .B1(_07830_),
    .Y(_07915_));
 sky130_fd_sc_hd__nand2_2 _17067_ (.A(_12061_[0]),
    .B(net3986),
    .Y(_07916_));
 sky130_fd_sc_hd__a21oi_1 _17068_ (.A1(_07761_),
    .A2(_07916_),
    .B1(net3995),
    .Y(_07917_));
 sky130_fd_sc_hd__nor2_4 _17069_ (.A(net3984),
    .B(net3985),
    .Y(_07918_));
 sky130_fd_sc_hd__o211ai_1 _17070_ (.A1(_07915_),
    .A2(_07917_),
    .B1(_07918_),
    .C1(_07906_),
    .Y(_07919_));
 sky130_fd_sc_hd__nand2_4 _17071_ (.A(_07704_),
    .B(_07718_),
    .Y(_07920_));
 sky130_fd_sc_hd__o21ai_0 _17072_ (.A1(net3986),
    .A2(_07847_),
    .B1(_07883_),
    .Y(_07921_));
 sky130_fd_sc_hd__a22oi_1 _17073_ (.A1(_12074_[0]),
    .A2(_07782_),
    .B1(_07921_),
    .B2(_07683_),
    .Y(_07922_));
 sky130_fd_sc_hd__nand2_1 _17074_ (.A(net3992),
    .B(net3988),
    .Y(_07923_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_753 ();
 sky130_fd_sc_hd__a21oi_1 _17076_ (.A1(_12061_[0]),
    .A2(_07718_),
    .B1(net3988),
    .Y(_07925_));
 sky130_fd_sc_hd__a21oi_1 _17077_ (.A1(_07718_),
    .A2(_07849_),
    .B1(_07925_),
    .Y(_07926_));
 sky130_fd_sc_hd__nand2_1 _17078_ (.A(_07718_),
    .B(net3986),
    .Y(_07927_));
 sky130_fd_sc_hd__o22ai_1 _17079_ (.A1(_07718_),
    .A2(_07766_),
    .B1(_07927_),
    .B2(net3995),
    .Y(_07928_));
 sky130_fd_sc_hd__a2bb2oi_1 _17080_ (.A1_N(_07684_),
    .A2_N(_07926_),
    .B1(_07928_),
    .B2(net3997),
    .Y(_07929_));
 sky130_fd_sc_hd__o21ai_0 _17081_ (.A1(_07807_),
    .A2(_07833_),
    .B1(_07668_),
    .Y(_07930_));
 sky130_fd_sc_hd__nor2_2 _17082_ (.A(_07791_),
    .B(_07871_),
    .Y(_07931_));
 sky130_fd_sc_hd__o2111ai_2 _17083_ (.A1(_07923_),
    .A2(_07889_),
    .B1(_07929_),
    .C1(_07930_),
    .D1(_07931_),
    .Y(_07932_));
 sky130_fd_sc_hd__a21oi_1 _17084_ (.A1(_12060_[0]),
    .A2(net3988),
    .B1(net3692),
    .Y(_07933_));
 sky130_fd_sc_hd__nand2_1 _17085_ (.A(_07916_),
    .B(_07933_),
    .Y(_07934_));
 sky130_fd_sc_hd__and2_4 _17086_ (.A(_12065_[0]),
    .B(net3986),
    .X(_07935_));
 sky130_fd_sc_hd__o21ai_0 _17087_ (.A1(_07744_),
    .A2(_07935_),
    .B1(net3693),
    .Y(_07936_));
 sky130_fd_sc_hd__a21oi_1 _17088_ (.A1(_07934_),
    .A2(_07936_),
    .B1(_07881_),
    .Y(_07937_));
 sky130_fd_sc_hd__and2_4 _17089_ (.A(_12074_[0]),
    .B(net3988),
    .X(_07938_));
 sky130_fd_sc_hd__o21ai_2 _17090_ (.A1(net3999),
    .A2(net3997),
    .B1(net3986),
    .Y(_07939_));
 sky130_fd_sc_hd__nand3_2 _17091_ (.A(net3692),
    .B(_07824_),
    .C(_07939_),
    .Y(_07940_));
 sky130_fd_sc_hd__o311a_1 _17092_ (.A1(net3693),
    .A2(_07841_),
    .A3(_07938_),
    .B1(_07940_),
    .C1(_07906_),
    .X(_07941_));
 sky130_fd_sc_hd__o21ai_0 _17093_ (.A1(_07937_),
    .A2(_07941_),
    .B1(_07840_),
    .Y(_07942_));
 sky130_fd_sc_hd__o311a_1 _17094_ (.A1(_07881_),
    .A2(_07920_),
    .A3(_07922_),
    .B1(_07932_),
    .C1(_07942_),
    .X(_07943_));
 sky130_fd_sc_hd__nand4_1 _17095_ (.A(_07905_),
    .B(_07914_),
    .C(_07919_),
    .D(_07943_),
    .Y(_00057_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_752 ();
 sky130_fd_sc_hd__nand2_1 _17097_ (.A(_07668_),
    .B(net3996),
    .Y(_07945_));
 sky130_fd_sc_hd__nor2_1 _17098_ (.A(_12084_[0]),
    .B(net3986),
    .Y(_07946_));
 sky130_fd_sc_hd__nand2_8 _17099_ (.A(net3984),
    .B(net3985),
    .Y(_07947_));
 sky130_fd_sc_hd__a311o_1 _17100_ (.A1(net3986),
    .A2(_07734_),
    .A3(_07945_),
    .B1(_07946_),
    .C1(_07947_),
    .X(_07948_));
 sky130_fd_sc_hd__nor2_4 _17101_ (.A(_07791_),
    .B(_07718_),
    .Y(_07949_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_751 ();
 sky130_fd_sc_hd__nor3_1 _17103_ (.A(net3989),
    .B(_07818_),
    .C(_07786_),
    .Y(_07951_));
 sky130_fd_sc_hd__a21oi_1 _17104_ (.A1(_12081_[0]),
    .A2(net3989),
    .B1(_07951_),
    .Y(_07952_));
 sky130_fd_sc_hd__a21oi_1 _17105_ (.A1(_07949_),
    .A2(_07952_),
    .B1(_07881_),
    .Y(_07953_));
 sky130_fd_sc_hd__o21ai_0 _17106_ (.A1(_07900_),
    .A2(_07788_),
    .B1(_12061_[0]),
    .Y(_07954_));
 sky130_fd_sc_hd__nor2_2 _17107_ (.A(net3999),
    .B(net3693),
    .Y(_07955_));
 sky130_fd_sc_hd__a22oi_1 _17108_ (.A1(_07732_),
    .A2(_07775_),
    .B1(_07955_),
    .B2(_07823_),
    .Y(_07956_));
 sky130_fd_sc_hd__nand3_1 _17109_ (.A(net3994),
    .B(_07954_),
    .C(_07956_),
    .Y(_07957_));
 sky130_fd_sc_hd__a21oi_1 _17110_ (.A1(_12060_[0]),
    .A2(net3989),
    .B1(_07841_),
    .Y(_07958_));
 sky130_fd_sc_hd__o31a_1 _17111_ (.A1(net3694),
    .A2(_07836_),
    .A3(_07900_),
    .B1(net3983),
    .X(_07959_));
 sky130_fd_sc_hd__o21ai_0 _17112_ (.A1(net3995),
    .A2(_07958_),
    .B1(_07959_),
    .Y(_07960_));
 sky130_fd_sc_hd__nand3_1 _17113_ (.A(net3991),
    .B(_07957_),
    .C(_07960_),
    .Y(_07961_));
 sky130_fd_sc_hd__nand3_1 _17114_ (.A(_07948_),
    .B(_07953_),
    .C(_07961_),
    .Y(_07962_));
 sky130_fd_sc_hd__nand2_2 _17115_ (.A(net3696),
    .B(net3997),
    .Y(_07963_));
 sky130_fd_sc_hd__nand2_1 _17116_ (.A(_12079_[0]),
    .B(net3986),
    .Y(_07964_));
 sky130_fd_sc_hd__o21ai_0 _17117_ (.A1(_07963_),
    .A2(_07781_),
    .B1(_07964_),
    .Y(_07965_));
 sky130_fd_sc_hd__nand2_2 _17118_ (.A(_07888_),
    .B(_07889_),
    .Y(_07966_));
 sky130_fd_sc_hd__o211ai_1 _17119_ (.A1(_12088_[0]),
    .A2(net3986),
    .B1(_07966_),
    .C1(net3992),
    .Y(_07967_));
 sky130_fd_sc_hd__o21ai_1 _17120_ (.A1(net3992),
    .A2(_07965_),
    .B1(_07967_),
    .Y(_07968_));
 sky130_fd_sc_hd__nor2_4 _17121_ (.A(_12062_[0]),
    .B(_12065_[0]),
    .Y(_07969_));
 sky130_fd_sc_hd__nand2_1 _17122_ (.A(net3996),
    .B(_07969_),
    .Y(_07970_));
 sky130_fd_sc_hd__nand2_2 _17123_ (.A(net3693),
    .B(_07847_),
    .Y(_07971_));
 sky130_fd_sc_hd__a311oi_1 _17124_ (.A1(net3986),
    .A2(_07970_),
    .A3(_07971_),
    .B1(_07894_),
    .C1(_07776_),
    .Y(_07972_));
 sky130_fd_sc_hd__a221oi_1 _17125_ (.A1(_12065_[0]),
    .A2(_07782_),
    .B1(_07958_),
    .B2(net3995),
    .C1(net3991),
    .Y(_07973_));
 sky130_fd_sc_hd__nor4_1 _17126_ (.A(net3983),
    .B(_07871_),
    .C(_07972_),
    .D(_07973_),
    .Y(_07974_));
 sky130_fd_sc_hd__a21oi_1 _17127_ (.A1(_07872_),
    .A2(_07968_),
    .B1(_07974_),
    .Y(_07975_));
 sky130_fd_sc_hd__nand2_4 _17128_ (.A(net3998),
    .B(net3989),
    .Y(_07976_));
 sky130_fd_sc_hd__nand2_4 _17129_ (.A(_12070_[0]),
    .B(net3989),
    .Y(_07977_));
 sky130_fd_sc_hd__a21oi_1 _17130_ (.A1(_07876_),
    .A2(_07977_),
    .B1(net3995),
    .Y(_07978_));
 sky130_fd_sc_hd__a31oi_1 _17131_ (.A1(net3995),
    .A2(_07876_),
    .A3(_07976_),
    .B1(_07978_),
    .Y(_07979_));
 sky130_fd_sc_hd__o21ai_2 _17132_ (.A1(_12074_[0]),
    .A2(net3986),
    .B1(net3692),
    .Y(_07980_));
 sky130_fd_sc_hd__nor2_1 _17133_ (.A(_07888_),
    .B(_07980_),
    .Y(_07981_));
 sky130_fd_sc_hd__nand2_2 _17134_ (.A(_12070_[0]),
    .B(net3986),
    .Y(_07982_));
 sky130_fd_sc_hd__a21oi_1 _17135_ (.A1(_07761_),
    .A2(_07982_),
    .B1(net3693),
    .Y(_07983_));
 sky130_fd_sc_hd__o21ai_0 _17136_ (.A1(_07981_),
    .A2(_07983_),
    .B1(net3991),
    .Y(_07984_));
 sky130_fd_sc_hd__o21ai_0 _17137_ (.A1(net3991),
    .A2(_07979_),
    .B1(_07984_),
    .Y(_07985_));
 sky130_fd_sc_hd__nand3_1 _17138_ (.A(net3996),
    .B(_07823_),
    .C(_07977_),
    .Y(_07986_));
 sky130_fd_sc_hd__o311ai_0 _17139_ (.A1(net3996),
    .A2(_07935_),
    .A3(_07938_),
    .B1(_07986_),
    .C1(net3993),
    .Y(_07987_));
 sky130_fd_sc_hd__a31oi_1 _17140_ (.A1(net3996),
    .A2(_07883_),
    .A3(_07977_),
    .B1(_07817_),
    .Y(_07988_));
 sky130_fd_sc_hd__a21oi_1 _17141_ (.A1(_07776_),
    .A2(_07988_),
    .B1(_07704_),
    .Y(_07989_));
 sky130_fd_sc_hd__a21oi_1 _17142_ (.A1(_07987_),
    .A2(_07989_),
    .B1(_07798_),
    .Y(_07990_));
 sky130_fd_sc_hd__o21ai_0 _17143_ (.A1(net3983),
    .A2(_07985_),
    .B1(_07990_),
    .Y(_07991_));
 sky130_fd_sc_hd__o21ai_2 _17144_ (.A1(net3989),
    .A2(_07819_),
    .B1(_07776_),
    .Y(_07992_));
 sky130_fd_sc_hd__nor2_1 _17145_ (.A(_07815_),
    .B(_07955_),
    .Y(_07993_));
 sky130_fd_sc_hd__nor2_1 _17146_ (.A(_12065_[0]),
    .B(net3693),
    .Y(_07994_));
 sky130_fd_sc_hd__nor2_1 _17147_ (.A(_12074_[0]),
    .B(net3995),
    .Y(_07995_));
 sky130_fd_sc_hd__o21ai_0 _17148_ (.A1(_07994_),
    .A2(_07995_),
    .B1(net3989),
    .Y(_07996_));
 sky130_fd_sc_hd__a31oi_1 _17149_ (.A1(net3992),
    .A2(_07966_),
    .A3(_07996_),
    .B1(_07704_),
    .Y(_07997_));
 sky130_fd_sc_hd__o21ai_0 _17150_ (.A1(_07992_),
    .A2(_07993_),
    .B1(_07997_),
    .Y(_07998_));
 sky130_fd_sc_hd__a21oi_1 _17151_ (.A1(_07823_),
    .A2(_07789_),
    .B1(net3693),
    .Y(_07999_));
 sky130_fd_sc_hd__a21oi_1 _17152_ (.A1(_07766_),
    .A2(_07855_),
    .B1(net3995),
    .Y(_08000_));
 sky130_fd_sc_hd__o21ai_0 _17153_ (.A1(_07999_),
    .A2(_08000_),
    .B1(net3992),
    .Y(_08001_));
 sky130_fd_sc_hd__nand2_4 _17154_ (.A(net3997),
    .B(net3986),
    .Y(_08002_));
 sky130_fd_sc_hd__nor2_2 _17155_ (.A(net3999),
    .B(net3995),
    .Y(_08003_));
 sky130_fd_sc_hd__nand3_1 _17156_ (.A(_08002_),
    .B(_07761_),
    .C(_08003_),
    .Y(_08004_));
 sky130_fd_sc_hd__o211ai_1 _17157_ (.A1(_12074_[0]),
    .A2(_07773_),
    .B1(_08004_),
    .C1(net3985),
    .Y(_08005_));
 sky130_fd_sc_hd__a31oi_1 _17158_ (.A1(_07704_),
    .A2(_08001_),
    .A3(_08005_),
    .B1(_07898_),
    .Y(_08006_));
 sky130_fd_sc_hd__nand2_2 _17159_ (.A(_07998_),
    .B(_08006_),
    .Y(_08007_));
 sky130_fd_sc_hd__nand4_1 _17160_ (.A(_07962_),
    .B(_07975_),
    .C(_07991_),
    .D(_08007_),
    .Y(_00058_));
 sky130_fd_sc_hd__nor2_4 _17161_ (.A(net3693),
    .B(net3989),
    .Y(_08008_));
 sky130_fd_sc_hd__a22oi_1 _17162_ (.A1(_12068_[0]),
    .A2(_08008_),
    .B1(_07786_),
    .B2(net3989),
    .Y(_08009_));
 sky130_fd_sc_hd__nor2_1 _17163_ (.A(net3986),
    .B(_07732_),
    .Y(_08010_));
 sky130_fd_sc_hd__o21ai_0 _17164_ (.A1(_07807_),
    .A2(_08010_),
    .B1(net3696),
    .Y(_08011_));
 sky130_fd_sc_hd__a31oi_1 _17165_ (.A1(_07949_),
    .A2(_08009_),
    .A3(_08011_),
    .B1(_07881_),
    .Y(_08012_));
 sky130_fd_sc_hd__a21oi_1 _17166_ (.A1(_07963_),
    .A2(_07732_),
    .B1(_08008_),
    .Y(_08013_));
 sky130_fd_sc_hd__nand3_1 _17167_ (.A(net3693),
    .B(_07768_),
    .C(_07977_),
    .Y(_08014_));
 sky130_fd_sc_hd__o311ai_0 _17168_ (.A1(net3693),
    .A2(_07749_),
    .A3(_07888_),
    .B1(_08014_),
    .C1(net3992),
    .Y(_08015_));
 sky130_fd_sc_hd__o21ai_0 _17169_ (.A1(net3992),
    .A2(_08013_),
    .B1(_08015_),
    .Y(_08016_));
 sky130_fd_sc_hd__nand3_2 _17170_ (.A(net3999),
    .B(net3997),
    .C(net3986),
    .Y(_08017_));
 sky130_fd_sc_hd__nand2_1 _17171_ (.A(_07918_),
    .B(_08017_),
    .Y(_08018_));
 sky130_fd_sc_hd__a211oi_1 _17172_ (.A1(_12068_[0]),
    .A2(_07908_),
    .B1(_07999_),
    .C1(_08018_),
    .Y(_08019_));
 sky130_fd_sc_hd__a21oi_1 _17173_ (.A1(_07791_),
    .A2(_08016_),
    .B1(_08019_),
    .Y(_08020_));
 sky130_fd_sc_hd__nor2_4 _17174_ (.A(_12061_[0]),
    .B(_07684_),
    .Y(_08021_));
 sky130_fd_sc_hd__nor2_1 _17175_ (.A(net3989),
    .B(_07866_),
    .Y(_08022_));
 sky130_fd_sc_hd__nor3_1 _17176_ (.A(net3996),
    .B(_07829_),
    .C(_07810_),
    .Y(_08023_));
 sky130_fd_sc_hd__a211oi_1 _17177_ (.A1(net3989),
    .A2(_08021_),
    .B1(_08022_),
    .C1(_08023_),
    .Y(_08024_));
 sky130_fd_sc_hd__o21ai_0 _17178_ (.A1(_07841_),
    .A2(_07810_),
    .B1(net3694),
    .Y(_08025_));
 sky130_fd_sc_hd__nand2_4 _17179_ (.A(net3997),
    .B(_07783_),
    .Y(_08026_));
 sky130_fd_sc_hd__a31oi_1 _17180_ (.A1(_07840_),
    .A2(_08025_),
    .A3(_08026_),
    .B1(_07871_),
    .Y(_08027_));
 sky130_fd_sc_hd__o31ai_1 _17181_ (.A1(net3983),
    .A2(net3993),
    .A3(_08024_),
    .B1(_08027_),
    .Y(_08028_));
 sky130_fd_sc_hd__a22oi_1 _17182_ (.A1(_07810_),
    .A2(_07732_),
    .B1(_08003_),
    .B2(_07976_),
    .Y(_08029_));
 sky130_fd_sc_hd__a21oi_1 _17183_ (.A1(_07764_),
    .A2(_08029_),
    .B1(_07947_),
    .Y(_08030_));
 sky130_fd_sc_hd__nand2_1 _17184_ (.A(_12068_[0]),
    .B(net3989),
    .Y(_08031_));
 sky130_fd_sc_hd__a21oi_1 _17185_ (.A1(_07743_),
    .A2(_08031_),
    .B1(net3694),
    .Y(_08032_));
 sky130_fd_sc_hd__a311oi_1 _17186_ (.A1(net3694),
    .A2(_07876_),
    .A3(_07761_),
    .B1(_07920_),
    .C1(_08032_),
    .Y(_08033_));
 sky130_fd_sc_hd__a21oi_1 _17187_ (.A1(_12070_[0]),
    .A2(_07784_),
    .B1(_08010_),
    .Y(_08034_));
 sky130_fd_sc_hd__nor2_1 _17188_ (.A(net3693),
    .B(_07749_),
    .Y(_08035_));
 sky130_fd_sc_hd__nand2_1 _17189_ (.A(net3986),
    .B(_07969_),
    .Y(_08036_));
 sky130_fd_sc_hd__a21oi_1 _17190_ (.A1(_07768_),
    .A2(_07761_),
    .B1(net3995),
    .Y(_08037_));
 sky130_fd_sc_hd__a211oi_1 _17191_ (.A1(_08035_),
    .A2(_08036_),
    .B1(_08037_),
    .C1(_07947_),
    .Y(_08038_));
 sky130_fd_sc_hd__o21ai_0 _17192_ (.A1(_07704_),
    .A2(_07766_),
    .B1(_07855_),
    .Y(_08039_));
 sky130_fd_sc_hd__nor3_1 _17193_ (.A(_12068_[0]),
    .B(net3994),
    .C(_07781_),
    .Y(_08040_));
 sky130_fd_sc_hd__nand3_1 _17194_ (.A(net3995),
    .B(_07704_),
    .C(net3989),
    .Y(_08041_));
 sky130_fd_sc_hd__nand3_1 _17195_ (.A(net3693),
    .B(_07791_),
    .C(net3986),
    .Y(_08042_));
 sky130_fd_sc_hd__a21oi_1 _17196_ (.A1(_08041_),
    .A2(_08042_),
    .B1(_12061_[0]),
    .Y(_08043_));
 sky130_fd_sc_hd__a2111oi_0 _17197_ (.A1(net3995),
    .A2(_08039_),
    .B1(_08040_),
    .C1(net3985),
    .D1(_08043_),
    .Y(_08044_));
 sky130_fd_sc_hd__a211oi_1 _17198_ (.A1(_07949_),
    .A2(_08034_),
    .B1(_08038_),
    .C1(_08044_),
    .Y(_08045_));
 sky130_fd_sc_hd__o32ai_1 _17199_ (.A1(_08028_),
    .A2(_08030_),
    .A3(_08033_),
    .B1(_08045_),
    .B2(_07898_),
    .Y(_08046_));
 sky130_fd_sc_hd__nor2_1 _17200_ (.A(_07791_),
    .B(_07823_),
    .Y(_08047_));
 sky130_fd_sc_hd__nand2_2 _17201_ (.A(_07791_),
    .B(net3988),
    .Y(_08048_));
 sky130_fd_sc_hd__nor2_4 _17202_ (.A(_12070_[0]),
    .B(net3988),
    .Y(_08049_));
 sky130_fd_sc_hd__nor2_1 _17203_ (.A(_07749_),
    .B(_08049_),
    .Y(_08050_));
 sky130_fd_sc_hd__o221ai_1 _17204_ (.A1(net3695),
    .A2(_08048_),
    .B1(_08050_),
    .B2(_07791_),
    .C1(net3995),
    .Y(_08051_));
 sky130_fd_sc_hd__o21ai_2 _17205_ (.A1(_07980_),
    .A2(_08047_),
    .B1(_08051_),
    .Y(_08052_));
 sky130_fd_sc_hd__o22ai_1 _17206_ (.A1(_12060_[0]),
    .A2(_07773_),
    .B1(_07781_),
    .B2(net3999),
    .Y(_08053_));
 sky130_fd_sc_hd__a21oi_1 _17207_ (.A1(net3996),
    .A2(_07766_),
    .B1(net3998),
    .Y(_08054_));
 sky130_fd_sc_hd__nor3_1 _17208_ (.A(net3983),
    .B(_08053_),
    .C(_08054_),
    .Y(_08055_));
 sky130_fd_sc_hd__nor2_2 _17209_ (.A(_12070_[0]),
    .B(net3996),
    .Y(_08056_));
 sky130_fd_sc_hd__a211oi_1 _17210_ (.A1(net3996),
    .A2(_07969_),
    .B1(_08056_),
    .C1(net3989),
    .Y(_08057_));
 sky130_fd_sc_hd__nor3_1 _17211_ (.A(_07704_),
    .B(_07894_),
    .C(_08057_),
    .Y(_08058_));
 sky130_fd_sc_hd__nor3_1 _17212_ (.A(net3993),
    .B(_08055_),
    .C(_08058_),
    .Y(_08059_));
 sky130_fd_sc_hd__a211oi_1 _17213_ (.A1(net3991),
    .A2(_08052_),
    .B1(_08059_),
    .C1(_07798_),
    .Y(_08060_));
 sky130_fd_sc_hd__a211oi_2 _17214_ (.A1(_08012_),
    .A2(_08020_),
    .B1(_08046_),
    .C1(_08060_),
    .Y(_00059_));
 sky130_fd_sc_hd__nand2_1 _17215_ (.A(net3995),
    .B(net3985),
    .Y(_08061_));
 sky130_fd_sc_hd__o22ai_1 _17216_ (.A1(net3985),
    .A2(_07890_),
    .B1(_08061_),
    .B2(net3999),
    .Y(_08062_));
 sky130_fd_sc_hd__a21oi_1 _17217_ (.A1(net3997),
    .A2(_07835_),
    .B1(net3999),
    .Y(_08063_));
 sky130_fd_sc_hd__nand2_1 _17218_ (.A(net3988),
    .B(_07732_),
    .Y(_08064_));
 sky130_fd_sc_hd__o22ai_1 _17219_ (.A1(net3988),
    .A2(_08062_),
    .B1(_08063_),
    .B2(_08064_),
    .Y(_08065_));
 sky130_fd_sc_hd__nand2_1 _17220_ (.A(net3995),
    .B(_07718_),
    .Y(_08066_));
 sky130_fd_sc_hd__o21ai_0 _17221_ (.A1(_07718_),
    .A2(_08002_),
    .B1(_08066_),
    .Y(_08067_));
 sky130_fd_sc_hd__a21oi_1 _17222_ (.A1(net3999),
    .A2(_08067_),
    .B1(net3994),
    .Y(_08068_));
 sky130_fd_sc_hd__a211oi_1 _17223_ (.A1(_07832_),
    .A2(_07883_),
    .B1(_07893_),
    .C1(_07718_),
    .Y(_08069_));
 sky130_fd_sc_hd__a311oi_1 _17224_ (.A1(_07718_),
    .A2(_07830_),
    .A3(_07982_),
    .B1(_08069_),
    .C1(net3983),
    .Y(_08070_));
 sky130_fd_sc_hd__a211oi_1 _17225_ (.A1(_08065_),
    .A2(_08068_),
    .B1(_08070_),
    .C1(_07881_),
    .Y(_08071_));
 sky130_fd_sc_hd__o21ai_1 _17226_ (.A1(_07822_),
    .A2(_08003_),
    .B1(net3986),
    .Y(_08072_));
 sky130_fd_sc_hd__o21ai_0 _17227_ (.A1(_07849_),
    .A2(_07860_),
    .B1(net3995),
    .Y(_08073_));
 sky130_fd_sc_hd__o31ai_1 _17228_ (.A1(net3995),
    .A2(_07888_),
    .A3(_07938_),
    .B1(_08073_),
    .Y(_08074_));
 sky130_fd_sc_hd__a221oi_2 _17229_ (.A1(_07820_),
    .A2(_08072_),
    .B1(_08074_),
    .B2(net3993),
    .C1(net3994),
    .Y(_08075_));
 sky130_fd_sc_hd__nor3_1 _17230_ (.A(net3989),
    .B(_07818_),
    .C(_08056_),
    .Y(_08076_));
 sky130_fd_sc_hd__a21oi_1 _17231_ (.A1(_07814_),
    .A2(_07866_),
    .B1(net3986),
    .Y(_08077_));
 sky130_fd_sc_hd__o21a_4 _17232_ (.A1(_08076_),
    .A2(_08077_),
    .B1(_07949_),
    .X(_08078_));
 sky130_fd_sc_hd__o21ai_0 _17233_ (.A1(_12070_[0]),
    .A2(net3691),
    .B1(_07918_),
    .Y(_08079_));
 sky130_fd_sc_hd__a31oi_1 _17234_ (.A1(net3691),
    .A2(_07878_),
    .A3(_07916_),
    .B1(_08079_),
    .Y(_08080_));
 sky130_fd_sc_hd__nor4_1 _17235_ (.A(_07871_),
    .B(_08075_),
    .C(_08078_),
    .D(_08080_),
    .Y(_08081_));
 sky130_fd_sc_hd__and4_1 _17236_ (.A(_07684_),
    .B(net3994),
    .C(_08002_),
    .D(_07789_),
    .X(_08082_));
 sky130_fd_sc_hd__a2111oi_0 _17237_ (.A1(net3986),
    .A2(_07847_),
    .B1(_07849_),
    .C1(_07684_),
    .D1(net3984),
    .Y(_08083_));
 sky130_fd_sc_hd__a21oi_1 _17238_ (.A1(_07980_),
    .A2(_08026_),
    .B1(net3994),
    .Y(_08084_));
 sky130_fd_sc_hd__o31ai_1 _17239_ (.A1(_08082_),
    .A2(_08083_),
    .A3(_08084_),
    .B1(net3985),
    .Y(_08085_));
 sky130_fd_sc_hd__o311ai_1 _17240_ (.A1(net3693),
    .A2(_07935_),
    .A3(_07911_),
    .B1(_07840_),
    .C1(_07901_),
    .Y(_08086_));
 sky130_fd_sc_hd__a21oi_1 _17241_ (.A1(_07918_),
    .A2(_07940_),
    .B1(_07798_),
    .Y(_08087_));
 sky130_fd_sc_hd__and3_1 _17242_ (.A(_08085_),
    .B(_08086_),
    .C(_08087_),
    .X(_08088_));
 sky130_fd_sc_hd__nand2_1 _17243_ (.A(_12072_[0]),
    .B(net3989),
    .Y(_08089_));
 sky130_fd_sc_hd__o21ai_2 _17244_ (.A1(net3989),
    .A2(_07814_),
    .B1(_08089_),
    .Y(_08090_));
 sky130_fd_sc_hd__o211ai_1 _17245_ (.A1(_12060_[0]),
    .A2(_07781_),
    .B1(_08017_),
    .C1(_07791_),
    .Y(_08091_));
 sky130_fd_sc_hd__a21oi_1 _17246_ (.A1(net3995),
    .A2(_07825_),
    .B1(_08091_),
    .Y(_08092_));
 sky130_fd_sc_hd__a211oi_2 _17247_ (.A1(net3994),
    .A2(_08090_),
    .B1(_08092_),
    .C1(net3992),
    .Y(_08093_));
 sky130_fd_sc_hd__nor2_1 _17248_ (.A(_07791_),
    .B(net3986),
    .Y(_08094_));
 sky130_fd_sc_hd__o21ai_0 _17249_ (.A1(_08094_),
    .A2(_08049_),
    .B1(_07684_),
    .Y(_08095_));
 sky130_fd_sc_hd__o21ai_2 _17250_ (.A1(_07856_),
    .A2(_07788_),
    .B1(net3989),
    .Y(_08096_));
 sky130_fd_sc_hd__nand2_1 _17251_ (.A(_07791_),
    .B(net3986),
    .Y(_08097_));
 sky130_fd_sc_hd__nor2_1 _17252_ (.A(_07732_),
    .B(_08097_),
    .Y(_08098_));
 sky130_fd_sc_hd__a31oi_1 _17253_ (.A1(net3999),
    .A2(net3994),
    .A3(_08008_),
    .B1(_08098_),
    .Y(_08099_));
 sky130_fd_sc_hd__nand4_1 _17254_ (.A(_07718_),
    .B(_08095_),
    .C(_08096_),
    .D(_08099_),
    .Y(_08100_));
 sky130_fd_sc_hd__nor3b_4 _17255_ (.A(_07898_),
    .B(_08093_),
    .C_N(_08100_),
    .Y(_08101_));
 sky130_fd_sc_hd__nor4_1 _17256_ (.A(_08071_),
    .B(_08081_),
    .C(_08088_),
    .D(_08101_),
    .Y(_00060_));
 sky130_fd_sc_hd__nor2_4 _17257_ (.A(net3992),
    .B(net3988),
    .Y(_08102_));
 sky130_fd_sc_hd__a21oi_1 _17258_ (.A1(net3992),
    .A2(_07773_),
    .B1(_08102_),
    .Y(_08103_));
 sky130_fd_sc_hd__nor2_1 _17259_ (.A(net3999),
    .B(_08103_),
    .Y(_08104_));
 sky130_fd_sc_hd__a211oi_1 _17260_ (.A1(net3999),
    .A2(_07923_),
    .B1(_08104_),
    .C1(net3997),
    .Y(_08105_));
 sky130_fd_sc_hd__nor2_1 _17261_ (.A(_07783_),
    .B(_08102_),
    .Y(_08106_));
 sky130_fd_sc_hd__nor2_1 _17262_ (.A(_07668_),
    .B(_08106_),
    .Y(_08107_));
 sky130_fd_sc_hd__nand2_1 _17263_ (.A(_12068_[0]),
    .B(_07782_),
    .Y(_08108_));
 sky130_fd_sc_hd__a21oi_1 _17264_ (.A1(_08026_),
    .A2(_08108_),
    .B1(net3985),
    .Y(_08109_));
 sky130_fd_sc_hd__nor2_1 _17265_ (.A(_07831_),
    .B(_07769_),
    .Y(_08110_));
 sky130_fd_sc_hd__a2111oi_0 _17266_ (.A1(_12070_[0]),
    .A2(_07908_),
    .B1(_07857_),
    .C1(_07935_),
    .D1(_07776_),
    .Y(_08111_));
 sky130_fd_sc_hd__a211o_1 _17267_ (.A1(_07776_),
    .A2(_08110_),
    .B1(_08111_),
    .C1(_07828_),
    .X(_08112_));
 sky130_fd_sc_hd__o41a_1 _17268_ (.A1(_07710_),
    .A2(_08105_),
    .A3(_08107_),
    .A4(_08109_),
    .B1(_08112_),
    .X(_08113_));
 sky130_fd_sc_hd__a21oi_1 _17269_ (.A1(net3995),
    .A2(_07878_),
    .B1(_07860_),
    .Y(_08114_));
 sky130_fd_sc_hd__nor2_1 _17270_ (.A(_07709_),
    .B(_08114_),
    .Y(_08115_));
 sky130_fd_sc_hd__a21oi_1 _17271_ (.A1(_07824_),
    .A2(_07916_),
    .B1(net3995),
    .Y(_08116_));
 sky130_fd_sc_hd__a211oi_1 _17272_ (.A1(net3999),
    .A2(_07783_),
    .B1(_08116_),
    .C1(_07758_),
    .Y(_08117_));
 sky130_fd_sc_hd__nor2_1 _17273_ (.A(_08115_),
    .B(_08117_),
    .Y(_08118_));
 sky130_fd_sc_hd__o22ai_1 _17274_ (.A1(net3988),
    .A2(_07889_),
    .B1(_08050_),
    .B2(net3692),
    .Y(_08119_));
 sky130_fd_sc_hd__nand2_1 _17275_ (.A(net3986),
    .B(_08021_),
    .Y(_08120_));
 sky130_fd_sc_hd__nor2_1 _17276_ (.A(_12060_[0]),
    .B(net3988),
    .Y(_08121_));
 sky130_fd_sc_hd__o21ai_0 _17277_ (.A1(_07938_),
    .A2(_08121_),
    .B1(net3692),
    .Y(_08122_));
 sky130_fd_sc_hd__a31o_1 _17278_ (.A1(_07709_),
    .A2(_08120_),
    .A3(_08122_),
    .B1(_07947_),
    .X(_08123_));
 sky130_fd_sc_hd__a21oi_1 _17279_ (.A1(_07758_),
    .A2(_08119_),
    .B1(_08123_),
    .Y(_08124_));
 sky130_fd_sc_hd__a211oi_1 _17280_ (.A1(_07840_),
    .A2(_08118_),
    .B1(_08124_),
    .C1(_07698_),
    .Y(_08125_));
 sky130_fd_sc_hd__a32oi_1 _17281_ (.A1(_07887_),
    .A2(_07900_),
    .A3(_07889_),
    .B1(_07969_),
    .B2(_08008_),
    .Y(_08126_));
 sky130_fd_sc_hd__nand3_1 _17282_ (.A(net3995),
    .B(_07876_),
    .C(_07789_),
    .Y(_08127_));
 sky130_fd_sc_hd__o21ai_2 _17283_ (.A1(_07836_),
    .A2(_07938_),
    .B1(net3692),
    .Y(_08128_));
 sky130_fd_sc_hd__o21ai_2 _17284_ (.A1(net3989),
    .A2(_07995_),
    .B1(_07704_),
    .Y(_08129_));
 sky130_fd_sc_hd__a21oi_2 _17285_ (.A1(_12065_[0]),
    .A2(_07908_),
    .B1(_08129_),
    .Y(_08130_));
 sky130_fd_sc_hd__a311oi_1 _17286_ (.A1(net3984),
    .A2(_08127_),
    .A3(_08128_),
    .B1(_08130_),
    .C1(net3985),
    .Y(_08131_));
 sky130_fd_sc_hd__a221oi_1 _17287_ (.A1(_12068_[0]),
    .A2(net3986),
    .B1(_07847_),
    .B2(_07783_),
    .C1(_07947_),
    .Y(_08132_));
 sky130_fd_sc_hd__a2111oi_0 _17288_ (.A1(_07949_),
    .A2(_08126_),
    .B1(_08131_),
    .C1(_07898_),
    .D1(_08132_),
    .Y(_08133_));
 sky130_fd_sc_hd__a31oi_1 _17289_ (.A1(net3997),
    .A2(net3994),
    .A3(_07809_),
    .B1(_07718_),
    .Y(_08134_));
 sky130_fd_sc_hd__a211oi_1 _17290_ (.A1(_07791_),
    .A2(_07888_),
    .B1(_08094_),
    .C1(net3997),
    .Y(_08135_));
 sky130_fd_sc_hd__a21oi_1 _17291_ (.A1(net3997),
    .A2(_08048_),
    .B1(_08135_),
    .Y(_08136_));
 sky130_fd_sc_hd__o211ai_1 _17292_ (.A1(_12065_[0]),
    .A2(_08048_),
    .B1(_08002_),
    .C1(_07684_),
    .Y(_08137_));
 sky130_fd_sc_hd__o21ai_1 _17293_ (.A1(_07684_),
    .A2(_08136_),
    .B1(_08137_),
    .Y(_08138_));
 sky130_fd_sc_hd__nand3_1 _17294_ (.A(net3995),
    .B(_07876_),
    .C(_07766_),
    .Y(_08139_));
 sky130_fd_sc_hd__o31ai_1 _17295_ (.A1(net3995),
    .A2(_07843_),
    .A3(_07860_),
    .B1(_08139_),
    .Y(_08140_));
 sky130_fd_sc_hd__o31ai_1 _17296_ (.A1(_07684_),
    .A2(net3986),
    .A3(_07847_),
    .B1(_08128_),
    .Y(_08141_));
 sky130_fd_sc_hd__a221o_1 _17297_ (.A1(_07918_),
    .A2(_08140_),
    .B1(_08141_),
    .B2(_07840_),
    .C1(_07798_),
    .X(_08142_));
 sky130_fd_sc_hd__a21oi_1 _17298_ (.A1(_08134_),
    .A2(_08138_),
    .B1(_08142_),
    .Y(_08143_));
 sky130_fd_sc_hd__a211oi_1 _17299_ (.A1(_08113_),
    .A2(_08125_),
    .B1(_08133_),
    .C1(_08143_),
    .Y(_00061_));
 sky130_fd_sc_hd__a21oi_1 _17300_ (.A1(net3999),
    .A2(net3995),
    .B1(_07939_),
    .Y(_08144_));
 sky130_fd_sc_hd__nor3_1 _17301_ (.A(_12077_[0]),
    .B(_12086_[0]),
    .C(net3986),
    .Y(_08145_));
 sky130_fd_sc_hd__nor3_1 _17302_ (.A(_07718_),
    .B(_08144_),
    .C(_08145_),
    .Y(_08146_));
 sky130_fd_sc_hd__o21ai_0 _17303_ (.A1(_12070_[0]),
    .A2(net3988),
    .B1(_07933_),
    .Y(_08147_));
 sky130_fd_sc_hd__a311oi_1 _17304_ (.A1(_12062_[0]),
    .A2(_07718_),
    .A3(_07782_),
    .B1(_07881_),
    .C1(net3983),
    .Y(_08148_));
 sky130_fd_sc_hd__o21ai_0 _17305_ (.A1(net3985),
    .A2(_08147_),
    .B1(_08148_),
    .Y(_08149_));
 sky130_fd_sc_hd__a21oi_1 _17306_ (.A1(_07789_),
    .A2(_08036_),
    .B1(net3995),
    .Y(_08150_));
 sky130_fd_sc_hd__a311oi_1 _17307_ (.A1(net3995),
    .A2(_07976_),
    .A3(_07982_),
    .B1(_08150_),
    .C1(net3985),
    .Y(_08151_));
 sky130_fd_sc_hd__nand2_2 _17308_ (.A(_12074_[0]),
    .B(net3989),
    .Y(_08152_));
 sky130_fd_sc_hd__a31o_4 _17309_ (.A1(net3996),
    .A2(_07855_),
    .A3(_08152_),
    .B1(net3993),
    .X(_08153_));
 sky130_fd_sc_hd__a31oi_1 _17310_ (.A1(net3694),
    .A2(_07939_),
    .A3(_07977_),
    .B1(_08153_),
    .Y(_08154_));
 sky130_fd_sc_hd__or4_1 _17311_ (.A(net3994),
    .B(_07881_),
    .C(_08151_),
    .D(_08154_),
    .X(_08155_));
 sky130_fd_sc_hd__a211oi_1 _17312_ (.A1(net3989),
    .A2(_07969_),
    .B1(_07860_),
    .C1(net3693),
    .Y(_08156_));
 sky130_fd_sc_hd__a311oi_1 _17313_ (.A1(net3693),
    .A2(_07823_),
    .A3(_07789_),
    .B1(_08156_),
    .C1(net3991),
    .Y(_08157_));
 sky130_fd_sc_hd__a21oi_1 _17314_ (.A1(_07668_),
    .A2(_07732_),
    .B1(net3990),
    .Y(_08158_));
 sky130_fd_sc_hd__nor2_1 _17315_ (.A(_07854_),
    .B(_08158_),
    .Y(_08159_));
 sky130_fd_sc_hd__o21ai_0 _17316_ (.A1(_08157_),
    .A2(_08159_),
    .B1(_07872_),
    .Y(_08160_));
 sky130_fd_sc_hd__o211ai_1 _17317_ (.A1(_08146_),
    .A2(_08149_),
    .B1(_08155_),
    .C1(_08160_),
    .Y(_08161_));
 sky130_fd_sc_hd__a31oi_1 _17318_ (.A1(net3999),
    .A2(net3997),
    .A3(net3995),
    .B1(_07744_),
    .Y(_08162_));
 sky130_fd_sc_hd__o211ai_1 _17319_ (.A1(_12074_[0]),
    .A2(_08162_),
    .B1(_08017_),
    .C1(_07889_),
    .Y(_08163_));
 sky130_fd_sc_hd__o21ai_0 _17320_ (.A1(_12074_[0]),
    .A2(_07803_),
    .B1(net3992),
    .Y(_08164_));
 sky130_fd_sc_hd__a21oi_1 _17321_ (.A1(net3695),
    .A2(_07684_),
    .B1(net3999),
    .Y(_08165_));
 sky130_fd_sc_hd__a221o_1 _17322_ (.A1(_07893_),
    .A2(_08102_),
    .B1(_08164_),
    .B2(_08165_),
    .C1(_07791_),
    .X(_08166_));
 sky130_fd_sc_hd__a21oi_1 _17323_ (.A1(net3992),
    .A2(_08163_),
    .B1(_08166_),
    .Y(_08167_));
 sky130_fd_sc_hd__nand2_1 _17324_ (.A(_07668_),
    .B(_07718_),
    .Y(_08168_));
 sky130_fd_sc_hd__nand2_1 _17325_ (.A(net3695),
    .B(net3985),
    .Y(_08169_));
 sky130_fd_sc_hd__a21oi_1 _17326_ (.A1(_08168_),
    .A2(_08169_),
    .B1(net3995),
    .Y(_08170_));
 sky130_fd_sc_hd__nor2_1 _17327_ (.A(_12070_[0]),
    .B(_08061_),
    .Y(_08171_));
 sky130_fd_sc_hd__o21ai_0 _17328_ (.A1(_07668_),
    .A2(net3995),
    .B1(net3997),
    .Y(_08172_));
 sky130_fd_sc_hd__a22oi_1 _17329_ (.A1(_12061_[0]),
    .A2(_07833_),
    .B1(_08172_),
    .B2(_07718_),
    .Y(_08173_));
 sky130_fd_sc_hd__o32ai_1 _17330_ (.A1(_08097_),
    .A2(_08170_),
    .A3(_08171_),
    .B1(_08048_),
    .B2(_08173_),
    .Y(_08174_));
 sky130_fd_sc_hd__nor3_1 _17331_ (.A(_07798_),
    .B(_08167_),
    .C(_08174_),
    .Y(_08175_));
 sky130_fd_sc_hd__a21oi_1 _17332_ (.A1(_12068_[0]),
    .A2(net3988),
    .B1(_08049_),
    .Y(_08176_));
 sky130_fd_sc_hd__o221ai_1 _17333_ (.A1(_07668_),
    .A2(_07773_),
    .B1(_08176_),
    .B2(net3995),
    .C1(net3992),
    .Y(_08177_));
 sky130_fd_sc_hd__a21oi_1 _17334_ (.A1(_07992_),
    .A2(_08177_),
    .B1(net3994),
    .Y(_08178_));
 sky130_fd_sc_hd__a2111oi_0 _17335_ (.A1(_12070_[0]),
    .A2(net3693),
    .B1(net3992),
    .C1(net3986),
    .D1(_07955_),
    .Y(_08179_));
 sky130_fd_sc_hd__a211oi_1 _17336_ (.A1(net3986),
    .A2(_08021_),
    .B1(_08037_),
    .C1(net3985),
    .Y(_08180_));
 sky130_fd_sc_hd__a2111oi_0 _17337_ (.A1(_12078_[0]),
    .A2(_08102_),
    .B1(_08179_),
    .C1(_08180_),
    .D1(_07791_),
    .Y(_08181_));
 sky130_fd_sc_hd__o21ai_1 _17338_ (.A1(_07859_),
    .A2(_07860_),
    .B1(net3694),
    .Y(_08182_));
 sky130_fd_sc_hd__o311ai_0 _17339_ (.A1(net3693),
    .A2(_07749_),
    .A3(_07888_),
    .B1(_08182_),
    .C1(net3985),
    .Y(_08183_));
 sky130_fd_sc_hd__a21oi_1 _17340_ (.A1(net3693),
    .A2(_07856_),
    .B1(_08021_),
    .Y(_08184_));
 sky130_fd_sc_hd__o211ai_1 _17341_ (.A1(net3986),
    .A2(_08184_),
    .B1(_07964_),
    .C1(net3992),
    .Y(_08185_));
 sky130_fd_sc_hd__nand3_1 _17342_ (.A(_07931_),
    .B(_08183_),
    .C(_08185_),
    .Y(_08186_));
 sky130_fd_sc_hd__o31ai_2 _17343_ (.A1(_07898_),
    .A2(_08178_),
    .A3(_08181_),
    .B1(_08186_),
    .Y(_08187_));
 sky130_fd_sc_hd__nor3_1 _17344_ (.A(_08161_),
    .B(_08175_),
    .C(_08187_),
    .Y(_00062_));
 sky130_fd_sc_hd__a21oi_1 _17345_ (.A1(_12068_[0]),
    .A2(net3986),
    .B1(net3995),
    .Y(_08188_));
 sky130_fd_sc_hd__nand2_1 _17346_ (.A(_07745_),
    .B(_08188_),
    .Y(_08189_));
 sky130_fd_sc_hd__a21oi_1 _17347_ (.A1(_07668_),
    .A2(_07774_),
    .B1(net3986),
    .Y(_08190_));
 sky130_fd_sc_hd__nor3_2 _17348_ (.A(_07920_),
    .B(_08057_),
    .C(_08190_),
    .Y(_08191_));
 sky130_fd_sc_hd__a31oi_1 _17349_ (.A1(_07934_),
    .A2(_07949_),
    .A3(_08189_),
    .B1(_08191_),
    .Y(_08192_));
 sky130_fd_sc_hd__nor3_1 _17350_ (.A(net3995),
    .B(_07859_),
    .C(_07888_),
    .Y(_08193_));
 sky130_fd_sc_hd__or3_4 _17351_ (.A(_07822_),
    .B(_07947_),
    .C(_08193_),
    .X(_08194_));
 sky130_fd_sc_hd__o21ai_0 _17352_ (.A1(_07849_),
    .A2(_08144_),
    .B1(_07840_),
    .Y(_08195_));
 sky130_fd_sc_hd__a31oi_2 _17353_ (.A1(_08192_),
    .A2(_08194_),
    .A3(_08195_),
    .B1(_07709_),
    .Y(_08196_));
 sky130_fd_sc_hd__nor2_1 _17354_ (.A(_12086_[0]),
    .B(net3988),
    .Y(_08197_));
 sky130_fd_sc_hd__a211oi_1 _17355_ (.A1(_12070_[0]),
    .A2(net3995),
    .B1(net3986),
    .C1(_07786_),
    .Y(_08198_));
 sky130_fd_sc_hd__a21oi_1 _17356_ (.A1(_07876_),
    .A2(_07809_),
    .B1(net3692),
    .Y(_08199_));
 sky130_fd_sc_hd__o21ai_0 _17357_ (.A1(_07917_),
    .A2(_08199_),
    .B1(_07840_),
    .Y(_08200_));
 sky130_fd_sc_hd__o31ai_1 _17358_ (.A1(_07947_),
    .A2(_08197_),
    .A3(_08198_),
    .B1(_08200_),
    .Y(_08201_));
 sky130_fd_sc_hd__o21ai_0 _17359_ (.A1(_07994_),
    .A2(_07788_),
    .B1(net3986),
    .Y(_08202_));
 sky130_fd_sc_hd__a21oi_1 _17360_ (.A1(_07732_),
    .A2(_07900_),
    .B1(_07920_),
    .Y(_08203_));
 sky130_fd_sc_hd__nand3_1 _17361_ (.A(_12062_[0]),
    .B(net3693),
    .C(net3989),
    .Y(_08204_));
 sky130_fd_sc_hd__o21ai_0 _17362_ (.A1(_12072_[0]),
    .A2(net3989),
    .B1(_08204_),
    .Y(_08205_));
 sky130_fd_sc_hd__a221o_4 _17363_ (.A1(_08202_),
    .A2(_08203_),
    .B1(_08205_),
    .B2(_07949_),
    .C1(_07758_),
    .X(_08206_));
 sky130_fd_sc_hd__o21ai_2 _17364_ (.A1(_08201_),
    .A2(_08206_),
    .B1(_07870_),
    .Y(_08207_));
 sky130_fd_sc_hd__o21ai_0 _17365_ (.A1(net3989),
    .A2(_07889_),
    .B1(_07976_),
    .Y(_08208_));
 sky130_fd_sc_hd__nand2_1 _17366_ (.A(_12060_[0]),
    .B(_08008_),
    .Y(_08209_));
 sky130_fd_sc_hd__nand4_1 _17367_ (.A(_07758_),
    .B(net3991),
    .C(_07909_),
    .D(_08209_),
    .Y(_08210_));
 sky130_fd_sc_hd__a21oi_1 _17368_ (.A1(net3696),
    .A2(_08208_),
    .B1(_08210_),
    .Y(_08211_));
 sky130_fd_sc_hd__nor3_1 _17369_ (.A(net3693),
    .B(_07888_),
    .C(_07938_),
    .Y(_08212_));
 sky130_fd_sc_hd__a2111oi_0 _17370_ (.A1(net3693),
    .A2(_08049_),
    .B1(_08212_),
    .C1(_07709_),
    .D1(net3991),
    .Y(_08213_));
 sky130_fd_sc_hd__nor2_1 _17371_ (.A(net3986),
    .B(_07963_),
    .Y(_08214_));
 sky130_fd_sc_hd__a21oi_1 _17372_ (.A1(_07823_),
    .A2(_07781_),
    .B1(net3696),
    .Y(_08215_));
 sky130_fd_sc_hd__o21ai_0 _17373_ (.A1(_08214_),
    .A2(_08215_),
    .B1(net3985),
    .Y(_08216_));
 sky130_fd_sc_hd__o21ai_0 _17374_ (.A1(net3695),
    .A2(_07773_),
    .B1(_07761_),
    .Y(_08217_));
 sky130_fd_sc_hd__nand2_1 _17375_ (.A(net3991),
    .B(_08217_),
    .Y(_08218_));
 sky130_fd_sc_hd__o21ai_0 _17376_ (.A1(_07782_),
    .A2(_08010_),
    .B1(net3696),
    .Y(_08219_));
 sky130_fd_sc_hd__a31oi_1 _17377_ (.A1(_08216_),
    .A2(_08218_),
    .A3(_08219_),
    .B1(_07758_),
    .Y(_08220_));
 sky130_fd_sc_hd__nor4_2 _17378_ (.A(net3983),
    .B(_08211_),
    .C(_08213_),
    .D(_08220_),
    .Y(_08221_));
 sky130_fd_sc_hd__o21ai_0 _17379_ (.A1(_07908_),
    .A2(_08102_),
    .B1(net3695),
    .Y(_08222_));
 sky130_fd_sc_hd__o21ai_0 _17380_ (.A1(_07887_),
    .A2(_07927_),
    .B1(_08222_),
    .Y(_08223_));
 sky130_fd_sc_hd__nand2_1 _17381_ (.A(_12061_[0]),
    .B(_07783_),
    .Y(_08224_));
 sky130_fd_sc_hd__nand2_1 _17382_ (.A(_07835_),
    .B(_08224_),
    .Y(_08225_));
 sky130_fd_sc_hd__a21oi_1 _17383_ (.A1(_07668_),
    .A2(_08223_),
    .B1(_08225_),
    .Y(_08226_));
 sky130_fd_sc_hd__o221ai_1 _17384_ (.A1(_12074_[0]),
    .A2(_07773_),
    .B1(_07784_),
    .B2(_12061_[0]),
    .C1(_07909_),
    .Y(_08227_));
 sky130_fd_sc_hd__nor2_1 _17385_ (.A(net3990),
    .B(_07732_),
    .Y(_08228_));
 sky130_fd_sc_hd__nor2_2 _17386_ (.A(_08152_),
    .B(_08056_),
    .Y(_08229_));
 sky130_fd_sc_hd__a21oi_1 _17387_ (.A1(_07883_),
    .A2(_07977_),
    .B1(net3996),
    .Y(_08230_));
 sky130_fd_sc_hd__o41ai_1 _17388_ (.A1(_07850_),
    .A2(_08228_),
    .A3(_08229_),
    .A4(_08230_),
    .B1(_07698_),
    .Y(_08231_));
 sky130_fd_sc_hd__a31oi_2 _17389_ (.A1(_07758_),
    .A2(_07840_),
    .A3(_08227_),
    .B1(_08231_),
    .Y(_08232_));
 sky130_fd_sc_hd__o21ai_2 _17390_ (.A1(_07794_),
    .A2(_08226_),
    .B1(_08232_),
    .Y(_08233_));
 sky130_fd_sc_hd__o22ai_4 _17391_ (.A1(_08196_),
    .A2(_08207_),
    .B1(_08221_),
    .B2(_08233_),
    .Y(_00063_));
 sky130_fd_sc_hd__xnor3_1 _17392_ (.A(\sa10_sr[7] ),
    .B(\sa00_sr[1] ),
    .C(net4207),
    .X(_08234_));
 sky130_fd_sc_hd__xnor3_1 _17393_ (.A(_05875_),
    .B(_05885_),
    .C(_08234_),
    .X(_08235_));
 sky130_fd_sc_hd__mux2i_2 _17394_ (.A0(\text_in_r[113] ),
    .A1(_08235_),
    .S(_05879_),
    .Y(_08236_));
 sky130_fd_sc_hd__xor2_4 _17395_ (.A(\u0.w[0][17] ),
    .B(_08236_),
    .X(_08237_));
 sky130_fd_sc_hd__clkinv_8 _17396_ (.A(_08237_),
    .Y(_08238_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_749 ();
 sky130_fd_sc_hd__xor2_1 _17399_ (.A(\sa00_sr[0] ),
    .B(\sa30_sr[0] ),
    .X(_08240_));
 sky130_fd_sc_hd__xnor3_1 _17400_ (.A(\sa20_sr[0] ),
    .B(_05970_),
    .C(_08240_),
    .X(_08241_));
 sky130_fd_sc_hd__mux2i_2 _17401_ (.A0(\text_in_r[112] ),
    .A1(_08241_),
    .S(_05879_),
    .Y(_08242_));
 sky130_fd_sc_hd__xor2_4 _17402_ (.A(\u0.w[0][16] ),
    .B(_08242_),
    .X(_08243_));
 sky130_fd_sc_hd__clkinv_16 _17403_ (.A(_08243_),
    .Y(_08244_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_747 ();
 sky130_fd_sc_hd__xnor3_1 _17406_ (.A(\sa20_sr[1] ),
    .B(\sa20_sr[2] ),
    .C(\sa00_sr[2] ),
    .X(_08246_));
 sky130_fd_sc_hd__xnor2_1 _17407_ (.A(_05895_),
    .B(_08246_),
    .Y(_08247_));
 sky130_fd_sc_hd__mux2i_2 _17408_ (.A0(\text_in_r[114] ),
    .A1(_08247_),
    .S(_05879_),
    .Y(_08248_));
 sky130_fd_sc_hd__xnor2_4 _17409_ (.A(\u0.w[0][18] ),
    .B(_08248_),
    .Y(_08249_));
 sky130_fd_sc_hd__clkinv_16 _17410_ (.A(_08249_),
    .Y(_08250_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_737 ();
 sky130_fd_sc_hd__nand2_2 _17421_ (.A(net4230),
    .B(\text_in_r[115] ),
    .Y(_08258_));
 sky130_fd_sc_hd__nand3_1 _17422_ (.A(\u0.w[0][19] ),
    .B(net4230),
    .C(_08258_),
    .Y(_08259_));
 sky130_fd_sc_hd__o21a_4 _17423_ (.A1(\u0.w[0][19] ),
    .A2(_08258_),
    .B1(_08259_),
    .X(_08260_));
 sky130_fd_sc_hd__and2_4 _17424_ (.A(\u0.w[0][19] ),
    .B(_08258_),
    .X(_08261_));
 sky130_fd_sc_hd__nor2_1 _17425_ (.A(\u0.w[0][19] ),
    .B(net4230),
    .Y(_08262_));
 sky130_fd_sc_hd__xnor3_1 _17426_ (.A(\sa20_sr[2] ),
    .B(\sa20_sr[3] ),
    .C(\sa00_sr[3] ),
    .X(_08263_));
 sky130_fd_sc_hd__xnor3_1 _17427_ (.A(_05929_),
    .B(net4109),
    .C(_08263_),
    .X(_08264_));
 sky130_fd_sc_hd__mux2i_4 _17428_ (.A0(_08261_),
    .A1(_08262_),
    .S(_08264_),
    .Y(_08265_));
 sky130_fd_sc_hd__nand2_8 _17429_ (.A(_08260_),
    .B(_08265_),
    .Y(_08266_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_736 ();
 sky130_fd_sc_hd__nand2_8 _17431_ (.A(net3978),
    .B(net3977),
    .Y(_08268_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_735 ();
 sky130_fd_sc_hd__nor2_4 _17433_ (.A(net3689),
    .B(net3978),
    .Y(_08270_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_733 ();
 sky130_fd_sc_hd__nand2_1 _17436_ (.A(net3982),
    .B(net3976),
    .Y(_08273_));
 sky130_fd_sc_hd__nand2_1 _17437_ (.A(_08270_),
    .B(_08273_),
    .Y(_08274_));
 sky130_fd_sc_hd__o21ai_0 _17438_ (.A1(_12097_[0]),
    .A2(_08268_),
    .B1(_08274_),
    .Y(_08275_));
 sky130_fd_sc_hd__xor2_1 _17439_ (.A(\sa20_sr[4] ),
    .B(\sa00_sr[5] ),
    .X(_08276_));
 sky130_fd_sc_hd__xnor2_2 _17440_ (.A(_05911_),
    .B(_08276_),
    .Y(_08277_));
 sky130_fd_sc_hd__mux2i_4 _17441_ (.A0(\text_in_r[117] ),
    .A1(_08277_),
    .S(_05879_),
    .Y(_08278_));
 sky130_fd_sc_hd__xor2_4 _17442_ (.A(net4172),
    .B(_08278_),
    .X(_08279_));
 sky130_fd_sc_hd__xnor3_1 _17443_ (.A(\sa20_sr[3] ),
    .B(\sa30_sr[4] ),
    .C(net4207),
    .X(_08280_));
 sky130_fd_sc_hd__xnor2_1 _17444_ (.A(\sa20_sr[4] ),
    .B(\sa00_sr[4] ),
    .Y(_08281_));
 sky130_fd_sc_hd__xnor3_1 _17445_ (.A(_05925_),
    .B(_08280_),
    .C(_08281_),
    .X(_08282_));
 sky130_fd_sc_hd__mux2i_4 _17446_ (.A0(\text_in_r[116] ),
    .A1(_08282_),
    .S(net4121),
    .Y(_08283_));
 sky130_fd_sc_hd__xnor2_4 _17447_ (.A(\u0.w[0][20] ),
    .B(_08283_),
    .Y(_08284_));
 sky130_fd_sc_hd__nor2_4 _17448_ (.A(_08279_),
    .B(_08284_),
    .Y(_08285_));
 sky130_fd_sc_hd__xnor2_4 _17449_ (.A(net4172),
    .B(_08278_),
    .Y(_08286_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_731 ();
 sky130_fd_sc_hd__nor3_2 _17452_ (.A(net3982),
    .B(net3980),
    .C(_08250_),
    .Y(_08289_));
 sky130_fd_sc_hd__and2_4 _17453_ (.A(_08265_),
    .B(_08260_),
    .X(_08290_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_729 ();
 sky130_fd_sc_hd__xor2_4 _17456_ (.A(\u0.w[0][20] ),
    .B(_08283_),
    .X(_08293_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_728 ();
 sky130_fd_sc_hd__o31ai_2 _17458_ (.A1(_08289_),
    .A2(net3965),
    .A3(_08270_),
    .B1(net3961),
    .Y(_08295_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_726 ();
 sky130_fd_sc_hd__nor2_1 _17461_ (.A(net3981),
    .B(net3978),
    .Y(_08298_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_724 ();
 sky130_fd_sc_hd__nor2_2 _17464_ (.A(_12094_[0]),
    .B(_08250_),
    .Y(_08301_));
 sky130_fd_sc_hd__nor3_1 _17465_ (.A(net3974),
    .B(_08298_),
    .C(_08301_),
    .Y(_08302_));
 sky130_fd_sc_hd__nor3_1 _17466_ (.A(net3968),
    .B(_08295_),
    .C(_08302_),
    .Y(_08303_));
 sky130_fd_sc_hd__a21oi_1 _17467_ (.A1(_08275_),
    .A2(_08285_),
    .B1(_08303_),
    .Y(_08304_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_722 ();
 sky130_fd_sc_hd__nand2_4 _17470_ (.A(net3596),
    .B(net3976),
    .Y(_08307_));
 sky130_fd_sc_hd__nand2_4 _17471_ (.A(net3690),
    .B(_08290_),
    .Y(_08308_));
 sky130_fd_sc_hd__nand2_8 _17472_ (.A(net3982),
    .B(_08290_),
    .Y(_08309_));
 sky130_fd_sc_hd__a32o_1 _17473_ (.A1(net3978),
    .A2(_08307_),
    .A3(_08308_),
    .B1(_08270_),
    .B2(_08309_),
    .X(_08310_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_721 ();
 sky130_fd_sc_hd__nor2_4 _17475_ (.A(net3981),
    .B(_08266_),
    .Y(_08312_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_720 ();
 sky130_fd_sc_hd__nor2_4 _17477_ (.A(_12106_[0]),
    .B(net3963),
    .Y(_08314_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_719 ();
 sky130_fd_sc_hd__nand2_2 _17479_ (.A(net3689),
    .B(net3963),
    .Y(_08316_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_716 ();
 sky130_fd_sc_hd__nand3_1 _17483_ (.A(net3632),
    .B(net3978),
    .C(_08266_),
    .Y(_08320_));
 sky130_fd_sc_hd__o311ai_0 _17484_ (.A1(net3978),
    .A2(_08312_),
    .A3(_08314_),
    .B1(_08316_),
    .C1(_08320_),
    .Y(_08321_));
 sky130_fd_sc_hd__nand2_1 _17485_ (.A(net3968),
    .B(_08321_),
    .Y(_08322_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_714 ();
 sky130_fd_sc_hd__o211ai_1 _17488_ (.A1(net3968),
    .A2(_08310_),
    .B1(_08322_),
    .C1(net3970),
    .Y(_08325_));
 sky130_fd_sc_hd__xnor2_1 _17489_ (.A(\sa20_sr[6] ),
    .B(net4207),
    .Y(_08326_));
 sky130_fd_sc_hd__xnor2_1 _17490_ (.A(_05974_),
    .B(_08326_),
    .Y(_08327_));
 sky130_fd_sc_hd__xnor2_1 _17491_ (.A(net4229),
    .B(_08327_),
    .Y(_08328_));
 sky130_fd_sc_hd__mux2i_2 _17492_ (.A0(\text_in_r[119] ),
    .A1(_08328_),
    .S(_05879_),
    .Y(_08329_));
 sky130_fd_sc_hd__xnor2_4 _17493_ (.A(\u0.w[0][23] ),
    .B(_08329_),
    .Y(_08330_));
 sky130_fd_sc_hd__xnor2_1 _17494_ (.A(net4208),
    .B(\sa00_sr[6] ),
    .Y(_08331_));
 sky130_fd_sc_hd__xnor2_2 _17495_ (.A(_05982_),
    .B(_08331_),
    .Y(_08332_));
 sky130_fd_sc_hd__nor2_2 _17496_ (.A(net398),
    .B(_08332_),
    .Y(_08333_));
 sky130_fd_sc_hd__a21oi_4 _17497_ (.A1(net398),
    .A2(\text_in_r[118] ),
    .B1(_08333_),
    .Y(_08334_));
 sky130_fd_sc_hd__xnor2_4 _17498_ (.A(net4171),
    .B(_08334_),
    .Y(_08335_));
 sky130_fd_sc_hd__nand2b_4 _17499_ (.A_N(_08330_),
    .B(_08335_),
    .Y(_08336_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_713 ();
 sky130_fd_sc_hd__a21oi_1 _17501_ (.A1(_08304_),
    .A2(_08325_),
    .B1(_08336_),
    .Y(_08338_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_711 ();
 sky130_fd_sc_hd__nor2_4 _17504_ (.A(_08250_),
    .B(_08266_),
    .Y(_08341_));
 sky130_fd_sc_hd__nor3_1 _17505_ (.A(net3982),
    .B(_08244_),
    .C(_08250_),
    .Y(_08342_));
 sky130_fd_sc_hd__o21ai_2 _17506_ (.A1(net3597),
    .A2(net3978),
    .B1(net3974),
    .Y(_08343_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_710 ();
 sky130_fd_sc_hd__o21ai_2 _17508_ (.A1(net3619),
    .A2(_08343_),
    .B1(net3961),
    .Y(_08345_));
 sky130_fd_sc_hd__a21oi_1 _17509_ (.A1(_12094_[0]),
    .A2(_08341_),
    .B1(_08345_),
    .Y(_08346_));
 sky130_fd_sc_hd__nor3_4 _17510_ (.A(net3981),
    .B(net3688),
    .C(net3973),
    .Y(_08347_));
 sky130_fd_sc_hd__o21ai_0 _17511_ (.A1(_12094_[0]),
    .A2(net3965),
    .B1(net3978),
    .Y(_08348_));
 sky130_fd_sc_hd__nor2_1 _17512_ (.A(_08347_),
    .B(_08348_),
    .Y(_08349_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_708 ();
 sky130_fd_sc_hd__nand2_8 _17515_ (.A(_08250_),
    .B(net3964),
    .Y(_08352_));
 sky130_fd_sc_hd__nor2_2 _17516_ (.A(_12100_[0]),
    .B(_08352_),
    .Y(_08353_));
 sky130_fd_sc_hd__nor3_1 _17517_ (.A(net3961),
    .B(_08349_),
    .C(_08353_),
    .Y(_08354_));
 sky130_fd_sc_hd__nor2_4 _17518_ (.A(_12097_[0]),
    .B(net3978),
    .Y(_08355_));
 sky130_fd_sc_hd__o31ai_2 _17519_ (.A1(net3974),
    .A2(net3619),
    .A3(_08355_),
    .B1(net3961),
    .Y(_08356_));
 sky130_fd_sc_hd__nor2_1 _17520_ (.A(net3633),
    .B(_08268_),
    .Y(_08357_));
 sky130_fd_sc_hd__nand2_8 _17521_ (.A(net3689),
    .B(net3977),
    .Y(_08358_));
 sky130_fd_sc_hd__nand2_1 _17522_ (.A(_12094_[0]),
    .B(net3964),
    .Y(_08359_));
 sky130_fd_sc_hd__a21oi_1 _17523_ (.A1(_08358_),
    .A2(_08359_),
    .B1(net3978),
    .Y(_08360_));
 sky130_fd_sc_hd__clkinvlp_2 _17524_ (.A(_12093_[0]),
    .Y(_08361_));
 sky130_fd_sc_hd__a21oi_1 _17525_ (.A1(_12113_[0]),
    .A2(net3975),
    .B1(net3961),
    .Y(_08362_));
 sky130_fd_sc_hd__o21ai_0 _17526_ (.A1(net3618),
    .A2(_08352_),
    .B1(_08362_),
    .Y(_08363_));
 sky130_fd_sc_hd__o311ai_0 _17527_ (.A1(_08356_),
    .A2(_08357_),
    .A3(_08360_),
    .B1(_08363_),
    .C1(net3971),
    .Y(_08364_));
 sky130_fd_sc_hd__xor2_4 _17528_ (.A(net4171),
    .B(_08334_),
    .X(_08365_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_707 ();
 sky130_fd_sc_hd__and2_4 _17530_ (.A(_08365_),
    .B(_08330_),
    .X(_08367_));
 sky130_fd_sc_hd__o311a_1 _17531_ (.A1(net3971),
    .A2(_08346_),
    .A3(_08354_),
    .B1(_08364_),
    .C1(_08367_),
    .X(_08368_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_705 ();
 sky130_fd_sc_hd__nand2_4 _17534_ (.A(net3690),
    .B(net3688),
    .Y(_08371_));
 sky130_fd_sc_hd__nor2_1 _17535_ (.A(_12100_[0]),
    .B(net3968),
    .Y(_08372_));
 sky130_fd_sc_hd__a21oi_2 _17536_ (.A1(net3968),
    .A2(_08371_),
    .B1(_08372_),
    .Y(_08373_));
 sky130_fd_sc_hd__xnor2_1 _17537_ (.A(net3968),
    .B(net3965),
    .Y(_08374_));
 sky130_fd_sc_hd__nor2_1 _17538_ (.A(_12100_[0]),
    .B(net3965),
    .Y(_08375_));
 sky130_fd_sc_hd__a22oi_1 _17539_ (.A1(net3632),
    .A2(_08374_),
    .B1(_08375_),
    .B2(net3968),
    .Y(_08376_));
 sky130_fd_sc_hd__nand2_8 _17540_ (.A(_08250_),
    .B(net3973),
    .Y(_08377_));
 sky130_fd_sc_hd__o21ai_0 _17541_ (.A1(net3632),
    .A2(net3971),
    .B1(_08341_),
    .Y(_08378_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_704 ();
 sky130_fd_sc_hd__a21o_1 _17543_ (.A1(_08377_),
    .A2(_08378_),
    .B1(net3633),
    .X(_08380_));
 sky130_fd_sc_hd__o221ai_1 _17544_ (.A1(_08352_),
    .A2(_08373_),
    .B1(_08376_),
    .B2(_08250_),
    .C1(_08380_),
    .Y(_08381_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_702 ();
 sky130_fd_sc_hd__a21oi_1 _17547_ (.A1(net3980),
    .A2(net3968),
    .B1(_08250_),
    .Y(_08384_));
 sky130_fd_sc_hd__nand2_2 _17548_ (.A(_08244_),
    .B(_08250_),
    .Y(_08385_));
 sky130_fd_sc_hd__nand3_1 _17549_ (.A(_12093_[0]),
    .B(net3978),
    .C(net3971),
    .Y(_08386_));
 sky130_fd_sc_hd__o221ai_1 _17550_ (.A1(net3982),
    .A2(_08384_),
    .B1(_08385_),
    .B2(net3971),
    .C1(_08386_),
    .Y(_08387_));
 sky130_fd_sc_hd__nand2_8 _17551_ (.A(_08244_),
    .B(net3978),
    .Y(_08388_));
 sky130_fd_sc_hd__nand2_4 _17552_ (.A(net3982),
    .B(net3980),
    .Y(_08389_));
 sky130_fd_sc_hd__a21oi_1 _17553_ (.A1(_08388_),
    .A2(_08389_),
    .B1(net3971),
    .Y(_08390_));
 sky130_fd_sc_hd__o31ai_1 _17554_ (.A1(net3632),
    .A2(net3978),
    .A3(net3968),
    .B1(net3974),
    .Y(_08391_));
 sky130_fd_sc_hd__o22ai_1 _17555_ (.A1(net3974),
    .A2(_08387_),
    .B1(_08390_),
    .B2(_08391_),
    .Y(_08392_));
 sky130_fd_sc_hd__nor2_4 _17556_ (.A(_08335_),
    .B(_08330_),
    .Y(_08393_));
 sky130_fd_sc_hd__o21ai_1 _17557_ (.A1(net3961),
    .A2(_08392_),
    .B1(_08393_),
    .Y(_08394_));
 sky130_fd_sc_hd__a21oi_1 _17558_ (.A1(net3961),
    .A2(_08381_),
    .B1(_08394_),
    .Y(_08395_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_700 ();
 sky130_fd_sc_hd__nor2_4 _17561_ (.A(net3632),
    .B(net3974),
    .Y(_08398_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_699 ();
 sky130_fd_sc_hd__nand3_1 _17563_ (.A(net3978),
    .B(_08309_),
    .C(_08358_),
    .Y(_08400_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_698 ();
 sky130_fd_sc_hd__o311ai_0 _17565_ (.A1(net3978),
    .A2(_08375_),
    .A3(_08398_),
    .B1(_08400_),
    .C1(net3961),
    .Y(_08402_));
 sky130_fd_sc_hd__nor2_4 _17566_ (.A(_12097_[0]),
    .B(net3963),
    .Y(_08403_));
 sky130_fd_sc_hd__nor2_4 _17567_ (.A(_12094_[0]),
    .B(_08266_),
    .Y(_08404_));
 sky130_fd_sc_hd__o21ai_2 _17568_ (.A1(_08403_),
    .A2(_08404_),
    .B1(net3978),
    .Y(_08405_));
 sky130_fd_sc_hd__nor2_4 _17569_ (.A(net3978),
    .B(_08266_),
    .Y(_08406_));
 sky130_fd_sc_hd__nand2_1 _17570_ (.A(net3633),
    .B(_08406_),
    .Y(_08407_));
 sky130_fd_sc_hd__nand3_1 _17571_ (.A(net3970),
    .B(_08405_),
    .C(_08407_),
    .Y(_08408_));
 sky130_fd_sc_hd__nand3_1 _17572_ (.A(net3968),
    .B(_08402_),
    .C(_08408_),
    .Y(_08409_));
 sky130_fd_sc_hd__nand2_4 _17573_ (.A(net3980),
    .B(net3974),
    .Y(_08410_));
 sky130_fd_sc_hd__nor2_2 _17574_ (.A(net3970),
    .B(_08410_),
    .Y(_08411_));
 sky130_fd_sc_hd__nor2_2 _17575_ (.A(_12097_[0]),
    .B(net3974),
    .Y(_08412_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_696 ();
 sky130_fd_sc_hd__nand2_2 _17578_ (.A(net3632),
    .B(net3974),
    .Y(_08415_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_695 ();
 sky130_fd_sc_hd__nand2_4 _17580_ (.A(net3597),
    .B(net397),
    .Y(_08417_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_694 ();
 sky130_fd_sc_hd__a21oi_1 _17582_ (.A1(_08415_),
    .A2(_08417_),
    .B1(_08250_),
    .Y(_08419_));
 sky130_fd_sc_hd__o21ai_0 _17583_ (.A1(net3961),
    .A2(_08419_),
    .B1(_08295_),
    .Y(_08420_));
 sky130_fd_sc_hd__o311ai_1 _17584_ (.A1(net3978),
    .A2(_08411_),
    .A3(_08412_),
    .B1(_08279_),
    .C1(_08420_),
    .Y(_08421_));
 sky130_fd_sc_hd__nand2_4 _17585_ (.A(_08335_),
    .B(_08330_),
    .Y(_08422_));
 sky130_fd_sc_hd__a21oi_1 _17586_ (.A1(_08409_),
    .A2(_08421_),
    .B1(_08422_),
    .Y(_08423_));
 sky130_fd_sc_hd__nor4_1 _17587_ (.A(_08338_),
    .B(_08368_),
    .C(_08395_),
    .D(_08423_),
    .Y(_00064_));
 sky130_fd_sc_hd__nor2_4 _17588_ (.A(_08244_),
    .B(_08290_),
    .Y(_08424_));
 sky130_fd_sc_hd__o21ai_0 _17589_ (.A1(net3978),
    .A2(_08424_),
    .B1(net3690),
    .Y(_08425_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_693 ();
 sky130_fd_sc_hd__nor2_4 _17591_ (.A(_08244_),
    .B(_08266_),
    .Y(_08426_));
 sky130_fd_sc_hd__nand2_1 _17592_ (.A(net3982),
    .B(_08426_),
    .Y(_08427_));
 sky130_fd_sc_hd__nand4_1 _17593_ (.A(_08268_),
    .B(_08285_),
    .C(_08425_),
    .D(_08427_),
    .Y(_08428_));
 sky130_fd_sc_hd__nand2_4 _17594_ (.A(_12097_[0]),
    .B(net3966),
    .Y(_08429_));
 sky130_fd_sc_hd__a21oi_1 _17595_ (.A1(_08415_),
    .A2(_08429_),
    .B1(_08250_),
    .Y(_08430_));
 sky130_fd_sc_hd__nor2_2 _17596_ (.A(net3980),
    .B(_08266_),
    .Y(_08431_));
 sky130_fd_sc_hd__nor3_1 _17597_ (.A(net3978),
    .B(_08431_),
    .C(_08424_),
    .Y(_08432_));
 sky130_fd_sc_hd__nor2_4 _17598_ (.A(_08279_),
    .B(net3960),
    .Y(_08433_));
 sky130_fd_sc_hd__o21ai_2 _17599_ (.A1(_08430_),
    .A2(_08432_),
    .B1(_08433_),
    .Y(_08434_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_692 ();
 sky130_fd_sc_hd__mux2i_1 _17601_ (.A0(net3632),
    .A1(_12106_[0]),
    .S(net3978),
    .Y(_08436_));
 sky130_fd_sc_hd__nor2_1 _17602_ (.A(net397),
    .B(_08436_),
    .Y(_08437_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_691 ();
 sky130_fd_sc_hd__xnor2_2 _17604_ (.A(_08250_),
    .B(net3964),
    .Y(_08439_));
 sky130_fd_sc_hd__o22ai_1 _17605_ (.A1(_12097_[0]),
    .A2(_08352_),
    .B1(_08439_),
    .B2(net3982),
    .Y(_08440_));
 sky130_fd_sc_hd__a21oi_1 _17606_ (.A1(net3970),
    .A2(_08440_),
    .B1(net3968),
    .Y(_08441_));
 sky130_fd_sc_hd__o21ai_2 _17607_ (.A1(_08356_),
    .A2(_08437_),
    .B1(_08441_),
    .Y(_08442_));
 sky130_fd_sc_hd__nand2_4 _17608_ (.A(net3690),
    .B(net3973),
    .Y(_08443_));
 sky130_fd_sc_hd__xnor2_1 _17609_ (.A(net3688),
    .B(_08250_),
    .Y(_08444_));
 sky130_fd_sc_hd__mux2i_1 _17610_ (.A0(_12092_[0]),
    .A1(net3980),
    .S(net3978),
    .Y(_08445_));
 sky130_fd_sc_hd__o22ai_1 _17611_ (.A1(_08443_),
    .A2(_08444_),
    .B1(_08445_),
    .B2(net3973),
    .Y(_08446_));
 sky130_fd_sc_hd__nand2_1 _17612_ (.A(_08286_),
    .B(_08446_),
    .Y(_08447_));
 sky130_fd_sc_hd__and2_4 _17613_ (.A(_12097_[0]),
    .B(_08266_),
    .X(_08448_));
 sky130_fd_sc_hd__o21ai_2 _17614_ (.A1(_08426_),
    .A2(_08448_),
    .B1(net3978),
    .Y(_08449_));
 sky130_fd_sc_hd__nor2_2 _17615_ (.A(net3690),
    .B(net3976),
    .Y(_08450_));
 sky130_fd_sc_hd__nor2_4 _17616_ (.A(net3982),
    .B(_08290_),
    .Y(_08451_));
 sky130_fd_sc_hd__o21ai_0 _17617_ (.A1(_08450_),
    .A2(_08451_),
    .B1(_08250_),
    .Y(_08452_));
 sky130_fd_sc_hd__a31oi_1 _17618_ (.A1(net3972),
    .A2(_08449_),
    .A3(_08452_),
    .B1(net3960),
    .Y(_08453_));
 sky130_fd_sc_hd__nand2_2 _17619_ (.A(_12100_[0]),
    .B(_08250_),
    .Y(_08454_));
 sky130_fd_sc_hd__nor3b_2 _17620_ (.A(_08289_),
    .B(net3975),
    .C_N(_08454_),
    .Y(_08455_));
 sky130_fd_sc_hd__nor3_1 _17621_ (.A(_12116_[0]),
    .B(_08286_),
    .C(net3964),
    .Y(_08456_));
 sky130_fd_sc_hd__or2_4 _17622_ (.A(_08455_),
    .B(_08456_),
    .X(_08457_));
 sky130_fd_sc_hd__a221oi_1 _17623_ (.A1(_08447_),
    .A2(_08453_),
    .B1(_08457_),
    .B2(net3960),
    .C1(_08330_),
    .Y(_08458_));
 sky130_fd_sc_hd__a41oi_2 _17624_ (.A1(_08330_),
    .A2(_08428_),
    .A3(_08434_),
    .A4(_08442_),
    .B1(_08458_),
    .Y(_08459_));
 sky130_fd_sc_hd__a21oi_1 _17625_ (.A1(net3690),
    .A2(_08244_),
    .B1(net3962),
    .Y(_08460_));
 sky130_fd_sc_hd__nand2_1 _17626_ (.A(_08361_),
    .B(net3976),
    .Y(_08461_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_690 ();
 sky130_fd_sc_hd__a21oi_1 _17628_ (.A1(net3588),
    .A2(_08429_),
    .B1(_08250_),
    .Y(_08463_));
 sky130_fd_sc_hd__a21o_1 _17629_ (.A1(_08250_),
    .A2(_08460_),
    .B1(_08463_),
    .X(_08464_));
 sky130_fd_sc_hd__nor2_1 _17630_ (.A(net3690),
    .B(_08358_),
    .Y(_08465_));
 sky130_fd_sc_hd__o22ai_2 _17631_ (.A1(net3618),
    .A2(_08352_),
    .B1(_08439_),
    .B2(_08244_),
    .Y(_08466_));
 sky130_fd_sc_hd__nor3_1 _17632_ (.A(_08286_),
    .B(_08465_),
    .C(_08466_),
    .Y(_08467_));
 sky130_fd_sc_hd__a21oi_1 _17633_ (.A1(_08286_),
    .A2(_08464_),
    .B1(_08467_),
    .Y(_08468_));
 sky130_fd_sc_hd__nor2_2 _17634_ (.A(_08371_),
    .B(net3976),
    .Y(_08469_));
 sky130_fd_sc_hd__nor2_2 _17635_ (.A(net3690),
    .B(_08268_),
    .Y(_08470_));
 sky130_fd_sc_hd__a2111oi_0 _17636_ (.A1(_08250_),
    .A2(_08307_),
    .B1(_08469_),
    .C1(_08470_),
    .D1(_08279_),
    .Y(_08471_));
 sky130_fd_sc_hd__nor2_2 _17637_ (.A(_12093_[0]),
    .B(_08290_),
    .Y(_08472_));
 sky130_fd_sc_hd__nor2_4 _17638_ (.A(_12092_[0]),
    .B(_08266_),
    .Y(_08473_));
 sky130_fd_sc_hd__o21ai_0 _17639_ (.A1(_08426_),
    .A2(_08403_),
    .B1(_08250_),
    .Y(_08474_));
 sky130_fd_sc_hd__o311a_1 _17640_ (.A1(_08250_),
    .A2(net3617),
    .A3(_08473_),
    .B1(_08474_),
    .C1(_08279_),
    .X(_08475_));
 sky130_fd_sc_hd__o21ai_0 _17641_ (.A1(_08471_),
    .A2(_08475_),
    .B1(net3969),
    .Y(_08476_));
 sky130_fd_sc_hd__and2_4 _17642_ (.A(_08335_),
    .B(_08330_),
    .X(_08477_));
 sky130_fd_sc_hd__o211ai_1 _17643_ (.A1(net3969),
    .A2(_08468_),
    .B1(_08476_),
    .C1(_08477_),
    .Y(_08478_));
 sky130_fd_sc_hd__nor3_1 _17644_ (.A(net3978),
    .B(_08426_),
    .C(net3617),
    .Y(_08479_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_689 ();
 sky130_fd_sc_hd__a211oi_1 _17646_ (.A1(_12092_[0]),
    .A2(net3973),
    .B1(_08404_),
    .C1(_08250_),
    .Y(_08481_));
 sky130_fd_sc_hd__o21ai_0 _17647_ (.A1(_08479_),
    .A2(_08481_),
    .B1(_08433_),
    .Y(_08482_));
 sky130_fd_sc_hd__o21ai_0 _17648_ (.A1(_08451_),
    .A2(_08473_),
    .B1(_08250_),
    .Y(_08483_));
 sky130_fd_sc_hd__nand2_1 _17649_ (.A(_08449_),
    .B(_08483_),
    .Y(_08484_));
 sky130_fd_sc_hd__a21oi_1 _17650_ (.A1(_08285_),
    .A2(_08484_),
    .B1(_08336_),
    .Y(_08485_));
 sky130_fd_sc_hd__nor3_4 _17651_ (.A(net3982),
    .B(net3980),
    .C(net3963),
    .Y(_08486_));
 sky130_fd_sc_hd__nor2_2 _17652_ (.A(_08404_),
    .B(_08486_),
    .Y(_08487_));
 sky130_fd_sc_hd__nor2_4 _17653_ (.A(_08286_),
    .B(net3960),
    .Y(_08488_));
 sky130_fd_sc_hd__nand2_8 _17654_ (.A(_12106_[0]),
    .B(_08290_),
    .Y(_08489_));
 sky130_fd_sc_hd__nand3_1 _17655_ (.A(net3978),
    .B(net3588),
    .C(_08489_),
    .Y(_08490_));
 sky130_fd_sc_hd__o211ai_1 _17656_ (.A1(net3978),
    .A2(_08487_),
    .B1(_08488_),
    .C1(_08490_),
    .Y(_08491_));
 sky130_fd_sc_hd__o21ai_0 _17657_ (.A1(net3617),
    .A2(_08469_),
    .B1(net3978),
    .Y(_08492_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_688 ();
 sky130_fd_sc_hd__nor2_4 _17659_ (.A(net3967),
    .B(net3969),
    .Y(_08494_));
 sky130_fd_sc_hd__nand2_4 _17660_ (.A(net3980),
    .B(_08406_),
    .Y(_08495_));
 sky130_fd_sc_hd__nand3_1 _17661_ (.A(_08492_),
    .B(_08494_),
    .C(_08495_),
    .Y(_08496_));
 sky130_fd_sc_hd__nand4_1 _17662_ (.A(_08482_),
    .B(_08485_),
    .C(_08491_),
    .D(_08496_),
    .Y(_08497_));
 sky130_fd_sc_hd__o211a_1 _17663_ (.A1(_08335_),
    .A2(_08459_),
    .B1(_08478_),
    .C1(_08497_),
    .X(_00065_));
 sky130_fd_sc_hd__nand2_2 _17664_ (.A(_12100_[0]),
    .B(_08266_),
    .Y(_08498_));
 sky130_fd_sc_hd__and3_4 _17665_ (.A(_12092_[0]),
    .B(_08260_),
    .C(_08265_),
    .X(_08499_));
 sky130_fd_sc_hd__nor3_1 _17666_ (.A(net3978),
    .B(net3616),
    .C(_08499_),
    .Y(_08500_));
 sky130_fd_sc_hd__a311oi_1 _17667_ (.A1(net3978),
    .A2(_08309_),
    .A3(_08498_),
    .B1(_08500_),
    .C1(_08286_),
    .Y(_08501_));
 sky130_fd_sc_hd__nor2_1 _17668_ (.A(net3690),
    .B(net3978),
    .Y(_08502_));
 sky130_fd_sc_hd__o21ai_0 _17669_ (.A1(_08312_),
    .A2(_08502_),
    .B1(_12093_[0]),
    .Y(_08503_));
 sky130_fd_sc_hd__nor2_1 _17670_ (.A(net3981),
    .B(_08250_),
    .Y(_08504_));
 sky130_fd_sc_hd__a32oi_1 _17671_ (.A1(net3981),
    .A2(_08388_),
    .A3(net3973),
    .B1(_08358_),
    .B2(_08504_),
    .Y(_08505_));
 sky130_fd_sc_hd__a21oi_1 _17672_ (.A1(_08503_),
    .A2(_08505_),
    .B1(net3972),
    .Y(_08506_));
 sky130_fd_sc_hd__or3_1 _17673_ (.A(net3960),
    .B(_08501_),
    .C(_08506_),
    .X(_08507_));
 sky130_fd_sc_hd__nand2_4 _17674_ (.A(net3690),
    .B(net3978),
    .Y(_08508_));
 sky130_fd_sc_hd__nand3_1 _17675_ (.A(net3974),
    .B(_08389_),
    .C(_08508_),
    .Y(_08509_));
 sky130_fd_sc_hd__o211ai_1 _17676_ (.A1(_12116_[0]),
    .A2(net3974),
    .B1(_08509_),
    .C1(_08279_),
    .Y(_08510_));
 sky130_fd_sc_hd__o21ai_0 _17677_ (.A1(net3632),
    .A2(net3978),
    .B1(net3974),
    .Y(_08511_));
 sky130_fd_sc_hd__a21oi_1 _17678_ (.A1(_12113_[0]),
    .A2(net397),
    .B1(net3971),
    .Y(_08512_));
 sky130_fd_sc_hd__o21ai_2 _17679_ (.A1(net3619),
    .A2(_08511_),
    .B1(_08512_),
    .Y(_08513_));
 sky130_fd_sc_hd__nand3_2 _17680_ (.A(net3961),
    .B(_08510_),
    .C(_08513_),
    .Y(_08514_));
 sky130_fd_sc_hd__a21oi_1 _17681_ (.A1(_08507_),
    .A2(_08514_),
    .B1(_08422_),
    .Y(_08515_));
 sky130_fd_sc_hd__nor3_1 _17682_ (.A(_08250_),
    .B(_08398_),
    .C(_08424_),
    .Y(_08516_));
 sky130_fd_sc_hd__nand2_2 _17683_ (.A(_12094_[0]),
    .B(net3974),
    .Y(_08517_));
 sky130_fd_sc_hd__a21oi_1 _17684_ (.A1(_08309_),
    .A2(_08517_),
    .B1(net3978),
    .Y(_08518_));
 sky130_fd_sc_hd__o21ai_0 _17685_ (.A1(_08516_),
    .A2(_08518_),
    .B1(net3970),
    .Y(_08519_));
 sky130_fd_sc_hd__nand2_1 _17686_ (.A(_08238_),
    .B(_08432_),
    .Y(_08520_));
 sky130_fd_sc_hd__o211ai_1 _17687_ (.A1(_12106_[0]),
    .A2(_08268_),
    .B1(_08520_),
    .C1(net3961),
    .Y(_08521_));
 sky130_fd_sc_hd__o21ai_1 _17688_ (.A1(_08342_),
    .A2(_08355_),
    .B1(net3974),
    .Y(_08522_));
 sky130_fd_sc_hd__o211ai_1 _17689_ (.A1(net3618),
    .A2(net3978),
    .B1(net3964),
    .C1(_08508_),
    .Y(_08523_));
 sky130_fd_sc_hd__a21oi_1 _17690_ (.A1(_12106_[0]),
    .A2(_08250_),
    .B1(net3974),
    .Y(_08524_));
 sky130_fd_sc_hd__nand2_1 _17691_ (.A(_12097_[0]),
    .B(net3978),
    .Y(_08525_));
 sky130_fd_sc_hd__a221oi_1 _17692_ (.A1(_08385_),
    .A2(_08451_),
    .B1(_08524_),
    .B2(_08525_),
    .C1(_08293_),
    .Y(_08526_));
 sky130_fd_sc_hd__a311oi_1 _17693_ (.A1(net3961),
    .A2(_08522_),
    .A3(_08523_),
    .B1(_08526_),
    .C1(net3968),
    .Y(_08527_));
 sky130_fd_sc_hd__or2_4 _17694_ (.A(_08335_),
    .B(_08330_),
    .X(_08528_));
 sky130_fd_sc_hd__a311oi_2 _17695_ (.A1(net3968),
    .A2(_08519_),
    .A3(_08521_),
    .B1(_08527_),
    .C1(_08528_),
    .Y(_08529_));
 sky130_fd_sc_hd__nor2_4 _17696_ (.A(_12094_[0]),
    .B(_12097_[0]),
    .Y(_08530_));
 sky130_fd_sc_hd__a21oi_1 _17697_ (.A1(net3976),
    .A2(_08530_),
    .B1(_08469_),
    .Y(_08531_));
 sky130_fd_sc_hd__a211oi_1 _17698_ (.A1(_12100_[0]),
    .A2(net3963),
    .B1(_08486_),
    .C1(net3979),
    .Y(_08532_));
 sky130_fd_sc_hd__a21oi_1 _17699_ (.A1(net3979),
    .A2(_08531_),
    .B1(_08532_),
    .Y(_08533_));
 sky130_fd_sc_hd__nor2_4 _17700_ (.A(net3978),
    .B(net3964),
    .Y(_08534_));
 sky130_fd_sc_hd__nand2_2 _17701_ (.A(_12097_[0]),
    .B(_08534_),
    .Y(_08535_));
 sky130_fd_sc_hd__o311ai_0 _17702_ (.A1(_08250_),
    .A2(net3617),
    .A3(_08499_),
    .B1(_08535_),
    .C1(_08285_),
    .Y(_08536_));
 sky130_fd_sc_hd__nand2_1 _17703_ (.A(_12111_[0]),
    .B(net3973),
    .Y(_08537_));
 sky130_fd_sc_hd__o41ai_1 _17704_ (.A1(net3981),
    .A2(_08244_),
    .A3(net3978),
    .A4(net3973),
    .B1(_08537_),
    .Y(_08538_));
 sky130_fd_sc_hd__nor2_2 _17705_ (.A(net3980),
    .B(net3978),
    .Y(_08539_));
 sky130_fd_sc_hd__o221ai_1 _17706_ (.A1(_12120_[0]),
    .A2(net3973),
    .B1(_08539_),
    .B2(_08443_),
    .C1(net3969),
    .Y(_08540_));
 sky130_fd_sc_hd__o211ai_1 _17707_ (.A1(net3969),
    .A2(_08538_),
    .B1(_08540_),
    .C1(_08279_),
    .Y(_08541_));
 sky130_fd_sc_hd__nand3_1 _17708_ (.A(_08367_),
    .B(_08536_),
    .C(_08541_),
    .Y(_08542_));
 sky130_fd_sc_hd__a21oi_1 _17709_ (.A1(_08433_),
    .A2(_08533_),
    .B1(_08542_),
    .Y(_08543_));
 sky130_fd_sc_hd__nor2_2 _17710_ (.A(net3597),
    .B(net3976),
    .Y(_08544_));
 sky130_fd_sc_hd__nor3_1 _17711_ (.A(_08250_),
    .B(_08424_),
    .C(_08544_),
    .Y(_08545_));
 sky130_fd_sc_hd__nor2_1 _17712_ (.A(net3596),
    .B(net3976),
    .Y(_08546_));
 sky130_fd_sc_hd__nor3_1 _17713_ (.A(net3978),
    .B(_08403_),
    .C(_08546_),
    .Y(_08547_));
 sky130_fd_sc_hd__o21ai_0 _17714_ (.A1(_08545_),
    .A2(_08547_),
    .B1(_08488_),
    .Y(_08548_));
 sky130_fd_sc_hd__nor2_1 _17715_ (.A(net3597),
    .B(_08250_),
    .Y(_08549_));
 sky130_fd_sc_hd__o21ai_1 _17716_ (.A1(_08298_),
    .A2(_08549_),
    .B1(net3974),
    .Y(_08550_));
 sky130_fd_sc_hd__nand2_1 _17717_ (.A(_08388_),
    .B(_08524_),
    .Y(_08551_));
 sky130_fd_sc_hd__nand3_2 _17718_ (.A(_08433_),
    .B(_08550_),
    .C(_08551_),
    .Y(_08552_));
 sky130_fd_sc_hd__nand3_1 _17719_ (.A(_08250_),
    .B(_08417_),
    .C(net3588),
    .Y(_08553_));
 sky130_fd_sc_hd__o21ai_0 _17720_ (.A1(_08426_),
    .A2(net3616),
    .B1(net3979),
    .Y(_08554_));
 sky130_fd_sc_hd__a21oi_1 _17721_ (.A1(_12102_[0]),
    .A2(_08290_),
    .B1(_08451_),
    .Y(_08555_));
 sky130_fd_sc_hd__nand2_4 _17722_ (.A(_08279_),
    .B(net3960),
    .Y(_08556_));
 sky130_fd_sc_hd__a211oi_2 _17723_ (.A1(net3978),
    .A2(_08555_),
    .B1(_08556_),
    .C1(_08355_),
    .Y(_08557_));
 sky130_fd_sc_hd__a31oi_1 _17724_ (.A1(_08285_),
    .A2(_08553_),
    .A3(_08554_),
    .B1(_08557_),
    .Y(_08558_));
 sky130_fd_sc_hd__a31oi_1 _17725_ (.A1(_08548_),
    .A2(_08552_),
    .A3(_08558_),
    .B1(_08336_),
    .Y(_08559_));
 sky130_fd_sc_hd__or4_4 _17726_ (.A(_08515_),
    .B(_08529_),
    .C(_08543_),
    .D(_08559_),
    .X(_00066_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_687 ();
 sky130_fd_sc_hd__nor2_1 _17728_ (.A(_12100_[0]),
    .B(_08266_),
    .Y(_08561_));
 sky130_fd_sc_hd__nor2_1 _17729_ (.A(net3633),
    .B(net3963),
    .Y(_08562_));
 sky130_fd_sc_hd__nor3_1 _17730_ (.A(_08250_),
    .B(_08561_),
    .C(_08562_),
    .Y(_08563_));
 sky130_fd_sc_hd__a31oi_1 _17731_ (.A1(_08250_),
    .A2(_08316_),
    .A3(net3588),
    .B1(_08563_),
    .Y(_08564_));
 sky130_fd_sc_hd__nand2_2 _17732_ (.A(_12093_[0]),
    .B(net3963),
    .Y(_08565_));
 sky130_fd_sc_hd__o211ai_1 _17733_ (.A1(net3596),
    .A2(net3963),
    .B1(_08565_),
    .C1(net3979),
    .Y(_08566_));
 sky130_fd_sc_hd__o311ai_0 _17734_ (.A1(net3979),
    .A2(_08450_),
    .A3(_08403_),
    .B1(_08566_),
    .C1(net3960),
    .Y(_08567_));
 sky130_fd_sc_hd__o21ai_0 _17735_ (.A1(net3960),
    .A2(_08564_),
    .B1(_08567_),
    .Y(_08568_));
 sky130_fd_sc_hd__nand2_1 _17736_ (.A(net3968),
    .B(_08367_),
    .Y(_08569_));
 sky130_fd_sc_hd__nand2_1 _17737_ (.A(net3972),
    .B(_08367_),
    .Y(_08570_));
 sky130_fd_sc_hd__nor2_2 _17738_ (.A(_08250_),
    .B(_08293_),
    .Y(_08571_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_686 ();
 sky130_fd_sc_hd__a211oi_1 _17740_ (.A1(net3980),
    .A2(net3960),
    .B1(net3978),
    .C1(net3982),
    .Y(_08573_));
 sky130_fd_sc_hd__a31oi_1 _17741_ (.A1(net3982),
    .A2(net3960),
    .A3(_08388_),
    .B1(_08573_),
    .Y(_08574_));
 sky130_fd_sc_hd__nand2_1 _17742_ (.A(_08250_),
    .B(_08293_),
    .Y(_08575_));
 sky130_fd_sc_hd__nor3_1 _17743_ (.A(net3982),
    .B(net3978),
    .C(_08284_),
    .Y(_08576_));
 sky130_fd_sc_hd__a2111oi_0 _17744_ (.A1(_12093_[0]),
    .A2(_08575_),
    .B1(_08576_),
    .C1(net397),
    .D1(_08571_),
    .Y(_08577_));
 sky130_fd_sc_hd__a21oi_1 _17745_ (.A1(net397),
    .A2(_08574_),
    .B1(_08577_),
    .Y(_08578_));
 sky130_fd_sc_hd__a21oi_2 _17746_ (.A1(net3688),
    .A2(_08571_),
    .B1(_08578_),
    .Y(_08579_));
 sky130_fd_sc_hd__o22a_1 _17747_ (.A1(_08568_),
    .A2(_08569_),
    .B1(_08570_),
    .B2(_08579_),
    .X(_08580_));
 sky130_fd_sc_hd__a21oi_1 _17748_ (.A1(net3978),
    .A2(_08530_),
    .B1(_08343_),
    .Y(_08581_));
 sky130_fd_sc_hd__a21oi_1 _17749_ (.A1(net3978),
    .A2(_08309_),
    .B1(net3980),
    .Y(_08582_));
 sky130_fd_sc_hd__o221ai_1 _17750_ (.A1(net3633),
    .A2(_08268_),
    .B1(_08352_),
    .B2(net3981),
    .C1(net3968),
    .Y(_08583_));
 sky130_fd_sc_hd__o32a_1 _17751_ (.A1(net3968),
    .A2(_08455_),
    .A3(_08581_),
    .B1(_08582_),
    .B2(_08583_),
    .X(_08584_));
 sky130_fd_sc_hd__nor2_1 _17752_ (.A(_12102_[0]),
    .B(net3964),
    .Y(_08585_));
 sky130_fd_sc_hd__o21ai_1 _17753_ (.A1(_08398_),
    .A2(net3586),
    .B1(net3978),
    .Y(_08586_));
 sky130_fd_sc_hd__nand3_1 _17754_ (.A(_08250_),
    .B(_08410_),
    .C(net3587),
    .Y(_08587_));
 sky130_fd_sc_hd__nand3_1 _17755_ (.A(net3968),
    .B(_08586_),
    .C(_08587_),
    .Y(_08588_));
 sky130_fd_sc_hd__a21oi_1 _17756_ (.A1(net3971),
    .A2(_08551_),
    .B1(net3961),
    .Y(_08589_));
 sky130_fd_sc_hd__a21oi_1 _17757_ (.A1(_08588_),
    .A2(_08589_),
    .B1(_08336_),
    .Y(_08590_));
 sky130_fd_sc_hd__o21ai_1 _17758_ (.A1(net3970),
    .A2(_08584_),
    .B1(_08590_),
    .Y(_08591_));
 sky130_fd_sc_hd__nor2_1 _17759_ (.A(net3970),
    .B(_08539_),
    .Y(_08592_));
 sky130_fd_sc_hd__a21o_1 _17760_ (.A1(_08273_),
    .A2(_08565_),
    .B1(_08250_),
    .X(_08593_));
 sky130_fd_sc_hd__o21ai_0 _17761_ (.A1(_08314_),
    .A2(_08544_),
    .B1(_08250_),
    .Y(_08594_));
 sky130_fd_sc_hd__a21oi_1 _17762_ (.A1(_08593_),
    .A2(_08594_),
    .B1(net3960),
    .Y(_08595_));
 sky130_fd_sc_hd__a311oi_1 _17763_ (.A1(_08268_),
    .A2(_08389_),
    .A3(_08592_),
    .B1(_08595_),
    .C1(_08286_),
    .Y(_08596_));
 sky130_fd_sc_hd__nor3_2 _17764_ (.A(net3980),
    .B(_08250_),
    .C(net3974),
    .Y(_08597_));
 sky130_fd_sc_hd__a21oi_1 _17765_ (.A1(_08266_),
    .A2(_08270_),
    .B1(_08597_),
    .Y(_08598_));
 sky130_fd_sc_hd__nor2_2 _17766_ (.A(_08250_),
    .B(net3965),
    .Y(_08599_));
 sky130_fd_sc_hd__nand2_1 _17767_ (.A(_12100_[0]),
    .B(_08599_),
    .Y(_08600_));
 sky130_fd_sc_hd__o211ai_1 _17768_ (.A1(net3981),
    .A2(_08598_),
    .B1(_08600_),
    .C1(_08285_),
    .Y(_08601_));
 sky130_fd_sc_hd__a21oi_1 _17769_ (.A1(net3618),
    .A2(_08406_),
    .B1(_08601_),
    .Y(_08602_));
 sky130_fd_sc_hd__nand2_2 _17770_ (.A(_08286_),
    .B(_08284_),
    .Y(_08603_));
 sky130_fd_sc_hd__o22ai_1 _17771_ (.A1(_08238_),
    .A2(_08410_),
    .B1(_08454_),
    .B2(net3975),
    .Y(_08604_));
 sky130_fd_sc_hd__nor3_1 _17772_ (.A(_08603_),
    .B(_08516_),
    .C(_08604_),
    .Y(_08605_));
 sky130_fd_sc_hd__o31ai_1 _17773_ (.A1(_08596_),
    .A2(_08602_),
    .A3(_08605_),
    .B1(_08477_),
    .Y(_08606_));
 sky130_fd_sc_hd__nand2_1 _17774_ (.A(net3978),
    .B(net3970),
    .Y(_08607_));
 sky130_fd_sc_hd__a21oi_1 _17775_ (.A1(_12094_[0]),
    .A2(net3975),
    .B1(_08398_),
    .Y(_08608_));
 sky130_fd_sc_hd__a21oi_1 _17776_ (.A1(net3597),
    .A2(_08439_),
    .B1(_08597_),
    .Y(_08609_));
 sky130_fd_sc_hd__o221ai_2 _17777_ (.A1(_08607_),
    .A2(_08608_),
    .B1(_08609_),
    .B2(net3970),
    .C1(net3968),
    .Y(_08610_));
 sky130_fd_sc_hd__nand2_1 _17778_ (.A(net3976),
    .B(_08530_),
    .Y(_08611_));
 sky130_fd_sc_hd__o211ai_1 _17779_ (.A1(_12093_[0]),
    .A2(net3976),
    .B1(_08611_),
    .C1(net3979),
    .Y(_08612_));
 sky130_fd_sc_hd__o311ai_0 _17780_ (.A1(net3979),
    .A2(_08314_),
    .A3(_08426_),
    .B1(_08494_),
    .C1(_08612_),
    .Y(_08613_));
 sky130_fd_sc_hd__nand3_1 _17781_ (.A(net3979),
    .B(_08309_),
    .C(_08517_),
    .Y(_08614_));
 sky130_fd_sc_hd__o31ai_1 _17782_ (.A1(net3979),
    .A2(net3616),
    .A3(_08561_),
    .B1(_08614_),
    .Y(_08615_));
 sky130_fd_sc_hd__a21oi_1 _17783_ (.A1(_08488_),
    .A2(_08615_),
    .B1(_08528_),
    .Y(_08616_));
 sky130_fd_sc_hd__nand3_1 _17784_ (.A(_08610_),
    .B(_08613_),
    .C(_08616_),
    .Y(_08617_));
 sky130_fd_sc_hd__nand4_1 _17785_ (.A(_08580_),
    .B(_08591_),
    .C(_08606_),
    .D(_08617_),
    .Y(_00067_));
 sky130_fd_sc_hd__nand2_1 _17786_ (.A(_08250_),
    .B(_08443_),
    .Y(_08618_));
 sky130_fd_sc_hd__o211ai_1 _17787_ (.A1(_08499_),
    .A2(_08618_),
    .B1(_08388_),
    .C1(_08285_),
    .Y(_08619_));
 sky130_fd_sc_hd__a21oi_2 _17788_ (.A1(_12102_[0]),
    .A2(net3973),
    .B1(net3978),
    .Y(_08620_));
 sky130_fd_sc_hd__o21ai_0 _17789_ (.A1(_08404_),
    .A2(_08620_),
    .B1(_08433_),
    .Y(_08621_));
 sky130_fd_sc_hd__nand3_2 _17790_ (.A(_08477_),
    .B(_08619_),
    .C(_08621_),
    .Y(_08622_));
 sky130_fd_sc_hd__nor2_1 _17791_ (.A(_08284_),
    .B(_08508_),
    .Y(_08623_));
 sky130_fd_sc_hd__a31oi_1 _17792_ (.A1(net3633),
    .A2(_08250_),
    .A3(_08284_),
    .B1(_08623_),
    .Y(_08624_));
 sky130_fd_sc_hd__nor2_4 _17793_ (.A(net3980),
    .B(_08250_),
    .Y(_08625_));
 sky130_fd_sc_hd__a21oi_1 _17794_ (.A1(net3980),
    .A2(_08575_),
    .B1(net3982),
    .Y(_08626_));
 sky130_fd_sc_hd__o21ai_0 _17795_ (.A1(_08625_),
    .A2(_08626_),
    .B1(net397),
    .Y(_08627_));
 sky130_fd_sc_hd__o21ai_0 _17796_ (.A1(_08411_),
    .A2(_08571_),
    .B1(net3982),
    .Y(_08628_));
 sky130_fd_sc_hd__o211ai_1 _17797_ (.A1(net397),
    .A2(_08624_),
    .B1(_08627_),
    .C1(_08628_),
    .Y(_08629_));
 sky130_fd_sc_hd__o311ai_1 _17798_ (.A1(_08250_),
    .A2(_08403_),
    .A3(_08499_),
    .B1(_08452_),
    .C1(net3969),
    .Y(_08630_));
 sky130_fd_sc_hd__o22ai_1 _17799_ (.A1(_08250_),
    .A2(_08426_),
    .B1(_08352_),
    .B2(net3596),
    .Y(_08631_));
 sky130_fd_sc_hd__a21oi_1 _17800_ (.A1(net3960),
    .A2(_08631_),
    .B1(_08336_),
    .Y(_08632_));
 sky130_fd_sc_hd__a21oi_1 _17801_ (.A1(_08630_),
    .A2(_08632_),
    .B1(_08286_),
    .Y(_08633_));
 sky130_fd_sc_hd__o21ai_0 _17802_ (.A1(_08622_),
    .A2(_08629_),
    .B1(_08633_),
    .Y(_08634_));
 sky130_fd_sc_hd__o21ai_0 _17803_ (.A1(net3632),
    .A2(net3978),
    .B1(_08525_),
    .Y(_08635_));
 sky130_fd_sc_hd__a21oi_1 _17804_ (.A1(net397),
    .A2(_08635_),
    .B1(_08295_),
    .Y(_08636_));
 sky130_fd_sc_hd__nor3_2 _17805_ (.A(net3978),
    .B(net3960),
    .C(_08487_),
    .Y(_08637_));
 sky130_fd_sc_hd__o311ai_0 _17806_ (.A1(_08336_),
    .A2(_08636_),
    .A3(_08637_),
    .B1(_08286_),
    .C1(_08622_),
    .Y(_08638_));
 sky130_fd_sc_hd__a21oi_1 _17807_ (.A1(net3633),
    .A2(_08250_),
    .B1(_08301_),
    .Y(_08639_));
 sky130_fd_sc_hd__nor3_1 _17808_ (.A(_08266_),
    .B(_08556_),
    .C(_08639_),
    .Y(_08640_));
 sky130_fd_sc_hd__a31oi_1 _17809_ (.A1(net3981),
    .A2(_08488_),
    .A3(_08620_),
    .B1(_08640_),
    .Y(_08641_));
 sky130_fd_sc_hd__nand3_1 _17810_ (.A(_12093_[0]),
    .B(_08250_),
    .C(net3973),
    .Y(_08642_));
 sky130_fd_sc_hd__a21oi_1 _17811_ (.A1(_12104_[0]),
    .A2(net3962),
    .B1(net3969),
    .Y(_08643_));
 sky130_fd_sc_hd__a21oi_1 _17812_ (.A1(_08642_),
    .A2(_08643_),
    .B1(net3972),
    .Y(_08644_));
 sky130_fd_sc_hd__o41ai_1 _17813_ (.A1(net3960),
    .A2(_08347_),
    .A3(_08470_),
    .A4(_08620_),
    .B1(_08644_),
    .Y(_08645_));
 sky130_fd_sc_hd__o211ai_1 _17814_ (.A1(net3960),
    .A2(net397),
    .B1(net3690),
    .C1(_08279_),
    .Y(_08646_));
 sky130_fd_sc_hd__a31oi_1 _17815_ (.A1(net3960),
    .A2(net397),
    .A3(_08639_),
    .B1(_08646_),
    .Y(_08647_));
 sky130_fd_sc_hd__nand2_1 _17816_ (.A(_08488_),
    .B(_08620_),
    .Y(_08648_));
 sky130_fd_sc_hd__nand2_1 _17817_ (.A(net3980),
    .B(_08648_),
    .Y(_08649_));
 sky130_fd_sc_hd__a21oi_1 _17818_ (.A1(_12102_[0]),
    .A2(_08250_),
    .B1(net3962),
    .Y(_08650_));
 sky130_fd_sc_hd__nand2_1 _17819_ (.A(_08488_),
    .B(_08650_),
    .Y(_08651_));
 sky130_fd_sc_hd__o311ai_0 _17820_ (.A1(net3978),
    .A2(_08473_),
    .A3(_08556_),
    .B1(_08651_),
    .C1(_08244_),
    .Y(_08652_));
 sky130_fd_sc_hd__o21ai_0 _17821_ (.A1(_08647_),
    .A2(_08649_),
    .B1(_08652_),
    .Y(_08653_));
 sky130_fd_sc_hd__a31oi_1 _17822_ (.A1(_08641_),
    .A2(_08645_),
    .A3(_08653_),
    .B1(net3687),
    .Y(_08654_));
 sky130_fd_sc_hd__nand2_2 _17823_ (.A(_08443_),
    .B(_08489_),
    .Y(_08655_));
 sky130_fd_sc_hd__nor3_4 _17824_ (.A(net3981),
    .B(_08244_),
    .C(_08290_),
    .Y(_08656_));
 sky130_fd_sc_hd__nor3_1 _17825_ (.A(_08250_),
    .B(_08412_),
    .C(_08656_),
    .Y(_08657_));
 sky130_fd_sc_hd__a211oi_1 _17826_ (.A1(_08250_),
    .A2(_08655_),
    .B1(_08657_),
    .C1(net3960),
    .Y(_08658_));
 sky130_fd_sc_hd__o21bai_1 _17827_ (.A1(net3633),
    .A2(_08250_),
    .B1_N(_08298_),
    .Y(_08659_));
 sky130_fd_sc_hd__a21oi_1 _17828_ (.A1(net3975),
    .A2(_08659_),
    .B1(_08356_),
    .Y(_08660_));
 sky130_fd_sc_hd__nor3_1 _17829_ (.A(net3968),
    .B(_08658_),
    .C(_08660_),
    .Y(_08661_));
 sky130_fd_sc_hd__a31oi_1 _17830_ (.A1(_08250_),
    .A2(_08415_),
    .A3(_08429_),
    .B1(_08549_),
    .Y(_08662_));
 sky130_fd_sc_hd__nor2_1 _17831_ (.A(net3974),
    .B(_08436_),
    .Y(_08663_));
 sky130_fd_sc_hd__o22ai_1 _17832_ (.A1(net3961),
    .A2(_08662_),
    .B1(_08663_),
    .B2(_08345_),
    .Y(_08664_));
 sky130_fd_sc_hd__o21ai_0 _17833_ (.A1(_08279_),
    .A2(_08664_),
    .B1(_08330_),
    .Y(_08665_));
 sky130_fd_sc_hd__o21ai_0 _17834_ (.A1(_08661_),
    .A2(_08665_),
    .B1(_08365_),
    .Y(_08666_));
 sky130_fd_sc_hd__o2bb2ai_1 _17835_ (.A1_N(_08634_),
    .A2_N(_08638_),
    .B1(_08654_),
    .B2(_08666_),
    .Y(_00068_));
 sky130_fd_sc_hd__o21ai_0 _17836_ (.A1(_12100_[0]),
    .A2(net3963),
    .B1(_08489_),
    .Y(_08667_));
 sky130_fd_sc_hd__nand2_1 _17837_ (.A(_08250_),
    .B(_08667_),
    .Y(_08668_));
 sky130_fd_sc_hd__nand3_1 _17838_ (.A(net3979),
    .B(net3588),
    .C(_08565_),
    .Y(_08669_));
 sky130_fd_sc_hd__a21oi_1 _17839_ (.A1(_08668_),
    .A2(_08669_),
    .B1(net3960),
    .Y(_08670_));
 sky130_fd_sc_hd__o311ai_0 _17840_ (.A1(_08250_),
    .A2(_08371_),
    .A3(net3976),
    .B1(_08498_),
    .C1(net3960),
    .Y(_08671_));
 sky130_fd_sc_hd__nand2_1 _17841_ (.A(net3972),
    .B(_08671_),
    .Y(_08672_));
 sky130_fd_sc_hd__a21oi_1 _17842_ (.A1(_12097_[0]),
    .A2(_08250_),
    .B1(net3976),
    .Y(_08673_));
 sky130_fd_sc_hd__nor2_1 _17843_ (.A(net3596),
    .B(_08377_),
    .Y(_08674_));
 sky130_fd_sc_hd__o221ai_1 _17844_ (.A1(_08308_),
    .A2(_08444_),
    .B1(_08611_),
    .B2(_08250_),
    .C1(net3960),
    .Y(_08675_));
 sky130_fd_sc_hd__o311ai_0 _17845_ (.A1(net3960),
    .A2(_08673_),
    .A3(_08674_),
    .B1(_08675_),
    .C1(_08286_),
    .Y(_08676_));
 sky130_fd_sc_hd__o211ai_1 _17846_ (.A1(_08670_),
    .A2(_08672_),
    .B1(_08393_),
    .C1(_08676_),
    .Y(_08677_));
 sky130_fd_sc_hd__a21oi_1 _17847_ (.A1(_12097_[0]),
    .A2(_08250_),
    .B1(_08625_),
    .Y(_08678_));
 sky130_fd_sc_hd__o21bai_1 _17848_ (.A1(net3975),
    .A2(_08678_),
    .B1_N(_08295_),
    .Y(_08679_));
 sky130_fd_sc_hd__nor2_1 _17849_ (.A(_08336_),
    .B(net3968),
    .Y(_08680_));
 sky130_fd_sc_hd__a21oi_1 _17850_ (.A1(_08371_),
    .A2(_08341_),
    .B1(net3960),
    .Y(_08681_));
 sky130_fd_sc_hd__nand2_1 _17851_ (.A(_08668_),
    .B(_08681_),
    .Y(_08682_));
 sky130_fd_sc_hd__a21oi_1 _17852_ (.A1(_08359_),
    .A2(_08415_),
    .B1(net3978),
    .Y(_08683_));
 sky130_fd_sc_hd__a211oi_2 _17853_ (.A1(net3981),
    .A2(_08341_),
    .B1(_08683_),
    .C1(net3961),
    .Y(_08684_));
 sky130_fd_sc_hd__o21ai_0 _17854_ (.A1(net3633),
    .A2(net3965),
    .B1(net3587),
    .Y(_08685_));
 sky130_fd_sc_hd__a221oi_1 _17855_ (.A1(net3618),
    .A2(_08599_),
    .B1(_08685_),
    .B2(_08250_),
    .C1(net3970),
    .Y(_08686_));
 sky130_fd_sc_hd__nor3_1 _17856_ (.A(_08570_),
    .B(_08684_),
    .C(_08686_),
    .Y(_08687_));
 sky130_fd_sc_hd__a31oi_1 _17857_ (.A1(_08679_),
    .A2(_08680_),
    .A3(_08682_),
    .B1(_08687_),
    .Y(_08688_));
 sky130_fd_sc_hd__nor2_2 _17858_ (.A(_08284_),
    .B(net3964),
    .Y(_08689_));
 sky130_fd_sc_hd__a21oi_2 _17859_ (.A1(net3970),
    .A2(_08312_),
    .B1(_08689_),
    .Y(_08690_));
 sky130_fd_sc_hd__o21ai_0 _17860_ (.A1(_08266_),
    .A2(_08285_),
    .B1(net3981),
    .Y(_08691_));
 sky130_fd_sc_hd__nand4_1 _17861_ (.A(net3689),
    .B(_08377_),
    .C(_08690_),
    .D(_08691_),
    .Y(_08692_));
 sky130_fd_sc_hd__a21oi_1 _17862_ (.A1(_08433_),
    .A2(_08454_),
    .B1(net3965),
    .Y(_08693_));
 sky130_fd_sc_hd__o21ai_0 _17863_ (.A1(_08341_),
    .A2(_08693_),
    .B1(net3981),
    .Y(_08694_));
 sky130_fd_sc_hd__a22o_1 _17864_ (.A1(net3980),
    .A2(_08341_),
    .B1(_08534_),
    .B2(_12100_[0]),
    .X(_08695_));
 sky130_fd_sc_hd__a21oi_1 _17865_ (.A1(net3970),
    .A2(_08695_),
    .B1(_08569_),
    .Y(_08696_));
 sky130_fd_sc_hd__a2111oi_0 _17866_ (.A1(net3597),
    .A2(_08406_),
    .B1(_08448_),
    .C1(net3961),
    .D1(_08349_),
    .Y(_08697_));
 sky130_fd_sc_hd__nand3_1 _17867_ (.A(_08250_),
    .B(_08309_),
    .C(_08307_),
    .Y(_08698_));
 sky130_fd_sc_hd__a21oi_1 _17868_ (.A1(_08405_),
    .A2(_08698_),
    .B1(net3970),
    .Y(_08699_));
 sky130_fd_sc_hd__nor4_1 _17869_ (.A(net3972),
    .B(_08422_),
    .C(_08697_),
    .D(_08699_),
    .Y(_08700_));
 sky130_fd_sc_hd__a31oi_1 _17870_ (.A1(_08692_),
    .A2(_08694_),
    .A3(_08696_),
    .B1(_08700_),
    .Y(_08701_));
 sky130_fd_sc_hd__a21oi_1 _17871_ (.A1(net3689),
    .A2(_08534_),
    .B1(net3970),
    .Y(_08702_));
 sky130_fd_sc_hd__o21ai_0 _17872_ (.A1(net3978),
    .A2(_08656_),
    .B1(_08429_),
    .Y(_08703_));
 sky130_fd_sc_hd__a22o_1 _17873_ (.A1(_08586_),
    .A2(_08702_),
    .B1(_08703_),
    .B2(net3970),
    .X(_08704_));
 sky130_fd_sc_hd__nor3_1 _17874_ (.A(net3978),
    .B(_08544_),
    .C(_08656_),
    .Y(_08705_));
 sky130_fd_sc_hd__a31oi_1 _17875_ (.A1(net3978),
    .A2(_08309_),
    .A3(net3588),
    .B1(_08705_),
    .Y(_08706_));
 sky130_fd_sc_hd__nor2_1 _17876_ (.A(net3980),
    .B(_08341_),
    .Y(_08707_));
 sky130_fd_sc_hd__nor3_1 _17877_ (.A(net3970),
    .B(_08347_),
    .C(_08707_),
    .Y(_08708_));
 sky130_fd_sc_hd__a2111oi_0 _17878_ (.A1(net3970),
    .A2(_08706_),
    .B1(_08708_),
    .C1(net3972),
    .D1(_08336_),
    .Y(_08709_));
 sky130_fd_sc_hd__a31oi_1 _17879_ (.A1(net3972),
    .A2(_08477_),
    .A3(_08704_),
    .B1(_08709_),
    .Y(_08710_));
 sky130_fd_sc_hd__nand4_1 _17880_ (.A(_08677_),
    .B(_08688_),
    .C(_08701_),
    .D(_08710_),
    .Y(_00069_));
 sky130_fd_sc_hd__a211oi_1 _17881_ (.A1(net3963),
    .A2(_08530_),
    .B1(_08656_),
    .C1(_08250_),
    .Y(_08711_));
 sky130_fd_sc_hd__a31oi_1 _17882_ (.A1(_08250_),
    .A2(_08358_),
    .A3(_08565_),
    .B1(_08711_),
    .Y(_08712_));
 sky130_fd_sc_hd__o21ai_0 _17883_ (.A1(_08404_),
    .A2(_08656_),
    .B1(_08250_),
    .Y(_08713_));
 sky130_fd_sc_hd__a21oi_1 _17884_ (.A1(_08593_),
    .A2(_08713_),
    .B1(net3972),
    .Y(_08714_));
 sky130_fd_sc_hd__a21oi_1 _17885_ (.A1(net3972),
    .A2(_08712_),
    .B1(_08714_),
    .Y(_08715_));
 sky130_fd_sc_hd__a21oi_1 _17886_ (.A1(_08238_),
    .A2(_08388_),
    .B1(net3963),
    .Y(_08716_));
 sky130_fd_sc_hd__o21ai_2 _17887_ (.A1(_12111_[0]),
    .A2(net3962),
    .B1(_08286_),
    .Y(_08717_));
 sky130_fd_sc_hd__o21ai_0 _17888_ (.A1(net3632),
    .A2(_08250_),
    .B1(net3963),
    .Y(_08718_));
 sky130_fd_sc_hd__a31oi_1 _17889_ (.A1(_08238_),
    .A2(net3980),
    .A3(_08250_),
    .B1(_08718_),
    .Y(_08719_));
 sky130_fd_sc_hd__o32ai_1 _17890_ (.A1(net3968),
    .A2(_08353_),
    .A3(_08716_),
    .B1(_08717_),
    .B2(_08719_),
    .Y(_08720_));
 sky130_fd_sc_hd__o21ai_0 _17891_ (.A1(net3960),
    .A2(_08720_),
    .B1(_08367_),
    .Y(_08721_));
 sky130_fd_sc_hd__a21oi_1 _17892_ (.A1(net3960),
    .A2(_08715_),
    .B1(_08721_),
    .Y(_08722_));
 sky130_fd_sc_hd__a31oi_1 _17893_ (.A1(net3982),
    .A2(net3980),
    .A3(net3978),
    .B1(_08431_),
    .Y(_08723_));
 sky130_fd_sc_hd__o221ai_2 _17894_ (.A1(_08238_),
    .A2(_08410_),
    .B1(_08723_),
    .B2(_12106_[0]),
    .C1(_08385_),
    .Y(_08724_));
 sky130_fd_sc_hd__nand2_1 _17895_ (.A(net3980),
    .B(net3960),
    .Y(_08725_));
 sky130_fd_sc_hd__o21ai_0 _17896_ (.A1(net3960),
    .A2(_08546_),
    .B1(net3978),
    .Y(_08726_));
 sky130_fd_sc_hd__a21oi_1 _17897_ (.A1(_08725_),
    .A2(_08726_),
    .B1(net3982),
    .Y(_08727_));
 sky130_fd_sc_hd__a221oi_1 _17898_ (.A1(_08625_),
    .A2(_08689_),
    .B1(_08724_),
    .B2(net3970),
    .C1(_08727_),
    .Y(_08728_));
 sky130_fd_sc_hd__nor3_1 _17899_ (.A(_08336_),
    .B(net3972),
    .C(_08728_),
    .Y(_08729_));
 sky130_fd_sc_hd__o32ai_1 _17900_ (.A1(net3978),
    .A2(_08314_),
    .A3(_08426_),
    .B1(_08268_),
    .B2(_12093_[0]),
    .Y(_08730_));
 sky130_fd_sc_hd__a21oi_1 _17901_ (.A1(_12102_[0]),
    .A2(_08250_),
    .B1(net3973),
    .Y(_08731_));
 sky130_fd_sc_hd__a221oi_1 _17902_ (.A1(_12110_[0]),
    .A2(net3973),
    .B1(_08508_),
    .B2(_08731_),
    .C1(net3969),
    .Y(_08732_));
 sky130_fd_sc_hd__a2111oi_0 _17903_ (.A1(net3970),
    .A2(_08730_),
    .B1(_08732_),
    .C1(_08528_),
    .D1(net3972),
    .Y(_08733_));
 sky130_fd_sc_hd__o21ai_0 _17904_ (.A1(net3597),
    .A2(net3970),
    .B1(net3974),
    .Y(_08734_));
 sky130_fd_sc_hd__nand3_1 _17905_ (.A(net3632),
    .B(net3961),
    .C(net3966),
    .Y(_08735_));
 sky130_fd_sc_hd__a211oi_1 _17906_ (.A1(net3982),
    .A2(net3970),
    .B1(_08411_),
    .C1(net3978),
    .Y(_08736_));
 sky130_fd_sc_hd__a31oi_1 _17907_ (.A1(net3978),
    .A2(_08734_),
    .A3(_08735_),
    .B1(_08736_),
    .Y(_08737_));
 sky130_fd_sc_hd__o21ai_0 _17908_ (.A1(net3960),
    .A2(_08316_),
    .B1(_08680_),
    .Y(_08738_));
 sky130_fd_sc_hd__o21ai_0 _17909_ (.A1(_08486_),
    .A2(_08544_),
    .B1(_08250_),
    .Y(_08739_));
 sky130_fd_sc_hd__nand3_1 _17910_ (.A(net3979),
    .B(_08517_),
    .C(_08489_),
    .Y(_08740_));
 sky130_fd_sc_hd__nand3_1 _17911_ (.A(_08494_),
    .B(_08739_),
    .C(_08740_),
    .Y(_08741_));
 sky130_fd_sc_hd__a21oi_1 _17912_ (.A1(net3974),
    .A2(_08530_),
    .B1(net3978),
    .Y(_08742_));
 sky130_fd_sc_hd__nor3_1 _17913_ (.A(_08250_),
    .B(_08431_),
    .C(net3586),
    .Y(_08743_));
 sky130_fd_sc_hd__o221ai_1 _17914_ (.A1(net3618),
    .A2(_08352_),
    .B1(_08742_),
    .B2(_08743_),
    .C1(_08488_),
    .Y(_08744_));
 sky130_fd_sc_hd__o21ai_1 _17915_ (.A1(net3690),
    .A2(_08250_),
    .B1(_08460_),
    .Y(_08745_));
 sky130_fd_sc_hd__o311ai_1 _17916_ (.A1(_12109_[0]),
    .A2(_12118_[0]),
    .A3(net3973),
    .B1(_08285_),
    .C1(_08745_),
    .Y(_08746_));
 sky130_fd_sc_hd__nor4_1 _17917_ (.A(_08250_),
    .B(_08603_),
    .C(_08499_),
    .D(net3586),
    .Y(_08747_));
 sky130_fd_sc_hd__a311oi_1 _17918_ (.A1(_12094_[0]),
    .A2(_08534_),
    .A3(_08433_),
    .B1(_08747_),
    .C1(_08422_),
    .Y(_08748_));
 sky130_fd_sc_hd__nand4_1 _17919_ (.A(_08741_),
    .B(_08744_),
    .C(_08746_),
    .D(_08748_),
    .Y(_08749_));
 sky130_fd_sc_hd__nand2_1 _17920_ (.A(net3961),
    .B(_08522_),
    .Y(_08750_));
 sky130_fd_sc_hd__a21oi_1 _17921_ (.A1(_12100_[0]),
    .A2(net3965),
    .B1(net3586),
    .Y(_08751_));
 sky130_fd_sc_hd__o221ai_1 _17922_ (.A1(_08238_),
    .A2(_08268_),
    .B1(_08751_),
    .B2(net3978),
    .C1(net3970),
    .Y(_08752_));
 sky130_fd_sc_hd__nand4_1 _17923_ (.A(net3971),
    .B(_08393_),
    .C(_08750_),
    .D(_08752_),
    .Y(_08753_));
 sky130_fd_sc_hd__o211ai_1 _17924_ (.A1(_08737_),
    .A2(_08738_),
    .B1(_08749_),
    .C1(_08753_),
    .Y(_08754_));
 sky130_fd_sc_hd__nor4_1 _17925_ (.A(_08722_),
    .B(_08729_),
    .C(_08733_),
    .D(_08754_),
    .Y(_00070_));
 sky130_fd_sc_hd__o221ai_1 _17926_ (.A1(net3596),
    .A2(_08268_),
    .B1(_08439_),
    .B2(_12093_[0]),
    .C1(_08495_),
    .Y(_08755_));
 sky130_fd_sc_hd__nor3_1 _17927_ (.A(_08365_),
    .B(net3960),
    .C(_08755_),
    .Y(_08756_));
 sky130_fd_sc_hd__and3_1 _17928_ (.A(net3978),
    .B(_08358_),
    .C(_08489_),
    .X(_08757_));
 sky130_fd_sc_hd__a2111oi_0 _17929_ (.A1(_08250_),
    .A2(_08555_),
    .B1(_08757_),
    .C1(_08365_),
    .D1(_08284_),
    .Y(_08758_));
 sky130_fd_sc_hd__o21ai_0 _17930_ (.A1(_08406_),
    .A2(_08689_),
    .B1(net3688),
    .Y(_08759_));
 sky130_fd_sc_hd__nor2_1 _17931_ (.A(net3978),
    .B(_08284_),
    .Y(_08760_));
 sky130_fd_sc_hd__a221oi_1 _17932_ (.A1(net3632),
    .A2(_08341_),
    .B1(_08571_),
    .B2(_08656_),
    .C1(_08760_),
    .Y(_08761_));
 sky130_fd_sc_hd__o21ai_1 _17933_ (.A1(net3982),
    .A2(_08759_),
    .B1(_08761_),
    .Y(_08762_));
 sky130_fd_sc_hd__nor2_1 _17934_ (.A(_08335_),
    .B(_08762_),
    .Y(_08763_));
 sky130_fd_sc_hd__nor3_2 _17935_ (.A(_08756_),
    .B(_08758_),
    .C(_08763_),
    .Y(_08764_));
 sky130_fd_sc_hd__nor3_1 _17936_ (.A(net3978),
    .B(_08431_),
    .C(_08585_),
    .Y(_08765_));
 sky130_fd_sc_hd__o21ai_1 _17937_ (.A1(_08268_),
    .A2(_08530_),
    .B1(_08309_),
    .Y(_08766_));
 sky130_fd_sc_hd__o21ai_2 _17938_ (.A1(_08765_),
    .A2(_08766_),
    .B1(_08286_),
    .Y(_08767_));
 sky130_fd_sc_hd__nor2_1 _17939_ (.A(_08286_),
    .B(_08412_),
    .Y(_08768_));
 sky130_fd_sc_hd__nand2_1 _17940_ (.A(_08745_),
    .B(_08768_),
    .Y(_08769_));
 sky130_fd_sc_hd__a21oi_1 _17941_ (.A1(_08767_),
    .A2(_08769_),
    .B1(net3960),
    .Y(_08770_));
 sky130_fd_sc_hd__o221ai_1 _17942_ (.A1(_12092_[0]),
    .A2(_08250_),
    .B1(_08404_),
    .B2(_08618_),
    .C1(_08279_),
    .Y(_08771_));
 sky130_fd_sc_hd__o21ai_0 _17943_ (.A1(_08371_),
    .A2(_08266_),
    .B1(_08498_),
    .Y(_08772_));
 sky130_fd_sc_hd__nor4_1 _17944_ (.A(_08250_),
    .B(_08279_),
    .C(_08472_),
    .D(_08473_),
    .Y(_08773_));
 sky130_fd_sc_hd__a31oi_1 _17945_ (.A1(_08250_),
    .A2(_08286_),
    .A3(_08772_),
    .B1(_08773_),
    .Y(_08774_));
 sky130_fd_sc_hd__and3_1 _17946_ (.A(net3960),
    .B(_08771_),
    .C(_08774_),
    .X(_08775_));
 sky130_fd_sc_hd__o21ai_0 _17947_ (.A1(_12093_[0]),
    .A2(net3978),
    .B1(net3962),
    .Y(_08776_));
 sky130_fd_sc_hd__a21oi_1 _17948_ (.A1(_12102_[0]),
    .A2(net3978),
    .B1(_08776_),
    .Y(_08777_));
 sky130_fd_sc_hd__nor2_1 _17949_ (.A(_12118_[0]),
    .B(net3962),
    .Y(_08778_));
 sky130_fd_sc_hd__a21oi_1 _17950_ (.A1(_08308_),
    .A2(_08461_),
    .B1(_08250_),
    .Y(_08779_));
 sky130_fd_sc_hd__o21ai_0 _17951_ (.A1(_08479_),
    .A2(_08779_),
    .B1(_08488_),
    .Y(_08780_));
 sky130_fd_sc_hd__nand3_1 _17952_ (.A(_12094_[0]),
    .B(_08250_),
    .C(net397),
    .Y(_08781_));
 sky130_fd_sc_hd__o21ai_0 _17953_ (.A1(_12104_[0]),
    .A2(_08290_),
    .B1(_08781_),
    .Y(_08782_));
 sky130_fd_sc_hd__nor2_1 _17954_ (.A(_12097_[0]),
    .B(_08250_),
    .Y(_08783_));
 sky130_fd_sc_hd__o21ai_0 _17955_ (.A1(_08502_),
    .A2(_08783_),
    .B1(net3976),
    .Y(_08784_));
 sky130_fd_sc_hd__a21oi_1 _17956_ (.A1(_08388_),
    .A2(_08312_),
    .B1(_08603_),
    .Y(_08785_));
 sky130_fd_sc_hd__a221oi_1 _17957_ (.A1(_08285_),
    .A2(_08782_),
    .B1(_08784_),
    .B2(_08785_),
    .C1(_08335_),
    .Y(_08786_));
 sky130_fd_sc_hd__o311ai_0 _17958_ (.A1(_08556_),
    .A2(_08777_),
    .A3(_08778_),
    .B1(_08780_),
    .C1(_08786_),
    .Y(_08787_));
 sky130_fd_sc_hd__o311ai_0 _17959_ (.A1(_08365_),
    .A2(_08770_),
    .A3(_08775_),
    .B1(_08787_),
    .C1(net3687),
    .Y(_08788_));
 sky130_fd_sc_hd__o21ai_0 _17960_ (.A1(_08534_),
    .A2(_08597_),
    .B1(_08238_),
    .Y(_08789_));
 sky130_fd_sc_hd__a21oi_1 _17961_ (.A1(_08352_),
    .A2(_08358_),
    .B1(_08238_),
    .Y(_08790_));
 sky130_fd_sc_hd__o21ai_0 _17962_ (.A1(_08347_),
    .A2(_08790_),
    .B1(net3960),
    .Y(_08791_));
 sky130_fd_sc_hd__o21ai_0 _17963_ (.A1(net3689),
    .A2(_08268_),
    .B1(_08316_),
    .Y(_08792_));
 sky130_fd_sc_hd__nand2_1 _17964_ (.A(net3970),
    .B(_08792_),
    .Y(_08793_));
 sky130_fd_sc_hd__a31oi_2 _17965_ (.A1(_08789_),
    .A2(_08791_),
    .A3(_08793_),
    .B1(_08528_),
    .Y(_08794_));
 sky130_fd_sc_hd__a21oi_1 _17966_ (.A1(net3688),
    .A2(_08534_),
    .B1(_08426_),
    .Y(_08795_));
 sky130_fd_sc_hd__nand2_1 _17967_ (.A(_12092_[0]),
    .B(_08599_),
    .Y(_08796_));
 sky130_fd_sc_hd__o2111ai_1 _17968_ (.A1(net3982),
    .A2(_08795_),
    .B1(_08796_),
    .C1(net3969),
    .D1(_08495_),
    .Y(_08797_));
 sky130_fd_sc_hd__o221ai_1 _17969_ (.A1(_12102_[0]),
    .A2(_08377_),
    .B1(_08655_),
    .B2(_08250_),
    .C1(net3960),
    .Y(_08798_));
 sky130_fd_sc_hd__a21oi_1 _17970_ (.A1(_08797_),
    .A2(_08798_),
    .B1(_08336_),
    .Y(_08799_));
 sky130_fd_sc_hd__o21ai_0 _17971_ (.A1(_08794_),
    .A2(_08799_),
    .B1(net3967),
    .Y(_08800_));
 sky130_fd_sc_hd__o311ai_2 _17972_ (.A1(net3687),
    .A2(net3967),
    .A3(_08764_),
    .B1(_08788_),
    .C1(_08800_),
    .Y(_00071_));
 sky130_fd_sc_hd__xnor2_2 _17973_ (.A(\sa11_sr[7] ),
    .B(\sa21_sr[7] ),
    .Y(_08801_));
 sky130_fd_sc_hd__xor3_1 _17974_ (.A(\sa21_sr[1] ),
    .B(\sa30_sub[1] ),
    .C(net4227),
    .X(_08802_));
 sky130_fd_sc_hd__xnor3_1 _17975_ (.A(_06489_),
    .B(_08801_),
    .C(_08802_),
    .X(_08803_));
 sky130_fd_sc_hd__mux2i_2 _17976_ (.A0(\text_in_r[81] ),
    .A1(_08803_),
    .S(net4117),
    .Y(_08804_));
 sky130_fd_sc_hd__xor2_4 _17977_ (.A(net4154),
    .B(_08804_),
    .X(_08805_));
 sky130_fd_sc_hd__inv_12 _17978_ (.A(_08805_),
    .Y(_08806_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_684 ();
 sky130_fd_sc_hd__xor2_1 _17981_ (.A(\sa01_sr[0] ),
    .B(\sa30_sub[0] ),
    .X(_08808_));
 sky130_fd_sc_hd__xnor3_1 _17982_ (.A(net4206),
    .B(_08801_),
    .C(_08808_),
    .X(_08809_));
 sky130_fd_sc_hd__mux2i_2 _17983_ (.A0(\text_in_r[80] ),
    .A1(_08809_),
    .S(_05879_),
    .Y(_08810_));
 sky130_fd_sc_hd__xor2_4 _17984_ (.A(net4155),
    .B(_08810_),
    .X(_08811_));
 sky130_fd_sc_hd__inv_16 _17985_ (.A(_08811_),
    .Y(_08812_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_682 ();
 sky130_fd_sc_hd__xnor3_1 _17988_ (.A(\sa21_sr[1] ),
    .B(\sa21_sr[2] ),
    .C(net4226),
    .X(_08814_));
 sky130_fd_sc_hd__xor2_1 _17989_ (.A(_06497_),
    .B(_08814_),
    .X(_08815_));
 sky130_fd_sc_hd__mux2i_2 _17990_ (.A0(\text_in_r[82] ),
    .A1(_08815_),
    .S(net4117),
    .Y(_08816_));
 sky130_fd_sc_hd__xnor2_4 _17991_ (.A(\u0.w[1][18] ),
    .B(_08816_),
    .Y(_08817_));
 sky130_fd_sc_hd__clkinv_16 _17992_ (.A(_08817_),
    .Y(_08818_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_675 ();
 sky130_fd_sc_hd__xnor3_1 _18000_ (.A(\sa21_sr[4] ),
    .B(\sa30_sub[5] ),
    .C(\sa01_sr[5] ),
    .X(_08823_));
 sky130_fd_sc_hd__xor2_1 _18001_ (.A(\sa11_sr[4] ),
    .B(net4203),
    .X(_08824_));
 sky130_fd_sc_hd__xnor2_2 _18002_ (.A(_08823_),
    .B(_08824_),
    .Y(_08825_));
 sky130_fd_sc_hd__mux2i_4 _18003_ (.A0(\text_in_r[85] ),
    .A1(_08825_),
    .S(net4120),
    .Y(_08826_));
 sky130_fd_sc_hd__xnor2_4 _18004_ (.A(\u0.w[1][21] ),
    .B(_08826_),
    .Y(_08827_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_674 ();
 sky130_fd_sc_hd__nor2b_1 _18006_ (.A(net4230),
    .B_N(\u0.w[1][19] ),
    .Y(_08829_));
 sky130_fd_sc_hd__nor2_1 _18007_ (.A(\u0.w[1][19] ),
    .B(net4230),
    .Y(_08830_));
 sky130_fd_sc_hd__xnor3_1 _18008_ (.A(\sa21_sr[2] ),
    .B(\sa30_sub[3] ),
    .C(\sa21_sr[7] ),
    .X(_08831_));
 sky130_fd_sc_hd__xnor2_1 _18009_ (.A(\sa21_sr[3] ),
    .B(net4225),
    .Y(_08832_));
 sky130_fd_sc_hd__xnor3_1 _18010_ (.A(_06528_),
    .B(_08831_),
    .C(_08832_),
    .X(_08833_));
 sky130_fd_sc_hd__mux2_8 _18011_ (.A0(_08829_),
    .A1(_08830_),
    .S(_08833_),
    .X(_08834_));
 sky130_fd_sc_hd__nand2_1 _18012_ (.A(\u0.w[1][19] ),
    .B(net4230),
    .Y(_08835_));
 sky130_fd_sc_hd__nand3b_1 _18013_ (.A_N(\u0.w[1][19] ),
    .B(net4230),
    .C(\text_in_r[83] ),
    .Y(_08836_));
 sky130_fd_sc_hd__o21ai_4 _18014_ (.A1(\text_in_r[83] ),
    .A2(_08835_),
    .B1(_08836_),
    .Y(_08837_));
 sky130_fd_sc_hd__or2_4 _18015_ (.A(_08834_),
    .B(_08837_),
    .X(_08838_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_673 ();
 sky130_fd_sc_hd__nor3_4 _18017_ (.A(net3958),
    .B(net3683),
    .C(_08838_),
    .Y(_08840_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_672 ();
 sky130_fd_sc_hd__nor2_4 _18019_ (.A(_08834_),
    .B(_08837_),
    .Y(_08842_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_671 ();
 sky130_fd_sc_hd__o21ai_0 _18021_ (.A1(_12126_[0]),
    .A2(net3947),
    .B1(net3956),
    .Y(_08844_));
 sky130_fd_sc_hd__xnor2_1 _18022_ (.A(\sa21_sr[3] ),
    .B(\sa30_sub[4] ),
    .Y(_08845_));
 sky130_fd_sc_hd__xnor3_1 _18023_ (.A(\sa11_sr[3] ),
    .B(net4204),
    .C(\sa01_sr[4] ),
    .X(_08846_));
 sky130_fd_sc_hd__xnor3_1 _18024_ (.A(_08801_),
    .B(_08845_),
    .C(_08846_),
    .X(_08847_));
 sky130_fd_sc_hd__mux2i_4 _18025_ (.A0(\text_in_r[84] ),
    .A1(_08847_),
    .S(net4120),
    .Y(_08848_));
 sky130_fd_sc_hd__xnor2_4 _18026_ (.A(\u0.w[1][20] ),
    .B(_08848_),
    .Y(_08849_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_670 ();
 sky130_fd_sc_hd__o21ai_0 _18028_ (.A1(_08840_),
    .A2(_08844_),
    .B1(_08849_),
    .Y(_08851_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_669 ();
 sky130_fd_sc_hd__nand2_8 _18030_ (.A(_08818_),
    .B(net3946),
    .Y(_08853_));
 sky130_fd_sc_hd__nor2_1 _18031_ (.A(_12132_[0]),
    .B(_08853_),
    .Y(_08854_));
 sky130_fd_sc_hd__nor2_4 _18032_ (.A(_12126_[0]),
    .B(_08838_),
    .Y(_08855_));
 sky130_fd_sc_hd__nor3_4 _18033_ (.A(net3958),
    .B(net3683),
    .C(net3946),
    .Y(_08856_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_668 ();
 sky130_fd_sc_hd__nor2_1 _18035_ (.A(net3956),
    .B(_08842_),
    .Y(_08858_));
 sky130_fd_sc_hd__nand2_1 _18036_ (.A(_12134_[0]),
    .B(net3681),
    .Y(_08859_));
 sky130_fd_sc_hd__xor2_4 _18037_ (.A(\u0.w[1][20] ),
    .B(_08848_),
    .X(_08860_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_667 ();
 sky130_fd_sc_hd__o311ai_0 _18039_ (.A1(_08818_),
    .A2(_08855_),
    .A3(_08856_),
    .B1(_08859_),
    .C1(net3941),
    .Y(_08862_));
 sky130_fd_sc_hd__o21ai_0 _18040_ (.A1(_08851_),
    .A2(_08854_),
    .B1(_08862_),
    .Y(_08863_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_663 ();
 sky130_fd_sc_hd__nand2_1 _18045_ (.A(_12124_[0]),
    .B(_08838_),
    .Y(_08868_));
 sky130_fd_sc_hd__nand2_1 _18046_ (.A(net3956),
    .B(_08868_),
    .Y(_08869_));
 sky130_fd_sc_hd__nor2_1 _18047_ (.A(_08840_),
    .B(_08869_),
    .Y(_08870_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_661 ();
 sky130_fd_sc_hd__nor2_4 _18050_ (.A(_12126_[0]),
    .B(_12129_[0]),
    .Y(_08873_));
 sky130_fd_sc_hd__nor2_2 _18051_ (.A(_08812_),
    .B(net3947),
    .Y(_08874_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_660 ();
 sky130_fd_sc_hd__a211oi_1 _18053_ (.A1(net3947),
    .A2(_08873_),
    .B1(_08874_),
    .C1(net3956),
    .Y(_08876_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_659 ();
 sky130_fd_sc_hd__o21ai_0 _18055_ (.A1(_08870_),
    .A2(_08876_),
    .B1(net3941),
    .Y(_08878_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_654 ();
 sky130_fd_sc_hd__nand2_4 _18061_ (.A(_12125_[0]),
    .B(_08818_),
    .Y(_08884_));
 sky130_fd_sc_hd__nor2_1 _18062_ (.A(_12145_[0]),
    .B(net3948),
    .Y(_08885_));
 sky130_fd_sc_hd__a21oi_1 _18063_ (.A1(net3948),
    .A2(_08884_),
    .B1(_08885_),
    .Y(_08886_));
 sky130_fd_sc_hd__a21oi_1 _18064_ (.A1(net3945),
    .A2(_08886_),
    .B1(net3955),
    .Y(_08887_));
 sky130_fd_sc_hd__xnor2_1 _18065_ (.A(\sa21_sr[6] ),
    .B(net4186),
    .Y(_08888_));
 sky130_fd_sc_hd__xnor3_1 _18066_ (.A(\sa01_sr[7] ),
    .B(\sa11_sr[6] ),
    .C(\sa21_sr[7] ),
    .X(_08889_));
 sky130_fd_sc_hd__xor2_1 _18067_ (.A(_08888_),
    .B(_08889_),
    .X(_08890_));
 sky130_fd_sc_hd__mux2i_4 _18068_ (.A0(\text_in_r[87] ),
    .A1(_08890_),
    .S(net4120),
    .Y(_08891_));
 sky130_fd_sc_hd__xnor2_4 _18069_ (.A(\u0.w[1][23] ),
    .B(_08891_),
    .Y(_08892_));
 sky130_fd_sc_hd__xor2_1 _18070_ (.A(net4203),
    .B(\sa01_sr[6] ),
    .X(_08893_));
 sky130_fd_sc_hd__xnor2_1 _18071_ (.A(_06596_),
    .B(_08893_),
    .Y(_08894_));
 sky130_fd_sc_hd__mux2i_4 _18072_ (.A0(\text_in_r[86] ),
    .A1(_08894_),
    .S(net4120),
    .Y(_08895_));
 sky130_fd_sc_hd__xor2_2 _18073_ (.A(net4152),
    .B(_08895_),
    .X(_08896_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_653 ();
 sky130_fd_sc_hd__nand2_2 _18075_ (.A(_08892_),
    .B(net3938),
    .Y(_08898_));
 sky130_fd_sc_hd__a221oi_1 _18076_ (.A1(net3955),
    .A2(_08863_),
    .B1(_08878_),
    .B2(_08887_),
    .C1(_08898_),
    .Y(_08899_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_652 ();
 sky130_fd_sc_hd__nand2_4 _18078_ (.A(net3959),
    .B(net3946),
    .Y(_08901_));
 sky130_fd_sc_hd__nand2_1 _18079_ (.A(_08812_),
    .B(_08838_),
    .Y(_08902_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_651 ();
 sky130_fd_sc_hd__nor2_1 _18081_ (.A(_12132_[0]),
    .B(net3947),
    .Y(_08904_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_650 ();
 sky130_fd_sc_hd__nor2_4 _18083_ (.A(_12125_[0]),
    .B(net3952),
    .Y(_08906_));
 sky130_fd_sc_hd__nor3_1 _18084_ (.A(net3956),
    .B(_08904_),
    .C(_08906_),
    .Y(_08907_));
 sky130_fd_sc_hd__a31oi_1 _18085_ (.A1(net3956),
    .A2(_08901_),
    .A3(net3615),
    .B1(_08907_),
    .Y(_08908_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_649 ();
 sky130_fd_sc_hd__o21ai_4 _18087_ (.A1(net3958),
    .A2(net3957),
    .B1(_08838_),
    .Y(_08910_));
 sky130_fd_sc_hd__nor2_2 _18088_ (.A(_12129_[0]),
    .B(_08838_),
    .Y(_08911_));
 sky130_fd_sc_hd__a221o_4 _18089_ (.A1(net3957),
    .A2(_08858_),
    .B1(_08910_),
    .B2(net3956),
    .C1(_08911_),
    .X(_08912_));
 sky130_fd_sc_hd__nor2_1 _18090_ (.A(net3955),
    .B(_08912_),
    .Y(_08913_));
 sky130_fd_sc_hd__a21oi_1 _18091_ (.A1(net3955),
    .A2(_08908_),
    .B1(_08913_),
    .Y(_08914_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_648 ();
 sky130_fd_sc_hd__xor2_4 _18093_ (.A(\u0.w[1][23] ),
    .B(_08891_),
    .X(_08916_));
 sky130_fd_sc_hd__nor2_4 _18094_ (.A(_08916_),
    .B(_08896_),
    .Y(_08917_));
 sky130_fd_sc_hd__nand2_2 _18095_ (.A(net3941),
    .B(_08917_),
    .Y(_08918_));
 sky130_fd_sc_hd__nor2_4 _18096_ (.A(net3957),
    .B(_08818_),
    .Y(_08919_));
 sky130_fd_sc_hd__a21oi_1 _18097_ (.A1(net3959),
    .A2(net3957),
    .B1(_08919_),
    .Y(_08920_));
 sky130_fd_sc_hd__xnor2_1 _18098_ (.A(net3946),
    .B(_08920_),
    .Y(_08921_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_647 ();
 sky130_fd_sc_hd__nand2_8 _18100_ (.A(_08806_),
    .B(_08812_),
    .Y(_08923_));
 sky130_fd_sc_hd__nand2_2 _18101_ (.A(net3946),
    .B(_08923_),
    .Y(_08924_));
 sky130_fd_sc_hd__nand2b_1 _18102_ (.A_N(_12124_[0]),
    .B(net3951),
    .Y(_08925_));
 sky130_fd_sc_hd__and2_4 _18103_ (.A(_12125_[0]),
    .B(net3950),
    .X(_08926_));
 sky130_fd_sc_hd__nor3_1 _18104_ (.A(_08818_),
    .B(_08904_),
    .C(_08926_),
    .Y(_08927_));
 sky130_fd_sc_hd__a311oi_1 _18105_ (.A1(_08818_),
    .A2(_08924_),
    .A3(_08925_),
    .B1(net3945),
    .C1(_08927_),
    .Y(_08928_));
 sky130_fd_sc_hd__a21oi_1 _18106_ (.A1(net3945),
    .A2(_08921_),
    .B1(_08928_),
    .Y(_08929_));
 sky130_fd_sc_hd__xor2_4 _18107_ (.A(\u0.w[1][21] ),
    .B(_08826_),
    .X(_08930_));
 sky130_fd_sc_hd__nor2_1 _18108_ (.A(_08892_),
    .B(_08930_),
    .Y(_08931_));
 sky130_fd_sc_hd__nand2_1 _18109_ (.A(net3938),
    .B(net3680),
    .Y(_08932_));
 sky130_fd_sc_hd__nor2_2 _18110_ (.A(net3684),
    .B(net3956),
    .Y(_08933_));
 sky130_fd_sc_hd__nand2_8 _18111_ (.A(net3958),
    .B(_08838_),
    .Y(_08934_));
 sky130_fd_sc_hd__nand2_8 _18112_ (.A(net3956),
    .B(_08838_),
    .Y(_08935_));
 sky130_fd_sc_hd__xnor2_4 _18113_ (.A(net4152),
    .B(_08895_),
    .Y(_08936_));
 sky130_fd_sc_hd__o311ai_0 _18114_ (.A1(_12129_[0]),
    .A2(_08849_),
    .A3(_08935_),
    .B1(_08931_),
    .C1(_08936_),
    .Y(_08937_));
 sky130_fd_sc_hd__a31oi_1 _18115_ (.A1(net3941),
    .A2(_08933_),
    .A3(_08934_),
    .B1(_08937_),
    .Y(_08938_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_646 ();
 sky130_fd_sc_hd__nor2_4 _18117_ (.A(_12138_[0]),
    .B(net3950),
    .Y(_08940_));
 sky130_fd_sc_hd__nand2_4 _18118_ (.A(net3685),
    .B(net3950),
    .Y(_08941_));
 sky130_fd_sc_hd__nand3b_1 _18119_ (.A_N(_08940_),
    .B(_08818_),
    .C(_08941_),
    .Y(_08942_));
 sky130_fd_sc_hd__nor2_4 _18120_ (.A(_08818_),
    .B(net3946),
    .Y(_08943_));
 sky130_fd_sc_hd__nand2_1 _18121_ (.A(_12125_[0]),
    .B(_08943_),
    .Y(_08944_));
 sky130_fd_sc_hd__nand2_8 _18122_ (.A(_08812_),
    .B(net3950),
    .Y(_08945_));
 sky130_fd_sc_hd__nand4_1 _18123_ (.A(_08849_),
    .B(_08942_),
    .C(_08944_),
    .D(_08945_),
    .Y(_08946_));
 sky130_fd_sc_hd__nand2_8 _18124_ (.A(_12125_[0]),
    .B(_08838_),
    .Y(_08947_));
 sky130_fd_sc_hd__nand2_4 _18125_ (.A(_12134_[0]),
    .B(net3950),
    .Y(_08948_));
 sky130_fd_sc_hd__and3_1 _18126_ (.A(net3956),
    .B(_08947_),
    .C(_08948_),
    .X(_08949_));
 sky130_fd_sc_hd__nor2_4 _18127_ (.A(_12129_[0]),
    .B(_08853_),
    .Y(_08950_));
 sky130_fd_sc_hd__nand2_4 _18128_ (.A(net3937),
    .B(_08917_),
    .Y(_08951_));
 sky130_fd_sc_hd__a2111oi_0 _18129_ (.A1(net3939),
    .A2(_08912_),
    .B1(_08949_),
    .C1(_08950_),
    .D1(_08951_),
    .Y(_08952_));
 sky130_fd_sc_hd__nor2_4 _18130_ (.A(_12129_[0]),
    .B(net3950),
    .Y(_08953_));
 sky130_fd_sc_hd__o21ai_0 _18131_ (.A1(_08855_),
    .A2(_08953_),
    .B1(net3956),
    .Y(_08954_));
 sky130_fd_sc_hd__nor2_4 _18132_ (.A(net3956),
    .B(_08838_),
    .Y(_08955_));
 sky130_fd_sc_hd__nand2_1 _18133_ (.A(_12124_[0]),
    .B(_08955_),
    .Y(_08956_));
 sky130_fd_sc_hd__nor2_4 _18134_ (.A(_08930_),
    .B(_08860_),
    .Y(_08957_));
 sky130_fd_sc_hd__and4_1 _18135_ (.A(_08917_),
    .B(_08954_),
    .C(_08956_),
    .D(_08957_),
    .X(_08958_));
 sky130_fd_sc_hd__a211oi_1 _18136_ (.A1(_08938_),
    .A2(_08946_),
    .B1(net3571),
    .C1(_08958_),
    .Y(_08959_));
 sky130_fd_sc_hd__o221ai_1 _18137_ (.A1(_08914_),
    .A2(_08918_),
    .B1(_08929_),
    .B2(_08932_),
    .C1(_08959_),
    .Y(_08960_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_645 ();
 sky130_fd_sc_hd__nand2_4 _18139_ (.A(_12138_[0]),
    .B(net3954),
    .Y(_08962_));
 sky130_fd_sc_hd__a32oi_1 _18140_ (.A1(net3956),
    .A2(_08941_),
    .A3(_08962_),
    .B1(_08901_),
    .B2(_08933_),
    .Y(_08963_));
 sky130_fd_sc_hd__nand2_1 _18141_ (.A(net3959),
    .B(_08818_),
    .Y(_08964_));
 sky130_fd_sc_hd__nor2_4 _18142_ (.A(_12125_[0]),
    .B(net3956),
    .Y(_08965_));
 sky130_fd_sc_hd__a221o_1 _18143_ (.A1(_08926_),
    .A2(_08964_),
    .B1(_08965_),
    .B2(_08901_),
    .C1(_08936_),
    .X(_08966_));
 sky130_fd_sc_hd__o21ai_0 _18144_ (.A1(net3938),
    .A2(_08963_),
    .B1(_08966_),
    .Y(_08967_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_644 ();
 sky130_fd_sc_hd__nand2_2 _18146_ (.A(_08916_),
    .B(net3937),
    .Y(_08969_));
 sky130_fd_sc_hd__nor2_4 _18147_ (.A(_08818_),
    .B(_08838_),
    .Y(_08970_));
 sky130_fd_sc_hd__o21ai_0 _18148_ (.A1(_08970_),
    .A2(net3681),
    .B1(_12124_[0]),
    .Y(_08971_));
 sky130_fd_sc_hd__nor2_2 _18149_ (.A(_12125_[0]),
    .B(_08935_),
    .Y(_08972_));
 sky130_fd_sc_hd__a21oi_1 _18150_ (.A1(_12132_[0]),
    .A2(_08955_),
    .B1(_08972_),
    .Y(_08973_));
 sky130_fd_sc_hd__nand3_1 _18151_ (.A(net3683),
    .B(net3956),
    .C(net3953),
    .Y(_08974_));
 sky130_fd_sc_hd__a21oi_1 _18152_ (.A1(_08853_),
    .A2(_08974_),
    .B1(net3958),
    .Y(_08975_));
 sky130_fd_sc_hd__nand2_2 _18153_ (.A(net3956),
    .B(net3946),
    .Y(_08976_));
 sky130_fd_sc_hd__nor2_2 _18154_ (.A(_12126_[0]),
    .B(_08976_),
    .Y(_08977_));
 sky130_fd_sc_hd__a2111oi_2 _18155_ (.A1(net3957),
    .A2(net3681),
    .B1(_08975_),
    .C1(_08977_),
    .D1(net3938),
    .Y(_08978_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_643 ();
 sky130_fd_sc_hd__a311oi_1 _18157_ (.A1(net3938),
    .A2(_08971_),
    .A3(_08973_),
    .B1(_08978_),
    .C1(net3945),
    .Y(_08980_));
 sky130_fd_sc_hd__a211oi_1 _18158_ (.A1(net3945),
    .A2(_08967_),
    .B1(_08969_),
    .C1(_08980_),
    .Y(_08981_));
 sky130_fd_sc_hd__or3_1 _18159_ (.A(_08899_),
    .B(_08960_),
    .C(_08981_),
    .X(_00072_));
 sky130_fd_sc_hd__nand2b_4 _18160_ (.A_N(_12125_[0]),
    .B(net3954),
    .Y(_08982_));
 sky130_fd_sc_hd__nand3_1 _18161_ (.A(_08806_),
    .B(_08812_),
    .C(net3946),
    .Y(_08983_));
 sky130_fd_sc_hd__a21oi_1 _18162_ (.A1(_08982_),
    .A2(net3614),
    .B1(net3682),
    .Y(_08984_));
 sky130_fd_sc_hd__nand2_1 _18163_ (.A(net3957),
    .B(_08955_),
    .Y(_08985_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_642 ();
 sky130_fd_sc_hd__nand3b_1 _18165_ (.A_N(_08984_),
    .B(_08985_),
    .C(net3939),
    .Y(_08987_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_639 ();
 sky130_fd_sc_hd__nand2_2 _18169_ (.A(_12126_[0]),
    .B(net3950),
    .Y(_08991_));
 sky130_fd_sc_hd__nand3_1 _18170_ (.A(net3682),
    .B(_08991_),
    .C(_08910_),
    .Y(_08992_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_638 ();
 sky130_fd_sc_hd__nand2_4 _18172_ (.A(_12138_[0]),
    .B(net3950),
    .Y(_08994_));
 sky130_fd_sc_hd__nand3_1 _18173_ (.A(net3956),
    .B(_08982_),
    .C(_08994_),
    .Y(_08995_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_636 ();
 sky130_fd_sc_hd__a311oi_1 _18176_ (.A1(net3943),
    .A2(_08992_),
    .A3(_08995_),
    .B1(_08827_),
    .C1(net3938),
    .Y(_08998_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_635 ();
 sky130_fd_sc_hd__nand2_8 _18178_ (.A(net3686),
    .B(net3952),
    .Y(_09000_));
 sky130_fd_sc_hd__nor2_2 _18179_ (.A(_08812_),
    .B(_08818_),
    .Y(_09001_));
 sky130_fd_sc_hd__nor2_4 _18180_ (.A(net3957),
    .B(net3956),
    .Y(_09002_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_634 ();
 sky130_fd_sc_hd__a21oi_1 _18182_ (.A1(_12124_[0]),
    .A2(_08818_),
    .B1(_09001_),
    .Y(_09004_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_632 ();
 sky130_fd_sc_hd__o32ai_1 _18185_ (.A1(_09000_),
    .A2(_09001_),
    .A3(_09002_),
    .B1(_09004_),
    .B2(net3951),
    .Y(_09007_));
 sky130_fd_sc_hd__a21oi_1 _18186_ (.A1(_12132_[0]),
    .A2(_08818_),
    .B1(net3951),
    .Y(_09008_));
 sky130_fd_sc_hd__o21ai_0 _18187_ (.A1(_08818_),
    .A2(_08923_),
    .B1(_09008_),
    .Y(_09009_));
 sky130_fd_sc_hd__o311a_1 _18188_ (.A1(_12148_[0]),
    .A2(net3955),
    .A3(net3948),
    .B1(_09009_),
    .C1(_08860_),
    .X(_09010_));
 sky130_fd_sc_hd__a21oi_2 _18189_ (.A1(_08957_),
    .A2(_09007_),
    .B1(_09010_),
    .Y(_09011_));
 sky130_fd_sc_hd__o2bb2ai_2 _18190_ (.A1_N(_08987_),
    .A2_N(_08998_),
    .B1(_08936_),
    .B2(_09011_),
    .Y(_09012_));
 sky130_fd_sc_hd__or3_4 _18191_ (.A(_12126_[0]),
    .B(_08834_),
    .C(_08837_),
    .X(_09013_));
 sky130_fd_sc_hd__a21oi_1 _18192_ (.A1(_08945_),
    .A2(_08947_),
    .B1(net3956),
    .Y(_09014_));
 sky130_fd_sc_hd__a31oi_1 _18193_ (.A1(net3956),
    .A2(_08868_),
    .A3(_09013_),
    .B1(_09014_),
    .Y(_09015_));
 sky130_fd_sc_hd__nor2_4 _18194_ (.A(net3957),
    .B(_08838_),
    .Y(_09016_));
 sky130_fd_sc_hd__o21ai_0 _18195_ (.A1(_08953_),
    .A2(_09016_),
    .B1(net3956),
    .Y(_09017_));
 sky130_fd_sc_hd__o211ai_1 _18196_ (.A1(_12124_[0]),
    .A2(_08838_),
    .B1(_09000_),
    .C1(_08818_),
    .Y(_09018_));
 sky130_fd_sc_hd__nand2_2 _18197_ (.A(_08827_),
    .B(net3939),
    .Y(_09019_));
 sky130_fd_sc_hd__a21oi_1 _18198_ (.A1(_09017_),
    .A2(_09018_),
    .B1(_09019_),
    .Y(_09020_));
 sky130_fd_sc_hd__a21oi_1 _18199_ (.A1(_08957_),
    .A2(_09015_),
    .B1(_09020_),
    .Y(_09021_));
 sky130_fd_sc_hd__nand3_2 _18200_ (.A(_08818_),
    .B(_08934_),
    .C(_08941_),
    .Y(_09022_));
 sky130_fd_sc_hd__or3_1 _18201_ (.A(_08818_),
    .B(_08953_),
    .C(_09016_),
    .X(_09023_));
 sky130_fd_sc_hd__nor2_4 _18202_ (.A(_08827_),
    .B(net3939),
    .Y(_09024_));
 sky130_fd_sc_hd__a41oi_1 _18203_ (.A1(net3938),
    .A2(_09022_),
    .A3(_09023_),
    .A4(_09024_),
    .B1(_08892_),
    .Y(_09025_));
 sky130_fd_sc_hd__o21ai_2 _18204_ (.A1(net3938),
    .A2(_09021_),
    .B1(_09025_),
    .Y(_09026_));
 sky130_fd_sc_hd__nand2_1 _18205_ (.A(net3682),
    .B(_08962_),
    .Y(_09027_));
 sky130_fd_sc_hd__o211ai_1 _18206_ (.A1(net3685),
    .A2(_08935_),
    .B1(net3614),
    .C1(_09027_),
    .Y(_09028_));
 sky130_fd_sc_hd__nand2_8 _18207_ (.A(_12124_[0]),
    .B(net3949),
    .Y(_09029_));
 sky130_fd_sc_hd__nor2_4 _18208_ (.A(net3684),
    .B(net3954),
    .Y(_09030_));
 sky130_fd_sc_hd__nor3_1 _18209_ (.A(net3956),
    .B(_09030_),
    .C(_08953_),
    .Y(_09031_));
 sky130_fd_sc_hd__a311oi_1 _18210_ (.A1(net3956),
    .A2(_08947_),
    .A3(_09029_),
    .B1(_09031_),
    .C1(_08827_),
    .Y(_09032_));
 sky130_fd_sc_hd__a211oi_1 _18211_ (.A1(_08827_),
    .A2(_09028_),
    .B1(_09032_),
    .C1(net3939),
    .Y(_09033_));
 sky130_fd_sc_hd__nand2_4 _18212_ (.A(_08930_),
    .B(net3939),
    .Y(_09034_));
 sky130_fd_sc_hd__xnor2_2 _18213_ (.A(_08818_),
    .B(net3949),
    .Y(_09035_));
 sky130_fd_sc_hd__nor2_2 _18214_ (.A(_08812_),
    .B(_09035_),
    .Y(_09036_));
 sky130_fd_sc_hd__o22ai_1 _18215_ (.A1(net3951),
    .A2(_08884_),
    .B1(net3615),
    .B2(net3685),
    .Y(_09037_));
 sky130_fd_sc_hd__a21oi_4 _18216_ (.A1(_08806_),
    .A2(_08812_),
    .B1(net3946),
    .Y(_09038_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_631 ();
 sky130_fd_sc_hd__nand2_1 _18218_ (.A(_12129_[0]),
    .B(net3946),
    .Y(_09040_));
 sky130_fd_sc_hd__a21oi_1 _18219_ (.A1(_08982_),
    .A2(_09040_),
    .B1(_08818_),
    .Y(_09041_));
 sky130_fd_sc_hd__a21oi_1 _18220_ (.A1(_08818_),
    .A2(_09038_),
    .B1(_09041_),
    .Y(_09042_));
 sky130_fd_sc_hd__o32ai_1 _18221_ (.A1(_09034_),
    .A2(_09036_),
    .A3(_09037_),
    .B1(_09042_),
    .B2(_09019_),
    .Y(_09043_));
 sky130_fd_sc_hd__nor3_2 _18222_ (.A(net3938),
    .B(_09033_),
    .C(_09043_),
    .Y(_09044_));
 sky130_fd_sc_hd__nor2_4 _18223_ (.A(net3685),
    .B(_08838_),
    .Y(_09045_));
 sky130_fd_sc_hd__o21ai_0 _18224_ (.A1(_12129_[0]),
    .A2(net3956),
    .B1(_09024_),
    .Y(_09046_));
 sky130_fd_sc_hd__a22oi_1 _18225_ (.A1(net3685),
    .A2(net3681),
    .B1(_09045_),
    .B2(_09046_),
    .Y(_09047_));
 sky130_fd_sc_hd__nand2_8 _18226_ (.A(_08930_),
    .B(net3943),
    .Y(_09048_));
 sky130_fd_sc_hd__o22ai_1 _18227_ (.A1(_08943_),
    .A2(_09019_),
    .B1(_09048_),
    .B2(_08950_),
    .Y(_09049_));
 sky130_fd_sc_hd__nor3_1 _18228_ (.A(net3956),
    .B(_08827_),
    .C(net3949),
    .Y(_09050_));
 sky130_fd_sc_hd__o21ai_0 _18229_ (.A1(_08970_),
    .A2(_09050_),
    .B1(net3685),
    .Y(_09051_));
 sky130_fd_sc_hd__o211ai_1 _18230_ (.A1(_08812_),
    .A2(_09047_),
    .B1(_09049_),
    .C1(_09051_),
    .Y(_09052_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_630 ();
 sky130_fd_sc_hd__nor3_1 _18232_ (.A(_08818_),
    .B(_08840_),
    .C(_08940_),
    .Y(_09054_));
 sky130_fd_sc_hd__nor2_4 _18233_ (.A(_12125_[0]),
    .B(net3946),
    .Y(_09055_));
 sky130_fd_sc_hd__nor3_1 _18234_ (.A(net3956),
    .B(net3585),
    .C(_09055_),
    .Y(_09056_));
 sky130_fd_sc_hd__nor2_2 _18235_ (.A(_08827_),
    .B(net3943),
    .Y(_09057_));
 sky130_fd_sc_hd__o21ai_0 _18236_ (.A1(_09054_),
    .A2(_09056_),
    .B1(_09057_),
    .Y(_09058_));
 sky130_fd_sc_hd__nor3_2 _18237_ (.A(net3956),
    .B(_08874_),
    .C(_09016_),
    .Y(_09059_));
 sky130_fd_sc_hd__nor3_1 _18238_ (.A(_08818_),
    .B(net3585),
    .C(_09055_),
    .Y(_09060_));
 sky130_fd_sc_hd__o21ai_0 _18239_ (.A1(_09059_),
    .A2(_09060_),
    .B1(_08957_),
    .Y(_09061_));
 sky130_fd_sc_hd__a41o_1 _18240_ (.A1(net3938),
    .A2(_09052_),
    .A3(_09058_),
    .A4(_09061_),
    .B1(_08916_),
    .X(_09062_));
 sky130_fd_sc_hd__o22ai_4 _18241_ (.A1(_09012_),
    .A2(_09026_),
    .B1(_09044_),
    .B2(_09062_),
    .Y(_00073_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_628 ();
 sky130_fd_sc_hd__nand2_2 _18244_ (.A(net3959),
    .B(net3957),
    .Y(_09064_));
 sky130_fd_sc_hd__nand2_2 _18245_ (.A(net3686),
    .B(net3956),
    .Y(_09065_));
 sky130_fd_sc_hd__a21oi_1 _18246_ (.A1(_09064_),
    .A2(_09065_),
    .B1(net3948),
    .Y(_09066_));
 sky130_fd_sc_hd__a21oi_1 _18247_ (.A1(_12148_[0]),
    .A2(net3948),
    .B1(_09066_),
    .Y(_09067_));
 sky130_fd_sc_hd__nor3_1 _18248_ (.A(net3959),
    .B(_08812_),
    .C(_08818_),
    .Y(_09068_));
 sky130_fd_sc_hd__nand2_1 _18249_ (.A(_12145_[0]),
    .B(net3948),
    .Y(_09069_));
 sky130_fd_sc_hd__o311ai_0 _18250_ (.A1(net3948),
    .A2(_08965_),
    .A3(_09068_),
    .B1(_09069_),
    .C1(net3955),
    .Y(_09070_));
 sky130_fd_sc_hd__o21ai_2 _18251_ (.A1(net3955),
    .A2(_09067_),
    .B1(_09070_),
    .Y(_09071_));
 sky130_fd_sc_hd__nand2_1 _18252_ (.A(_08941_),
    .B(_08964_),
    .Y(_09072_));
 sky130_fd_sc_hd__a32oi_1 _18253_ (.A1(net3685),
    .A2(net3956),
    .A3(net3615),
    .B1(_09072_),
    .B2(_12125_[0]),
    .Y(_09073_));
 sky130_fd_sc_hd__o2111ai_1 _18254_ (.A1(_08934_),
    .A2(_08919_),
    .B1(_09073_),
    .C1(_08957_),
    .D1(_08917_),
    .Y(_09074_));
 sky130_fd_sc_hd__nand2_2 _18255_ (.A(_08982_),
    .B(_09029_),
    .Y(_09075_));
 sky130_fd_sc_hd__nand2_4 _18256_ (.A(_12132_[0]),
    .B(net3951),
    .Y(_09076_));
 sky130_fd_sc_hd__nand3_1 _18257_ (.A(net3956),
    .B(_08901_),
    .C(_09076_),
    .Y(_09077_));
 sky130_fd_sc_hd__o21ai_0 _18258_ (.A1(net3956),
    .A2(_09075_),
    .B1(_09077_),
    .Y(_09078_));
 sky130_fd_sc_hd__nand3_1 _18259_ (.A(_08917_),
    .B(_09024_),
    .C(_09078_),
    .Y(_09079_));
 sky130_fd_sc_hd__o211ai_1 _18260_ (.A1(_08918_),
    .A2(_09071_),
    .B1(_09074_),
    .C1(_09079_),
    .Y(_09080_));
 sky130_fd_sc_hd__a21oi_2 _18261_ (.A1(_12126_[0]),
    .A2(net3954),
    .B1(_09045_),
    .Y(_09081_));
 sky130_fd_sc_hd__nor2_1 _18262_ (.A(net3957),
    .B(net3950),
    .Y(_09082_));
 sky130_fd_sc_hd__o21ai_1 _18263_ (.A1(_09082_),
    .A2(_08926_),
    .B1(net3956),
    .Y(_09083_));
 sky130_fd_sc_hd__o21ai_0 _18264_ (.A1(net3956),
    .A2(_09081_),
    .B1(_09083_),
    .Y(_09084_));
 sky130_fd_sc_hd__nor2_1 _18265_ (.A(_12138_[0]),
    .B(_08935_),
    .Y(_09085_));
 sky130_fd_sc_hd__a211oi_2 _18266_ (.A1(net3685),
    .A2(_09059_),
    .B1(_09085_),
    .C1(net3943),
    .Y(_09086_));
 sky130_fd_sc_hd__a211oi_1 _18267_ (.A1(net3944),
    .A2(_09084_),
    .B1(_09086_),
    .C1(net3937),
    .Y(_09087_));
 sky130_fd_sc_hd__nor2_1 _18268_ (.A(_09000_),
    .B(_09002_),
    .Y(_09088_));
 sky130_fd_sc_hd__nand2_1 _18269_ (.A(_12138_[0]),
    .B(_08818_),
    .Y(_09089_));
 sky130_fd_sc_hd__nand2_1 _18270_ (.A(net3948),
    .B(_09089_),
    .Y(_09090_));
 sky130_fd_sc_hd__a21oi_1 _18271_ (.A1(_12129_[0]),
    .A2(net3956),
    .B1(_09090_),
    .Y(_09091_));
 sky130_fd_sc_hd__nand3_1 _18272_ (.A(net3948),
    .B(_08884_),
    .C(_09065_),
    .Y(_09092_));
 sky130_fd_sc_hd__o21ai_0 _18273_ (.A1(_12129_[0]),
    .A2(net3956),
    .B1(_08860_),
    .Y(_09093_));
 sky130_fd_sc_hd__nand2_2 _18274_ (.A(_08860_),
    .B(net3946),
    .Y(_09094_));
 sky130_fd_sc_hd__o21ai_0 _18275_ (.A1(_09068_),
    .A2(_09093_),
    .B1(_09094_),
    .Y(_09095_));
 sky130_fd_sc_hd__nand2_1 _18276_ (.A(_09092_),
    .B(_09095_),
    .Y(_09096_));
 sky130_fd_sc_hd__o311a_1 _18277_ (.A1(_08860_),
    .A2(_09088_),
    .A3(_09091_),
    .B1(_09096_),
    .C1(net3937),
    .X(_09097_));
 sky130_fd_sc_hd__or4_1 _18278_ (.A(_08892_),
    .B(_08936_),
    .C(_09087_),
    .D(_09097_),
    .X(_09098_));
 sky130_fd_sc_hd__nand3_1 _18279_ (.A(net3956),
    .B(_08945_),
    .C(_08947_),
    .Y(_09099_));
 sky130_fd_sc_hd__nand3_1 _18280_ (.A(net3682),
    .B(_08982_),
    .C(_08948_),
    .Y(_09100_));
 sky130_fd_sc_hd__nor2_4 _18281_ (.A(_12134_[0]),
    .B(net3950),
    .Y(_09101_));
 sky130_fd_sc_hd__or3_1 _18282_ (.A(net3682),
    .B(_09030_),
    .C(_09101_),
    .X(_09102_));
 sky130_fd_sc_hd__or3_4 _18283_ (.A(_12138_[0]),
    .B(_08834_),
    .C(_08837_),
    .X(_09103_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_627 ();
 sky130_fd_sc_hd__nand3_1 _18285_ (.A(net3682),
    .B(_09000_),
    .C(_09103_),
    .Y(_09105_));
 sky130_fd_sc_hd__a21oi_1 _18286_ (.A1(_09102_),
    .A2(_09105_),
    .B1(net3940),
    .Y(_09106_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_626 ();
 sky130_fd_sc_hd__a311o_1 _18288_ (.A1(net3940),
    .A2(_09099_),
    .A3(_09100_),
    .B1(_09106_),
    .C1(net3937),
    .X(_09108_));
 sky130_fd_sc_hd__nor2_1 _18289_ (.A(net3957),
    .B(net3940),
    .Y(_09109_));
 sky130_fd_sc_hd__a211oi_1 _18290_ (.A1(net3685),
    .A2(net3940),
    .B1(net3950),
    .C1(_09109_),
    .Y(_09110_));
 sky130_fd_sc_hd__o21ai_0 _18291_ (.A1(_12134_[0]),
    .A2(net3954),
    .B1(net3956),
    .Y(_09111_));
 sky130_fd_sc_hd__nor2_4 _18292_ (.A(_08860_),
    .B(net3952),
    .Y(_09112_));
 sky130_fd_sc_hd__mux2i_1 _18293_ (.A0(_12129_[0]),
    .A1(_12138_[0]),
    .S(_09112_),
    .Y(_09113_));
 sky130_fd_sc_hd__o221ai_1 _18294_ (.A1(_09110_),
    .A2(_09111_),
    .B1(_09113_),
    .B2(net3956),
    .C1(net3937),
    .Y(_09114_));
 sky130_fd_sc_hd__nand4_1 _18295_ (.A(_08916_),
    .B(_08936_),
    .C(_09108_),
    .D(_09114_),
    .Y(_09115_));
 sky130_fd_sc_hd__nor2_4 _18296_ (.A(_08916_),
    .B(_08936_),
    .Y(_09116_));
 sky130_fd_sc_hd__nand2_4 _18297_ (.A(net3951),
    .B(_08873_),
    .Y(_09117_));
 sky130_fd_sc_hd__a21oi_1 _18298_ (.A1(net3614),
    .A2(_09117_),
    .B1(_08818_),
    .Y(_09118_));
 sky130_fd_sc_hd__nor2_2 _18299_ (.A(_12132_[0]),
    .B(net3951),
    .Y(_09119_));
 sky130_fd_sc_hd__nor3_1 _18300_ (.A(net3956),
    .B(_09038_),
    .C(_09119_),
    .Y(_09120_));
 sky130_fd_sc_hd__o221ai_1 _18301_ (.A1(_12152_[0]),
    .A2(net3952),
    .B1(_09000_),
    .B2(_09002_),
    .C1(net3937),
    .Y(_09121_));
 sky130_fd_sc_hd__o311ai_0 _18302_ (.A1(net3937),
    .A2(_09118_),
    .A3(_09120_),
    .B1(net3945),
    .C1(_09121_),
    .Y(_09122_));
 sky130_fd_sc_hd__nand2_1 _18303_ (.A(_12129_[0]),
    .B(_08818_),
    .Y(_09123_));
 sky130_fd_sc_hd__o22ai_1 _18304_ (.A1(net3946),
    .A2(_09123_),
    .B1(_09075_),
    .B2(_08818_),
    .Y(_09124_));
 sky130_fd_sc_hd__nor2_2 _18305_ (.A(net3958),
    .B(_08812_),
    .Y(_09125_));
 sky130_fd_sc_hd__nand3_1 _18306_ (.A(_08818_),
    .B(net3946),
    .C(_09125_),
    .Y(_09126_));
 sky130_fd_sc_hd__a21oi_1 _18307_ (.A1(_12143_[0]),
    .A2(net3952),
    .B1(_08827_),
    .Y(_09127_));
 sky130_fd_sc_hd__a221o_1 _18308_ (.A1(net3955),
    .A2(_09124_),
    .B1(_09126_),
    .B2(_09127_),
    .C1(net3945),
    .X(_09128_));
 sky130_fd_sc_hd__nand3_2 _18309_ (.A(_09116_),
    .B(_09122_),
    .C(_09128_),
    .Y(_09129_));
 sky130_fd_sc_hd__nand4b_1 _18310_ (.A_N(_09080_),
    .B(_09098_),
    .C(_09115_),
    .D(_09129_),
    .Y(_00074_));
 sky130_fd_sc_hd__nor3_1 _18311_ (.A(net3956),
    .B(_09055_),
    .C(_09119_),
    .Y(_09130_));
 sky130_fd_sc_hd__a21oi_1 _18312_ (.A1(net3956),
    .A2(_09081_),
    .B1(_09130_),
    .Y(_09131_));
 sky130_fd_sc_hd__a21oi_1 _18313_ (.A1(_12126_[0]),
    .A2(net3954),
    .B1(_08906_),
    .Y(_09132_));
 sky130_fd_sc_hd__o31ai_1 _18314_ (.A1(net3682),
    .A2(net3940),
    .A3(_09132_),
    .B1(_08827_),
    .Y(_09133_));
 sky130_fd_sc_hd__nand3_4 _18315_ (.A(_08812_),
    .B(net3956),
    .C(net3947),
    .Y(_09134_));
 sky130_fd_sc_hd__nand3_1 _18316_ (.A(_12134_[0]),
    .B(net3939),
    .C(_09035_),
    .Y(_09135_));
 sky130_fd_sc_hd__o21ai_0 _18317_ (.A1(net3943),
    .A2(_09134_),
    .B1(_09135_),
    .Y(_09136_));
 sky130_fd_sc_hd__o22ai_1 _18318_ (.A1(_09048_),
    .A2(_09131_),
    .B1(_09133_),
    .B2(_09136_),
    .Y(_09137_));
 sky130_fd_sc_hd__a21oi_2 _18319_ (.A1(_08945_),
    .A2(_08962_),
    .B1(net3956),
    .Y(_09138_));
 sky130_fd_sc_hd__nor3_1 _18320_ (.A(_12126_[0]),
    .B(_12129_[0]),
    .C(net3950),
    .Y(_09139_));
 sky130_fd_sc_hd__nor3_1 _18321_ (.A(net3682),
    .B(_08906_),
    .C(_09139_),
    .Y(_09140_));
 sky130_fd_sc_hd__nor3_1 _18322_ (.A(_09034_),
    .B(_09138_),
    .C(_09140_),
    .Y(_09141_));
 sky130_fd_sc_hd__nor3_1 _18323_ (.A(_08936_),
    .B(_09137_),
    .C(_09141_),
    .Y(_09142_));
 sky130_fd_sc_hd__a211oi_1 _18324_ (.A1(_12132_[0]),
    .A2(net3946),
    .B1(_09101_),
    .C1(net3956),
    .Y(_09143_));
 sky130_fd_sc_hd__a311oi_1 _18325_ (.A1(net3956),
    .A2(net3614),
    .A3(_09117_),
    .B1(_09143_),
    .C1(net3945),
    .Y(_09144_));
 sky130_fd_sc_hd__nor3_1 _18326_ (.A(_08860_),
    .B(_08919_),
    .C(_09090_),
    .Y(_09145_));
 sky130_fd_sc_hd__o21ai_1 _18327_ (.A1(_09144_),
    .A2(_09145_),
    .B1(net3937),
    .Y(_09146_));
 sky130_fd_sc_hd__nor2_4 _18328_ (.A(_08930_),
    .B(net3943),
    .Y(_09147_));
 sky130_fd_sc_hd__nand2_1 _18329_ (.A(net3685),
    .B(_08955_),
    .Y(_09148_));
 sky130_fd_sc_hd__o21ai_0 _18330_ (.A1(net3682),
    .A2(_09045_),
    .B1(net3684),
    .Y(_09149_));
 sky130_fd_sc_hd__o2111ai_1 _18331_ (.A1(_12124_[0]),
    .A2(_08935_),
    .B1(_09147_),
    .C1(_09148_),
    .D1(_09149_),
    .Y(_09150_));
 sky130_fd_sc_hd__nand2_4 _18332_ (.A(_12125_[0]),
    .B(net3946),
    .Y(_09151_));
 sky130_fd_sc_hd__nand2_2 _18333_ (.A(_12134_[0]),
    .B(net3952),
    .Y(_09152_));
 sky130_fd_sc_hd__nand2_4 _18334_ (.A(_09151_),
    .B(_09152_),
    .Y(_09153_));
 sky130_fd_sc_hd__nand2_1 _18335_ (.A(net3956),
    .B(_09153_),
    .Y(_09154_));
 sky130_fd_sc_hd__nand3_1 _18336_ (.A(_08818_),
    .B(net3615),
    .C(_09103_),
    .Y(_09155_));
 sky130_fd_sc_hd__a31oi_1 _18337_ (.A1(_08957_),
    .A2(_09154_),
    .A3(_09155_),
    .B1(net3938),
    .Y(_09156_));
 sky130_fd_sc_hd__and3_1 _18338_ (.A(_09146_),
    .B(_09150_),
    .C(_09156_),
    .X(_09157_));
 sky130_fd_sc_hd__nor2_1 _18339_ (.A(_12124_[0]),
    .B(net3950),
    .Y(_09158_));
 sky130_fd_sc_hd__nor3_1 _18340_ (.A(net3682),
    .B(_09158_),
    .C(_09119_),
    .Y(_09159_));
 sky130_fd_sc_hd__a31oi_1 _18341_ (.A1(net3682),
    .A2(_08945_),
    .A3(_08982_),
    .B1(_09159_),
    .Y(_09160_));
 sky130_fd_sc_hd__or3_1 _18342_ (.A(net3682),
    .B(_08940_),
    .C(_08926_),
    .X(_09161_));
 sky130_fd_sc_hd__o311ai_0 _18343_ (.A1(net3956),
    .A2(_09045_),
    .A3(_08953_),
    .B1(_09161_),
    .C1(net3940),
    .Y(_09162_));
 sky130_fd_sc_hd__o21ai_0 _18344_ (.A1(net3940),
    .A2(_09160_),
    .B1(_09162_),
    .Y(_09163_));
 sky130_fd_sc_hd__o31ai_1 _18345_ (.A1(net3944),
    .A2(_08901_),
    .A3(_08919_),
    .B1(_09116_),
    .Y(_09164_));
 sky130_fd_sc_hd__a311oi_1 _18346_ (.A1(net3685),
    .A2(net3944),
    .A3(_08955_),
    .B1(_09164_),
    .C1(net3955),
    .Y(_09165_));
 sky130_fd_sc_hd__nor2_4 _18347_ (.A(_08860_),
    .B(net3950),
    .Y(_09166_));
 sky130_fd_sc_hd__nor2_1 _18348_ (.A(_08818_),
    .B(net3944),
    .Y(_09167_));
 sky130_fd_sc_hd__a21oi_1 _18349_ (.A1(_08818_),
    .A2(_09166_),
    .B1(_09167_),
    .Y(_09168_));
 sky130_fd_sc_hd__o21ai_0 _18350_ (.A1(net3957),
    .A2(_09167_),
    .B1(net3950),
    .Y(_09169_));
 sky130_fd_sc_hd__o221ai_1 _18351_ (.A1(_08964_),
    .A2(_09166_),
    .B1(_09168_),
    .B2(_12125_[0]),
    .C1(_09169_),
    .Y(_09170_));
 sky130_fd_sc_hd__a32oi_1 _18352_ (.A1(_09116_),
    .A2(net3955),
    .A3(_09163_),
    .B1(_09165_),
    .B2(_09170_),
    .Y(_09171_));
 sky130_fd_sc_hd__a21oi_2 _18353_ (.A1(_08934_),
    .A2(_09151_),
    .B1(_08818_),
    .Y(_09172_));
 sky130_fd_sc_hd__a31oi_1 _18354_ (.A1(_08818_),
    .A2(_08948_),
    .A3(_08962_),
    .B1(_09172_),
    .Y(_09173_));
 sky130_fd_sc_hd__nor2_1 _18355_ (.A(net3944),
    .B(_09002_),
    .Y(_09174_));
 sky130_fd_sc_hd__a31oi_1 _18356_ (.A1(_08935_),
    .A2(_09064_),
    .A3(_09174_),
    .B1(net3955),
    .Y(_09175_));
 sky130_fd_sc_hd__o21ai_0 _18357_ (.A1(_08860_),
    .A2(_09173_),
    .B1(_09175_),
    .Y(_09176_));
 sky130_fd_sc_hd__nand2_1 _18358_ (.A(_12132_[0]),
    .B(_08943_),
    .Y(_09177_));
 sky130_fd_sc_hd__nand2_2 _18359_ (.A(_08818_),
    .B(_08838_),
    .Y(_09178_));
 sky130_fd_sc_hd__o21ai_0 _18360_ (.A1(net3684),
    .A2(_09178_),
    .B1(_09134_),
    .Y(_09179_));
 sky130_fd_sc_hd__nand2_1 _18361_ (.A(net3685),
    .B(_09179_),
    .Y(_09180_));
 sky130_fd_sc_hd__o2111ai_2 _18362_ (.A1(_12125_[0]),
    .A2(_08853_),
    .B1(_09147_),
    .C1(_09177_),
    .D1(_09180_),
    .Y(_09181_));
 sky130_fd_sc_hd__nor2_4 _18363_ (.A(net3684),
    .B(_08934_),
    .Y(_09182_));
 sky130_fd_sc_hd__a21oi_1 _18364_ (.A1(_12132_[0]),
    .A2(_08955_),
    .B1(_09182_),
    .Y(_09183_));
 sky130_fd_sc_hd__nand3_1 _18365_ (.A(_08957_),
    .B(_09083_),
    .C(_09183_),
    .Y(_09184_));
 sky130_fd_sc_hd__nand4_1 _18366_ (.A(_08917_),
    .B(_09176_),
    .C(_09181_),
    .D(_09184_),
    .Y(_09185_));
 sky130_fd_sc_hd__o311a_1 _18367_ (.A1(_08892_),
    .A2(_09142_),
    .A3(_09157_),
    .B1(_09171_),
    .C1(_09185_),
    .X(_00075_));
 sky130_fd_sc_hd__a211oi_1 _18368_ (.A1(_12134_[0]),
    .A2(net3956),
    .B1(_08930_),
    .C1(_09056_),
    .Y(_09186_));
 sky130_fd_sc_hd__and2_4 _18369_ (.A(_08934_),
    .B(_09103_),
    .X(_09187_));
 sky130_fd_sc_hd__nor3_1 _18370_ (.A(_08818_),
    .B(_08856_),
    .C(net3585),
    .Y(_09188_));
 sky130_fd_sc_hd__a211oi_1 _18371_ (.A1(_08818_),
    .A2(_09187_),
    .B1(_09188_),
    .C1(_08827_),
    .Y(_09189_));
 sky130_fd_sc_hd__nor3_1 _18372_ (.A(net3939),
    .B(_09186_),
    .C(_09189_),
    .Y(_09190_));
 sky130_fd_sc_hd__nand2_1 _18373_ (.A(net3956),
    .B(_09103_),
    .Y(_09191_));
 sky130_fd_sc_hd__a2bb2oi_1 _18374_ (.A1_N(_08856_),
    .A2_N(_09191_),
    .B1(_09153_),
    .B2(_08818_),
    .Y(_09192_));
 sky130_fd_sc_hd__a21oi_1 _18375_ (.A1(_08827_),
    .A2(_09192_),
    .B1(net3943),
    .Y(_09193_));
 sky130_fd_sc_hd__nor3_1 _18376_ (.A(_08936_),
    .B(_09190_),
    .C(_09193_),
    .Y(_09194_));
 sky130_fd_sc_hd__a221oi_1 _18377_ (.A1(net3958),
    .A2(net3956),
    .B1(net3681),
    .B2(_12124_[0]),
    .C1(_09048_),
    .Y(_09195_));
 sky130_fd_sc_hd__a21oi_1 _18378_ (.A1(_12134_[0]),
    .A2(_08838_),
    .B1(net3956),
    .Y(_09196_));
 sky130_fd_sc_hd__nor2_1 _18379_ (.A(_08855_),
    .B(_09196_),
    .Y(_09197_));
 sky130_fd_sc_hd__nor2_1 _18380_ (.A(net3939),
    .B(_09197_),
    .Y(_09198_));
 sky130_fd_sc_hd__a311oi_1 _18381_ (.A1(_08818_),
    .A2(_09000_),
    .A3(_09029_),
    .B1(net3943),
    .C1(_08919_),
    .Y(_09199_));
 sky130_fd_sc_hd__nor3_1 _18382_ (.A(_08930_),
    .B(_09198_),
    .C(_09199_),
    .Y(_09200_));
 sky130_fd_sc_hd__nand2_1 _18383_ (.A(_09057_),
    .B(_09134_),
    .Y(_09201_));
 sky130_fd_sc_hd__a211oi_1 _18384_ (.A1(net3685),
    .A2(_09035_),
    .B1(_09182_),
    .C1(_09201_),
    .Y(_09202_));
 sky130_fd_sc_hd__a2111oi_0 _18385_ (.A1(net3614),
    .A2(_09195_),
    .B1(_09200_),
    .C1(net3938),
    .D1(_09202_),
    .Y(_09203_));
 sky130_fd_sc_hd__a21oi_1 _18386_ (.A1(_09000_),
    .A2(_09040_),
    .B1(net3956),
    .Y(_09204_));
 sky130_fd_sc_hd__nor4_1 _18387_ (.A(_08936_),
    .B(_08870_),
    .C(_09034_),
    .D(_09204_),
    .Y(_09205_));
 sky130_fd_sc_hd__nand4_1 _18388_ (.A(_08818_),
    .B(_08991_),
    .C(_08910_),
    .D(_08957_),
    .Y(_09206_));
 sky130_fd_sc_hd__nor2_1 _18389_ (.A(net3949),
    .B(_08923_),
    .Y(_09207_));
 sky130_fd_sc_hd__o21ai_1 _18390_ (.A1(_09082_),
    .A2(_08906_),
    .B1(net3682),
    .Y(_09208_));
 sky130_fd_sc_hd__o311ai_1 _18391_ (.A1(_08818_),
    .A2(_08911_),
    .A3(_09207_),
    .B1(_09147_),
    .C1(_09208_),
    .Y(_09209_));
 sky130_fd_sc_hd__o211ai_1 _18392_ (.A1(_12129_[0]),
    .A2(net3949),
    .B1(_09029_),
    .C1(net3956),
    .Y(_09210_));
 sky130_fd_sc_hd__o22ai_1 _18393_ (.A1(net3682),
    .A2(_09030_),
    .B1(_08853_),
    .B2(_12138_[0]),
    .Y(_09211_));
 sky130_fd_sc_hd__a32oi_1 _18394_ (.A1(_09022_),
    .A2(_09024_),
    .A3(_09210_),
    .B1(_09211_),
    .B2(_09057_),
    .Y(_09212_));
 sky130_fd_sc_hd__a31oi_2 _18395_ (.A1(_09206_),
    .A2(_09209_),
    .A3(_09212_),
    .B1(net3938),
    .Y(_09213_));
 sky130_fd_sc_hd__nand2_4 _18396_ (.A(_08827_),
    .B(_08849_),
    .Y(_09214_));
 sky130_fd_sc_hd__a2111oi_0 _18397_ (.A1(net3958),
    .A2(_08943_),
    .B1(_09214_),
    .C1(_09196_),
    .D1(_08840_),
    .Y(_09215_));
 sky130_fd_sc_hd__o21ai_0 _18398_ (.A1(_08874_),
    .A2(_09045_),
    .B1(net3956),
    .Y(_09216_));
 sky130_fd_sc_hd__a31oi_1 _18399_ (.A1(_08859_),
    .A2(net3614),
    .A3(_09216_),
    .B1(_09048_),
    .Y(_09217_));
 sky130_fd_sc_hd__a21oi_1 _18400_ (.A1(net3615),
    .A2(_09029_),
    .B1(net3956),
    .Y(_09218_));
 sky130_fd_sc_hd__nor4_1 _18401_ (.A(_08856_),
    .B(_08977_),
    .C(_09034_),
    .D(_09218_),
    .Y(_09219_));
 sky130_fd_sc_hd__nor2_2 _18402_ (.A(_12136_[0]),
    .B(net3953),
    .Y(_09220_));
 sky130_fd_sc_hd__a21oi_2 _18403_ (.A1(net3951),
    .A2(_08884_),
    .B1(_09220_),
    .Y(_09221_));
 sky130_fd_sc_hd__o21ai_0 _18404_ (.A1(_09019_),
    .A2(_09221_),
    .B1(net3938),
    .Y(_09222_));
 sky130_fd_sc_hd__nor4_1 _18405_ (.A(_09215_),
    .B(_09217_),
    .C(_09219_),
    .D(_09222_),
    .Y(_09223_));
 sky130_fd_sc_hd__or3_1 _18406_ (.A(_08892_),
    .B(_09213_),
    .C(_09223_),
    .X(_09224_));
 sky130_fd_sc_hd__o41ai_1 _18407_ (.A1(_08916_),
    .A2(_09194_),
    .A3(_09203_),
    .A4(_09205_),
    .B1(_09224_),
    .Y(_00076_));
 sky130_fd_sc_hd__a21oi_1 _18408_ (.A1(net3683),
    .A2(_08976_),
    .B1(_08840_),
    .Y(_09225_));
 sky130_fd_sc_hd__o21ai_0 _18409_ (.A1(_12134_[0]),
    .A2(_08838_),
    .B1(_08818_),
    .Y(_09226_));
 sky130_fd_sc_hd__o32ai_1 _18410_ (.A1(_08818_),
    .A2(_09045_),
    .A3(_09055_),
    .B1(_09226_),
    .B2(_08856_),
    .Y(_09227_));
 sky130_fd_sc_hd__nand2_1 _18411_ (.A(net3943),
    .B(_09227_),
    .Y(_09228_));
 sky130_fd_sc_hd__o211ai_1 _18412_ (.A1(net3943),
    .A2(_09225_),
    .B1(_09228_),
    .C1(_08936_),
    .Y(_09229_));
 sky130_fd_sc_hd__o32ai_1 _18413_ (.A1(_08941_),
    .A2(_09001_),
    .A3(_09002_),
    .B1(_09117_),
    .B2(_08818_),
    .Y(_09230_));
 sky130_fd_sc_hd__a21oi_2 _18414_ (.A1(net3948),
    .A2(_09123_),
    .B1(_08860_),
    .Y(_09231_));
 sky130_fd_sc_hd__o21ai_0 _18415_ (.A1(_12138_[0]),
    .A2(_09178_),
    .B1(_09231_),
    .Y(_09232_));
 sky130_fd_sc_hd__o211ai_1 _18416_ (.A1(_08849_),
    .A2(_09230_),
    .B1(_09232_),
    .C1(net3938),
    .Y(_09233_));
 sky130_fd_sc_hd__nand3_1 _18417_ (.A(net3680),
    .B(_09229_),
    .C(_09233_),
    .Y(_09234_));
 sky130_fd_sc_hd__nor2_1 _18418_ (.A(_08935_),
    .B(_08923_),
    .Y(_09235_));
 sky130_fd_sc_hd__o21a_1 _18419_ (.A1(_08976_),
    .A2(_08923_),
    .B1(_09076_),
    .X(_09236_));
 sky130_fd_sc_hd__a21oi_1 _18420_ (.A1(net3938),
    .A2(_09236_),
    .B1(net3943),
    .Y(_09237_));
 sky130_fd_sc_hd__o41ai_1 _18421_ (.A1(net3938),
    .A2(_08950_),
    .A3(_09036_),
    .A4(_09235_),
    .B1(_09237_),
    .Y(_09238_));
 sky130_fd_sc_hd__a21oi_1 _18422_ (.A1(_08982_),
    .A2(_09151_),
    .B1(_08936_),
    .Y(_09239_));
 sky130_fd_sc_hd__a211oi_1 _18423_ (.A1(_08936_),
    .A2(_08924_),
    .B1(_09239_),
    .C1(_08818_),
    .Y(_09240_));
 sky130_fd_sc_hd__a311o_1 _18424_ (.A1(_08818_),
    .A2(_09076_),
    .A3(_09103_),
    .B1(_09240_),
    .C1(net3942),
    .X(_09241_));
 sky130_fd_sc_hd__nand4_1 _18425_ (.A(_08916_),
    .B(_08930_),
    .C(_09238_),
    .D(_09241_),
    .Y(_09242_));
 sky130_fd_sc_hd__a221o_1 _18426_ (.A1(_12129_[0]),
    .A2(net3951),
    .B1(_08955_),
    .B2(_12134_[0]),
    .C1(_08851_),
    .X(_09243_));
 sky130_fd_sc_hd__o311ai_0 _18427_ (.A1(_08818_),
    .A2(_08855_),
    .A3(_08953_),
    .B1(_08942_),
    .C1(net3941),
    .Y(_09244_));
 sky130_fd_sc_hd__nand4_1 _18428_ (.A(net3955),
    .B(_08917_),
    .C(_09243_),
    .D(_09244_),
    .Y(_09245_));
 sky130_fd_sc_hd__a21oi_2 _18429_ (.A1(_08991_),
    .A2(_08947_),
    .B1(net3956),
    .Y(_09246_));
 sky130_fd_sc_hd__a21oi_1 _18430_ (.A1(net3959),
    .A2(_08970_),
    .B1(_09246_),
    .Y(_09247_));
 sky130_fd_sc_hd__a21oi_1 _18431_ (.A1(_08925_),
    .A2(_08994_),
    .B1(net3956),
    .Y(_09248_));
 sky130_fd_sc_hd__nor3_1 _18432_ (.A(net3945),
    .B(_08972_),
    .C(_09248_),
    .Y(_09249_));
 sky130_fd_sc_hd__a21oi_2 _18433_ (.A1(net3945),
    .A2(_09247_),
    .B1(_09249_),
    .Y(_09250_));
 sky130_fd_sc_hd__nand2_1 _18434_ (.A(_08849_),
    .B(_08943_),
    .Y(_09251_));
 sky130_fd_sc_hd__o21ai_0 _18435_ (.A1(net3686),
    .A2(_09112_),
    .B1(_08812_),
    .Y(_09252_));
 sky130_fd_sc_hd__a31oi_1 _18436_ (.A1(net3686),
    .A2(_09094_),
    .A3(_09251_),
    .B1(_09252_),
    .Y(_09253_));
 sky130_fd_sc_hd__a22oi_1 _18437_ (.A1(net3957),
    .A2(_08970_),
    .B1(net3681),
    .B2(_12132_[0]),
    .Y(_09254_));
 sky130_fd_sc_hd__o32ai_1 _18438_ (.A1(net3686),
    .A2(_08955_),
    .A3(_09166_),
    .B1(_09254_),
    .B2(net3942),
    .Y(_09255_));
 sky130_fd_sc_hd__nor4_1 _18439_ (.A(_08898_),
    .B(net3937),
    .C(_09253_),
    .D(_09255_),
    .Y(_09256_));
 sky130_fd_sc_hd__a221oi_1 _18440_ (.A1(_12129_[0]),
    .A2(_09112_),
    .B1(_09153_),
    .B2(net3942),
    .C1(_08818_),
    .Y(_09257_));
 sky130_fd_sc_hd__nand2_1 _18441_ (.A(_08849_),
    .B(_09125_),
    .Y(_09258_));
 sky130_fd_sc_hd__nand2_1 _18442_ (.A(net3942),
    .B(_09002_),
    .Y(_09259_));
 sky130_fd_sc_hd__a21oi_1 _18443_ (.A1(_09258_),
    .A2(_09259_),
    .B1(net3946),
    .Y(_09260_));
 sky130_fd_sc_hd__nor3_1 _18444_ (.A(_08951_),
    .B(_09257_),
    .C(_09260_),
    .Y(_09261_));
 sky130_fd_sc_hd__a311oi_2 _18445_ (.A1(_09116_),
    .A2(net3937),
    .A3(_09250_),
    .B1(_09256_),
    .C1(_09261_),
    .Y(_09262_));
 sky130_fd_sc_hd__nand4_1 _18446_ (.A(_09234_),
    .B(_09242_),
    .C(_09245_),
    .D(_09262_),
    .Y(_00077_));
 sky130_fd_sc_hd__nor2_1 _18447_ (.A(_08855_),
    .B(_08856_),
    .Y(_09263_));
 sky130_fd_sc_hd__nor2_1 _18448_ (.A(net3956),
    .B(_09263_),
    .Y(_09264_));
 sky130_fd_sc_hd__o21ai_2 _18449_ (.A1(_08806_),
    .A2(_08818_),
    .B1(_09038_),
    .Y(_09265_));
 sky130_fd_sc_hd__o311ai_0 _18450_ (.A1(_12141_[0]),
    .A2(_12150_[0]),
    .A3(net3952),
    .B1(_09265_),
    .C1(_08936_),
    .Y(_09266_));
 sky130_fd_sc_hd__o31ai_1 _18451_ (.A1(_08936_),
    .A2(_09172_),
    .A3(_09264_),
    .B1(_09266_),
    .Y(_09267_));
 sky130_fd_sc_hd__o21a_1 _18452_ (.A1(_12124_[0]),
    .A2(net3952),
    .B1(_09152_),
    .X(_09268_));
 sky130_fd_sc_hd__nand2_1 _18453_ (.A(_12126_[0]),
    .B(net3681),
    .Y(_09269_));
 sky130_fd_sc_hd__o21ai_0 _18454_ (.A1(_08818_),
    .A2(_09268_),
    .B1(_09269_),
    .Y(_09270_));
 sky130_fd_sc_hd__o21ai_0 _18455_ (.A1(_12125_[0]),
    .A2(_08818_),
    .B1(net3946),
    .Y(_09271_));
 sky130_fd_sc_hd__a21oi_1 _18456_ (.A1(_08818_),
    .A2(_09125_),
    .B1(_09271_),
    .Y(_09272_));
 sky130_fd_sc_hd__o21ai_0 _18457_ (.A1(_12143_[0]),
    .A2(net3946),
    .B1(net3938),
    .Y(_09273_));
 sky130_fd_sc_hd__o221a_1 _18458_ (.A1(net3938),
    .A2(_09270_),
    .B1(_09272_),
    .B2(_09273_),
    .C1(_08849_),
    .X(_09274_));
 sky130_fd_sc_hd__a2111oi_0 _18459_ (.A1(net3942),
    .A2(_09267_),
    .B1(_09274_),
    .C1(net3937),
    .D1(_08916_),
    .Y(_09275_));
 sky130_fd_sc_hd__a21oi_1 _18460_ (.A1(net3942),
    .A2(_09153_),
    .B1(_09166_),
    .Y(_09276_));
 sky130_fd_sc_hd__nor2_1 _18461_ (.A(_08849_),
    .B(net3946),
    .Y(_09277_));
 sky130_fd_sc_hd__a22o_1 _18462_ (.A1(net3958),
    .A2(_08849_),
    .B1(_09277_),
    .B2(net3957),
    .X(_09278_));
 sky130_fd_sc_hd__a221oi_1 _18463_ (.A1(_08812_),
    .A2(_09112_),
    .B1(_09278_),
    .B2(_08818_),
    .C1(net3938),
    .Y(_09279_));
 sky130_fd_sc_hd__o21ai_0 _18464_ (.A1(_08818_),
    .A2(_09276_),
    .B1(_09279_),
    .Y(_09280_));
 sky130_fd_sc_hd__a21oi_1 _18465_ (.A1(net3959),
    .A2(net3951),
    .B1(_08818_),
    .Y(_09281_));
 sky130_fd_sc_hd__o21ai_0 _18466_ (.A1(_09143_),
    .A2(_09281_),
    .B1(net3945),
    .Y(_09282_));
 sky130_fd_sc_hd__nand3b_1 _18467_ (.A_N(_09095_),
    .B(_09282_),
    .C(net3938),
    .Y(_09283_));
 sky130_fd_sc_hd__a21oi_1 _18468_ (.A1(_09280_),
    .A2(_09283_),
    .B1(_08969_),
    .Y(_09284_));
 sky130_fd_sc_hd__o21ai_0 _18469_ (.A1(net3958),
    .A2(_08919_),
    .B1(net3952),
    .Y(_09285_));
 sky130_fd_sc_hd__nor2_1 _18470_ (.A(_08854_),
    .B(_09048_),
    .Y(_09286_));
 sky130_fd_sc_hd__a211oi_1 _18471_ (.A1(net3947),
    .A2(_08873_),
    .B1(_08856_),
    .C1(_08818_),
    .Y(_09287_));
 sky130_fd_sc_hd__a311oi_1 _18472_ (.A1(_08818_),
    .A2(net3615),
    .A3(_09151_),
    .B1(_09034_),
    .C1(_09287_),
    .Y(_09288_));
 sky130_fd_sc_hd__a21oi_1 _18473_ (.A1(_09285_),
    .A2(_09286_),
    .B1(_09288_),
    .Y(_09289_));
 sky130_fd_sc_hd__nand2_1 _18474_ (.A(_12126_[0]),
    .B(_08838_),
    .Y(_09290_));
 sky130_fd_sc_hd__nand3_1 _18475_ (.A(net3956),
    .B(_08994_),
    .C(_09290_),
    .Y(_09291_));
 sky130_fd_sc_hd__nand3_1 _18476_ (.A(net3682),
    .B(_08910_),
    .C(_08948_),
    .Y(_09292_));
 sky130_fd_sc_hd__nand2_1 _18477_ (.A(_09291_),
    .B(_09292_),
    .Y(_09293_));
 sky130_fd_sc_hd__nor3_1 _18478_ (.A(net3956),
    .B(_08926_),
    .C(_09139_),
    .Y(_09294_));
 sky130_fd_sc_hd__nor3_1 _18479_ (.A(_08818_),
    .B(net3679),
    .C(_09101_),
    .Y(_09295_));
 sky130_fd_sc_hd__o21ai_0 _18480_ (.A1(_09294_),
    .A2(_09295_),
    .B1(net3944),
    .Y(_09296_));
 sky130_fd_sc_hd__o21ai_2 _18481_ (.A1(net3944),
    .A2(_09293_),
    .B1(_09296_),
    .Y(_09297_));
 sky130_fd_sc_hd__o22ai_1 _18482_ (.A1(_08898_),
    .A2(_09289_),
    .B1(_09297_),
    .B2(_08951_),
    .Y(_09298_));
 sky130_fd_sc_hd__a21oi_1 _18483_ (.A1(net3959),
    .A2(_09001_),
    .B1(net3679),
    .Y(_09299_));
 sky130_fd_sc_hd__nor2_1 _18484_ (.A(_12138_[0]),
    .B(_09299_),
    .Y(_09300_));
 sky130_fd_sc_hd__o31ai_1 _18485_ (.A1(_09002_),
    .A2(_09182_),
    .A3(_09300_),
    .B1(_08849_),
    .Y(_09301_));
 sky130_fd_sc_hd__o22ai_1 _18486_ (.A1(_08849_),
    .A2(_09002_),
    .B1(_09103_),
    .B2(_08818_),
    .Y(_09302_));
 sky130_fd_sc_hd__a221oi_1 _18487_ (.A1(_08919_),
    .A2(_09277_),
    .B1(_09302_),
    .B2(net3686),
    .C1(net3938),
    .Y(_09303_));
 sky130_fd_sc_hd__nand2_1 _18488_ (.A(_12142_[0]),
    .B(net3952),
    .Y(_09304_));
 sky130_fd_sc_hd__nand2_1 _18489_ (.A(_12134_[0]),
    .B(_08818_),
    .Y(_09305_));
 sky130_fd_sc_hd__nand3_1 _18490_ (.A(net3948),
    .B(_09065_),
    .C(_09305_),
    .Y(_09306_));
 sky130_fd_sc_hd__a21oi_1 _18491_ (.A1(_09304_),
    .A2(_09306_),
    .B1(_08849_),
    .Y(_09307_));
 sky130_fd_sc_hd__o31ai_1 _18492_ (.A1(_08860_),
    .A2(_08972_),
    .A3(_09138_),
    .B1(net3938),
    .Y(_09308_));
 sky130_fd_sc_hd__o21ai_0 _18493_ (.A1(_09307_),
    .A2(_09308_),
    .B1(net3680),
    .Y(_09309_));
 sky130_fd_sc_hd__a21oi_1 _18494_ (.A1(_09301_),
    .A2(_09303_),
    .B1(_09309_),
    .Y(_09310_));
 sky130_fd_sc_hd__nor4_1 _18495_ (.A(_09275_),
    .B(_09284_),
    .C(_09298_),
    .D(_09310_),
    .Y(_00078_));
 sky130_fd_sc_hd__o21ai_0 _18496_ (.A1(_08812_),
    .A2(_08935_),
    .B1(_08945_),
    .Y(_09311_));
 sky130_fd_sc_hd__a21oi_1 _18497_ (.A1(_09178_),
    .A2(_09134_),
    .B1(net3958),
    .Y(_09312_));
 sky130_fd_sc_hd__a21oi_1 _18498_ (.A1(net3957),
    .A2(net3946),
    .B1(net3958),
    .Y(_09313_));
 sky130_fd_sc_hd__a311oi_1 _18499_ (.A1(net3958),
    .A2(_08853_),
    .A3(_08902_),
    .B1(_09313_),
    .C1(_08849_),
    .Y(_09314_));
 sky130_fd_sc_hd__a211o_4 _18500_ (.A1(_08849_),
    .A2(_09311_),
    .B1(_09312_),
    .C1(_09314_),
    .X(_09315_));
 sky130_fd_sc_hd__a21oi_1 _18501_ (.A1(_08818_),
    .A2(_08923_),
    .B1(net3953),
    .Y(_09316_));
 sky130_fd_sc_hd__o21ai_0 _18502_ (.A1(_08906_),
    .A2(_09038_),
    .B1(net3956),
    .Y(_09317_));
 sky130_fd_sc_hd__o21ai_0 _18503_ (.A1(net3942),
    .A2(_09316_),
    .B1(_09317_),
    .Y(_09318_));
 sky130_fd_sc_hd__a31oi_2 _18504_ (.A1(_08849_),
    .A2(_09125_),
    .A3(_08943_),
    .B1(_08969_),
    .Y(_09319_));
 sky130_fd_sc_hd__a22o_4 _18505_ (.A1(net3680),
    .A2(_09315_),
    .B1(_09318_),
    .B2(_09319_),
    .X(_09320_));
 sky130_fd_sc_hd__a21oi_2 _18506_ (.A1(_08916_),
    .A2(_08936_),
    .B1(_09320_),
    .Y(_09321_));
 sky130_fd_sc_hd__a21oi_1 _18507_ (.A1(net3684),
    .A2(net3681),
    .B1(_09030_),
    .Y(_09322_));
 sky130_fd_sc_hd__nor2_1 _18508_ (.A(net3958),
    .B(_09322_),
    .Y(_09323_));
 sky130_fd_sc_hd__a221oi_1 _18509_ (.A1(_12124_[0]),
    .A2(_08943_),
    .B1(_08955_),
    .B2(net3957),
    .C1(_09323_),
    .Y(_09324_));
 sky130_fd_sc_hd__o221ai_2 _18510_ (.A1(_12138_[0]),
    .A2(_08935_),
    .B1(_09035_),
    .B2(_12125_[0]),
    .C1(_08985_),
    .Y(_09325_));
 sky130_fd_sc_hd__a21oi_2 _18511_ (.A1(_08930_),
    .A2(_09325_),
    .B1(net3939),
    .Y(_09326_));
 sky130_fd_sc_hd__nand3_1 _18512_ (.A(net3682),
    .B(_08948_),
    .C(_09000_),
    .Y(_09327_));
 sky130_fd_sc_hd__nand3_1 _18513_ (.A(net3956),
    .B(net3615),
    .C(_08994_),
    .Y(_09328_));
 sky130_fd_sc_hd__nand3_1 _18514_ (.A(_09057_),
    .B(_09327_),
    .C(_09328_),
    .Y(_09329_));
 sky130_fd_sc_hd__o221ai_1 _18515_ (.A1(_12134_[0]),
    .A2(_09178_),
    .B1(_09187_),
    .B2(_08818_),
    .C1(_09147_),
    .Y(_09330_));
 sky130_fd_sc_hd__nand2_2 _18516_ (.A(_09329_),
    .B(_09330_),
    .Y(_09331_));
 sky130_fd_sc_hd__o22ai_4 _18517_ (.A1(_09214_),
    .A2(_09324_),
    .B1(_09326_),
    .B2(_09331_),
    .Y(_09332_));
 sky130_fd_sc_hd__a21oi_1 _18518_ (.A1(_12134_[0]),
    .A2(net3956),
    .B1(_08965_),
    .Y(_09333_));
 sky130_fd_sc_hd__nand2_1 _18519_ (.A(_12150_[0]),
    .B(net3952),
    .Y(_09334_));
 sky130_fd_sc_hd__o21ai_1 _18520_ (.A1(net3952),
    .A2(_09333_),
    .B1(_09334_),
    .Y(_09335_));
 sky130_fd_sc_hd__nand3_1 _18521_ (.A(_12126_[0]),
    .B(_08818_),
    .C(net3946),
    .Y(_09336_));
 sky130_fd_sc_hd__o211ai_1 _18522_ (.A1(_12136_[0]),
    .A2(net3946),
    .B1(_09336_),
    .C1(_08827_),
    .Y(_09337_));
 sky130_fd_sc_hd__o2111a_1 _18523_ (.A1(_08827_),
    .A2(_09335_),
    .B1(_09337_),
    .C1(net3942),
    .D1(_09116_),
    .X(_09338_));
 sky130_fd_sc_hd__nor2_1 _18524_ (.A(_12124_[0]),
    .B(_08818_),
    .Y(_09339_));
 sky130_fd_sc_hd__a31oi_1 _18525_ (.A1(_08818_),
    .A2(_09013_),
    .A3(_09000_),
    .B1(_09339_),
    .Y(_09340_));
 sky130_fd_sc_hd__nor2_1 _18526_ (.A(net3942),
    .B(net3585),
    .Y(_09341_));
 sky130_fd_sc_hd__a2bb2oi_1 _18527_ (.A1_N(_08849_),
    .A2_N(_09340_),
    .B1(_09341_),
    .B2(_09265_),
    .Y(_09342_));
 sky130_fd_sc_hd__nor2_1 _18528_ (.A(_08951_),
    .B(_09342_),
    .Y(_09343_));
 sky130_fd_sc_hd__nand2_1 _18529_ (.A(_09116_),
    .B(_09112_),
    .Y(_09344_));
 sky130_fd_sc_hd__a21oi_1 _18530_ (.A1(_08818_),
    .A2(_08827_),
    .B1(net3957),
    .Y(_09345_));
 sky130_fd_sc_hd__o21ai_0 _18531_ (.A1(_08818_),
    .A2(_08827_),
    .B1(net3686),
    .Y(_09346_));
 sky130_fd_sc_hd__o32ai_1 _18532_ (.A1(net3686),
    .A2(_08827_),
    .A3(_09002_),
    .B1(_09345_),
    .B2(_09346_),
    .Y(_09347_));
 sky130_fd_sc_hd__a31o_1 _18533_ (.A1(_08818_),
    .A2(_08983_),
    .A3(_09076_),
    .B1(net3945),
    .X(_09348_));
 sky130_fd_sc_hd__a31oi_1 _18534_ (.A1(net3956),
    .A2(_08947_),
    .A3(_09029_),
    .B1(_09348_),
    .Y(_09349_));
 sky130_fd_sc_hd__a211o_1 _18535_ (.A1(_08941_),
    .A2(_09117_),
    .B1(_08818_),
    .C1(net3941),
    .X(_09350_));
 sky130_fd_sc_hd__o2111ai_1 _18536_ (.A1(_09016_),
    .A2(_09101_),
    .B1(_08818_),
    .C1(_08849_),
    .D1(_08901_),
    .Y(_09351_));
 sky130_fd_sc_hd__nand4_1 _18537_ (.A(net3955),
    .B(_08917_),
    .C(_09350_),
    .D(_09351_),
    .Y(_09352_));
 sky130_fd_sc_hd__nand2_1 _18538_ (.A(_12125_[0]),
    .B(net3937),
    .Y(_09353_));
 sky130_fd_sc_hd__o211ai_1 _18539_ (.A1(net3958),
    .A2(net3937),
    .B1(_09353_),
    .C1(_08818_),
    .Y(_09354_));
 sky130_fd_sc_hd__nand2_1 _18540_ (.A(_12129_[0]),
    .B(_08827_),
    .Y(_09355_));
 sky130_fd_sc_hd__o211ai_1 _18541_ (.A1(_12125_[0]),
    .A2(_08827_),
    .B1(_09355_),
    .C1(net3956),
    .Y(_09356_));
 sky130_fd_sc_hd__nand4_1 _18542_ (.A(_09116_),
    .B(_09166_),
    .C(_09354_),
    .D(_09356_),
    .Y(_09357_));
 sky130_fd_sc_hd__o221ai_2 _18543_ (.A1(_09344_),
    .A2(_09347_),
    .B1(_09349_),
    .B2(_09352_),
    .C1(_09357_),
    .Y(_09358_));
 sky130_fd_sc_hd__a2111oi_2 _18544_ (.A1(net3938),
    .A2(_09320_),
    .B1(_09338_),
    .C1(_09343_),
    .D1(_09358_),
    .Y(_09359_));
 sky130_fd_sc_hd__o21ai_4 _18545_ (.A1(_09321_),
    .A2(_09332_),
    .B1(_09359_),
    .Y(_00079_));
 sky130_fd_sc_hd__xnor3_1 _18546_ (.A(\sa12_sr[0] ),
    .B(net4201),
    .C(\sa02_sr[1] ),
    .X(_09360_));
 sky130_fd_sc_hd__xnor3_1 _18547_ (.A(_07075_),
    .B(_07108_),
    .C(_09360_),
    .X(_09361_));
 sky130_fd_sc_hd__mux2i_2 _18548_ (.A0(\text_in_r[49] ),
    .A1(_09361_),
    .S(net4111),
    .Y(_09362_));
 sky130_fd_sc_hd__xor2_4 _18549_ (.A(net4139),
    .B(_09362_),
    .X(_09363_));
 sky130_fd_sc_hd__inv_12 _18550_ (.A(_09363_),
    .Y(_09364_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_624 ();
 sky130_fd_sc_hd__xor2_1 _18553_ (.A(\sa02_sr[0] ),
    .B(\sa31_sub[0] ),
    .X(_09366_));
 sky130_fd_sc_hd__xor3_1 _18554_ (.A(net4201),
    .B(_07108_),
    .C(_09366_),
    .X(_09367_));
 sky130_fd_sc_hd__mux2i_1 _18555_ (.A0(\text_in_r[48] ),
    .A1(_09367_),
    .S(net4111),
    .Y(_09368_));
 sky130_fd_sc_hd__xor2_1 _18556_ (.A(\u0.w[2][16] ),
    .B(_09368_),
    .X(_09369_));
 sky130_fd_sc_hd__clkinv_16 _18557_ (.A(net3932),
    .Y(_09370_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_623 ();
 sky130_fd_sc_hd__xnor3_1 _18559_ (.A(\sa20_sub[1] ),
    .B(net4200),
    .C(net4224),
    .X(_09371_));
 sky130_fd_sc_hd__xor2_1 _18560_ (.A(_07096_),
    .B(_09371_),
    .X(_09372_));
 sky130_fd_sc_hd__mux2i_2 _18561_ (.A0(\text_in_r[50] ),
    .A1(_09372_),
    .S(net4111),
    .Y(_09373_));
 sky130_fd_sc_hd__xnor2_4 _18562_ (.A(\u0.w[2][18] ),
    .B(_09373_),
    .Y(_09374_));
 sky130_fd_sc_hd__clkinv_16 _18563_ (.A(_09374_),
    .Y(_09375_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_615 ();
 sky130_fd_sc_hd__xnor3_1 _18572_ (.A(net4199),
    .B(\sa20_sub[4] ),
    .C(\sa02_sr[4] ),
    .X(_09381_));
 sky130_fd_sc_hd__xnor3_1 _18573_ (.A(_07108_),
    .B(_07136_),
    .C(_09381_),
    .X(_09382_));
 sky130_fd_sc_hd__nand2_1 _18574_ (.A(net398),
    .B(\text_in_r[52] ),
    .Y(_09383_));
 sky130_fd_sc_hd__o21a_4 _18575_ (.A1(net398),
    .A2(_09382_),
    .B1(_09383_),
    .X(_09384_));
 sky130_fd_sc_hd__xor2_4 _18576_ (.A(net4138),
    .B(_09384_),
    .X(_09385_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_613 ();
 sky130_fd_sc_hd__xor2_1 _18579_ (.A(net4198),
    .B(\sa02_sr[5] ),
    .X(_09388_));
 sky130_fd_sc_hd__xnor2_1 _18580_ (.A(_07126_),
    .B(_09388_),
    .Y(_09389_));
 sky130_fd_sc_hd__mux2i_4 _18581_ (.A0(\text_in_r[53] ),
    .A1(_09389_),
    .S(net4112),
    .Y(_09390_));
 sky130_fd_sc_hd__xnor2_4 _18582_ (.A(\u0.w[2][21] ),
    .B(_09390_),
    .Y(_09391_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_609 ();
 sky130_fd_sc_hd__nor2b_1 _18587_ (.A(net4230),
    .B_N(\u0.w[2][19] ),
    .Y(_09396_));
 sky130_fd_sc_hd__nor2_1 _18588_ (.A(\u0.w[2][19] ),
    .B(net4230),
    .Y(_09397_));
 sky130_fd_sc_hd__xor2_1 _18589_ (.A(\sa20_sub[3] ),
    .B(net4196),
    .X(_09398_));
 sky130_fd_sc_hd__xor2_1 _18590_ (.A(net4200),
    .B(net4183),
    .X(_09399_));
 sky130_fd_sc_hd__xnor3_1 _18591_ (.A(\sa12_sr[7] ),
    .B(net4213),
    .C(\sa02_sr[3] ),
    .X(_09400_));
 sky130_fd_sc_hd__xnor3_1 _18592_ (.A(_09398_),
    .B(_09399_),
    .C(_09400_),
    .X(_09401_));
 sky130_fd_sc_hd__mux2_8 _18593_ (.A0(_09396_),
    .A1(_09397_),
    .S(_09401_),
    .X(_09402_));
 sky130_fd_sc_hd__nand2_1 _18594_ (.A(\u0.w[2][19] ),
    .B(net4230),
    .Y(_09403_));
 sky130_fd_sc_hd__nand3b_1 _18595_ (.A_N(\u0.w[2][19] ),
    .B(net4230),
    .C(\text_in_r[51] ),
    .Y(_09404_));
 sky130_fd_sc_hd__o21ai_2 _18596_ (.A1(\text_in_r[51] ),
    .A2(_09403_),
    .B1(_09404_),
    .Y(_09405_));
 sky130_fd_sc_hd__nor2_4 _18597_ (.A(_09402_),
    .B(_09405_),
    .Y(_09406_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_608 ();
 sky130_fd_sc_hd__nand2_8 _18599_ (.A(_09375_),
    .B(net3926),
    .Y(_09408_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_607 ();
 sky130_fd_sc_hd__nor2_4 _18601_ (.A(_12157_[0]),
    .B(_09406_),
    .Y(_09410_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_606 ();
 sky130_fd_sc_hd__or2_4 _18603_ (.A(_09402_),
    .B(_09405_),
    .X(_09412_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_604 ();
 sky130_fd_sc_hd__nor2_4 _18606_ (.A(_12166_[0]),
    .B(_09412_),
    .Y(_09415_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_603 ();
 sky130_fd_sc_hd__o21ai_0 _18608_ (.A1(_09410_),
    .A2(_09415_),
    .B1(net3931),
    .Y(_09417_));
 sky130_fd_sc_hd__o21ai_0 _18609_ (.A1(_12161_[0]),
    .A2(_09408_),
    .B1(_09417_),
    .Y(_09418_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_602 ();
 sky130_fd_sc_hd__nor2_4 _18611_ (.A(_12158_[0]),
    .B(_09412_),
    .Y(_09420_));
 sky130_fd_sc_hd__nor2_1 _18612_ (.A(_12161_[0]),
    .B(_09406_),
    .Y(_09421_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_600 ();
 sky130_fd_sc_hd__o21ai_2 _18615_ (.A1(_09420_),
    .A2(net3584),
    .B1(net3931),
    .Y(_09424_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_598 ();
 sky130_fd_sc_hd__nor2_4 _18618_ (.A(net3931),
    .B(_09412_),
    .Y(_09427_));
 sky130_fd_sc_hd__nand2_1 _18619_ (.A(_12156_[0]),
    .B(_09427_),
    .Y(_09428_));
 sky130_fd_sc_hd__nand3_1 _18620_ (.A(net3927),
    .B(_09424_),
    .C(_09428_),
    .Y(_09429_));
 sky130_fd_sc_hd__o21ai_0 _18621_ (.A1(net3927),
    .A2(_09418_),
    .B1(_09429_),
    .Y(_09430_));
 sky130_fd_sc_hd__xnor2_4 _18622_ (.A(net4138),
    .B(_09384_),
    .Y(_09431_));
 sky130_fd_sc_hd__xor2_4 _18623_ (.A(\u0.w[2][21] ),
    .B(_09390_),
    .X(_09432_));
 sky130_fd_sc_hd__nor2_4 _18624_ (.A(_09431_),
    .B(_09432_),
    .Y(_09433_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_596 ();
 sky130_fd_sc_hd__nor2_4 _18627_ (.A(net3936),
    .B(_09375_),
    .Y(_09436_));
 sky130_fd_sc_hd__a211o_1 _18628_ (.A1(_12157_[0]),
    .A2(_09375_),
    .B1(net3917),
    .C1(_09436_),
    .X(_09437_));
 sky130_fd_sc_hd__nor2_4 _18629_ (.A(net3934),
    .B(_09375_),
    .Y(_09438_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_595 ();
 sky130_fd_sc_hd__nor2_1 _18631_ (.A(_12164_[0]),
    .B(net3931),
    .Y(_09440_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_593 ();
 sky130_fd_sc_hd__o21ai_0 _18634_ (.A1(_09438_),
    .A2(_09440_),
    .B1(net3917),
    .Y(_09443_));
 sky130_fd_sc_hd__nand3_2 _18635_ (.A(_09433_),
    .B(_09437_),
    .C(_09443_),
    .Y(_09444_));
 sky130_fd_sc_hd__o21ai_4 _18636_ (.A1(net3936),
    .A2(net3934),
    .B1(net3917),
    .Y(_09445_));
 sky130_fd_sc_hd__nand2_8 _18637_ (.A(_09370_),
    .B(net3915),
    .Y(_09446_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_592 ();
 sky130_fd_sc_hd__nand2_1 _18639_ (.A(_12161_[0]),
    .B(net3926),
    .Y(_09448_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_590 ();
 sky130_fd_sc_hd__a21o_1 _18642_ (.A1(_09446_),
    .A2(_09448_),
    .B1(net3931),
    .X(_09451_));
 sky130_fd_sc_hd__nor2_4 _18643_ (.A(_09431_),
    .B(_09391_),
    .Y(_09452_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_589 ();
 sky130_fd_sc_hd__o211ai_1 _18645_ (.A1(_09375_),
    .A2(_09445_),
    .B1(_09451_),
    .C1(_09452_),
    .Y(_09454_));
 sky130_fd_sc_hd__xor2_2 _18646_ (.A(\sa31_sub[6] ),
    .B(\sa02_sr[6] ),
    .X(_09455_));
 sky130_fd_sc_hd__xnor3_1 _18647_ (.A(\sa12_sr[5] ),
    .B(net4197),
    .C(\sa20_sub[6] ),
    .X(_09456_));
 sky130_fd_sc_hd__xnor2_1 _18648_ (.A(_09455_),
    .B(_09456_),
    .Y(_09457_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_588 ();
 sky130_fd_sc_hd__mux2i_4 _18650_ (.A0(\text_in_r[54] ),
    .A1(_09457_),
    .S(net4112),
    .Y(_09459_));
 sky130_fd_sc_hd__xnor2_4 _18651_ (.A(\u0.w[2][22] ),
    .B(_09459_),
    .Y(_09460_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_587 ();
 sky130_fd_sc_hd__o2111ai_1 _18653_ (.A1(net3929),
    .A2(_09430_),
    .B1(_09444_),
    .C1(_09454_),
    .D1(_09460_),
    .Y(_09462_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_585 ();
 sky130_fd_sc_hd__nor3_1 _18656_ (.A(net3935),
    .B(_09370_),
    .C(net3923),
    .Y(_09465_));
 sky130_fd_sc_hd__nor2_4 _18657_ (.A(net3931),
    .B(net3920),
    .Y(_09466_));
 sky130_fd_sc_hd__nand2_2 _18658_ (.A(_12166_[0]),
    .B(_09466_),
    .Y(_09467_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_583 ();
 sky130_fd_sc_hd__o311ai_0 _18661_ (.A1(net3677),
    .A2(net3613),
    .A3(_09420_),
    .B1(_09467_),
    .C1(net3930),
    .Y(_09470_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_581 ();
 sky130_fd_sc_hd__nor2_4 _18664_ (.A(_12164_[0]),
    .B(_09408_),
    .Y(_09473_));
 sky130_fd_sc_hd__nor3_4 _18665_ (.A(net3936),
    .B(_09370_),
    .C(_09412_),
    .Y(_09474_));
 sky130_fd_sc_hd__nor2_2 _18666_ (.A(_12158_[0]),
    .B(net3925),
    .Y(_09475_));
 sky130_fd_sc_hd__nor3_1 _18667_ (.A(_09375_),
    .B(_09474_),
    .C(_09475_),
    .Y(_09476_));
 sky130_fd_sc_hd__nor3_1 _18668_ (.A(net3929),
    .B(_09473_),
    .C(_09476_),
    .Y(_09477_));
 sky130_fd_sc_hd__nor3_1 _18669_ (.A(_09460_),
    .B(_09432_),
    .C(_09477_),
    .Y(_09478_));
 sky130_fd_sc_hd__nor2_4 _18670_ (.A(net3933),
    .B(net3931),
    .Y(_09479_));
 sky130_fd_sc_hd__nor2_1 _18671_ (.A(_12156_[0]),
    .B(_09375_),
    .Y(_09480_));
 sky130_fd_sc_hd__o21ai_2 _18672_ (.A1(_09479_),
    .A2(_09480_),
    .B1(net3914),
    .Y(_09481_));
 sky130_fd_sc_hd__nor2_4 _18673_ (.A(_12158_[0]),
    .B(_12161_[0]),
    .Y(_09482_));
 sky130_fd_sc_hd__nor3_2 _18674_ (.A(net3936),
    .B(_09370_),
    .C(_09375_),
    .Y(_09483_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_580 ();
 sky130_fd_sc_hd__a211o_1 _18676_ (.A1(_09375_),
    .A2(_09482_),
    .B1(_09483_),
    .C1(net3917),
    .X(_09485_));
 sky130_fd_sc_hd__xor2_4 _18677_ (.A(\u0.w[2][22] ),
    .B(_09459_),
    .X(_09486_));
 sky130_fd_sc_hd__nand2_1 _18678_ (.A(_09486_),
    .B(_09432_),
    .Y(_09487_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_579 ();
 sky130_fd_sc_hd__a221oi_1 _18680_ (.A1(_12177_[0]),
    .A2(net3917),
    .B1(_09427_),
    .B2(_12157_[0]),
    .C1(net3929),
    .Y(_09489_));
 sky130_fd_sc_hd__a311oi_1 _18681_ (.A1(net3929),
    .A2(_09481_),
    .A3(_09485_),
    .B1(_09487_),
    .C1(_09489_),
    .Y(_09490_));
 sky130_fd_sc_hd__xor2_1 _18682_ (.A(\sa20_sub[6] ),
    .B(\sa31_sub[7] ),
    .X(_09491_));
 sky130_fd_sc_hd__xnor2_1 _18683_ (.A(\sa12_sr[6] ),
    .B(net4196),
    .Y(_09492_));
 sky130_fd_sc_hd__xnor2_1 _18684_ (.A(_09491_),
    .B(_09492_),
    .Y(_09493_));
 sky130_fd_sc_hd__xnor2_1 _18685_ (.A(net4223),
    .B(_09493_),
    .Y(_09494_));
 sky130_fd_sc_hd__nor2_1 _18686_ (.A(net398),
    .B(_09494_),
    .Y(_09495_));
 sky130_fd_sc_hd__a21oi_4 _18687_ (.A1(net398),
    .A2(\text_in_r[55] ),
    .B1(_09495_),
    .Y(_09496_));
 sky130_fd_sc_hd__xor2_4 _18688_ (.A(\u0.w[2][23] ),
    .B(_09496_),
    .X(_09497_));
 sky130_fd_sc_hd__a211oi_1 _18689_ (.A1(_09470_),
    .A2(_09478_),
    .B1(_09490_),
    .C1(_09497_),
    .Y(_09498_));
 sky130_fd_sc_hd__nand2_4 _18690_ (.A(_09486_),
    .B(net3912),
    .Y(_09499_));
 sky130_fd_sc_hd__nor3_1 _18691_ (.A(net3934),
    .B(net3931),
    .C(_09412_),
    .Y(_09500_));
 sky130_fd_sc_hd__nand3_1 _18692_ (.A(_09364_),
    .B(_09499_),
    .C(_09500_),
    .Y(_09501_));
 sky130_fd_sc_hd__xnor2_2 _18693_ (.A(_09375_),
    .B(net3926),
    .Y(_09502_));
 sky130_fd_sc_hd__nor2_1 _18694_ (.A(net3934),
    .B(_09502_),
    .Y(_09503_));
 sky130_fd_sc_hd__nand2_4 _18695_ (.A(net3933),
    .B(net3925),
    .Y(_09504_));
 sky130_fd_sc_hd__nor2_2 _18696_ (.A(_09364_),
    .B(_09504_),
    .Y(_09505_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_578 ();
 sky130_fd_sc_hd__nor2_1 _18698_ (.A(_12157_[0]),
    .B(_09412_),
    .Y(_09507_));
 sky130_fd_sc_hd__a21oi_1 _18699_ (.A1(_12164_[0]),
    .A2(_09412_),
    .B1(_09507_),
    .Y(_09508_));
 sky130_fd_sc_hd__nand2_4 _18700_ (.A(_09486_),
    .B(net3929),
    .Y(_09509_));
 sky130_fd_sc_hd__a21oi_1 _18701_ (.A1(_12156_[0]),
    .A2(_09466_),
    .B1(_09509_),
    .Y(_09510_));
 sky130_fd_sc_hd__o21ai_0 _18702_ (.A1(_09375_),
    .A2(_09508_),
    .B1(_09510_),
    .Y(_09511_));
 sky130_fd_sc_hd__o41ai_1 _18703_ (.A1(_09499_),
    .A2(_09503_),
    .A3(_09505_),
    .A4(net3613),
    .B1(_09511_),
    .Y(_09512_));
 sky130_fd_sc_hd__nand2_4 _18704_ (.A(net3931),
    .B(net3917),
    .Y(_09513_));
 sky130_fd_sc_hd__nor2_4 _18705_ (.A(_09364_),
    .B(net3919),
    .Y(_09514_));
 sky130_fd_sc_hd__nand2_1 _18706_ (.A(net3934),
    .B(_09375_),
    .Y(_09515_));
 sky130_fd_sc_hd__o22ai_1 _18707_ (.A1(_12161_[0]),
    .A2(_09513_),
    .B1(_09514_),
    .B2(_09515_),
    .Y(_09516_));
 sky130_fd_sc_hd__nor2_1 _18708_ (.A(_09364_),
    .B(_09412_),
    .Y(_09517_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_577 ();
 sky130_fd_sc_hd__and2_4 _18710_ (.A(_12170_[0]),
    .B(_09412_),
    .X(_09519_));
 sky130_fd_sc_hd__o21ai_0 _18711_ (.A1(_09517_),
    .A2(_09519_),
    .B1(_09375_),
    .Y(_09520_));
 sky130_fd_sc_hd__and3_4 _18712_ (.A(_12157_[0]),
    .B(net3931),
    .C(_09412_),
    .X(_09521_));
 sky130_fd_sc_hd__nor2_4 _18713_ (.A(net3933),
    .B(_09412_),
    .Y(_09522_));
 sky130_fd_sc_hd__nor3_1 _18714_ (.A(net3929),
    .B(_09521_),
    .C(_09522_),
    .Y(_09523_));
 sky130_fd_sc_hd__a221oi_1 _18715_ (.A1(net3929),
    .A2(_09516_),
    .B1(_09520_),
    .B2(_09523_),
    .C1(_09486_),
    .Y(_09524_));
 sky130_fd_sc_hd__xnor2_4 _18716_ (.A(\u0.w[2][23] ),
    .B(_09496_),
    .Y(_09525_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_576 ();
 sky130_fd_sc_hd__a2111oi_0 _18718_ (.A1(_09501_),
    .A2(_09512_),
    .B1(_09524_),
    .C1(_09432_),
    .D1(_09525_),
    .Y(_09527_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_573 ();
 sky130_fd_sc_hd__nor2_4 _18722_ (.A(net3935),
    .B(_09412_),
    .Y(_09531_));
 sky130_fd_sc_hd__o32ai_1 _18723_ (.A1(_09375_),
    .A2(_09519_),
    .A3(_09531_),
    .B1(_09515_),
    .B2(net3612),
    .Y(_09532_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_572 ();
 sky130_fd_sc_hd__nand2_4 _18725_ (.A(net3935),
    .B(net3921),
    .Y(_09534_));
 sky130_fd_sc_hd__nor2_2 _18726_ (.A(_12157_[0]),
    .B(net3931),
    .Y(_09535_));
 sky130_fd_sc_hd__nor2_2 _18727_ (.A(net3678),
    .B(net3931),
    .Y(_09536_));
 sky130_fd_sc_hd__nand2_8 _18728_ (.A(_12157_[0]),
    .B(net3920),
    .Y(_09537_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_571 ();
 sky130_fd_sc_hd__o2bb2ai_1 _18730_ (.A1_N(_09534_),
    .A2_N(_09535_),
    .B1(_09536_),
    .B2(_09537_),
    .Y(_09539_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_569 ();
 sky130_fd_sc_hd__o21ai_0 _18733_ (.A1(_09460_),
    .A2(_09539_),
    .B1(net3912),
    .Y(_09542_));
 sky130_fd_sc_hd__a21oi_1 _18734_ (.A1(_09460_),
    .A2(_09532_),
    .B1(_09542_),
    .Y(_09543_));
 sky130_fd_sc_hd__nand2_4 _18735_ (.A(_09460_),
    .B(net3929),
    .Y(_09544_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_568 ();
 sky130_fd_sc_hd__nand2_2 _18737_ (.A(net3931),
    .B(net3919),
    .Y(_09546_));
 sky130_fd_sc_hd__nand2_1 _18738_ (.A(net3934),
    .B(_09466_),
    .Y(_09547_));
 sky130_fd_sc_hd__o21ai_0 _18739_ (.A1(_12158_[0]),
    .A2(_09546_),
    .B1(_09547_),
    .Y(_09548_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_566 ();
 sky130_fd_sc_hd__a21oi_1 _18742_ (.A1(_09412_),
    .A2(_09438_),
    .B1(_09427_),
    .Y(_09550_));
 sky130_fd_sc_hd__nor2_1 _18743_ (.A(net3936),
    .B(_09550_),
    .Y(_09551_));
 sky130_fd_sc_hd__nor2_1 _18744_ (.A(_12156_[0]),
    .B(_09502_),
    .Y(_09552_));
 sky130_fd_sc_hd__nor3_1 _18745_ (.A(_09521_),
    .B(_09473_),
    .C(_09552_),
    .Y(_09553_));
 sky130_fd_sc_hd__o32ai_1 _18746_ (.A1(_09544_),
    .A2(_09548_),
    .A3(_09551_),
    .B1(_09553_),
    .B2(_09509_),
    .Y(_09554_));
 sky130_fd_sc_hd__nor4_1 _18747_ (.A(net3927),
    .B(_09525_),
    .C(_09543_),
    .D(_09554_),
    .Y(_09555_));
 sky130_fd_sc_hd__a211oi_1 _18748_ (.A1(_09462_),
    .A2(_09498_),
    .B1(_09527_),
    .C1(_09555_),
    .Y(_00080_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_565 ();
 sky130_fd_sc_hd__nor2_1 _18750_ (.A(_09522_),
    .B(_09421_),
    .Y(_09557_));
 sky130_fd_sc_hd__nor2_1 _18751_ (.A(_12156_[0]),
    .B(_09412_),
    .Y(_09558_));
 sky130_fd_sc_hd__nand2_8 _18752_ (.A(net3678),
    .B(_09412_),
    .Y(_09559_));
 sky130_fd_sc_hd__nand3b_1 _18753_ (.A_N(_09558_),
    .B(net3677),
    .C(_09559_),
    .Y(_09560_));
 sky130_fd_sc_hd__o21ai_0 _18754_ (.A1(net3677),
    .A2(_09557_),
    .B1(_09560_),
    .Y(_09561_));
 sky130_fd_sc_hd__a21oi_1 _18755_ (.A1(net3678),
    .A2(_09522_),
    .B1(_09410_),
    .Y(_09562_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_564 ();
 sky130_fd_sc_hd__nand3_1 _18757_ (.A(net3933),
    .B(_09375_),
    .C(net3926),
    .Y(_09564_));
 sky130_fd_sc_hd__o21ai_1 _18758_ (.A1(_09375_),
    .A2(_09562_),
    .B1(_09564_),
    .Y(_09565_));
 sky130_fd_sc_hd__nor2_4 _18759_ (.A(_09370_),
    .B(_09412_),
    .Y(_09566_));
 sky130_fd_sc_hd__and2_0 _18760_ (.A(_12156_[0]),
    .B(_09412_),
    .X(_09567_));
 sky130_fd_sc_hd__o21ai_0 _18761_ (.A1(_12158_[0]),
    .A2(_09412_),
    .B1(net3931),
    .Y(_09568_));
 sky130_fd_sc_hd__o32ai_1 _18762_ (.A1(net3931),
    .A2(_09566_),
    .A3(_09410_),
    .B1(_09567_),
    .B2(_09568_),
    .Y(_09569_));
 sky130_fd_sc_hd__nor3_2 _18763_ (.A(net3935),
    .B(net3933),
    .C(net3923),
    .Y(_09570_));
 sky130_fd_sc_hd__o21ai_1 _18764_ (.A1(_09420_),
    .A2(_09570_),
    .B1(net3677),
    .Y(_09571_));
 sky130_fd_sc_hd__nand2b_4 _18765_ (.A_N(_12157_[0]),
    .B(_09412_),
    .Y(_09572_));
 sky130_fd_sc_hd__nand2_4 _18766_ (.A(_12170_[0]),
    .B(net3922),
    .Y(_09573_));
 sky130_fd_sc_hd__a31oi_1 _18767_ (.A1(net3931),
    .A2(_09572_),
    .A3(_09573_),
    .B1(_09391_),
    .Y(_09574_));
 sky130_fd_sc_hd__a221oi_1 _18768_ (.A1(_09391_),
    .A2(_09569_),
    .B1(_09571_),
    .B2(_09574_),
    .C1(net3930),
    .Y(_09575_));
 sky130_fd_sc_hd__a221oi_1 _18769_ (.A1(_09433_),
    .A2(_09561_),
    .B1(_09565_),
    .B2(_09452_),
    .C1(_09575_),
    .Y(_09576_));
 sky130_fd_sc_hd__nor3_1 _18770_ (.A(_09486_),
    .B(_09525_),
    .C(_09576_),
    .Y(_09577_));
 sky130_fd_sc_hd__nor2_4 _18771_ (.A(net3929),
    .B(net3910),
    .Y(_09578_));
 sky130_fd_sc_hd__o21ai_0 _18772_ (.A1(_12161_[0]),
    .A2(_09412_),
    .B1(_09572_),
    .Y(_09579_));
 sky130_fd_sc_hd__nor2_4 _18773_ (.A(_09370_),
    .B(_09406_),
    .Y(_09580_));
 sky130_fd_sc_hd__or3_4 _18774_ (.A(net3931),
    .B(_09580_),
    .C(_09522_),
    .X(_09581_));
 sky130_fd_sc_hd__o21ai_0 _18775_ (.A1(net3677),
    .A2(_09579_),
    .B1(_09581_),
    .Y(_09582_));
 sky130_fd_sc_hd__nor2_4 _18776_ (.A(_09375_),
    .B(net3918),
    .Y(_09583_));
 sky130_fd_sc_hd__nand2_2 _18777_ (.A(_09385_),
    .B(_09391_),
    .Y(_09584_));
 sky130_fd_sc_hd__nand2_1 _18778_ (.A(net3933),
    .B(_09412_),
    .Y(_09585_));
 sky130_fd_sc_hd__a21oi_1 _18779_ (.A1(net3677),
    .A2(_09585_),
    .B1(net3935),
    .Y(_09586_));
 sky130_fd_sc_hd__nor4_1 _18780_ (.A(_09505_),
    .B(_09583_),
    .C(_09584_),
    .D(_09586_),
    .Y(_09587_));
 sky130_fd_sc_hd__nand2_2 _18781_ (.A(_09486_),
    .B(_09525_),
    .Y(_09588_));
 sky130_fd_sc_hd__nor2_4 _18782_ (.A(_12170_[0]),
    .B(net3926),
    .Y(_09589_));
 sky130_fd_sc_hd__nor3_1 _18783_ (.A(_09375_),
    .B(_09589_),
    .C(_09474_),
    .Y(_09590_));
 sky130_fd_sc_hd__nor2_2 _18784_ (.A(_12161_[0]),
    .B(_09412_),
    .Y(_09591_));
 sky130_fd_sc_hd__nor3_1 _18785_ (.A(net3931),
    .B(_09410_),
    .C(_09591_),
    .Y(_09592_));
 sky130_fd_sc_hd__o21ai_0 _18786_ (.A1(_09590_),
    .A2(_09592_),
    .B1(net3929),
    .Y(_09593_));
 sky130_fd_sc_hd__o221ai_1 _18787_ (.A1(net3936),
    .A2(_09502_),
    .B1(_09408_),
    .B2(_12161_[0]),
    .C1(net3912),
    .Y(_09594_));
 sky130_fd_sc_hd__a21oi_1 _18788_ (.A1(_09593_),
    .A2(_09594_),
    .B1(net3927),
    .Y(_09595_));
 sky130_fd_sc_hd__a2111oi_0 _18789_ (.A1(_09578_),
    .A2(_09582_),
    .B1(_09587_),
    .C1(_09588_),
    .D1(_09595_),
    .Y(_09596_));
 sky130_fd_sc_hd__and3_1 _18790_ (.A(net3931),
    .B(_09572_),
    .C(_09448_),
    .X(_09597_));
 sky130_fd_sc_hd__a21oi_1 _18791_ (.A1(_09375_),
    .A2(_09445_),
    .B1(_09597_),
    .Y(_09598_));
 sky130_fd_sc_hd__o22ai_1 _18792_ (.A1(_09370_),
    .A2(_09502_),
    .B1(_09446_),
    .B2(_09364_),
    .Y(_09599_));
 sky130_fd_sc_hd__a211oi_1 _18793_ (.A1(_12157_[0]),
    .A2(_09427_),
    .B1(net3927),
    .C1(_09599_),
    .Y(_09600_));
 sky130_fd_sc_hd__a211o_1 _18794_ (.A1(net3927),
    .A2(_09598_),
    .B1(_09600_),
    .C1(_09544_),
    .X(_09601_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_563 ();
 sky130_fd_sc_hd__o21ai_0 _18796_ (.A1(_09566_),
    .A2(net3584),
    .B1(_09375_),
    .Y(_09603_));
 sky130_fd_sc_hd__a31oi_1 _18797_ (.A1(_12156_[0]),
    .A2(net3931),
    .A3(net3926),
    .B1(_09521_),
    .Y(_09604_));
 sky130_fd_sc_hd__nand3_1 _18798_ (.A(net3910),
    .B(_09603_),
    .C(_09604_),
    .Y(_09605_));
 sky130_fd_sc_hd__nand3_4 _18799_ (.A(net3678),
    .B(_09370_),
    .C(_09406_),
    .Y(_09606_));
 sky130_fd_sc_hd__a2bb2oi_1 _18800_ (.A1_N(net3931),
    .A2_N(_09519_),
    .B1(_09583_),
    .B2(net3936),
    .Y(_09607_));
 sky130_fd_sc_hd__nand2_4 _18801_ (.A(_09460_),
    .B(net3912),
    .Y(_09608_));
 sky130_fd_sc_hd__a31oi_1 _18802_ (.A1(net3927),
    .A2(_09606_),
    .A3(_09607_),
    .B1(_09608_),
    .Y(_09609_));
 sky130_fd_sc_hd__nand2_1 _18803_ (.A(_09605_),
    .B(_09609_),
    .Y(_09610_));
 sky130_fd_sc_hd__a21oi_1 _18804_ (.A1(_09601_),
    .A2(_09610_),
    .B1(_09497_),
    .Y(_09611_));
 sky130_fd_sc_hd__nand2_4 _18805_ (.A(_09486_),
    .B(_09497_),
    .Y(_09612_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_562 ();
 sky130_fd_sc_hd__nor2_1 _18807_ (.A(net3935),
    .B(net3933),
    .Y(_09614_));
 sky130_fd_sc_hd__nand2_1 _18808_ (.A(net3931),
    .B(_09614_),
    .Y(_09615_));
 sky130_fd_sc_hd__nand2_2 _18809_ (.A(_12164_[0]),
    .B(_09375_),
    .Y(_09616_));
 sky130_fd_sc_hd__nor3_1 _18810_ (.A(_12180_[0]),
    .B(net3920),
    .C(_09391_),
    .Y(_09617_));
 sky130_fd_sc_hd__a31oi_1 _18811_ (.A1(net3921),
    .A2(_09615_),
    .A3(_09616_),
    .B1(_09617_),
    .Y(_09618_));
 sky130_fd_sc_hd__nor2_1 _18812_ (.A(net3911),
    .B(_09618_),
    .Y(_09619_));
 sky130_fd_sc_hd__nor2_4 _18813_ (.A(_09370_),
    .B(_09375_),
    .Y(_09620_));
 sky130_fd_sc_hd__a21oi_1 _18814_ (.A1(_12156_[0]),
    .A2(_09375_),
    .B1(_09620_),
    .Y(_09621_));
 sky130_fd_sc_hd__o32ai_2 _18815_ (.A1(_09479_),
    .A2(_09559_),
    .A3(_09620_),
    .B1(_09621_),
    .B2(net3913),
    .Y(_09622_));
 sky130_fd_sc_hd__nor3_1 _18816_ (.A(net3931),
    .B(_09514_),
    .C(_09531_),
    .Y(_09623_));
 sky130_fd_sc_hd__a211oi_1 _18817_ (.A1(net3931),
    .A2(_09557_),
    .B1(_09623_),
    .C1(net3928),
    .Y(_09624_));
 sky130_fd_sc_hd__a211oi_1 _18818_ (.A1(net3928),
    .A2(_09622_),
    .B1(_09624_),
    .C1(net3930),
    .Y(_09625_));
 sky130_fd_sc_hd__nor3_1 _18819_ (.A(_09612_),
    .B(_09619_),
    .C(_09625_),
    .Y(_09626_));
 sky130_fd_sc_hd__nor4_1 _18820_ (.A(_09577_),
    .B(_09596_),
    .C(_09611_),
    .D(_09626_),
    .Y(_00081_));
 sky130_fd_sc_hd__nor3_1 _18821_ (.A(_09375_),
    .B(_09580_),
    .C(_09415_),
    .Y(_09627_));
 sky130_fd_sc_hd__nor2_4 _18822_ (.A(_12170_[0]),
    .B(_09412_),
    .Y(_09628_));
 sky130_fd_sc_hd__nor3_1 _18823_ (.A(net3931),
    .B(net3584),
    .C(_09628_),
    .Y(_09629_));
 sky130_fd_sc_hd__nor2_2 _18824_ (.A(net3930),
    .B(net3928),
    .Y(_09630_));
 sky130_fd_sc_hd__o21ai_0 _18825_ (.A1(_09627_),
    .A2(_09629_),
    .B1(_09630_),
    .Y(_09631_));
 sky130_fd_sc_hd__nand2_1 _18826_ (.A(_12166_[0]),
    .B(net3924),
    .Y(_09632_));
 sky130_fd_sc_hd__nand3_1 _18827_ (.A(net3931),
    .B(_09559_),
    .C(_09632_),
    .Y(_09633_));
 sky130_fd_sc_hd__o211ai_1 _18828_ (.A1(_12161_[0]),
    .A2(net3931),
    .B1(_09452_),
    .C1(_09633_),
    .Y(_09634_));
 sky130_fd_sc_hd__o21ai_0 _18829_ (.A1(_09566_),
    .A2(_09410_),
    .B1(net3931),
    .Y(_09635_));
 sky130_fd_sc_hd__nand3_1 _18830_ (.A(_09375_),
    .B(_09572_),
    .C(_09632_),
    .Y(_09636_));
 sky130_fd_sc_hd__nand2_1 _18831_ (.A(net3678),
    .B(_09375_),
    .Y(_09637_));
 sky130_fd_sc_hd__o21ai_0 _18832_ (.A1(_12166_[0]),
    .A2(_09375_),
    .B1(_09637_),
    .Y(_09638_));
 sky130_fd_sc_hd__a211oi_1 _18833_ (.A1(_12170_[0]),
    .A2(_09375_),
    .B1(_09412_),
    .C1(_09438_),
    .Y(_09639_));
 sky130_fd_sc_hd__a21oi_1 _18834_ (.A1(_09412_),
    .A2(_09638_),
    .B1(_09639_),
    .Y(_09640_));
 sky130_fd_sc_hd__a32oi_1 _18835_ (.A1(_09433_),
    .A2(_09635_),
    .A3(_09636_),
    .B1(_09640_),
    .B2(_09578_),
    .Y(_09641_));
 sky130_fd_sc_hd__a41o_4 _18836_ (.A1(_09460_),
    .A2(_09631_),
    .A3(_09634_),
    .A4(_09641_),
    .B1(_09525_),
    .X(_09642_));
 sky130_fd_sc_hd__nor2_4 _18837_ (.A(_09375_),
    .B(_09412_),
    .Y(_09643_));
 sky130_fd_sc_hd__nand2_1 _18838_ (.A(_09446_),
    .B(_09573_),
    .Y(_09644_));
 sky130_fd_sc_hd__a221oi_1 _18839_ (.A1(_12161_[0]),
    .A2(_09643_),
    .B1(_09644_),
    .B2(_09375_),
    .C1(_09514_),
    .Y(_09645_));
 sky130_fd_sc_hd__a21oi_1 _18840_ (.A1(_09537_),
    .A2(_09446_),
    .B1(_09375_),
    .Y(_09646_));
 sky130_fd_sc_hd__nor3_1 _18841_ (.A(net3931),
    .B(_09531_),
    .C(_09475_),
    .Y(_09647_));
 sky130_fd_sc_hd__o21ai_0 _18842_ (.A1(_09646_),
    .A2(_09647_),
    .B1(net3927),
    .Y(_09648_));
 sky130_fd_sc_hd__o21ai_2 _18843_ (.A1(net3927),
    .A2(_09645_),
    .B1(_09648_),
    .Y(_09649_));
 sky130_fd_sc_hd__o21ai_0 _18844_ (.A1(_12161_[0]),
    .A2(net3931),
    .B1(net3929),
    .Y(_09650_));
 sky130_fd_sc_hd__o22ai_2 _18845_ (.A1(net3917),
    .A2(net3912),
    .B1(_09483_),
    .B2(_09650_),
    .Y(_09651_));
 sky130_fd_sc_hd__o221a_1 _18846_ (.A1(_12170_[0]),
    .A2(_09513_),
    .B1(_09581_),
    .B2(net3936),
    .C1(_09433_),
    .X(_09652_));
 sky130_fd_sc_hd__a311o_1 _18847_ (.A1(_09432_),
    .A2(_09437_),
    .A3(_09651_),
    .B1(_09652_),
    .C1(_09460_),
    .X(_09653_));
 sky130_fd_sc_hd__a21oi_1 _18848_ (.A1(net3912),
    .A2(_09649_),
    .B1(_09653_),
    .Y(_09654_));
 sky130_fd_sc_hd__nor3_1 _18849_ (.A(net3918),
    .B(_09535_),
    .C(_09483_),
    .Y(_09655_));
 sky130_fd_sc_hd__a21oi_1 _18850_ (.A1(_12177_[0]),
    .A2(net3918),
    .B1(_09486_),
    .Y(_09656_));
 sky130_fd_sc_hd__nand2_1 _18851_ (.A(_09433_),
    .B(_09656_),
    .Y(_09657_));
 sky130_fd_sc_hd__o21ai_0 _18852_ (.A1(_09655_),
    .A2(_09657_),
    .B1(_09525_),
    .Y(_09658_));
 sky130_fd_sc_hd__nor2_2 _18853_ (.A(net3935),
    .B(_09370_),
    .Y(_09659_));
 sky130_fd_sc_hd__o21ai_0 _18854_ (.A1(_12184_[0]),
    .A2(_09385_),
    .B1(net3919),
    .Y(_09660_));
 sky130_fd_sc_hd__a31oi_1 _18855_ (.A1(_09375_),
    .A2(_09385_),
    .A3(_09659_),
    .B1(_09660_),
    .Y(_09661_));
 sky130_fd_sc_hd__a21oi_1 _18856_ (.A1(_12175_[0]),
    .A2(_09385_),
    .B1(net3919),
    .Y(_09662_));
 sky130_fd_sc_hd__o31a_1 _18857_ (.A1(net3935),
    .A2(_09385_),
    .A3(_09479_),
    .B1(_09662_),
    .X(_09663_));
 sky130_fd_sc_hd__nor2_1 _18858_ (.A(_09364_),
    .B(_09370_),
    .Y(_09664_));
 sky130_fd_sc_hd__or3_1 _18859_ (.A(net3919),
    .B(_09436_),
    .C(_09664_),
    .X(_09665_));
 sky130_fd_sc_hd__o21ai_0 _18860_ (.A1(_12180_[0]),
    .A2(net3913),
    .B1(_09665_),
    .Y(_09666_));
 sky130_fd_sc_hd__o32a_1 _18861_ (.A1(_09460_),
    .A2(_09661_),
    .A3(_09663_),
    .B1(_09666_),
    .B2(_09544_),
    .X(_09667_));
 sky130_fd_sc_hd__nand2_4 _18862_ (.A(_12164_[0]),
    .B(net3914),
    .Y(_09668_));
 sky130_fd_sc_hd__nand3_1 _18863_ (.A(net3931),
    .B(_09668_),
    .C(_09534_),
    .Y(_09669_));
 sky130_fd_sc_hd__a21oi_2 _18864_ (.A1(_12156_[0]),
    .A2(net3924),
    .B1(net3931),
    .Y(_09670_));
 sky130_fd_sc_hd__a21oi_1 _18865_ (.A1(_09572_),
    .A2(_09670_),
    .B1(_09608_),
    .Y(_09671_));
 sky130_fd_sc_hd__nand2_2 _18866_ (.A(_09669_),
    .B(_09671_),
    .Y(_09672_));
 sky130_fd_sc_hd__nand2_4 _18867_ (.A(net3917),
    .B(_09482_),
    .Y(_09673_));
 sky130_fd_sc_hd__a21oi_2 _18868_ (.A1(_09606_),
    .A2(_09673_),
    .B1(_09375_),
    .Y(_09674_));
 sky130_fd_sc_hd__or3_4 _18869_ (.A(_12164_[0]),
    .B(_09402_),
    .C(_09405_),
    .X(_09675_));
 sky130_fd_sc_hd__and3_1 _18870_ (.A(_09375_),
    .B(_09445_),
    .C(_09675_),
    .X(_09676_));
 sky130_fd_sc_hd__o21bai_1 _18871_ (.A1(_09674_),
    .A2(_09676_),
    .B1_N(_09499_),
    .Y(_09677_));
 sky130_fd_sc_hd__nor3_1 _18872_ (.A(_12157_[0]),
    .B(_09514_),
    .C(_09436_),
    .Y(_09678_));
 sky130_fd_sc_hd__o32ai_1 _18873_ (.A1(_09364_),
    .A2(_09375_),
    .A3(_09580_),
    .B1(_09559_),
    .B2(_09620_),
    .Y(_09679_));
 sky130_fd_sc_hd__nor3_1 _18874_ (.A(_09608_),
    .B(_09678_),
    .C(_09679_),
    .Y(_09680_));
 sky130_fd_sc_hd__nand2_1 _18875_ (.A(_12157_[0]),
    .B(net3917),
    .Y(_09681_));
 sky130_fd_sc_hd__o21ai_0 _18876_ (.A1(_12156_[0]),
    .A2(net3917),
    .B1(_09681_),
    .Y(_09682_));
 sky130_fd_sc_hd__a221oi_1 _18877_ (.A1(_12161_[0]),
    .A2(_09466_),
    .B1(_09682_),
    .B2(net3931),
    .C1(_09509_),
    .Y(_09683_));
 sky130_fd_sc_hd__nor3_1 _18878_ (.A(_09432_),
    .B(_09680_),
    .C(_09683_),
    .Y(_09684_));
 sky130_fd_sc_hd__a32oi_1 _18879_ (.A1(_09432_),
    .A2(_09667_),
    .A3(_09672_),
    .B1(_09677_),
    .B2(_09684_),
    .Y(_09685_));
 sky130_fd_sc_hd__o22ai_2 _18880_ (.A1(_09642_),
    .A2(_09654_),
    .B1(_09658_),
    .B2(_09685_),
    .Y(_00082_));
 sky130_fd_sc_hd__nand2_1 _18881_ (.A(_12158_[0]),
    .B(net3917),
    .Y(_09686_));
 sky130_fd_sc_hd__nand2_1 _18882_ (.A(_12157_[0]),
    .B(net3927),
    .Y(_09687_));
 sky130_fd_sc_hd__o211ai_1 _18883_ (.A1(net3936),
    .A2(net3927),
    .B1(_09687_),
    .C1(net3925),
    .Y(_09688_));
 sky130_fd_sc_hd__a21oi_1 _18884_ (.A1(_12164_[0]),
    .A2(net3925),
    .B1(net3927),
    .Y(_09689_));
 sky130_fd_sc_hd__a21oi_1 _18885_ (.A1(_09681_),
    .A2(_09689_),
    .B1(net3931),
    .Y(_09690_));
 sky130_fd_sc_hd__a311oi_1 _18886_ (.A1(net3931),
    .A2(_09686_),
    .A3(_09688_),
    .B1(_09690_),
    .C1(net3930),
    .Y(_09691_));
 sky130_fd_sc_hd__nor3b_1 _18887_ (.A(_09375_),
    .B(_09507_),
    .C_N(_09673_),
    .Y(_09692_));
 sky130_fd_sc_hd__nor3_2 _18888_ (.A(net3931),
    .B(_09566_),
    .C(_09589_),
    .Y(_09693_));
 sky130_fd_sc_hd__nand2_2 _18889_ (.A(_09370_),
    .B(net3931),
    .Y(_09694_));
 sky130_fd_sc_hd__nor2_1 _18890_ (.A(_09412_),
    .B(_09694_),
    .Y(_09695_));
 sky130_fd_sc_hd__a211o_1 _18891_ (.A1(_12166_[0]),
    .A2(_09502_),
    .B1(_09432_),
    .C1(_09695_),
    .X(_09696_));
 sky130_fd_sc_hd__o311a_4 _18892_ (.A1(net3927),
    .A2(_09692_),
    .A3(_09693_),
    .B1(_09696_),
    .C1(net3929),
    .X(_09697_));
 sky130_fd_sc_hd__o211ai_1 _18893_ (.A1(_12156_[0]),
    .A2(net3925),
    .B1(_09675_),
    .C1(net3931),
    .Y(_09698_));
 sky130_fd_sc_hd__o311ai_0 _18894_ (.A1(net3931),
    .A2(_09522_),
    .A3(_09410_),
    .B1(_09578_),
    .C1(_09698_),
    .Y(_09699_));
 sky130_fd_sc_hd__o21ai_0 _18895_ (.A1(net3612),
    .A2(_09410_),
    .B1(_09375_),
    .Y(_09700_));
 sky130_fd_sc_hd__nand2_2 _18896_ (.A(net3933),
    .B(_09643_),
    .Y(_09701_));
 sky130_fd_sc_hd__a31oi_1 _18897_ (.A1(_09630_),
    .A2(_09700_),
    .A3(_09701_),
    .B1(_09588_),
    .Y(_09702_));
 sky130_fd_sc_hd__o22ai_1 _18898_ (.A1(_09534_),
    .A2(_09438_),
    .B1(_09637_),
    .B2(_09566_),
    .Y(_09703_));
 sky130_fd_sc_hd__o21ai_0 _18899_ (.A1(_09521_),
    .A2(_09703_),
    .B1(_09452_),
    .Y(_09704_));
 sky130_fd_sc_hd__nor3b_1 _18900_ (.A(_09375_),
    .B(_09589_),
    .C_N(_09537_),
    .Y(_09705_));
 sky130_fd_sc_hd__nor3_1 _18901_ (.A(net3931),
    .B(net3612),
    .C(net3584),
    .Y(_09706_));
 sky130_fd_sc_hd__o21ai_0 _18902_ (.A1(_09705_),
    .A2(_09706_),
    .B1(_09433_),
    .Y(_09707_));
 sky130_fd_sc_hd__nand4_1 _18903_ (.A(_09699_),
    .B(_09702_),
    .C(_09704_),
    .D(_09707_),
    .Y(_09708_));
 sky130_fd_sc_hd__nand2_1 _18904_ (.A(net3933),
    .B(_09391_),
    .Y(_09709_));
 sky130_fd_sc_hd__a21oi_1 _18905_ (.A1(net3677),
    .A2(_09537_),
    .B1(_09709_),
    .Y(_09710_));
 sky130_fd_sc_hd__nor2_2 _18906_ (.A(net3936),
    .B(net3911),
    .Y(_09711_));
 sky130_fd_sc_hd__nand2_1 _18907_ (.A(_09513_),
    .B(_09711_),
    .Y(_09712_));
 sky130_fd_sc_hd__nor3_1 _18908_ (.A(_09479_),
    .B(_09710_),
    .C(_09712_),
    .Y(_09713_));
 sky130_fd_sc_hd__nand2_2 _18909_ (.A(net3921),
    .B(_09432_),
    .Y(_09714_));
 sky130_fd_sc_hd__o22ai_1 _18910_ (.A1(_09668_),
    .A2(_09432_),
    .B1(_09714_),
    .B2(net3933),
    .Y(_09715_));
 sky130_fd_sc_hd__nand3_1 _18911_ (.A(net3931),
    .B(net3930),
    .C(_09715_),
    .Y(_09716_));
 sky130_fd_sc_hd__o311ai_0 _18912_ (.A1(_12157_[0]),
    .A2(_09408_),
    .A3(_09584_),
    .B1(_09716_),
    .C1(_09525_),
    .Y(_09717_));
 sky130_fd_sc_hd__o211ai_1 _18913_ (.A1(net3678),
    .A2(net3922),
    .B1(_09537_),
    .C1(net3931),
    .Y(_09718_));
 sky130_fd_sc_hd__o31ai_1 _18914_ (.A1(net3931),
    .A2(_09589_),
    .A3(_09415_),
    .B1(_09718_),
    .Y(_09719_));
 sky130_fd_sc_hd__o22ai_1 _18915_ (.A1(net3678),
    .A2(_09585_),
    .B1(_09616_),
    .B2(net3916),
    .Y(_09720_));
 sky130_fd_sc_hd__nor3_1 _18916_ (.A(net3910),
    .B(_09646_),
    .C(_09720_),
    .Y(_09721_));
 sky130_fd_sc_hd__a211oi_1 _18917_ (.A1(net3910),
    .A2(_09719_),
    .B1(_09721_),
    .C1(net3930),
    .Y(_09722_));
 sky130_fd_sc_hd__nand2_8 _18918_ (.A(_12166_[0]),
    .B(net3916),
    .Y(_09723_));
 sky130_fd_sc_hd__and3_1 _18919_ (.A(_09375_),
    .B(_09723_),
    .C(_09675_),
    .X(_09724_));
 sky130_fd_sc_hd__o21ai_0 _18920_ (.A1(_09674_),
    .A2(_09724_),
    .B1(_09452_),
    .Y(_09725_));
 sky130_fd_sc_hd__nand4_1 _18921_ (.A(net3931),
    .B(_09391_),
    .C(_09537_),
    .D(_09723_),
    .Y(_09726_));
 sky130_fd_sc_hd__nand3_1 _18922_ (.A(net3920),
    .B(net3910),
    .C(_09620_),
    .Y(_09727_));
 sky130_fd_sc_hd__nor3_1 _18923_ (.A(net3934),
    .B(net3920),
    .C(net3910),
    .Y(_09728_));
 sky130_fd_sc_hd__o21ai_0 _18924_ (.A1(_09628_),
    .A2(_09728_),
    .B1(_09375_),
    .Y(_09729_));
 sky130_fd_sc_hd__a31o_1 _18925_ (.A1(_09726_),
    .A2(_09727_),
    .A3(_09729_),
    .B1(net3930),
    .X(_09730_));
 sky130_fd_sc_hd__or3_1 _18926_ (.A(net3913),
    .B(_09436_),
    .C(_09664_),
    .X(_09731_));
 sky130_fd_sc_hd__nand4_1 _18927_ (.A(net3930),
    .B(_09391_),
    .C(_09481_),
    .D(_09731_),
    .Y(_09732_));
 sky130_fd_sc_hd__nand4_1 _18928_ (.A(_09497_),
    .B(_09725_),
    .C(_09730_),
    .D(_09732_),
    .Y(_09733_));
 sky130_fd_sc_hd__o311ai_0 _18929_ (.A1(_09713_),
    .A2(_09717_),
    .A3(_09722_),
    .B1(_09733_),
    .C1(_09460_),
    .Y(_09734_));
 sky130_fd_sc_hd__o311a_4 _18930_ (.A1(_09612_),
    .A2(_09691_),
    .A3(_09697_),
    .B1(_09708_),
    .C1(_09734_),
    .X(_00083_));
 sky130_fd_sc_hd__nand3_1 _18931_ (.A(net3677),
    .B(_09585_),
    .C(_09537_),
    .Y(_09735_));
 sky130_fd_sc_hd__o311ai_0 _18932_ (.A1(net3677),
    .A2(_09570_),
    .A3(net3583),
    .B1(_09735_),
    .C1(net3930),
    .Y(_09736_));
 sky130_fd_sc_hd__o211ai_1 _18933_ (.A1(net3930),
    .A2(_09571_),
    .B1(_09736_),
    .C1(net3928),
    .Y(_09737_));
 sky130_fd_sc_hd__o21ai_0 _18934_ (.A1(net3931),
    .A2(_09628_),
    .B1(_09701_),
    .Y(_09738_));
 sky130_fd_sc_hd__a21oi_1 _18935_ (.A1(_09452_),
    .A2(_09738_),
    .B1(_09486_),
    .Y(_09739_));
 sky130_fd_sc_hd__a21oi_1 _18936_ (.A1(_12161_[0]),
    .A2(_09412_),
    .B1(_09558_),
    .Y(_09740_));
 sky130_fd_sc_hd__nor2_1 _18937_ (.A(net3677),
    .B(_09740_),
    .Y(_09741_));
 sky130_fd_sc_hd__o21ai_0 _18938_ (.A1(_09623_),
    .A2(_09741_),
    .B1(_09630_),
    .Y(_09742_));
 sky130_fd_sc_hd__a31oi_2 _18939_ (.A1(_09737_),
    .A2(_09739_),
    .A3(_09742_),
    .B1(_09525_),
    .Y(_09743_));
 sky130_fd_sc_hd__nand2_2 _18940_ (.A(net3911),
    .B(net3928),
    .Y(_09744_));
 sky130_fd_sc_hd__o21ai_0 _18941_ (.A1(net3916),
    .A2(_09659_),
    .B1(_09559_),
    .Y(_09745_));
 sky130_fd_sc_hd__a21boi_0 _18942_ (.A1(net3931),
    .A2(_09745_),
    .B1_N(_09467_),
    .Y(_09746_));
 sky130_fd_sc_hd__nand2_1 _18943_ (.A(_12168_[0]),
    .B(net3923),
    .Y(_09747_));
 sky130_fd_sc_hd__nand3_1 _18944_ (.A(_12157_[0]),
    .B(net3677),
    .C(_09412_),
    .Y(_09748_));
 sky130_fd_sc_hd__o21ai_0 _18945_ (.A1(_09580_),
    .A2(net3612),
    .B1(net3931),
    .Y(_09749_));
 sky130_fd_sc_hd__nand2_8 _18946_ (.A(_09431_),
    .B(_09432_),
    .Y(_09750_));
 sky130_fd_sc_hd__a31oi_1 _18947_ (.A1(_09467_),
    .A2(_09606_),
    .A3(_09749_),
    .B1(_09750_),
    .Y(_09751_));
 sky130_fd_sc_hd__a311oi_1 _18948_ (.A1(_09433_),
    .A2(_09747_),
    .A3(_09748_),
    .B1(_09751_),
    .C1(_09460_),
    .Y(_09752_));
 sky130_fd_sc_hd__nand2_2 _18949_ (.A(net3678),
    .B(_09580_),
    .Y(_09753_));
 sky130_fd_sc_hd__nand2_1 _18950_ (.A(_09446_),
    .B(_09670_),
    .Y(_09754_));
 sky130_fd_sc_hd__nand2_1 _18951_ (.A(_09568_),
    .B(_09754_),
    .Y(_09755_));
 sky130_fd_sc_hd__nand3_2 _18952_ (.A(_09753_),
    .B(_09452_),
    .C(_09755_),
    .Y(_09756_));
 sky130_fd_sc_hd__o211ai_1 _18953_ (.A1(_09744_),
    .A2(_09746_),
    .B1(_09752_),
    .C1(_09756_),
    .Y(_09757_));
 sky130_fd_sc_hd__a21oi_1 _18954_ (.A1(net3677),
    .A2(net3930),
    .B1(_09370_),
    .Y(_09758_));
 sky130_fd_sc_hd__o21ai_0 _18955_ (.A1(_09536_),
    .A2(_09758_),
    .B1(_09406_),
    .Y(_09759_));
 sky130_fd_sc_hd__nand2_1 _18956_ (.A(net3931),
    .B(_09711_),
    .Y(_09760_));
 sky130_fd_sc_hd__a31oi_1 _18957_ (.A1(_12156_[0]),
    .A2(net3677),
    .A3(net3911),
    .B1(_09406_),
    .Y(_09761_));
 sky130_fd_sc_hd__a21oi_1 _18958_ (.A1(_09760_),
    .A2(_09761_),
    .B1(net3928),
    .Y(_09762_));
 sky130_fd_sc_hd__a211oi_1 _18959_ (.A1(_09559_),
    .A2(_09670_),
    .B1(_09438_),
    .C1(_09584_),
    .Y(_09763_));
 sky130_fd_sc_hd__nand3_1 _18960_ (.A(net3934),
    .B(net3913),
    .C(_09385_),
    .Y(_09764_));
 sky130_fd_sc_hd__a21boi_0 _18961_ (.A1(net3931),
    .A2(net3911),
    .B1_N(_09764_),
    .Y(_09765_));
 sky130_fd_sc_hd__a21oi_1 _18962_ (.A1(net3677),
    .A2(_09723_),
    .B1(_09420_),
    .Y(_09766_));
 sky130_fd_sc_hd__o32ai_1 _18963_ (.A1(net3678),
    .A2(net3928),
    .A3(_09765_),
    .B1(_09766_),
    .B2(_09744_),
    .Y(_09767_));
 sky130_fd_sc_hd__a211oi_1 _18964_ (.A1(_09759_),
    .A2(_09762_),
    .B1(_09763_),
    .C1(_09767_),
    .Y(_09768_));
 sky130_fd_sc_hd__o21ai_0 _18965_ (.A1(_09486_),
    .A2(_09768_),
    .B1(_09525_),
    .Y(_09769_));
 sky130_fd_sc_hd__o21ai_0 _18966_ (.A1(_12166_[0]),
    .A2(net3677),
    .B1(_09578_),
    .Y(_09770_));
 sky130_fd_sc_hd__a21oi_1 _18967_ (.A1(net3677),
    .A2(_09579_),
    .B1(_09770_),
    .Y(_09771_));
 sky130_fd_sc_hd__nor4_1 _18968_ (.A(net3677),
    .B(net3613),
    .C(net3583),
    .D(_09750_),
    .Y(_09772_));
 sky130_fd_sc_hd__o41ai_1 _18969_ (.A1(net3931),
    .A2(_09514_),
    .A3(_09750_),
    .A4(_09628_),
    .B1(_09486_),
    .Y(_09773_));
 sky130_fd_sc_hd__nor3_1 _18970_ (.A(_09375_),
    .B(_09474_),
    .C(_09567_),
    .Y(_09774_));
 sky130_fd_sc_hd__nor3_1 _18971_ (.A(net3931),
    .B(_09514_),
    .C(net3583),
    .Y(_09775_));
 sky130_fd_sc_hd__o21ai_0 _18972_ (.A1(_09774_),
    .A2(_09775_),
    .B1(_09452_),
    .Y(_09776_));
 sky130_fd_sc_hd__a21oi_1 _18973_ (.A1(_09537_),
    .A2(_09723_),
    .B1(net3931),
    .Y(_09777_));
 sky130_fd_sc_hd__nor3_1 _18974_ (.A(net3677),
    .B(net3613),
    .C(_09628_),
    .Y(_09778_));
 sky130_fd_sc_hd__o21ai_0 _18975_ (.A1(_09777_),
    .A2(_09778_),
    .B1(_09433_),
    .Y(_09779_));
 sky130_fd_sc_hd__nand2_1 _18976_ (.A(_09776_),
    .B(_09779_),
    .Y(_09780_));
 sky130_fd_sc_hd__nor4_2 _18977_ (.A(_09771_),
    .B(_09772_),
    .C(_09773_),
    .D(_09780_),
    .Y(_09781_));
 sky130_fd_sc_hd__o2bb2ai_2 _18978_ (.A1_N(_09743_),
    .A2_N(_09757_),
    .B1(_09769_),
    .B2(_09781_),
    .Y(_00084_));
 sky130_fd_sc_hd__nor3_1 _18979_ (.A(net3931),
    .B(net3913),
    .C(net3911),
    .Y(_09782_));
 sky130_fd_sc_hd__a31oi_1 _18980_ (.A1(net3913),
    .A2(net3911),
    .A3(_09616_),
    .B1(_09782_),
    .Y(_09783_));
 sky130_fd_sc_hd__nand2_1 _18981_ (.A(_12164_[0]),
    .B(_09466_),
    .Y(_09784_));
 sky130_fd_sc_hd__a31oi_1 _18982_ (.A1(net3911),
    .A2(_09546_),
    .A3(_09784_),
    .B1(_09711_),
    .Y(_09785_));
 sky130_fd_sc_hd__o21ai_0 _18983_ (.A1(net3929),
    .A2(_09620_),
    .B1(net3919),
    .Y(_09786_));
 sky130_fd_sc_hd__o311ai_0 _18984_ (.A1(net3919),
    .A2(net3929),
    .A3(_09440_),
    .B1(_09786_),
    .C1(_09364_),
    .Y(_09787_));
 sky130_fd_sc_hd__o221ai_1 _18985_ (.A1(_09364_),
    .A2(_09783_),
    .B1(_09785_),
    .B2(_09370_),
    .C1(_09787_),
    .Y(_09788_));
 sky130_fd_sc_hd__nand2_1 _18986_ (.A(_12158_[0]),
    .B(net3926),
    .Y(_09789_));
 sky130_fd_sc_hd__a21oi_1 _18987_ (.A1(_09789_),
    .A2(_09681_),
    .B1(net3931),
    .Y(_09790_));
 sky130_fd_sc_hd__a211oi_1 _18988_ (.A1(net3936),
    .A2(_09643_),
    .B1(_09790_),
    .C1(net3930),
    .Y(_09791_));
 sky130_fd_sc_hd__o21ai_0 _18989_ (.A1(_12156_[0]),
    .A2(net3925),
    .B1(_09573_),
    .Y(_09792_));
 sky130_fd_sc_hd__nor2_1 _18990_ (.A(_12157_[0]),
    .B(_09513_),
    .Y(_09793_));
 sky130_fd_sc_hd__a211oi_1 _18991_ (.A1(_09375_),
    .A2(_09792_),
    .B1(_09793_),
    .C1(net3912),
    .Y(_09794_));
 sky130_fd_sc_hd__nor3_1 _18992_ (.A(net3927),
    .B(_09791_),
    .C(_09794_),
    .Y(_09795_));
 sky130_fd_sc_hd__a211oi_1 _18993_ (.A1(net3927),
    .A2(_09788_),
    .B1(_09795_),
    .C1(_09497_),
    .Y(_09796_));
 sky130_fd_sc_hd__nor4_1 _18994_ (.A(net3935),
    .B(net3913),
    .C(_09479_),
    .D(_09620_),
    .Y(_09797_));
 sky130_fd_sc_hd__o21ai_0 _18995_ (.A1(net3677),
    .A2(_09673_),
    .B1(_09433_),
    .Y(_09798_));
 sky130_fd_sc_hd__o211ai_1 _18996_ (.A1(net3913),
    .A2(_09615_),
    .B1(_09452_),
    .C1(_09668_),
    .Y(_09799_));
 sky130_fd_sc_hd__o21ai_0 _18997_ (.A1(_09797_),
    .A2(_09798_),
    .B1(_09799_),
    .Y(_09800_));
 sky130_fd_sc_hd__nand2_2 _18998_ (.A(_12161_[0]),
    .B(_09427_),
    .Y(_09801_));
 sky130_fd_sc_hd__o21ai_0 _18999_ (.A1(_12170_[0]),
    .A2(net3931),
    .B1(net3913),
    .Y(_09802_));
 sky130_fd_sc_hd__nor3b_1 _19000_ (.A(_09628_),
    .B(net3931),
    .C_N(_09668_),
    .Y(_09803_));
 sky130_fd_sc_hd__a311oi_1 _19001_ (.A1(net3931),
    .A2(_09537_),
    .A3(_09572_),
    .B1(_09803_),
    .C1(_09391_),
    .Y(_09804_));
 sky130_fd_sc_hd__a311oi_1 _19002_ (.A1(_09391_),
    .A2(_09801_),
    .A3(_09802_),
    .B1(_09804_),
    .C1(net3930),
    .Y(_09805_));
 sky130_fd_sc_hd__nor3_2 _19003_ (.A(_09525_),
    .B(_09800_),
    .C(_09805_),
    .Y(_09806_));
 sky130_fd_sc_hd__nand2_1 _19004_ (.A(net3923),
    .B(_09391_),
    .Y(_09807_));
 sky130_fd_sc_hd__o21ai_0 _19005_ (.A1(_09391_),
    .A2(_09559_),
    .B1(_09807_),
    .Y(_09808_));
 sky130_fd_sc_hd__o32ai_1 _19006_ (.A1(_12161_[0]),
    .A2(net3931),
    .A3(_09714_),
    .B1(_09709_),
    .B2(_09531_),
    .Y(_09809_));
 sky130_fd_sc_hd__a211oi_1 _19007_ (.A1(_09438_),
    .A2(_09808_),
    .B1(_09809_),
    .C1(net3911),
    .Y(_09810_));
 sky130_fd_sc_hd__nor2_1 _19008_ (.A(net3677),
    .B(_09714_),
    .Y(_09811_));
 sky130_fd_sc_hd__o21ai_0 _19009_ (.A1(_09466_),
    .A2(_09811_),
    .B1(net3933),
    .Y(_09812_));
 sky130_fd_sc_hd__nor2_1 _19010_ (.A(net3913),
    .B(_09614_),
    .Y(_09813_));
 sky130_fd_sc_hd__a21oi_1 _19011_ (.A1(net3931),
    .A2(_09813_),
    .B1(_09803_),
    .Y(_09814_));
 sky130_fd_sc_hd__nor3_1 _19012_ (.A(net3931),
    .B(_09465_),
    .C(_09415_),
    .Y(_09815_));
 sky130_fd_sc_hd__a311oi_1 _19013_ (.A1(net3931),
    .A2(_09534_),
    .A3(_09572_),
    .B1(_09815_),
    .C1(_09432_),
    .Y(_09816_));
 sky130_fd_sc_hd__a21oi_1 _19014_ (.A1(_09432_),
    .A2(_09814_),
    .B1(_09816_),
    .Y(_09817_));
 sky130_fd_sc_hd__a221oi_2 _19015_ (.A1(_09810_),
    .A2(_09812_),
    .B1(_09817_),
    .B2(net3911),
    .C1(_09525_),
    .Y(_09818_));
 sky130_fd_sc_hd__nand2_1 _19016_ (.A(net3931),
    .B(_09448_),
    .Y(_09819_));
 sky130_fd_sc_hd__a21oi_1 _19017_ (.A1(_09753_),
    .A2(_09819_),
    .B1(net3927),
    .Y(_09820_));
 sky130_fd_sc_hd__a221oi_1 _19018_ (.A1(_12161_[0]),
    .A2(_09412_),
    .B1(_09427_),
    .B2(_12166_[0]),
    .C1(net3910),
    .Y(_09821_));
 sky130_fd_sc_hd__o31a_1 _19019_ (.A1(_09375_),
    .A2(_09474_),
    .A3(_09475_),
    .B1(_09821_),
    .X(_09822_));
 sky130_fd_sc_hd__nand3_1 _19020_ (.A(net3931),
    .B(_09537_),
    .C(_09723_),
    .Y(_09823_));
 sky130_fd_sc_hd__nand3_1 _19021_ (.A(_09370_),
    .B(_09375_),
    .C(_09412_),
    .Y(_09824_));
 sky130_fd_sc_hd__a31oi_1 _19022_ (.A1(_09452_),
    .A2(_09823_),
    .A3(_09824_),
    .B1(_09497_),
    .Y(_09825_));
 sky130_fd_sc_hd__o311ai_0 _19023_ (.A1(net3931),
    .A2(net3612),
    .A3(_09519_),
    .B1(_09424_),
    .C1(_09433_),
    .Y(_09826_));
 sky130_fd_sc_hd__o311ai_1 _19024_ (.A1(net3929),
    .A2(_09820_),
    .A3(_09822_),
    .B1(_09825_),
    .C1(_09826_),
    .Y(_09827_));
 sky130_fd_sc_hd__nand2_1 _19025_ (.A(_09460_),
    .B(_09827_),
    .Y(_09828_));
 sky130_fd_sc_hd__o32ai_1 _19026_ (.A1(_09460_),
    .A2(_09796_),
    .A3(_09806_),
    .B1(_09818_),
    .B2(_09828_),
    .Y(_00085_));
 sky130_fd_sc_hd__o21ai_0 _19027_ (.A1(_12156_[0]),
    .A2(net3917),
    .B1(_09723_),
    .Y(_09829_));
 sky130_fd_sc_hd__a22oi_1 _19028_ (.A1(_12158_[0]),
    .A2(_09466_),
    .B1(_09829_),
    .B2(net3931),
    .Y(_09830_));
 sky130_fd_sc_hd__nor2_1 _19029_ (.A(net3925),
    .B(_09482_),
    .Y(_09831_));
 sky130_fd_sc_hd__nand3_1 _19030_ (.A(net3931),
    .B(_09504_),
    .C(_09723_),
    .Y(_09832_));
 sky130_fd_sc_hd__o311ai_0 _19031_ (.A1(net3931),
    .A2(_09507_),
    .A3(_09831_),
    .B1(_09832_),
    .C1(_09432_),
    .Y(_09833_));
 sky130_fd_sc_hd__o21ai_0 _19032_ (.A1(_09432_),
    .A2(_09830_),
    .B1(_09833_),
    .Y(_09834_));
 sky130_fd_sc_hd__a21o_1 _19033_ (.A1(net3936),
    .A2(net3931),
    .B1(_09445_),
    .X(_09835_));
 sky130_fd_sc_hd__o311ai_0 _19034_ (.A1(_12173_[0]),
    .A2(_12182_[0]),
    .A3(net3917),
    .B1(_09433_),
    .C1(_09835_),
    .Y(_09836_));
 sky130_fd_sc_hd__a21oi_1 _19035_ (.A1(_09686_),
    .A2(_09573_),
    .B1(_09375_),
    .Y(_09837_));
 sky130_fd_sc_hd__nor3_2 _19036_ (.A(net3931),
    .B(_09415_),
    .C(_09570_),
    .Y(_09838_));
 sky130_fd_sc_hd__o21ai_0 _19037_ (.A1(_09837_),
    .A2(_09838_),
    .B1(_09452_),
    .Y(_09839_));
 sky130_fd_sc_hd__nand2_1 _19038_ (.A(_09836_),
    .B(_09839_),
    .Y(_09840_));
 sky130_fd_sc_hd__a21oi_1 _19039_ (.A1(net3912),
    .A2(_09834_),
    .B1(_09840_),
    .Y(_09841_));
 sky130_fd_sc_hd__nor2_2 _19040_ (.A(_12175_[0]),
    .B(net3919),
    .Y(_09842_));
 sky130_fd_sc_hd__nor2_1 _19041_ (.A(_12157_[0]),
    .B(net3677),
    .Y(_09843_));
 sky130_fd_sc_hd__a211oi_1 _19042_ (.A1(net3677),
    .A2(_09659_),
    .B1(_09843_),
    .C1(net3916),
    .Y(_09844_));
 sky130_fd_sc_hd__o311ai_0 _19043_ (.A1(net3931),
    .A2(net3613),
    .A3(_09420_),
    .B1(_09433_),
    .C1(_09718_),
    .Y(_09845_));
 sky130_fd_sc_hd__a21oi_1 _19044_ (.A1(net3926),
    .A2(_09482_),
    .B1(_09375_),
    .Y(_09846_));
 sky130_fd_sc_hd__a32oi_1 _19045_ (.A1(_09375_),
    .A2(_09537_),
    .A3(_09446_),
    .B1(_09846_),
    .B2(_09753_),
    .Y(_09847_));
 sky130_fd_sc_hd__a21oi_1 _19046_ (.A1(net3678),
    .A2(_09694_),
    .B1(net3926),
    .Y(_09848_));
 sky130_fd_sc_hd__nor3_2 _19047_ (.A(_09473_),
    .B(_09750_),
    .C(_09848_),
    .Y(_09849_));
 sky130_fd_sc_hd__a211oi_2 _19048_ (.A1(_09452_),
    .A2(_09847_),
    .B1(_09849_),
    .C1(_09588_),
    .Y(_09850_));
 sky130_fd_sc_hd__o311ai_2 _19049_ (.A1(_09744_),
    .A2(_09842_),
    .A3(_09844_),
    .B1(_09845_),
    .C1(_09850_),
    .Y(_09851_));
 sky130_fd_sc_hd__nor2_1 _19050_ (.A(_09693_),
    .B(_09793_),
    .Y(_09852_));
 sky130_fd_sc_hd__a211o_1 _19051_ (.A1(_12166_[0]),
    .A2(_09375_),
    .B1(_09412_),
    .C1(_09436_),
    .X(_09853_));
 sky130_fd_sc_hd__a21oi_1 _19052_ (.A1(_12174_[0]),
    .A2(_09412_),
    .B1(_09509_),
    .Y(_09854_));
 sky130_fd_sc_hd__a21oi_1 _19053_ (.A1(_09853_),
    .A2(_09854_),
    .B1(_09432_),
    .Y(_09855_));
 sky130_fd_sc_hd__o21ai_0 _19054_ (.A1(_09499_),
    .A2(_09852_),
    .B1(_09855_),
    .Y(_09856_));
 sky130_fd_sc_hd__a21oi_1 _19055_ (.A1(net3936),
    .A2(_09620_),
    .B1(_09522_),
    .Y(_09857_));
 sky130_fd_sc_hd__a21oi_1 _19056_ (.A1(net3936),
    .A2(_09580_),
    .B1(_09479_),
    .Y(_09858_));
 sky130_fd_sc_hd__o21ai_0 _19057_ (.A1(_12170_[0]),
    .A2(_09857_),
    .B1(_09858_),
    .Y(_09859_));
 sky130_fd_sc_hd__a21oi_1 _19058_ (.A1(net3913),
    .A2(_09438_),
    .B1(_09659_),
    .Y(_09860_));
 sky130_fd_sc_hd__o21ai_0 _19059_ (.A1(_09385_),
    .A2(_09628_),
    .B1(_09436_),
    .Y(_09861_));
 sky130_fd_sc_hd__o211ai_1 _19060_ (.A1(net3911),
    .A2(_09860_),
    .B1(_09861_),
    .C1(_09460_),
    .Y(_09862_));
 sky130_fd_sc_hd__a21oi_2 _19061_ (.A1(net3911),
    .A2(_09859_),
    .B1(_09862_),
    .Y(_09863_));
 sky130_fd_sc_hd__a211oi_1 _19062_ (.A1(net3936),
    .A2(_09583_),
    .B1(_09724_),
    .C1(net3929),
    .Y(_09864_));
 sky130_fd_sc_hd__o211ai_1 _19063_ (.A1(_09364_),
    .A2(net3929),
    .B1(_09764_),
    .C1(_09375_),
    .Y(_09865_));
 sky130_fd_sc_hd__o21ai_0 _19064_ (.A1(_12166_[0]),
    .A2(net3912),
    .B1(net3917),
    .Y(_09866_));
 sky130_fd_sc_hd__o211ai_1 _19065_ (.A1(net3912),
    .A2(_09537_),
    .B1(_09866_),
    .C1(net3931),
    .Y(_09867_));
 sky130_fd_sc_hd__nand2_1 _19066_ (.A(_09460_),
    .B(_09432_),
    .Y(_09868_));
 sky130_fd_sc_hd__a221o_1 _19067_ (.A1(net3912),
    .A2(_09522_),
    .B1(_09865_),
    .B2(_09867_),
    .C1(_09868_),
    .X(_09869_));
 sky130_fd_sc_hd__o311a_1 _19068_ (.A1(_09487_),
    .A2(_09651_),
    .A3(_09864_),
    .B1(_09869_),
    .C1(_09497_),
    .X(_09870_));
 sky130_fd_sc_hd__o21ai_0 _19069_ (.A1(_09856_),
    .A2(_09863_),
    .B1(_09870_),
    .Y(_09871_));
 sky130_fd_sc_hd__o311ai_0 _19070_ (.A1(_09486_),
    .A2(_09497_),
    .A3(_09841_),
    .B1(_09851_),
    .C1(_09871_),
    .Y(_00086_));
 sky130_fd_sc_hd__nor2_1 _19071_ (.A(_12182_[0]),
    .B(net3925),
    .Y(_09872_));
 sky130_fd_sc_hd__a211oi_1 _19072_ (.A1(_12166_[0]),
    .A2(net3931),
    .B1(net3917),
    .C1(_09535_),
    .Y(_09873_));
 sky130_fd_sc_hd__nor3_1 _19073_ (.A(net3927),
    .B(_09872_),
    .C(_09873_),
    .Y(_09874_));
 sky130_fd_sc_hd__a21oi_1 _19074_ (.A1(_12158_[0]),
    .A2(_09375_),
    .B1(_09412_),
    .Y(_09875_));
 sky130_fd_sc_hd__a211oi_1 _19075_ (.A1(_12168_[0]),
    .A2(_09412_),
    .B1(net3910),
    .C1(_09875_),
    .Y(_09876_));
 sky130_fd_sc_hd__o21ai_0 _19076_ (.A1(_09566_),
    .A2(_09410_),
    .B1(_09375_),
    .Y(_09877_));
 sky130_fd_sc_hd__o311ai_0 _19077_ (.A1(_09375_),
    .A2(_09531_),
    .A3(_09410_),
    .B1(_09877_),
    .C1(net3910),
    .Y(_09878_));
 sky130_fd_sc_hd__nor2_1 _19078_ (.A(_12161_[0]),
    .B(_09375_),
    .Y(_09879_));
 sky130_fd_sc_hd__o21ai_0 _19079_ (.A1(_09536_),
    .A2(_09879_),
    .B1(net3917),
    .Y(_09880_));
 sky130_fd_sc_hd__a21oi_1 _19080_ (.A1(_09531_),
    .A2(_09694_),
    .B1(_09432_),
    .Y(_09881_));
 sky130_fd_sc_hd__nand2_1 _19081_ (.A(_09880_),
    .B(_09881_),
    .Y(_09882_));
 sky130_fd_sc_hd__nand3_1 _19082_ (.A(net3912),
    .B(_09878_),
    .C(_09882_),
    .Y(_09883_));
 sky130_fd_sc_hd__nor3b_1 _19083_ (.A(net3931),
    .B(_09420_),
    .C_N(_09559_),
    .Y(_09884_));
 sky130_fd_sc_hd__o21ai_0 _19084_ (.A1(_09480_),
    .A2(_09884_),
    .B1(_09452_),
    .Y(_09885_));
 sky130_fd_sc_hd__a21o_1 _19085_ (.A1(_09668_),
    .A2(_09606_),
    .B1(net3931),
    .X(_09886_));
 sky130_fd_sc_hd__nand3_1 _19086_ (.A(_09433_),
    .B(_09604_),
    .C(_09886_),
    .Y(_09887_));
 sky130_fd_sc_hd__nor2_2 _19087_ (.A(_09591_),
    .B(_09750_),
    .Y(_09888_));
 sky130_fd_sc_hd__a21oi_1 _19088_ (.A1(_09888_),
    .A2(_09835_),
    .B1(_09486_),
    .Y(_09889_));
 sky130_fd_sc_hd__a21oi_1 _19089_ (.A1(_09504_),
    .A2(_09723_),
    .B1(net3931),
    .Y(_09890_));
 sky130_fd_sc_hd__o21ai_0 _19090_ (.A1(_09513_),
    .A2(_09482_),
    .B1(_09534_),
    .Y(_09891_));
 sky130_fd_sc_hd__o21ai_0 _19091_ (.A1(_09890_),
    .A2(_09891_),
    .B1(_09578_),
    .Y(_09892_));
 sky130_fd_sc_hd__a41oi_1 _19092_ (.A1(_09885_),
    .A2(_09887_),
    .A3(_09889_),
    .A4(_09892_),
    .B1(_09497_),
    .Y(_09893_));
 sky130_fd_sc_hd__o311ai_0 _19093_ (.A1(net3912),
    .A2(_09874_),
    .A3(_09876_),
    .B1(_09883_),
    .C1(_09893_),
    .Y(_09894_));
 sky130_fd_sc_hd__o21ai_0 _19094_ (.A1(_09375_),
    .A2(net3930),
    .B1(net3934),
    .Y(_09895_));
 sky130_fd_sc_hd__o21ai_0 _19095_ (.A1(net3934),
    .A2(net3930),
    .B1(_09895_),
    .Y(_09896_));
 sky130_fd_sc_hd__o21ai_0 _19096_ (.A1(net3914),
    .A2(_09479_),
    .B1(net3678),
    .Y(_09897_));
 sky130_fd_sc_hd__a21oi_1 _19097_ (.A1(net3914),
    .A2(_09896_),
    .B1(_09897_),
    .Y(_09898_));
 sky130_fd_sc_hd__a221oi_1 _19098_ (.A1(_09375_),
    .A2(net3930),
    .B1(_09643_),
    .B2(_12157_[0]),
    .C1(_09898_),
    .Y(_09899_));
 sky130_fd_sc_hd__a21oi_1 _19099_ (.A1(net3934),
    .A2(_09583_),
    .B1(_09522_),
    .Y(_09900_));
 sky130_fd_sc_hd__o21ai_0 _19100_ (.A1(_09466_),
    .A2(_09695_),
    .B1(_09364_),
    .Y(_09901_));
 sky130_fd_sc_hd__a21oi_1 _19101_ (.A1(_09408_),
    .A2(_09446_),
    .B1(_09364_),
    .Y(_09902_));
 sky130_fd_sc_hd__o21ai_0 _19102_ (.A1(_09474_),
    .A2(_09902_),
    .B1(net3929),
    .Y(_09903_));
 sky130_fd_sc_hd__o2111ai_1 _19103_ (.A1(net3929),
    .A2(_09900_),
    .B1(_09901_),
    .C1(net3927),
    .D1(_09903_),
    .Y(_09904_));
 sky130_fd_sc_hd__xnor2_1 _19104_ (.A(net3931),
    .B(net3925),
    .Y(_09905_));
 sky130_fd_sc_hd__a221oi_1 _19105_ (.A1(_12157_[0]),
    .A2(_09905_),
    .B1(_09583_),
    .B2(_12170_[0]),
    .C1(_09500_),
    .Y(_09906_));
 sky130_fd_sc_hd__nand3_1 _19106_ (.A(_12156_[0]),
    .B(net3931),
    .C(_09412_),
    .Y(_09907_));
 sky130_fd_sc_hd__nand3_1 _19107_ (.A(_09564_),
    .B(_09578_),
    .C(_09907_),
    .Y(_09908_));
 sky130_fd_sc_hd__a21oi_1 _19108_ (.A1(_09504_),
    .A2(_09824_),
    .B1(net3936),
    .Y(_09909_));
 sky130_fd_sc_hd__o22a_1 _19109_ (.A1(_09750_),
    .A2(_09906_),
    .B1(_09908_),
    .B2(_09909_),
    .X(_09910_));
 sky130_fd_sc_hd__nand3_1 _19110_ (.A(_09375_),
    .B(_09559_),
    .C(_09632_),
    .Y(_09911_));
 sky130_fd_sc_hd__o211ai_1 _19111_ (.A1(_09375_),
    .A2(_09644_),
    .B1(_09911_),
    .C1(_09452_),
    .Y(_09912_));
 sky130_fd_sc_hd__nor3_1 _19112_ (.A(_12166_[0]),
    .B(net3931),
    .C(net3924),
    .Y(_09913_));
 sky130_fd_sc_hd__a31oi_1 _19113_ (.A1(net3931),
    .A2(_09573_),
    .A3(_09559_),
    .B1(_09913_),
    .Y(_09914_));
 sky130_fd_sc_hd__a21oi_1 _19114_ (.A1(_09433_),
    .A2(_09914_),
    .B1(_09486_),
    .Y(_09915_));
 sky130_fd_sc_hd__a31oi_2 _19115_ (.A1(_09910_),
    .A2(_09912_),
    .A3(_09915_),
    .B1(_09525_),
    .Y(_09916_));
 sky130_fd_sc_hd__o211ai_1 _19116_ (.A1(net3927),
    .A2(_09899_),
    .B1(_09904_),
    .C1(_09916_),
    .Y(_09917_));
 sky130_fd_sc_hd__o21ai_0 _19117_ (.A1(_09893_),
    .A2(_09916_),
    .B1(_09460_),
    .Y(_09918_));
 sky130_fd_sc_hd__nand3_1 _19118_ (.A(_09894_),
    .B(_09917_),
    .C(_09918_),
    .Y(_00087_));
 sky130_fd_sc_hd__xnor3_1 _19119_ (.A(net4211),
    .B(net4195),
    .C(\sa03_sr[1] ),
    .X(_09919_));
 sky130_fd_sc_hd__xnor3_1 _19120_ (.A(_07660_),
    .B(_07692_),
    .C(_09919_),
    .X(_09920_));
 sky130_fd_sc_hd__mux2i_2 _19121_ (.A0(\text_in_r[17] ),
    .A1(_09920_),
    .S(_05879_),
    .Y(_09921_));
 sky130_fd_sc_hd__xor2_4 _19122_ (.A(\u0.tmp_w[17] ),
    .B(_09921_),
    .X(_09922_));
 sky130_fd_sc_hd__clkinv_16 _19123_ (.A(net3907),
    .Y(_09923_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_560 ();
 sky130_fd_sc_hd__xor2_1 _19126_ (.A(\sa03_sr[0] ),
    .B(\sa32_sub[0] ),
    .X(_09925_));
 sky130_fd_sc_hd__xnor3_1 _19127_ (.A(net4195),
    .B(_07692_),
    .C(_09925_),
    .X(_09926_));
 sky130_fd_sc_hd__mux2i_2 _19128_ (.A0(\text_in_r[16] ),
    .A1(_09926_),
    .S(_05879_),
    .Y(_09927_));
 sky130_fd_sc_hd__xor2_4 _19129_ (.A(\u0.tmp_w[16] ),
    .B(_09927_),
    .X(_09928_));
 sky130_fd_sc_hd__clkinv_16 _19130_ (.A(net408),
    .Y(_09929_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_558 ();
 sky130_fd_sc_hd__xor2_1 _19133_ (.A(\sa32_sub[2] ),
    .B(net4222),
    .X(_09931_));
 sky130_fd_sc_hd__xnor3_1 _19134_ (.A(net4210),
    .B(\sa21_sub[1] ),
    .C(net4193),
    .X(_09932_));
 sky130_fd_sc_hd__xnor2_1 _19135_ (.A(_09931_),
    .B(_09932_),
    .Y(_09933_));
 sky130_fd_sc_hd__mux2i_2 _19136_ (.A0(\text_in_r[18] ),
    .A1(_09933_),
    .S(_05879_),
    .Y(_09934_));
 sky130_fd_sc_hd__xnor2_4 _19137_ (.A(\u0.tmp_w[18] ),
    .B(_09934_),
    .Y(_09935_));
 sky130_fd_sc_hd__clkinv_16 _19138_ (.A(_09935_),
    .Y(_09936_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_551 ();
 sky130_fd_sc_hd__xnor2_1 _19146_ (.A(\sa32_sub[6] ),
    .B(\sa03_sr[6] ),
    .Y(_09941_));
 sky130_fd_sc_hd__xor3_1 _19147_ (.A(\sa21_sub[6] ),
    .B(_07700_),
    .C(_09941_),
    .X(_09942_));
 sky130_fd_sc_hd__mux2i_4 _19148_ (.A0(\text_in_r[22] ),
    .A1(_09942_),
    .S(_05879_),
    .Y(_09943_));
 sky130_fd_sc_hd__xor2_4 _19149_ (.A(\u0.tmp_w[22] ),
    .B(_09943_),
    .X(_09944_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_550 ();
 sky130_fd_sc_hd__xnor2_1 _19151_ (.A(\sa21_sub[6] ),
    .B(net4179),
    .Y(_09946_));
 sky130_fd_sc_hd__xnor3_1 _19152_ (.A(\sa03_sr[7] ),
    .B(\sa10_sub[6] ),
    .C(\sa21_sub[7] ),
    .X(_09947_));
 sky130_fd_sc_hd__xor2_2 _19153_ (.A(_09946_),
    .B(_09947_),
    .X(_09948_));
 sky130_fd_sc_hd__mux2i_4 _19154_ (.A0(\text_in_r[23] ),
    .A1(_09948_),
    .S(_05879_),
    .Y(_09949_));
 sky130_fd_sc_hd__xnor2_4 _19155_ (.A(\u0.tmp_w[23] ),
    .B(_09949_),
    .Y(_09950_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_549 ();
 sky130_fd_sc_hd__nor2_1 _19157_ (.A(net3903),
    .B(_09950_),
    .Y(_09952_));
 sky130_fd_sc_hd__xnor3_1 _19158_ (.A(\sa21_sub[4] ),
    .B(\sa32_sub[5] ),
    .C(\sa03_sr[5] ),
    .X(_09953_));
 sky130_fd_sc_hd__xor2_1 _19159_ (.A(\sa10_sub[4] ),
    .B(\sa21_sub[5] ),
    .X(_09954_));
 sky130_fd_sc_hd__xnor2_2 _19160_ (.A(_09953_),
    .B(_09954_),
    .Y(_09955_));
 sky130_fd_sc_hd__mux2i_4 _19161_ (.A0(\text_in_r[21] ),
    .A1(_09955_),
    .S(net4115),
    .Y(_09956_));
 sky130_fd_sc_hd__xnor2_4 _19162_ (.A(net4133),
    .B(_09956_),
    .Y(_09957_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_546 ();
 sky130_fd_sc_hd__nor2b_2 _19166_ (.A(net4230),
    .B_N(\u0.tmp_w[19] ),
    .Y(_09961_));
 sky130_fd_sc_hd__nor2_1 _19167_ (.A(\u0.tmp_w[19] ),
    .B(net4230),
    .Y(_09962_));
 sky130_fd_sc_hd__xnor2_1 _19168_ (.A(\sa10_sub[7] ),
    .B(\sa10_sub[2] ),
    .Y(_09963_));
 sky130_fd_sc_hd__xnor3_1 _19169_ (.A(\sa21_sub[2] ),
    .B(\sa32_sub[3] ),
    .C(\sa21_sub[7] ),
    .X(_09964_));
 sky130_fd_sc_hd__xnor2_1 _19170_ (.A(net4192),
    .B(\sa03_sr[3] ),
    .Y(_09965_));
 sky130_fd_sc_hd__xnor3_1 _19171_ (.A(_09963_),
    .B(_09964_),
    .C(_09965_),
    .X(_09966_));
 sky130_fd_sc_hd__mux2i_4 _19172_ (.A0(_09961_),
    .A1(_09962_),
    .S(_09966_),
    .Y(_09967_));
 sky130_fd_sc_hd__nor2_2 _19173_ (.A(\u0.tmp_w[19] ),
    .B(net4115),
    .Y(_09968_));
 sky130_fd_sc_hd__nand2_1 _19174_ (.A(\u0.tmp_w[19] ),
    .B(net398),
    .Y(_09969_));
 sky130_fd_sc_hd__nor2_2 _19175_ (.A(\text_in_r[19] ),
    .B(_09969_),
    .Y(_09970_));
 sky130_fd_sc_hd__a21oi_4 _19176_ (.A1(\text_in_r[19] ),
    .A2(_09968_),
    .B1(_09970_),
    .Y(_09971_));
 sky130_fd_sc_hd__and2_4 _19177_ (.A(_09967_),
    .B(_09971_),
    .X(_09972_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_544 ();
 sky130_fd_sc_hd__nand2_8 _19180_ (.A(net3908),
    .B(net3900),
    .Y(_09975_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_543 ();
 sky130_fd_sc_hd__nand2_8 _19182_ (.A(_09967_),
    .B(_09971_),
    .Y(_09977_));
 sky130_fd_sc_hd__nand2_4 _19183_ (.A(_12202_[0]),
    .B(_09977_),
    .Y(_09978_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_541 ();
 sky130_fd_sc_hd__a21oi_1 _19186_ (.A1(_09975_),
    .A2(_09978_),
    .B1(net3904),
    .Y(_09981_));
 sky130_fd_sc_hd__inv_6 _19187_ (.A(_12189_[0]),
    .Y(_09982_));
 sky130_fd_sc_hd__nand2_8 _19188_ (.A(net3904),
    .B(_09977_),
    .Y(_09983_));
 sky130_fd_sc_hd__nand2_8 _19189_ (.A(_09929_),
    .B(net3899),
    .Y(_09984_));
 sky130_fd_sc_hd__o21ai_0 _19190_ (.A1(_09982_),
    .A2(_09983_),
    .B1(_09984_),
    .Y(_09985_));
 sky130_fd_sc_hd__xnor2_1 _19191_ (.A(net4192),
    .B(\sa32_sub[4] ),
    .Y(_09986_));
 sky130_fd_sc_hd__xnor3_1 _19192_ (.A(\sa10_sub[3] ),
    .B(\sa21_sub[4] ),
    .C(\sa03_sr[4] ),
    .X(_09987_));
 sky130_fd_sc_hd__xnor3_1 _19193_ (.A(_07692_),
    .B(_09986_),
    .C(_09987_),
    .X(_09988_));
 sky130_fd_sc_hd__mux2i_4 _19194_ (.A0(\text_in_r[20] ),
    .A1(_09988_),
    .S(net4115),
    .Y(_09989_));
 sky130_fd_sc_hd__xnor2_4 _19195_ (.A(\u0.tmp_w[20] ),
    .B(_09989_),
    .Y(_09990_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_540 ();
 sky130_fd_sc_hd__o21ai_0 _19197_ (.A1(_09981_),
    .A2(_09985_),
    .B1(net3895),
    .Y(_09992_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_539 ();
 sky130_fd_sc_hd__nor2_2 _19199_ (.A(_09923_),
    .B(_09972_),
    .Y(_09994_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_537 ();
 sky130_fd_sc_hd__nand2_2 _19202_ (.A(net3906),
    .B(_09936_),
    .Y(_09997_));
 sky130_fd_sc_hd__xor2_4 _19203_ (.A(\u0.tmp_w[20] ),
    .B(_09989_),
    .X(_09998_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_534 ();
 sky130_fd_sc_hd__o221ai_1 _19207_ (.A1(_12193_[0]),
    .A2(_09983_),
    .B1(_09994_),
    .B2(_09997_),
    .C1(net3893),
    .Y(_10002_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_533 ();
 sky130_fd_sc_hd__nand2_4 _19209_ (.A(_09936_),
    .B(net3900),
    .Y(_10004_));
 sky130_fd_sc_hd__o21ai_0 _19210_ (.A1(net3906),
    .A2(_09983_),
    .B1(_10004_),
    .Y(_10005_));
 sky130_fd_sc_hd__nor2_4 _19211_ (.A(net3904),
    .B(_09972_),
    .Y(_10006_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_532 ();
 sky130_fd_sc_hd__nand2_1 _19213_ (.A(net3904),
    .B(net3899),
    .Y(_10008_));
 sky130_fd_sc_hd__nor2_1 _19214_ (.A(_12190_[0]),
    .B(_10008_),
    .Y(_10009_));
 sky130_fd_sc_hd__a221oi_1 _19215_ (.A1(_09923_),
    .A2(_10005_),
    .B1(_10006_),
    .B2(net3906),
    .C1(_10009_),
    .Y(_10010_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_531 ();
 sky130_fd_sc_hd__nand2_2 _19217_ (.A(_09923_),
    .B(_09972_),
    .Y(_10012_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_530 ();
 sky130_fd_sc_hd__nor2_2 _19219_ (.A(_09923_),
    .B(_09977_),
    .Y(_10014_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_529 ();
 sky130_fd_sc_hd__o21ai_0 _19221_ (.A1(_10014_),
    .A2(_09997_),
    .B1(net3895),
    .Y(_10016_));
 sky130_fd_sc_hd__a31oi_1 _19222_ (.A1(net3904),
    .A2(_09978_),
    .A3(_10012_),
    .B1(_10016_),
    .Y(_10017_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_528 ();
 sky130_fd_sc_hd__a211oi_1 _19224_ (.A1(_09998_),
    .A2(_10010_),
    .B1(_10017_),
    .C1(net3902),
    .Y(_10019_));
 sky130_fd_sc_hd__a31oi_1 _19225_ (.A1(net3902),
    .A2(_09992_),
    .A3(_10002_),
    .B1(_10019_),
    .Y(_10020_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_526 ();
 sky130_fd_sc_hd__nand2_8 _19228_ (.A(_09929_),
    .B(_09977_),
    .Y(_10023_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_524 ();
 sky130_fd_sc_hd__nor2_4 _19231_ (.A(_12189_[0]),
    .B(_09977_),
    .Y(_10026_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_523 ();
 sky130_fd_sc_hd__nor2_1 _19233_ (.A(_12196_[0]),
    .B(net3899),
    .Y(_10028_));
 sky130_fd_sc_hd__nor3_1 _19234_ (.A(net3904),
    .B(_10026_),
    .C(_10028_),
    .Y(_10029_));
 sky130_fd_sc_hd__a31oi_1 _19235_ (.A1(net3904),
    .A2(_09975_),
    .A3(_10023_),
    .B1(_10029_),
    .Y(_10030_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_522 ();
 sky130_fd_sc_hd__nor2_2 _19237_ (.A(_12193_[0]),
    .B(_09972_),
    .Y(_10032_));
 sky130_fd_sc_hd__nor2_4 _19238_ (.A(_12190_[0]),
    .B(_09977_),
    .Y(_10033_));
 sky130_fd_sc_hd__o21ai_2 _19239_ (.A1(_10032_),
    .A2(_10033_),
    .B1(net3904),
    .Y(_10034_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_521 ();
 sky130_fd_sc_hd__nor2_4 _19241_ (.A(net3904),
    .B(_09977_),
    .Y(_10036_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_520 ();
 sky130_fd_sc_hd__a21oi_1 _19243_ (.A1(_12188_[0]),
    .A2(_10036_),
    .B1(net3892),
    .Y(_10038_));
 sky130_fd_sc_hd__a221oi_1 _19244_ (.A1(net3892),
    .A2(_10030_),
    .B1(_10034_),
    .B2(_10038_),
    .C1(net3903),
    .Y(_10039_));
 sky130_fd_sc_hd__xnor2_4 _19245_ (.A(net4132),
    .B(_09943_),
    .Y(_10040_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_518 ();
 sky130_fd_sc_hd__clkinvlp_2 _19248_ (.A(_12198_[0]),
    .Y(_10043_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_517 ();
 sky130_fd_sc_hd__nand2_2 _19250_ (.A(_09936_),
    .B(net3894),
    .Y(_10045_));
 sky130_fd_sc_hd__nor2_1 _19251_ (.A(_10043_),
    .B(_10045_),
    .Y(_10046_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_516 ();
 sky130_fd_sc_hd__nand2_1 _19253_ (.A(_12190_[0]),
    .B(net3895),
    .Y(_10048_));
 sky130_fd_sc_hd__nand2_2 _19254_ (.A(_09923_),
    .B(net3905),
    .Y(_10049_));
 sky130_fd_sc_hd__nand2_1 _19255_ (.A(_09998_),
    .B(_10049_),
    .Y(_10050_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_514 ();
 sky130_fd_sc_hd__a21oi_1 _19258_ (.A1(_10048_),
    .A2(_10050_),
    .B1(_09936_),
    .Y(_10053_));
 sky130_fd_sc_hd__nor4_1 _19259_ (.A(_10040_),
    .B(_09972_),
    .C(_10046_),
    .D(_10053_),
    .Y(_10054_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_512 ();
 sky130_fd_sc_hd__a21oi_1 _19262_ (.A1(_09923_),
    .A2(net3905),
    .B1(_09998_),
    .Y(_10057_));
 sky130_fd_sc_hd__a21oi_1 _19263_ (.A1(_12190_[0]),
    .A2(_09998_),
    .B1(_10057_),
    .Y(_10058_));
 sky130_fd_sc_hd__nand2_2 _19264_ (.A(_09936_),
    .B(_09990_),
    .Y(_10059_));
 sky130_fd_sc_hd__o22ai_1 _19265_ (.A1(_09936_),
    .A2(_10058_),
    .B1(_10059_),
    .B2(_12196_[0]),
    .Y(_10060_));
 sky130_fd_sc_hd__o311ai_0 _19266_ (.A1(_10040_),
    .A2(_09977_),
    .A3(_10060_),
    .B1(_09950_),
    .C1(net3901),
    .Y(_10061_));
 sky130_fd_sc_hd__nor3_1 _19267_ (.A(_10039_),
    .B(_10054_),
    .C(_10061_),
    .Y(_10062_));
 sky130_fd_sc_hd__xnor2_4 _19268_ (.A(net3904),
    .B(net3900),
    .Y(_10063_));
 sky130_fd_sc_hd__nor2_2 _19269_ (.A(_12189_[0]),
    .B(_09983_),
    .Y(_10064_));
 sky130_fd_sc_hd__a221oi_1 _19270_ (.A1(_12196_[0]),
    .A2(_10036_),
    .B1(_10063_),
    .B2(_12188_[0]),
    .C1(_10064_),
    .Y(_10065_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_510 ();
 sky130_fd_sc_hd__nand2_2 _19273_ (.A(net3908),
    .B(_09936_),
    .Y(_10068_));
 sky130_fd_sc_hd__nor2_4 _19274_ (.A(_12189_[0]),
    .B(net3904),
    .Y(_10069_));
 sky130_fd_sc_hd__a32oi_1 _19275_ (.A1(_12189_[0]),
    .A2(_09972_),
    .A3(_10068_),
    .B1(_10069_),
    .B2(_09975_),
    .Y(_10070_));
 sky130_fd_sc_hd__nand2_1 _19276_ (.A(net3895),
    .B(_10070_),
    .Y(_10071_));
 sky130_fd_sc_hd__o21ai_0 _19277_ (.A1(net3895),
    .A2(_10065_),
    .B1(_10071_),
    .Y(_10072_));
 sky130_fd_sc_hd__xor2_4 _19278_ (.A(net4133),
    .B(_09956_),
    .X(_10073_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_508 ();
 sky130_fd_sc_hd__nor2_4 _19281_ (.A(_10040_),
    .B(_09950_),
    .Y(_10076_));
 sky130_fd_sc_hd__nand2_2 _19282_ (.A(net3890),
    .B(_10076_),
    .Y(_10077_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_507 ();
 sky130_fd_sc_hd__nand2_1 _19284_ (.A(net3908),
    .B(net3906),
    .Y(_10079_));
 sky130_fd_sc_hd__nand2_8 _19285_ (.A(_09929_),
    .B(net3904),
    .Y(_10080_));
 sky130_fd_sc_hd__nand2_1 _19286_ (.A(_10079_),
    .B(_10080_),
    .Y(_10081_));
 sky130_fd_sc_hd__xnor2_1 _19287_ (.A(net3897),
    .B(_10081_),
    .Y(_10082_));
 sky130_fd_sc_hd__nor2_4 _19288_ (.A(net3906),
    .B(_09977_),
    .Y(_10083_));
 sky130_fd_sc_hd__a221oi_1 _19289_ (.A1(_12188_[0]),
    .A2(_09977_),
    .B1(_10083_),
    .B2(_09923_),
    .C1(net3904),
    .Y(_10084_));
 sky130_fd_sc_hd__nand2_8 _19290_ (.A(_09982_),
    .B(net3899),
    .Y(_10085_));
 sky130_fd_sc_hd__nand2_8 _19291_ (.A(_12196_[0]),
    .B(_09977_),
    .Y(_10086_));
 sky130_fd_sc_hd__nand3_1 _19292_ (.A(net3904),
    .B(_10085_),
    .C(_10086_),
    .Y(_10087_));
 sky130_fd_sc_hd__nand2_1 _19293_ (.A(net3893),
    .B(_10087_),
    .Y(_10088_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_506 ();
 sky130_fd_sc_hd__xor2_4 _19295_ (.A(\u0.tmp_w[23] ),
    .B(_09949_),
    .X(_10090_));
 sky130_fd_sc_hd__nand2_4 _19296_ (.A(net3903),
    .B(_10090_),
    .Y(_10091_));
 sky130_fd_sc_hd__nor2_4 _19297_ (.A(net3890),
    .B(_10091_),
    .Y(_10092_));
 sky130_fd_sc_hd__o221ai_1 _19298_ (.A1(net3893),
    .A2(_10082_),
    .B1(_10084_),
    .B2(_10088_),
    .C1(_10092_),
    .Y(_10093_));
 sky130_fd_sc_hd__nor3_2 _19299_ (.A(net3908),
    .B(_09929_),
    .C(_09936_),
    .Y(_10094_));
 sky130_fd_sc_hd__nor2_2 _19300_ (.A(_12193_[0]),
    .B(net3904),
    .Y(_10095_));
 sky130_fd_sc_hd__o31ai_2 _19301_ (.A1(_09977_),
    .A2(_10094_),
    .A3(_10095_),
    .B1(_09998_),
    .Y(_10096_));
 sky130_fd_sc_hd__nor2_1 _19302_ (.A(_12188_[0]),
    .B(_09983_),
    .Y(_10097_));
 sky130_fd_sc_hd__nand2_2 _19303_ (.A(_12190_[0]),
    .B(_09972_),
    .Y(_10098_));
 sky130_fd_sc_hd__a21oi_1 _19304_ (.A1(_10023_),
    .A2(_10098_),
    .B1(net3904),
    .Y(_10099_));
 sky130_fd_sc_hd__nand2_4 _19305_ (.A(_12189_[0]),
    .B(_09936_),
    .Y(_10100_));
 sky130_fd_sc_hd__nand2_1 _19306_ (.A(_12209_[0]),
    .B(net3896),
    .Y(_10101_));
 sky130_fd_sc_hd__o211ai_1 _19307_ (.A1(net3896),
    .A2(_10100_),
    .B1(_10101_),
    .C1(net3895),
    .Y(_10102_));
 sky130_fd_sc_hd__nand2_1 _19308_ (.A(_09944_),
    .B(_09950_),
    .Y(_10103_));
 sky130_fd_sc_hd__nor2_2 _19309_ (.A(_09957_),
    .B(_10103_),
    .Y(_10104_));
 sky130_fd_sc_hd__o311ai_0 _19310_ (.A1(_10096_),
    .A2(_10097_),
    .A3(_10099_),
    .B1(_10102_),
    .C1(_10104_),
    .Y(_10105_));
 sky130_fd_sc_hd__nor2_4 _19311_ (.A(net3908),
    .B(net3905),
    .Y(_10106_));
 sky130_fd_sc_hd__nor2_2 _19312_ (.A(net3899),
    .B(_10106_),
    .Y(_10107_));
 sky130_fd_sc_hd__nand2_4 _19313_ (.A(_12198_[0]),
    .B(net3899),
    .Y(_10108_));
 sky130_fd_sc_hd__nand2_8 _19314_ (.A(_12189_[0]),
    .B(net3898),
    .Y(_10109_));
 sky130_fd_sc_hd__nor2_4 _19315_ (.A(_09944_),
    .B(_10090_),
    .Y(_10110_));
 sky130_fd_sc_hd__nand2_1 _19316_ (.A(net3891),
    .B(_10110_),
    .Y(_10111_));
 sky130_fd_sc_hd__a41oi_1 _19317_ (.A1(net3904),
    .A2(net3895),
    .A3(_10108_),
    .A4(_10109_),
    .B1(_10111_),
    .Y(_10112_));
 sky130_fd_sc_hd__nor2_2 _19318_ (.A(_12193_[0]),
    .B(_09977_),
    .Y(_10113_));
 sky130_fd_sc_hd__nand2_8 _19319_ (.A(net3906),
    .B(_09977_),
    .Y(_10114_));
 sky130_fd_sc_hd__nor2_1 _19320_ (.A(net3895),
    .B(_10114_),
    .Y(_10115_));
 sky130_fd_sc_hd__o21ai_0 _19321_ (.A1(_10113_),
    .A2(_10115_),
    .B1(net3676),
    .Y(_10116_));
 sky130_fd_sc_hd__o311ai_2 _19322_ (.A1(net3676),
    .A2(net3895),
    .A3(_10107_),
    .B1(_10112_),
    .C1(_10116_),
    .Y(_10117_));
 sky130_fd_sc_hd__o2111ai_2 _19323_ (.A1(_10072_),
    .A2(_10077_),
    .B1(_10093_),
    .C1(_10105_),
    .D1(_10117_),
    .Y(_10118_));
 sky130_fd_sc_hd__a211o_1 _19324_ (.A1(_09952_),
    .A2(_10020_),
    .B1(_10062_),
    .C1(_10118_),
    .X(_00088_));
 sky130_fd_sc_hd__nand2_4 _19325_ (.A(_09923_),
    .B(_10083_),
    .Y(_10119_));
 sky130_fd_sc_hd__nand2_8 _19326_ (.A(_09982_),
    .B(net3898),
    .Y(_10120_));
 sky130_fd_sc_hd__a21oi_1 _19327_ (.A1(_10119_),
    .A2(_10120_),
    .B1(net3676),
    .Y(_10121_));
 sky130_fd_sc_hd__nand2_4 _19328_ (.A(net3891),
    .B(net3892),
    .Y(_10122_));
 sky130_fd_sc_hd__a211oi_1 _19329_ (.A1(net3905),
    .A2(_10036_),
    .B1(_10121_),
    .C1(_10122_),
    .Y(_10123_));
 sky130_fd_sc_hd__nor2_1 _19330_ (.A(net3908),
    .B(net3899),
    .Y(_10124_));
 sky130_fd_sc_hd__nor2_2 _19331_ (.A(_12188_[0]),
    .B(_09977_),
    .Y(_10125_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_505 ();
 sky130_fd_sc_hd__nand2_2 _19333_ (.A(_12193_[0]),
    .B(_09977_),
    .Y(_10127_));
 sky130_fd_sc_hd__nand2_8 _19334_ (.A(net3906),
    .B(net3900),
    .Y(_10128_));
 sky130_fd_sc_hd__nand3_1 _19335_ (.A(net3904),
    .B(_10127_),
    .C(_10128_),
    .Y(_10129_));
 sky130_fd_sc_hd__nor2_2 _19336_ (.A(net3891),
    .B(_09990_),
    .Y(_10130_));
 sky130_fd_sc_hd__o311a_1 _19337_ (.A1(net3904),
    .A2(_10124_),
    .A3(_10125_),
    .B1(_10129_),
    .C1(_10130_),
    .X(_10131_));
 sky130_fd_sc_hd__a21oi_1 _19338_ (.A1(net3898),
    .A2(_10106_),
    .B1(_10033_),
    .Y(_10132_));
 sky130_fd_sc_hd__nand2_8 _19339_ (.A(_12202_[0]),
    .B(_09972_),
    .Y(_10133_));
 sky130_fd_sc_hd__a21oi_1 _19340_ (.A1(_10120_),
    .A2(_10133_),
    .B1(_09936_),
    .Y(_10134_));
 sky130_fd_sc_hd__a21oi_1 _19341_ (.A1(net3676),
    .A2(_10132_),
    .B1(_10134_),
    .Y(_10135_));
 sky130_fd_sc_hd__nand2_8 _19342_ (.A(net3891),
    .B(net3895),
    .Y(_10136_));
 sky130_fd_sc_hd__nand2_4 _19343_ (.A(net3902),
    .B(net3895),
    .Y(_10137_));
 sky130_fd_sc_hd__nand2b_2 _19344_ (.A_N(_12188_[0]),
    .B(net3896),
    .Y(_10138_));
 sky130_fd_sc_hd__a21oi_1 _19345_ (.A1(_10098_),
    .A2(_10138_),
    .B1(_09936_),
    .Y(_10139_));
 sky130_fd_sc_hd__a31oi_1 _19346_ (.A1(_09936_),
    .A2(_10120_),
    .A3(_10128_),
    .B1(_10139_),
    .Y(_10140_));
 sky130_fd_sc_hd__o22ai_1 _19347_ (.A1(_10135_),
    .A2(_10136_),
    .B1(_10137_),
    .B2(_10140_),
    .Y(_10141_));
 sky130_fd_sc_hd__nor4_1 _19348_ (.A(_09950_),
    .B(_10123_),
    .C(_10131_),
    .D(_10141_),
    .Y(_10142_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_504 ();
 sky130_fd_sc_hd__nand2_4 _19350_ (.A(_12193_[0]),
    .B(net3899),
    .Y(_10144_));
 sky130_fd_sc_hd__a21oi_1 _19351_ (.A1(_10120_),
    .A2(_10144_),
    .B1(net3676),
    .Y(_10145_));
 sky130_fd_sc_hd__a21oi_1 _19352_ (.A1(net3676),
    .A2(_10107_),
    .B1(_10145_),
    .Y(_10146_));
 sky130_fd_sc_hd__nand2_1 _19353_ (.A(net3676),
    .B(_09978_),
    .Y(_10147_));
 sky130_fd_sc_hd__nor2_4 _19354_ (.A(_09936_),
    .B(_09972_),
    .Y(_10148_));
 sky130_fd_sc_hd__a21oi_4 _19355_ (.A1(net3908),
    .A2(_10148_),
    .B1(_09998_),
    .Y(_10149_));
 sky130_fd_sc_hd__nand3_1 _19356_ (.A(_10119_),
    .B(_10147_),
    .C(_10149_),
    .Y(_10150_));
 sky130_fd_sc_hd__o21ai_0 _19357_ (.A1(net3895),
    .A2(_10146_),
    .B1(_10150_),
    .Y(_10151_));
 sky130_fd_sc_hd__nand2_8 _19358_ (.A(_09923_),
    .B(_09977_),
    .Y(_10152_));
 sky130_fd_sc_hd__a21oi_1 _19359_ (.A1(_10008_),
    .A2(_10152_),
    .B1(net3905),
    .Y(_10153_));
 sky130_fd_sc_hd__a221oi_2 _19360_ (.A1(net3905),
    .A2(_10148_),
    .B1(_10036_),
    .B2(_09982_),
    .C1(_10153_),
    .Y(_10154_));
 sky130_fd_sc_hd__nand2_4 _19361_ (.A(_12188_[0]),
    .B(net3899),
    .Y(_10155_));
 sky130_fd_sc_hd__and3_1 _19362_ (.A(net3904),
    .B(_10109_),
    .C(_10155_),
    .X(_10156_));
 sky130_fd_sc_hd__a21oi_1 _19363_ (.A1(_09984_),
    .A2(_10127_),
    .B1(net3904),
    .Y(_10157_));
 sky130_fd_sc_hd__nor2_1 _19364_ (.A(_10156_),
    .B(_10157_),
    .Y(_10158_));
 sky130_fd_sc_hd__o221ai_1 _19365_ (.A1(_10122_),
    .A2(_10154_),
    .B1(_10158_),
    .B2(_10136_),
    .C1(_09950_),
    .Y(_10159_));
 sky130_fd_sc_hd__a21oi_1 _19366_ (.A1(net3901),
    .A2(_10151_),
    .B1(_10159_),
    .Y(_10160_));
 sky130_fd_sc_hd__a21oi_1 _19367_ (.A1(_10109_),
    .A2(_10144_),
    .B1(net3676),
    .Y(_10161_));
 sky130_fd_sc_hd__a31oi_1 _19368_ (.A1(net3676),
    .A2(_09984_),
    .A3(_10114_),
    .B1(_10161_),
    .Y(_10162_));
 sky130_fd_sc_hd__nor2_4 _19369_ (.A(_09929_),
    .B(_09972_),
    .Y(_10163_));
 sky130_fd_sc_hd__o21ai_0 _19370_ (.A1(net3904),
    .A2(_10163_),
    .B1(_09923_),
    .Y(_10164_));
 sky130_fd_sc_hd__o2111ai_1 _19371_ (.A1(_09923_),
    .A2(_10128_),
    .B1(_10164_),
    .C1(_09983_),
    .D1(_10130_),
    .Y(_10165_));
 sky130_fd_sc_hd__o21ai_0 _19372_ (.A1(_10137_),
    .A2(_10162_),
    .B1(_10165_),
    .Y(_10166_));
 sky130_fd_sc_hd__nand2_1 _19373_ (.A(_09923_),
    .B(_10063_),
    .Y(_10167_));
 sky130_fd_sc_hd__o21ai_0 _19374_ (.A1(_12193_[0]),
    .A2(_10004_),
    .B1(_10167_),
    .Y(_10168_));
 sky130_fd_sc_hd__nand2_1 _19375_ (.A(_12202_[0]),
    .B(net3904),
    .Y(_10169_));
 sky130_fd_sc_hd__a21oi_1 _19376_ (.A1(_10100_),
    .A2(_10169_),
    .B1(net3899),
    .Y(_10170_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_503 ();
 sky130_fd_sc_hd__o21ai_0 _19378_ (.A1(_10096_),
    .A2(_10170_),
    .B1(net3890),
    .Y(_10172_));
 sky130_fd_sc_hd__a21oi_1 _19379_ (.A1(net3895),
    .A2(_10168_),
    .B1(_10172_),
    .Y(_10173_));
 sky130_fd_sc_hd__nor2_4 _19380_ (.A(_10040_),
    .B(_10090_),
    .Y(_10174_));
 sky130_fd_sc_hd__o21ai_0 _19381_ (.A1(_10166_),
    .A2(_10173_),
    .B1(_10174_),
    .Y(_10175_));
 sky130_fd_sc_hd__and2_4 _19382_ (.A(_12196_[0]),
    .B(_09936_),
    .X(_10176_));
 sky130_fd_sc_hd__nor3_1 _19383_ (.A(net3908),
    .B(net3906),
    .C(_09936_),
    .Y(_10177_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_502 ();
 sky130_fd_sc_hd__o31ai_2 _19385_ (.A1(_09977_),
    .A2(_10176_),
    .A3(_10177_),
    .B1(net3893),
    .Y(_10179_));
 sky130_fd_sc_hd__nor3_1 _19386_ (.A(_12212_[0]),
    .B(net3902),
    .C(net3899),
    .Y(_10180_));
 sky130_fd_sc_hd__nor2_4 _19387_ (.A(_09929_),
    .B(_09936_),
    .Y(_10181_));
 sky130_fd_sc_hd__nor2_1 _19388_ (.A(net3906),
    .B(net3904),
    .Y(_10182_));
 sky130_fd_sc_hd__a21oi_1 _19389_ (.A1(_12188_[0]),
    .A2(_09936_),
    .B1(_10181_),
    .Y(_10183_));
 sky130_fd_sc_hd__o32ai_1 _19390_ (.A1(_10181_),
    .A2(_10152_),
    .A3(_10182_),
    .B1(_10183_),
    .B2(net3897),
    .Y(_10184_));
 sky130_fd_sc_hd__nand3_2 _19391_ (.A(_09936_),
    .B(_09975_),
    .C(_10152_),
    .Y(_10185_));
 sky130_fd_sc_hd__a21oi_1 _19392_ (.A1(_10129_),
    .A2(_10185_),
    .B1(net3901),
    .Y(_10186_));
 sky130_fd_sc_hd__a21oi_1 _19393_ (.A1(net3902),
    .A2(_10184_),
    .B1(_10186_),
    .Y(_10187_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_501 ();
 sky130_fd_sc_hd__o221ai_1 _19395_ (.A1(_10179_),
    .A2(_10180_),
    .B1(_10187_),
    .B2(_09998_),
    .C1(_10076_),
    .Y(_10189_));
 sky130_fd_sc_hd__o311ai_0 _19396_ (.A1(_09944_),
    .A2(_10142_),
    .A3(_10160_),
    .B1(_10175_),
    .C1(_10189_),
    .Y(_00089_));
 sky130_fd_sc_hd__nand2_2 _19397_ (.A(_09923_),
    .B(net3904),
    .Y(_10190_));
 sky130_fd_sc_hd__a21oi_1 _19398_ (.A1(_10079_),
    .A2(_10190_),
    .B1(net3899),
    .Y(_10191_));
 sky130_fd_sc_hd__a21oi_1 _19399_ (.A1(_12212_[0]),
    .A2(net3899),
    .B1(_10191_),
    .Y(_10192_));
 sky130_fd_sc_hd__a21oi_1 _19400_ (.A1(_10120_),
    .A2(_10155_),
    .B1(net3904),
    .Y(_10193_));
 sky130_fd_sc_hd__a21oi_1 _19401_ (.A1(_09975_),
    .A2(_10086_),
    .B1(net3676),
    .Y(_10194_));
 sky130_fd_sc_hd__o21ai_0 _19402_ (.A1(_10193_),
    .A2(_10194_),
    .B1(net3895),
    .Y(_10195_));
 sky130_fd_sc_hd__o21ai_0 _19403_ (.A1(net3895),
    .A2(_10192_),
    .B1(_10195_),
    .Y(_10196_));
 sky130_fd_sc_hd__nand2_2 _19404_ (.A(net3902),
    .B(_10110_),
    .Y(_10197_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_500 ();
 sky130_fd_sc_hd__nor2_2 _19406_ (.A(net3909),
    .B(_09936_),
    .Y(_10199_));
 sky130_fd_sc_hd__nand2_1 _19407_ (.A(_10012_),
    .B(_10068_),
    .Y(_10200_));
 sky130_fd_sc_hd__a222oi_1 _19408_ (.A1(_09994_),
    .A2(_10080_),
    .B1(_10199_),
    .B2(_10023_),
    .C1(_10200_),
    .C2(_12189_[0]),
    .Y(_10201_));
 sky130_fd_sc_hd__nand2_1 _19409_ (.A(_12209_[0]),
    .B(_09972_),
    .Y(_10202_));
 sky130_fd_sc_hd__o311ai_0 _19410_ (.A1(_09972_),
    .A2(_10094_),
    .A3(_10069_),
    .B1(_10202_),
    .C1(net3893),
    .Y(_10203_));
 sky130_fd_sc_hd__o21ai_2 _19411_ (.A1(net3893),
    .A2(_10201_),
    .B1(_10203_),
    .Y(_10204_));
 sky130_fd_sc_hd__o22ai_1 _19412_ (.A1(_10111_),
    .A2(_10196_),
    .B1(_10197_),
    .B2(_10204_),
    .Y(_10205_));
 sky130_fd_sc_hd__nand2_4 _19413_ (.A(_10040_),
    .B(net3889),
    .Y(_10206_));
 sky130_fd_sc_hd__nand3_1 _19414_ (.A(net3676),
    .B(_10127_),
    .C(_10133_),
    .Y(_10207_));
 sky130_fd_sc_hd__nand3_1 _19415_ (.A(net3904),
    .B(_10023_),
    .C(_10108_),
    .Y(_10208_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_499 ();
 sky130_fd_sc_hd__nand2_4 _19417_ (.A(_12198_[0]),
    .B(_09977_),
    .Y(_10210_));
 sky130_fd_sc_hd__nor2_1 _19418_ (.A(_12202_[0]),
    .B(_09977_),
    .Y(_10211_));
 sky130_fd_sc_hd__o21a_1 _19419_ (.A1(_10124_),
    .A2(_10211_),
    .B1(_09936_),
    .X(_10212_));
 sky130_fd_sc_hd__a311oi_2 _19420_ (.A1(net3904),
    .A2(_09984_),
    .A3(_10210_),
    .B1(_10212_),
    .C1(_10073_),
    .Y(_10213_));
 sky130_fd_sc_hd__a311oi_1 _19421_ (.A1(net3891),
    .A2(_10207_),
    .A3(_10208_),
    .B1(_10213_),
    .C1(net3892),
    .Y(_10214_));
 sky130_fd_sc_hd__nand3_1 _19422_ (.A(net3676),
    .B(_10108_),
    .C(_10120_),
    .Y(_10215_));
 sky130_fd_sc_hd__nor2_4 _19423_ (.A(_12189_[0]),
    .B(_09972_),
    .Y(_10216_));
 sky130_fd_sc_hd__nor2_4 _19424_ (.A(_09929_),
    .B(_09977_),
    .Y(_10217_));
 sky130_fd_sc_hd__o21ai_0 _19425_ (.A1(_10216_),
    .A2(_10217_),
    .B1(net3904),
    .Y(_10218_));
 sky130_fd_sc_hd__a311oi_1 _19426_ (.A1(net3904),
    .A2(_10108_),
    .A3(_10152_),
    .B1(_10095_),
    .C1(net3902),
    .Y(_10219_));
 sky130_fd_sc_hd__a311oi_1 _19427_ (.A1(net3902),
    .A2(_10215_),
    .A3(_10218_),
    .B1(_10219_),
    .C1(net3895),
    .Y(_10220_));
 sky130_fd_sc_hd__a32oi_1 _19428_ (.A1(net3904),
    .A2(_10120_),
    .A3(_10155_),
    .B1(_10006_),
    .B2(_12193_[0]),
    .Y(_10221_));
 sky130_fd_sc_hd__a21oi_1 _19429_ (.A1(_12207_[0]),
    .A2(_09977_),
    .B1(_09957_),
    .Y(_10222_));
 sky130_fd_sc_hd__o31ai_1 _19430_ (.A1(net3904),
    .A2(_09977_),
    .A3(_10049_),
    .B1(_10222_),
    .Y(_10223_));
 sky130_fd_sc_hd__o211ai_1 _19431_ (.A1(net3890),
    .A2(_10221_),
    .B1(_10223_),
    .C1(_09998_),
    .Y(_10224_));
 sky130_fd_sc_hd__nor2_4 _19432_ (.A(_12190_[0]),
    .B(_12193_[0]),
    .Y(_10225_));
 sky130_fd_sc_hd__xnor2_1 _19433_ (.A(_09929_),
    .B(_10073_),
    .Y(_10226_));
 sky130_fd_sc_hd__a21oi_1 _19434_ (.A1(net3904),
    .A2(_09957_),
    .B1(_09923_),
    .Y(_10227_));
 sky130_fd_sc_hd__a21oi_1 _19435_ (.A1(_09936_),
    .A2(_10226_),
    .B1(_10227_),
    .Y(_10228_));
 sky130_fd_sc_hd__nor2_1 _19436_ (.A(net3894),
    .B(net3900),
    .Y(_10229_));
 sky130_fd_sc_hd__o311ai_0 _19437_ (.A1(_09936_),
    .A2(net3890),
    .A3(_10225_),
    .B1(_10228_),
    .C1(_10229_),
    .Y(_10230_));
 sky130_fd_sc_hd__nand2_1 _19438_ (.A(_09990_),
    .B(net3900),
    .Y(_10231_));
 sky130_fd_sc_hd__a21oi_1 _19439_ (.A1(_12216_[0]),
    .A2(net3890),
    .B1(_10231_),
    .Y(_10232_));
 sky130_fd_sc_hd__o31ai_1 _19440_ (.A1(net3890),
    .A2(_10176_),
    .A3(_10177_),
    .B1(_10232_),
    .Y(_10233_));
 sky130_fd_sc_hd__nand4_1 _19441_ (.A(_10174_),
    .B(_10224_),
    .C(_10230_),
    .D(_10233_),
    .Y(_10234_));
 sky130_fd_sc_hd__o31ai_1 _19442_ (.A1(_10206_),
    .A2(_10214_),
    .A3(_10220_),
    .B1(_10234_),
    .Y(_10235_));
 sky130_fd_sc_hd__and3_1 _19443_ (.A(_09972_),
    .B(_10100_),
    .C(_10190_),
    .X(_10236_));
 sky130_fd_sc_hd__o21ai_2 _19444_ (.A1(_10094_),
    .A2(_10095_),
    .B1(net3897),
    .Y(_10237_));
 sky130_fd_sc_hd__nand2_4 _19445_ (.A(net3893),
    .B(_10237_),
    .Y(_10238_));
 sky130_fd_sc_hd__nor2_4 _19446_ (.A(_09936_),
    .B(_09977_),
    .Y(_10239_));
 sky130_fd_sc_hd__a21oi_1 _19447_ (.A1(_10023_),
    .A2(_10133_),
    .B1(net3904),
    .Y(_10240_));
 sky130_fd_sc_hd__a211oi_1 _19448_ (.A1(_12193_[0]),
    .A2(_10239_),
    .B1(_10240_),
    .C1(_09994_),
    .Y(_10241_));
 sky130_fd_sc_hd__o22a_1 _19449_ (.A1(_10236_),
    .A2(_10238_),
    .B1(_10241_),
    .B2(net3893),
    .X(_10242_));
 sky130_fd_sc_hd__a21oi_2 _19450_ (.A1(_12190_[0]),
    .A2(net3897),
    .B1(_10014_),
    .Y(_10243_));
 sky130_fd_sc_hd__nand3_1 _19451_ (.A(net3904),
    .B(_10085_),
    .C(_10114_),
    .Y(_10244_));
 sky130_fd_sc_hd__o211ai_1 _19452_ (.A1(net3904),
    .A2(_10243_),
    .B1(_10244_),
    .C1(net3895),
    .Y(_10245_));
 sky130_fd_sc_hd__nand2_1 _19453_ (.A(_09923_),
    .B(_09936_),
    .Y(_10246_));
 sky130_fd_sc_hd__o32ai_1 _19454_ (.A1(_10083_),
    .A2(_10163_),
    .A3(_10246_),
    .B1(_09983_),
    .B2(_12202_[0]),
    .Y(_10247_));
 sky130_fd_sc_hd__nand2_1 _19455_ (.A(net3893),
    .B(_10247_),
    .Y(_10248_));
 sky130_fd_sc_hd__nand3_1 _19456_ (.A(_10092_),
    .B(_10245_),
    .C(_10248_),
    .Y(_10249_));
 sky130_fd_sc_hd__o21ai_2 _19457_ (.A1(_10077_),
    .A2(_10242_),
    .B1(_10249_),
    .Y(_10250_));
 sky130_fd_sc_hd__or3_1 _19458_ (.A(_10205_),
    .B(_10235_),
    .C(_10250_),
    .X(_00090_));
 sky130_fd_sc_hd__nand2_2 _19459_ (.A(_09929_),
    .B(_09936_),
    .Y(_10251_));
 sky130_fd_sc_hd__o2111ai_2 _19460_ (.A1(net3890),
    .A2(_10128_),
    .B1(_10251_),
    .C1(_09983_),
    .D1(_09923_),
    .Y(_10252_));
 sky130_fd_sc_hd__nand2_1 _19461_ (.A(net3890),
    .B(_10083_),
    .Y(_10253_));
 sky130_fd_sc_hd__o21ai_0 _19462_ (.A1(net3890),
    .A2(_10086_),
    .B1(_10253_),
    .Y(_10254_));
 sky130_fd_sc_hd__a32oi_1 _19463_ (.A1(net3902),
    .A2(_09972_),
    .A3(_10069_),
    .B1(_10254_),
    .B2(net3904),
    .Y(_10255_));
 sky130_fd_sc_hd__nand3_1 _19464_ (.A(net3893),
    .B(_10252_),
    .C(_10255_),
    .Y(_10256_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_498 ();
 sky130_fd_sc_hd__a221oi_1 _19466_ (.A1(_12196_[0]),
    .A2(_10036_),
    .B1(_10163_),
    .B2(net3908),
    .C1(_10137_),
    .Y(_10257_));
 sky130_fd_sc_hd__a21oi_4 _19467_ (.A1(_10085_),
    .A2(_10152_),
    .B1(_09936_),
    .Y(_10258_));
 sky130_fd_sc_hd__a21oi_1 _19468_ (.A1(_09978_),
    .A2(_10108_),
    .B1(net3904),
    .Y(_10259_));
 sky130_fd_sc_hd__nor2_1 _19469_ (.A(_10258_),
    .B(_10259_),
    .Y(_10260_));
 sky130_fd_sc_hd__nor2_1 _19470_ (.A(_10136_),
    .B(_10260_),
    .Y(_10261_));
 sky130_fd_sc_hd__a21oi_1 _19471_ (.A1(_10244_),
    .A2(_10257_),
    .B1(_10261_),
    .Y(_10262_));
 sky130_fd_sc_hd__o21ai_0 _19472_ (.A1(_12198_[0]),
    .A2(net3904),
    .B1(net3897),
    .Y(_10263_));
 sky130_fd_sc_hd__a21oi_1 _19473_ (.A1(net3904),
    .A2(_10225_),
    .B1(_10263_),
    .Y(_10264_));
 sky130_fd_sc_hd__nor3_1 _19474_ (.A(net3902),
    .B(_10179_),
    .C(_10264_),
    .Y(_10265_));
 sky130_fd_sc_hd__nand2_2 _19475_ (.A(_09957_),
    .B(net3892),
    .Y(_10266_));
 sky130_fd_sc_hd__a21oi_1 _19476_ (.A1(net3904),
    .A2(_09975_),
    .B1(net3906),
    .Y(_10267_));
 sky130_fd_sc_hd__a2111oi_0 _19477_ (.A1(_09923_),
    .A2(_10036_),
    .B1(_10097_),
    .C1(_10266_),
    .D1(_10267_),
    .Y(_10268_));
 sky130_fd_sc_hd__a21oi_4 _19478_ (.A1(_09967_),
    .A2(_09971_),
    .B1(_10043_),
    .Y(_10269_));
 sky130_fd_sc_hd__a21oi_4 _19479_ (.A1(_12189_[0]),
    .A2(net3900),
    .B1(_10269_),
    .Y(_10270_));
 sky130_fd_sc_hd__nand2_1 _19480_ (.A(net3902),
    .B(_10270_),
    .Y(_10271_));
 sky130_fd_sc_hd__nand2_1 _19481_ (.A(net3890),
    .B(_10217_),
    .Y(_10272_));
 sky130_fd_sc_hd__nor2_2 _19482_ (.A(net3905),
    .B(net3899),
    .Y(_10273_));
 sky130_fd_sc_hd__a211oi_1 _19483_ (.A1(net3902),
    .A2(_10273_),
    .B1(net3582),
    .C1(net3904),
    .Y(_10274_));
 sky130_fd_sc_hd__a311oi_1 _19484_ (.A1(net3904),
    .A2(_10271_),
    .A3(_10272_),
    .B1(_09998_),
    .C1(_10274_),
    .Y(_10275_));
 sky130_fd_sc_hd__nor3_2 _19485_ (.A(_10265_),
    .B(_10268_),
    .C(_10275_),
    .Y(_10276_));
 sky130_fd_sc_hd__nor2_1 _19486_ (.A(_10206_),
    .B(_10276_),
    .Y(_10277_));
 sky130_fd_sc_hd__nor2_1 _19487_ (.A(net3909),
    .B(_10251_),
    .Y(_10278_));
 sky130_fd_sc_hd__a311oi_1 _19488_ (.A1(net3909),
    .A2(net3900),
    .A3(_10080_),
    .B1(_10278_),
    .C1(_09990_),
    .Y(_10279_));
 sky130_fd_sc_hd__nor2_1 _19489_ (.A(net3906),
    .B(_09936_),
    .Y(_10280_));
 sky130_fd_sc_hd__a211oi_1 _19490_ (.A1(_09923_),
    .A2(_10036_),
    .B1(_10280_),
    .C1(net3894),
    .Y(_10281_));
 sky130_fd_sc_hd__xnor2_1 _19491_ (.A(_09936_),
    .B(net3894),
    .Y(_10282_));
 sky130_fd_sc_hd__o221ai_1 _19492_ (.A1(_09923_),
    .A2(_10045_),
    .B1(_10282_),
    .B2(_12189_[0]),
    .C1(_09977_),
    .Y(_10283_));
 sky130_fd_sc_hd__o211ai_1 _19493_ (.A1(_10279_),
    .A2(_10281_),
    .B1(_10104_),
    .C1(_10283_),
    .Y(_10284_));
 sky130_fd_sc_hd__nand2_2 _19494_ (.A(_12189_[0]),
    .B(net3900),
    .Y(_10285_));
 sky130_fd_sc_hd__o211ai_1 _19495_ (.A1(_12202_[0]),
    .A2(net3900),
    .B1(_10285_),
    .C1(net3904),
    .Y(_10286_));
 sky130_fd_sc_hd__o31a_1 _19496_ (.A1(net3904),
    .A2(_10014_),
    .A3(_10032_),
    .B1(_10286_),
    .X(_10287_));
 sky130_fd_sc_hd__o211ai_1 _19497_ (.A1(_12196_[0]),
    .A2(net3896),
    .B1(_10138_),
    .C1(net3904),
    .Y(_10288_));
 sky130_fd_sc_hd__o311ai_0 _19498_ (.A1(net3904),
    .A2(_10083_),
    .A3(_10216_),
    .B1(_10288_),
    .C1(_09990_),
    .Y(_10289_));
 sky130_fd_sc_hd__o2111ai_1 _19499_ (.A1(_09990_),
    .A2(_10287_),
    .B1(_10289_),
    .C1(_10174_),
    .D1(_09957_),
    .Y(_10290_));
 sky130_fd_sc_hd__nand2_1 _19500_ (.A(_12198_[0]),
    .B(net3894),
    .Y(_10291_));
 sky130_fd_sc_hd__nor2_4 _19501_ (.A(_09990_),
    .B(_09977_),
    .Y(_10292_));
 sky130_fd_sc_hd__nand2_1 _19502_ (.A(_12190_[0]),
    .B(_09977_),
    .Y(_10293_));
 sky130_fd_sc_hd__a21oi_1 _19503_ (.A1(_10085_),
    .A2(_10293_),
    .B1(net3893),
    .Y(_10294_));
 sky130_fd_sc_hd__a21oi_1 _19504_ (.A1(_09929_),
    .A2(_10292_),
    .B1(_10294_),
    .Y(_10295_));
 sky130_fd_sc_hd__o221ai_1 _19505_ (.A1(_10291_),
    .A2(_10063_),
    .B1(_10295_),
    .B2(_09936_),
    .C1(_10092_),
    .Y(_10296_));
 sky130_fd_sc_hd__nor2_1 _19506_ (.A(_12196_[0]),
    .B(net3896),
    .Y(_10297_));
 sky130_fd_sc_hd__nor3_1 _19507_ (.A(net3904),
    .B(_10216_),
    .C(_10297_),
    .Y(_10298_));
 sky130_fd_sc_hd__a21o_1 _19508_ (.A1(net3904),
    .A2(_10243_),
    .B1(_10298_),
    .X(_10299_));
 sky130_fd_sc_hd__a21oi_1 _19509_ (.A1(_09978_),
    .A2(_09984_),
    .B1(net3904),
    .Y(_10300_));
 sky130_fd_sc_hd__a211oi_1 _19510_ (.A1(net3896),
    .A2(_10225_),
    .B1(_10026_),
    .C1(_09936_),
    .Y(_10301_));
 sky130_fd_sc_hd__o21ai_0 _19511_ (.A1(_10300_),
    .A2(_10301_),
    .B1(net3893),
    .Y(_10302_));
 sky130_fd_sc_hd__o2111ai_1 _19512_ (.A1(net3893),
    .A2(_10299_),
    .B1(_10302_),
    .C1(_10076_),
    .D1(net3890),
    .Y(_10303_));
 sky130_fd_sc_hd__nand4_1 _19513_ (.A(_10284_),
    .B(_10290_),
    .C(_10296_),
    .D(_10303_),
    .Y(_10304_));
 sky130_fd_sc_hd__a311oi_1 _19514_ (.A1(_10110_),
    .A2(_10256_),
    .A3(_10262_),
    .B1(_10277_),
    .C1(_10304_),
    .Y(_00091_));
 sky130_fd_sc_hd__o22ai_1 _19515_ (.A1(_12202_[0]),
    .A2(_10004_),
    .B1(_10217_),
    .B2(_09936_),
    .Y(_10305_));
 sky130_fd_sc_hd__and2_4 _19516_ (.A(_12193_[0]),
    .B(_09977_),
    .X(_10306_));
 sky130_fd_sc_hd__o311ai_0 _19517_ (.A1(_09936_),
    .A2(_10306_),
    .A3(_10125_),
    .B1(_10185_),
    .C1(_09990_),
    .Y(_10307_));
 sky130_fd_sc_hd__o21ai_0 _19518_ (.A1(_09990_),
    .A2(_10305_),
    .B1(_10307_),
    .Y(_10308_));
 sky130_fd_sc_hd__a21oi_1 _19519_ (.A1(_09977_),
    .A2(_10106_),
    .B1(_10113_),
    .Y(_10309_));
 sky130_fd_sc_hd__nand2_1 _19520_ (.A(net3904),
    .B(_10309_),
    .Y(_10310_));
 sky130_fd_sc_hd__o21ai_0 _19521_ (.A1(_10273_),
    .A2(_10026_),
    .B1(_09936_),
    .Y(_10311_));
 sky130_fd_sc_hd__o21ai_0 _19522_ (.A1(_10059_),
    .A2(_10132_),
    .B1(net3901),
    .Y(_10312_));
 sky130_fd_sc_hd__a31oi_1 _19523_ (.A1(net3892),
    .A2(_10310_),
    .A3(_10311_),
    .B1(_10312_),
    .Y(_10313_));
 sky130_fd_sc_hd__a21oi_1 _19524_ (.A1(net3891),
    .A2(_10308_),
    .B1(_10313_),
    .Y(_10314_));
 sky130_fd_sc_hd__nor2_4 _19525_ (.A(_12190_[0]),
    .B(_09936_),
    .Y(_10315_));
 sky130_fd_sc_hd__a21oi_1 _19526_ (.A1(_12188_[0]),
    .A2(_09936_),
    .B1(_10315_),
    .Y(_10316_));
 sky130_fd_sc_hd__o21ai_0 _19527_ (.A1(_10163_),
    .A2(_10182_),
    .B1(_12198_[0]),
    .Y(_10317_));
 sky130_fd_sc_hd__a21oi_1 _19528_ (.A1(_10012_),
    .A2(_10181_),
    .B1(_10083_),
    .Y(_10318_));
 sky130_fd_sc_hd__a21oi_2 _19529_ (.A1(_10317_),
    .A2(_10318_),
    .B1(_09998_),
    .Y(_10319_));
 sky130_fd_sc_hd__o21ai_0 _19530_ (.A1(_09998_),
    .A2(net3899),
    .B1(net3904),
    .Y(_10320_));
 sky130_fd_sc_hd__o21ai_0 _19531_ (.A1(_10059_),
    .A2(_10269_),
    .B1(_10049_),
    .Y(_10321_));
 sky130_fd_sc_hd__a21oi_1 _19532_ (.A1(_09929_),
    .A2(_10320_),
    .B1(_10321_),
    .Y(_10322_));
 sky130_fd_sc_hd__a2111oi_0 _19533_ (.A1(_10292_),
    .A2(_10316_),
    .B1(_10319_),
    .C1(_10322_),
    .D1(net3901),
    .Y(_10323_));
 sky130_fd_sc_hd__nor2_1 _19534_ (.A(_12200_[0]),
    .B(net3897),
    .Y(_10324_));
 sky130_fd_sc_hd__a21oi_2 _19535_ (.A1(net3897),
    .A2(_10100_),
    .B1(_10324_),
    .Y(_10325_));
 sky130_fd_sc_hd__o221ai_1 _19536_ (.A1(net3908),
    .A2(_10128_),
    .B1(_10269_),
    .B2(net3904),
    .C1(_10149_),
    .Y(_10326_));
 sky130_fd_sc_hd__o21ai_0 _19537_ (.A1(net3895),
    .A2(_10325_),
    .B1(_10326_),
    .Y(_10327_));
 sky130_fd_sc_hd__nand2_1 _19538_ (.A(net3908),
    .B(_09990_),
    .Y(_10328_));
 sky130_fd_sc_hd__a21boi_0 _19539_ (.A1(_12188_[0]),
    .A2(_10292_),
    .B1_N(_10328_),
    .Y(_10329_));
 sky130_fd_sc_hd__o2bb2ai_1 _19540_ (.A1_N(_10292_),
    .A2_N(_10315_),
    .B1(_10329_),
    .B2(net3904),
    .Y(_10330_));
 sky130_fd_sc_hd__a31oi_1 _19541_ (.A1(_10073_),
    .A2(_10210_),
    .A3(_10330_),
    .B1(_10091_),
    .Y(_10331_));
 sky130_fd_sc_hd__o21ai_1 _19542_ (.A1(_10073_),
    .A2(_10327_),
    .B1(_10331_),
    .Y(_10332_));
 sky130_fd_sc_hd__nand3_1 _19543_ (.A(_09936_),
    .B(_10152_),
    .C(_10155_),
    .Y(_10333_));
 sky130_fd_sc_hd__a21oi_1 _19544_ (.A1(_09936_),
    .A2(_10210_),
    .B1(_10033_),
    .Y(_10334_));
 sky130_fd_sc_hd__nor2_1 _19545_ (.A(net3892),
    .B(_10334_),
    .Y(_10335_));
 sky130_fd_sc_hd__a311oi_1 _19546_ (.A1(net3892),
    .A2(_10080_),
    .A3(_10333_),
    .B1(_10335_),
    .C1(net3891),
    .Y(_10336_));
 sky130_fd_sc_hd__nand2_1 _19547_ (.A(net3909),
    .B(_10163_),
    .Y(_10337_));
 sky130_fd_sc_hd__nand2_1 _19548_ (.A(_09929_),
    .B(_10239_),
    .Y(_10338_));
 sky130_fd_sc_hd__o211ai_1 _19549_ (.A1(net3908),
    .A2(_10063_),
    .B1(_10337_),
    .C1(_10338_),
    .Y(_10339_));
 sky130_fd_sc_hd__a221oi_1 _19550_ (.A1(net3908),
    .A2(net3904),
    .B1(_10006_),
    .B2(_12188_[0]),
    .C1(_10136_),
    .Y(_10340_));
 sky130_fd_sc_hd__a21oi_1 _19551_ (.A1(_10119_),
    .A2(_10340_),
    .B1(_09944_),
    .Y(_10341_));
 sky130_fd_sc_hd__o21ai_0 _19552_ (.A1(_10122_),
    .A2(_10339_),
    .B1(_10341_),
    .Y(_10342_));
 sky130_fd_sc_hd__nor3_4 _19553_ (.A(net3907),
    .B(_09929_),
    .C(net3899),
    .Y(_10343_));
 sky130_fd_sc_hd__nor3_1 _19554_ (.A(_09990_),
    .B(net3582),
    .C(_10343_),
    .Y(_10344_));
 sky130_fd_sc_hd__a211oi_1 _19555_ (.A1(_12198_[0]),
    .A2(_09990_),
    .B1(_10344_),
    .C1(_09936_),
    .Y(_10345_));
 sky130_fd_sc_hd__nand2_1 _19556_ (.A(_09998_),
    .B(_10270_),
    .Y(_10346_));
 sky130_fd_sc_hd__nand3_1 _19557_ (.A(net3895),
    .B(_10109_),
    .C(_10144_),
    .Y(_10347_));
 sky130_fd_sc_hd__a21oi_1 _19558_ (.A1(_10346_),
    .A2(_10347_),
    .B1(net3904),
    .Y(_10348_));
 sky130_fd_sc_hd__nor3_1 _19559_ (.A(net3891),
    .B(_10345_),
    .C(_10348_),
    .Y(_10349_));
 sky130_fd_sc_hd__o21ai_0 _19560_ (.A1(_12188_[0]),
    .A2(_09936_),
    .B1(_10246_),
    .Y(_10350_));
 sky130_fd_sc_hd__a21oi_2 _19561_ (.A1(_09977_),
    .A2(_10350_),
    .B1(_10096_),
    .Y(_10351_));
 sky130_fd_sc_hd__nand2_1 _19562_ (.A(_10152_),
    .B(_10133_),
    .Y(_10352_));
 sky130_fd_sc_hd__nor3_1 _19563_ (.A(_09936_),
    .B(_10113_),
    .C(_10343_),
    .Y(_10353_));
 sky130_fd_sc_hd__a211oi_1 _19564_ (.A1(_09936_),
    .A2(_10352_),
    .B1(_10353_),
    .C1(net3892),
    .Y(_10354_));
 sky130_fd_sc_hd__o31ai_1 _19565_ (.A1(net3901),
    .A2(_10351_),
    .A3(_10354_),
    .B1(net3903),
    .Y(_10355_));
 sky130_fd_sc_hd__o221ai_1 _19566_ (.A1(_10336_),
    .A2(_10342_),
    .B1(_10349_),
    .B2(_10355_),
    .C1(_09950_),
    .Y(_10356_));
 sky130_fd_sc_hd__o221ai_1 _19567_ (.A1(_10206_),
    .A2(_10314_),
    .B1(_10323_),
    .B2(_10332_),
    .C1(_10356_),
    .Y(_00092_));
 sky130_fd_sc_hd__nor2_4 _19568_ (.A(net3909),
    .B(_09977_),
    .Y(_10357_));
 sky130_fd_sc_hd__o21ai_0 _19569_ (.A1(_09929_),
    .A2(_10357_),
    .B1(_10338_),
    .Y(_10358_));
 sky130_fd_sc_hd__a211oi_1 _19570_ (.A1(_10043_),
    .A2(net3900),
    .B1(_10343_),
    .C1(net3904),
    .Y(_10359_));
 sky130_fd_sc_hd__a311oi_1 _19571_ (.A1(net3904),
    .A2(_09975_),
    .A3(_10120_),
    .B1(_10359_),
    .C1(_09998_),
    .Y(_10360_));
 sky130_fd_sc_hd__a21oi_1 _19572_ (.A1(net3894),
    .A2(_10358_),
    .B1(_10360_),
    .Y(_10361_));
 sky130_fd_sc_hd__o21ai_0 _19573_ (.A1(net3909),
    .A2(_09929_),
    .B1(net3900),
    .Y(_10362_));
 sky130_fd_sc_hd__a21oi_1 _19574_ (.A1(_10293_),
    .A2(_10362_),
    .B1(_09936_),
    .Y(_10363_));
 sky130_fd_sc_hd__a211oi_1 _19575_ (.A1(_12198_[0]),
    .A2(_10036_),
    .B1(_10306_),
    .C1(_10363_),
    .Y(_10364_));
 sky130_fd_sc_hd__nand3_1 _19576_ (.A(_09936_),
    .B(_09975_),
    .C(_09978_),
    .Y(_10365_));
 sky130_fd_sc_hd__a31oi_1 _19577_ (.A1(net3893),
    .A2(_10034_),
    .A3(_10365_),
    .B1(_10197_),
    .Y(_10366_));
 sky130_fd_sc_hd__o21ai_0 _19578_ (.A1(net3894),
    .A2(_10364_),
    .B1(_10366_),
    .Y(_10367_));
 sky130_fd_sc_hd__o41ai_1 _19579_ (.A1(_09944_),
    .A2(_09950_),
    .A3(net3890),
    .A4(_10361_),
    .B1(_10367_),
    .Y(_10368_));
 sky130_fd_sc_hd__nand2_1 _19580_ (.A(_09923_),
    .B(_09929_),
    .Y(_10369_));
 sky130_fd_sc_hd__nor3b_2 _19581_ (.A(net3582),
    .B(net3904),
    .C_N(_10086_),
    .Y(_10370_));
 sky130_fd_sc_hd__a21oi_1 _19582_ (.A1(_10239_),
    .A2(_10369_),
    .B1(_10370_),
    .Y(_10371_));
 sky130_fd_sc_hd__a221oi_1 _19583_ (.A1(_10148_),
    .A2(_10106_),
    .B1(_10063_),
    .B2(net3905),
    .C1(net3895),
    .Y(_10372_));
 sky130_fd_sc_hd__o21ai_0 _19584_ (.A1(_12193_[0]),
    .A2(_10004_),
    .B1(_10372_),
    .Y(_10373_));
 sky130_fd_sc_hd__o2111ai_1 _19585_ (.A1(net3894),
    .A2(_10371_),
    .B1(_10373_),
    .C1(_10040_),
    .D1(net3890),
    .Y(_10374_));
 sky130_fd_sc_hd__a21oi_1 _19586_ (.A1(_10138_),
    .A2(_10133_),
    .B1(net3904),
    .Y(_10375_));
 sky130_fd_sc_hd__o21ai_0 _19587_ (.A1(_10064_),
    .A2(_10375_),
    .B1(_09944_),
    .Y(_10376_));
 sky130_fd_sc_hd__a221oi_1 _19588_ (.A1(_09929_),
    .A2(_10006_),
    .B1(_10270_),
    .B2(net3904),
    .C1(_09944_),
    .Y(_10377_));
 sky130_fd_sc_hd__nor2_1 _19589_ (.A(_10122_),
    .B(_10377_),
    .Y(_10378_));
 sky130_fd_sc_hd__a21oi_1 _19590_ (.A1(net3904),
    .A2(_10144_),
    .B1(_10343_),
    .Y(_10379_));
 sky130_fd_sc_hd__nor3_1 _19591_ (.A(_09944_),
    .B(_10136_),
    .C(_10379_),
    .Y(_10380_));
 sky130_fd_sc_hd__a21oi_1 _19592_ (.A1(_10098_),
    .A2(_10109_),
    .B1(net3904),
    .Y(_10381_));
 sky130_fd_sc_hd__a2111oi_0 _19593_ (.A1(net3908),
    .A2(_10239_),
    .B1(_10136_),
    .C1(_10381_),
    .D1(_10040_),
    .Y(_10382_));
 sky130_fd_sc_hd__a211oi_1 _19594_ (.A1(_10376_),
    .A2(_10378_),
    .B1(_10380_),
    .C1(_10382_),
    .Y(_10383_));
 sky130_fd_sc_hd__mux2i_1 _19595_ (.A0(_10374_),
    .A1(_10383_),
    .S(_09950_),
    .Y(_10384_));
 sky130_fd_sc_hd__a211oi_1 _19596_ (.A1(_09990_),
    .A2(_10148_),
    .B1(_10292_),
    .C1(net3908),
    .Y(_10385_));
 sky130_fd_sc_hd__a21oi_1 _19597_ (.A1(net3908),
    .A2(_10231_),
    .B1(_10385_),
    .Y(_10386_));
 sky130_fd_sc_hd__a22oi_1 _19598_ (.A1(net3906),
    .A2(_10239_),
    .B1(_10006_),
    .B2(_12196_[0]),
    .Y(_10387_));
 sky130_fd_sc_hd__nor2_1 _19599_ (.A(_09990_),
    .B(net3900),
    .Y(_10388_));
 sky130_fd_sc_hd__o21ai_0 _19600_ (.A1(_10239_),
    .A2(_10388_),
    .B1(net3908),
    .Y(_10389_));
 sky130_fd_sc_hd__o21ai_0 _19601_ (.A1(net3894),
    .A2(_10387_),
    .B1(_10389_),
    .Y(_10390_));
 sky130_fd_sc_hd__a21oi_1 _19602_ (.A1(_09929_),
    .A2(_10386_),
    .B1(_10390_),
    .Y(_10391_));
 sky130_fd_sc_hd__nor3_1 _19603_ (.A(net3890),
    .B(_10103_),
    .C(_10391_),
    .Y(_10392_));
 sky130_fd_sc_hd__o21ai_0 _19604_ (.A1(net3890),
    .A2(_09997_),
    .B1(_10080_),
    .Y(_10393_));
 sky130_fd_sc_hd__nand3_1 _19605_ (.A(net3904),
    .B(_09957_),
    .C(_10225_),
    .Y(_10394_));
 sky130_fd_sc_hd__nand2_1 _19606_ (.A(_12196_[0]),
    .B(net3890),
    .Y(_10395_));
 sky130_fd_sc_hd__a21oi_1 _19607_ (.A1(_10394_),
    .A2(_10395_),
    .B1(net3900),
    .Y(_10396_));
 sky130_fd_sc_hd__a21oi_1 _19608_ (.A1(_10357_),
    .A2(_10393_),
    .B1(_10396_),
    .Y(_10397_));
 sky130_fd_sc_hd__a311o_1 _19609_ (.A1(net3904),
    .A2(_10285_),
    .A3(_10120_),
    .B1(_10370_),
    .C1(_09957_),
    .X(_10398_));
 sky130_fd_sc_hd__nand2_1 _19610_ (.A(_12193_[0]),
    .B(_10036_),
    .Y(_10399_));
 sky130_fd_sc_hd__o21ai_0 _19611_ (.A1(_12202_[0]),
    .A2(net3904),
    .B1(_09977_),
    .Y(_10400_));
 sky130_fd_sc_hd__a31oi_1 _19612_ (.A1(_09957_),
    .A2(_10399_),
    .A3(_10400_),
    .B1(net3894),
    .Y(_10401_));
 sky130_fd_sc_hd__a221oi_1 _19613_ (.A1(net3894),
    .A2(_10397_),
    .B1(_10398_),
    .B2(_10401_),
    .C1(_10091_),
    .Y(_10402_));
 sky130_fd_sc_hd__nor4_1 _19614_ (.A(_10368_),
    .B(_10384_),
    .C(_10392_),
    .D(_10402_),
    .Y(_00093_));
 sky130_fd_sc_hd__a211oi_1 _19615_ (.A1(_09972_),
    .A2(_10225_),
    .B1(_10343_),
    .C1(_09936_),
    .Y(_10403_));
 sky130_fd_sc_hd__a21oi_1 _19616_ (.A1(_10085_),
    .A2(_10114_),
    .B1(net3904),
    .Y(_10404_));
 sky130_fd_sc_hd__o21ai_0 _19617_ (.A1(net3908),
    .A2(_10280_),
    .B1(_09977_),
    .Y(_10405_));
 sky130_fd_sc_hd__o211ai_1 _19618_ (.A1(_12196_[0]),
    .A2(_10004_),
    .B1(_10405_),
    .C1(net3895),
    .Y(_10406_));
 sky130_fd_sc_hd__o311ai_0 _19619_ (.A1(net3895),
    .A2(_10403_),
    .A3(_10404_),
    .B1(_10406_),
    .C1(net3890),
    .Y(_10407_));
 sky130_fd_sc_hd__nor3_1 _19620_ (.A(net3904),
    .B(_10033_),
    .C(_10343_),
    .Y(_10408_));
 sky130_fd_sc_hd__nor2_1 _19621_ (.A(net3904),
    .B(_10049_),
    .Y(_10409_));
 sky130_fd_sc_hd__o21ai_0 _19622_ (.A1(_12189_[0]),
    .A2(_09936_),
    .B1(_09972_),
    .Y(_10410_));
 sky130_fd_sc_hd__o221ai_1 _19623_ (.A1(_12207_[0]),
    .A2(_09972_),
    .B1(_10409_),
    .B2(_10410_),
    .C1(net3895),
    .Y(_10411_));
 sky130_fd_sc_hd__o311ai_0 _19624_ (.A1(net3895),
    .A2(_10258_),
    .A3(_10408_),
    .B1(_10411_),
    .C1(_09957_),
    .Y(_10412_));
 sky130_fd_sc_hd__nor3_1 _19625_ (.A(_09936_),
    .B(_10217_),
    .C(_10269_),
    .Y(_10413_));
 sky130_fd_sc_hd__nor2_1 _19626_ (.A(_09972_),
    .B(_10225_),
    .Y(_10414_));
 sky130_fd_sc_hd__nor3_1 _19627_ (.A(net3904),
    .B(_10026_),
    .C(_10414_),
    .Y(_10415_));
 sky130_fd_sc_hd__o21ai_0 _19628_ (.A1(_10413_),
    .A2(_10415_),
    .B1(net3890),
    .Y(_10416_));
 sky130_fd_sc_hd__o21ai_0 _19629_ (.A1(_10125_),
    .A2(_10269_),
    .B1(net3904),
    .Y(_10417_));
 sky130_fd_sc_hd__a21oi_1 _19630_ (.A1(_12190_[0]),
    .A2(_10006_),
    .B1(net3890),
    .Y(_10418_));
 sky130_fd_sc_hd__a21oi_1 _19631_ (.A1(_10417_),
    .A2(_10418_),
    .B1(net3892),
    .Y(_10419_));
 sky130_fd_sc_hd__a21oi_1 _19632_ (.A1(_10416_),
    .A2(_10419_),
    .B1(net3903),
    .Y(_10420_));
 sky130_fd_sc_hd__o21ai_2 _19633_ (.A1(_09923_),
    .A2(_09936_),
    .B1(_10107_),
    .Y(_10421_));
 sky130_fd_sc_hd__or3_4 _19634_ (.A(_12205_[0]),
    .B(_12214_[0]),
    .C(net3897),
    .X(_10422_));
 sky130_fd_sc_hd__a21oi_2 _19635_ (.A1(_12198_[0]),
    .A2(_09936_),
    .B1(net3897),
    .Y(_10423_));
 sky130_fd_sc_hd__a21oi_2 _19636_ (.A1(_10169_),
    .A2(_10423_),
    .B1(_10122_),
    .Y(_10424_));
 sky130_fd_sc_hd__a32oi_1 _19637_ (.A1(net3676),
    .A2(_10106_),
    .A3(_10108_),
    .B1(_10133_),
    .B2(_10315_),
    .Y(_10425_));
 sky130_fd_sc_hd__a32oi_2 _19638_ (.A1(_10130_),
    .A2(_10421_),
    .A3(_10422_),
    .B1(_10424_),
    .B2(_10425_),
    .Y(_10426_));
 sky130_fd_sc_hd__a32o_1 _19639_ (.A1(_09944_),
    .A2(_10407_),
    .A3(_10412_),
    .B1(_10420_),
    .B2(_10426_),
    .X(_10427_));
 sky130_fd_sc_hd__a21oi_1 _19640_ (.A1(net3909),
    .A2(_10181_),
    .B1(_10083_),
    .Y(_10428_));
 sky130_fd_sc_hd__o2111a_1 _19641_ (.A1(_12202_[0]),
    .A2(_10428_),
    .B1(_10337_),
    .C1(_10251_),
    .D1(_09990_),
    .X(_10429_));
 sky130_fd_sc_hd__a21oi_2 _19642_ (.A1(_09929_),
    .A2(_10148_),
    .B1(_10050_),
    .Y(_10430_));
 sky130_fd_sc_hd__o21ai_0 _19643_ (.A1(net3894),
    .A2(net3582),
    .B1(_10199_),
    .Y(_10431_));
 sky130_fd_sc_hd__o211ai_1 _19644_ (.A1(_10429_),
    .A2(_10430_),
    .B1(_10431_),
    .C1(_10040_),
    .Y(_10432_));
 sky130_fd_sc_hd__a22oi_1 _19645_ (.A1(_12206_[0]),
    .A2(net3897),
    .B1(_10190_),
    .B2(_10423_),
    .Y(_10433_));
 sky130_fd_sc_hd__o31a_1 _19646_ (.A1(net3893),
    .A2(_10064_),
    .A3(_10300_),
    .B1(_09944_),
    .X(_10434_));
 sky130_fd_sc_hd__o21ai_0 _19647_ (.A1(net3895),
    .A2(_10433_),
    .B1(_10434_),
    .Y(_10435_));
 sky130_fd_sc_hd__nor2_1 _19648_ (.A(_12198_[0]),
    .B(net3900),
    .Y(_10436_));
 sky130_fd_sc_hd__a21oi_1 _19649_ (.A1(_12196_[0]),
    .A2(net3900),
    .B1(_10436_),
    .Y(_10437_));
 sky130_fd_sc_hd__o21ai_0 _19650_ (.A1(net3904),
    .A2(_10437_),
    .B1(_10149_),
    .Y(_10438_));
 sky130_fd_sc_hd__o21ai_0 _19651_ (.A1(_09990_),
    .A2(_10114_),
    .B1(_10328_),
    .Y(_10439_));
 sky130_fd_sc_hd__o21ai_0 _19652_ (.A1(_09998_),
    .A2(_09977_),
    .B1(net3904),
    .Y(_10440_));
 sky130_fd_sc_hd__a21oi_1 _19653_ (.A1(_09998_),
    .A2(_10270_),
    .B1(_10440_),
    .Y(_10441_));
 sky130_fd_sc_hd__o211ai_1 _19654_ (.A1(net3906),
    .A2(_10231_),
    .B1(net3890),
    .C1(_10040_),
    .Y(_10442_));
 sky130_fd_sc_hd__a211oi_1 _19655_ (.A1(_09936_),
    .A2(_10439_),
    .B1(_10441_),
    .C1(_10442_),
    .Y(_10443_));
 sky130_fd_sc_hd__a41o_1 _19656_ (.A1(_09944_),
    .A2(net3890),
    .A3(_10238_),
    .A4(_10438_),
    .B1(_10443_),
    .X(_10444_));
 sky130_fd_sc_hd__a311o_1 _19657_ (.A1(_09957_),
    .A2(_10432_),
    .A3(_10435_),
    .B1(_10444_),
    .C1(_09950_),
    .X(_10445_));
 sky130_fd_sc_hd__o21ai_1 _19658_ (.A1(net3889),
    .A2(_10427_),
    .B1(_10445_),
    .Y(_00094_));
 sky130_fd_sc_hd__o21ai_0 _19659_ (.A1(_10217_),
    .A2(_10269_),
    .B1(_09936_),
    .Y(_10446_));
 sky130_fd_sc_hd__o211ai_1 _19660_ (.A1(_09983_),
    .A2(_10225_),
    .B1(_10446_),
    .C1(_09975_),
    .Y(_10447_));
 sky130_fd_sc_hd__nor2_1 _19661_ (.A(net3901),
    .B(_10113_),
    .Y(_10448_));
 sky130_fd_sc_hd__a221o_1 _19662_ (.A1(net3901),
    .A2(_10447_),
    .B1(_10448_),
    .B2(_10421_),
    .C1(net3892),
    .X(_10449_));
 sky130_fd_sc_hd__o21ai_0 _19663_ (.A1(net3903),
    .A2(_10449_),
    .B1(_09950_),
    .Y(_10450_));
 sky130_fd_sc_hd__a211o_1 _19664_ (.A1(_12198_[0]),
    .A2(net3904),
    .B1(_09977_),
    .C1(_10069_),
    .X(_10451_));
 sky130_fd_sc_hd__o21ai_0 _19665_ (.A1(_12214_[0]),
    .A2(net3899),
    .B1(_10451_),
    .Y(_10452_));
 sky130_fd_sc_hd__nand3_1 _19666_ (.A(_12190_[0]),
    .B(_09936_),
    .C(_09972_),
    .Y(_10453_));
 sky130_fd_sc_hd__o21ai_0 _19667_ (.A1(_12200_[0]),
    .A2(_09972_),
    .B1(_10453_),
    .Y(_10454_));
 sky130_fd_sc_hd__o21ai_0 _19668_ (.A1(net3890),
    .A2(_10454_),
    .B1(net3893),
    .Y(_10455_));
 sky130_fd_sc_hd__a21oi_1 _19669_ (.A1(net3890),
    .A2(_10452_),
    .B1(_10455_),
    .Y(_10456_));
 sky130_fd_sc_hd__nor3_1 _19670_ (.A(_09936_),
    .B(_10357_),
    .C(_10216_),
    .Y(_10457_));
 sky130_fd_sc_hd__a311oi_1 _19671_ (.A1(_09936_),
    .A2(_09984_),
    .A3(_10109_),
    .B1(_10136_),
    .C1(_10457_),
    .Y(_10458_));
 sky130_fd_sc_hd__o21ai_0 _19672_ (.A1(_12193_[0]),
    .A2(_09936_),
    .B1(_10068_),
    .Y(_10459_));
 sky130_fd_sc_hd__a221oi_1 _19673_ (.A1(_10357_),
    .A2(_10080_),
    .B1(_10459_),
    .B2(net3897),
    .C1(_10137_),
    .Y(_10460_));
 sky130_fd_sc_hd__nor4_2 _19674_ (.A(_10040_),
    .B(_10456_),
    .C(_10458_),
    .D(_10460_),
    .Y(_10461_));
 sky130_fd_sc_hd__nand2_1 _19675_ (.A(_09936_),
    .B(_10152_),
    .Y(_10462_));
 sky130_fd_sc_hd__o22ai_1 _19676_ (.A1(_12188_[0]),
    .A2(_09936_),
    .B1(_10033_),
    .B2(_10462_),
    .Y(_10463_));
 sky130_fd_sc_hd__a31oi_1 _19677_ (.A1(net3676),
    .A2(_10119_),
    .A3(_10086_),
    .B1(_10156_),
    .Y(_10464_));
 sky130_fd_sc_hd__nor2_1 _19678_ (.A(net3891),
    .B(_10464_),
    .Y(_10465_));
 sky130_fd_sc_hd__a2111oi_0 _19679_ (.A1(net3891),
    .A2(_10463_),
    .B1(_09990_),
    .C1(net3903),
    .D1(_10465_),
    .Y(_10466_));
 sky130_fd_sc_hd__nor3_1 _19680_ (.A(_12198_[0]),
    .B(net3904),
    .C(net3899),
    .Y(_10467_));
 sky130_fd_sc_hd__nor2_1 _19681_ (.A(_09936_),
    .B(_10352_),
    .Y(_10468_));
 sky130_fd_sc_hd__nor2_1 _19682_ (.A(net3905),
    .B(_10004_),
    .Y(_10469_));
 sky130_fd_sc_hd__a221oi_1 _19683_ (.A1(_12202_[0]),
    .A2(_10148_),
    .B1(_10063_),
    .B2(_12189_[0]),
    .C1(_10469_),
    .Y(_10470_));
 sky130_fd_sc_hd__o32ai_1 _19684_ (.A1(_10266_),
    .A2(_10467_),
    .A3(_10468_),
    .B1(_10136_),
    .B2(_10470_),
    .Y(_10471_));
 sky130_fd_sc_hd__a32oi_1 _19685_ (.A1(net3908),
    .A2(_09936_),
    .A3(_10108_),
    .B1(_10181_),
    .B2(_10133_),
    .Y(_10472_));
 sky130_fd_sc_hd__a21oi_1 _19686_ (.A1(_10424_),
    .A2(_10472_),
    .B1(_09944_),
    .Y(_10473_));
 sky130_fd_sc_hd__a21oi_1 _19687_ (.A1(net3676),
    .A2(_10273_),
    .B1(_10217_),
    .Y(_10474_));
 sky130_fd_sc_hd__a221oi_1 _19688_ (.A1(_12188_[0]),
    .A2(_10148_),
    .B1(_10036_),
    .B2(net3905),
    .C1(_10137_),
    .Y(_10475_));
 sky130_fd_sc_hd__o21ai_0 _19689_ (.A1(net3908),
    .A2(_10474_),
    .B1(_10475_),
    .Y(_10476_));
 sky130_fd_sc_hd__nand2_1 _19690_ (.A(_10473_),
    .B(_10476_),
    .Y(_10477_));
 sky130_fd_sc_hd__o21ai_0 _19691_ (.A1(_10471_),
    .A2(_10477_),
    .B1(net3889),
    .Y(_10478_));
 sky130_fd_sc_hd__a21oi_1 _19692_ (.A1(_09929_),
    .A2(_10239_),
    .B1(_10006_),
    .Y(_10479_));
 sky130_fd_sc_hd__a21oi_1 _19693_ (.A1(_10004_),
    .A2(_10023_),
    .B1(_09923_),
    .Y(_10480_));
 sky130_fd_sc_hd__a211oi_1 _19694_ (.A1(_09923_),
    .A2(_10217_),
    .B1(_10480_),
    .C1(net3895),
    .Y(_10481_));
 sky130_fd_sc_hd__a211oi_1 _19695_ (.A1(net3906),
    .A2(_10148_),
    .B1(_10083_),
    .C1(_09998_),
    .Y(_10482_));
 sky130_fd_sc_hd__o22ai_2 _19696_ (.A1(net3908),
    .A2(_10479_),
    .B1(_10481_),
    .B2(_10482_),
    .Y(_10483_));
 sky130_fd_sc_hd__o21ai_0 _19697_ (.A1(_10036_),
    .A2(_10388_),
    .B1(_09929_),
    .Y(_10484_));
 sky130_fd_sc_hd__o31ai_1 _19698_ (.A1(_09929_),
    .A2(net3894),
    .A3(_09983_),
    .B1(_10484_),
    .Y(_10485_));
 sky130_fd_sc_hd__o2111ai_1 _19699_ (.A1(_09936_),
    .A2(_10285_),
    .B1(_10045_),
    .C1(net3890),
    .D1(_10090_),
    .Y(_10486_));
 sky130_fd_sc_hd__a21oi_2 _19700_ (.A1(_09923_),
    .A2(_10485_),
    .B1(_10486_),
    .Y(_10487_));
 sky130_fd_sc_hd__a211oi_4 _19701_ (.A1(_09957_),
    .A2(_10483_),
    .B1(_10487_),
    .C1(_10040_),
    .Y(_10488_));
 sky130_fd_sc_hd__o32ai_1 _19702_ (.A1(_10450_),
    .A2(_10461_),
    .A3(_10466_),
    .B1(_10478_),
    .B2(_10488_),
    .Y(_00095_));
 sky130_fd_sc_hd__xnor2_1 _19703_ (.A(\sa00_sr[1] ),
    .B(\sa30_sr[7] ),
    .Y(_10489_));
 sky130_fd_sc_hd__xnor2_1 _19704_ (.A(\sa10_sr[1] ),
    .B(\sa30_sr[0] ),
    .Y(_10490_));
 sky130_fd_sc_hd__xnor3_1 _19705_ (.A(\sa30_sr[1] ),
    .B(\sa20_sr[0] ),
    .C(net4207),
    .X(_10491_));
 sky130_fd_sc_hd__xnor3_1 _19706_ (.A(_10489_),
    .B(_10490_),
    .C(_10491_),
    .X(_10492_));
 sky130_fd_sc_hd__mux2i_2 _19707_ (.A0(\text_in_r[105] ),
    .A1(_10492_),
    .S(_05879_),
    .Y(_10493_));
 sky130_fd_sc_hd__xor2_4 _19708_ (.A(net4158),
    .B(_10493_),
    .X(_10494_));
 sky130_fd_sc_hd__inv_16 _19709_ (.A(net389),
    .Y(_10495_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_497 ();
 sky130_fd_sc_hd__xnor3_1 _19711_ (.A(net4220),
    .B(net4207),
    .C(net4189),
    .X(_10496_));
 sky130_fd_sc_hd__xnor2_1 _19712_ (.A(_08240_),
    .B(_10496_),
    .Y(_10497_));
 sky130_fd_sc_hd__mux2i_1 _19713_ (.A0(\text_in_r[104] ),
    .A1(_10497_),
    .S(_05879_),
    .Y(_10498_));
 sky130_fd_sc_hd__xor2_2 _19714_ (.A(\u0.w[0][8] ),
    .B(_10498_),
    .X(_10499_));
 sky130_fd_sc_hd__clkinv_16 _19715_ (.A(net3885),
    .Y(_10500_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_496 ();
 sky130_fd_sc_hd__xnor3_1 _19717_ (.A(net4219),
    .B(\sa30_sr[2] ),
    .C(\sa00_sr[2] ),
    .X(_10501_));
 sky130_fd_sc_hd__xnor2_2 _19718_ (.A(net4122),
    .B(_10501_),
    .Y(_10502_));
 sky130_fd_sc_hd__a21oi_1 _19719_ (.A1(net4230),
    .A2(\text_in_r[106] ),
    .B1(\u0.w[0][10] ),
    .Y(_10503_));
 sky130_fd_sc_hd__a21bo_4 _19720_ (.A1(net4117),
    .A2(_10502_),
    .B1_N(_10503_),
    .X(_10504_));
 sky130_fd_sc_hd__and3_4 _19721_ (.A(\u0.w[0][10] ),
    .B(net4230),
    .C(\text_in_r[106] ),
    .X(_10505_));
 sky130_fd_sc_hd__a31oi_4 _19722_ (.A1(\u0.w[0][10] ),
    .A2(net4117),
    .A3(_10502_),
    .B1(_10505_),
    .Y(_10506_));
 sky130_fd_sc_hd__and2_4 _19723_ (.A(_10504_),
    .B(_10506_),
    .X(_10507_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_495 ();
 sky130_fd_sc_hd__clkinv_16 _19725_ (.A(_10507_),
    .Y(_10509_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_487 ();
 sky130_fd_sc_hd__xnor3_1 _19734_ (.A(\sa30_sr[4] ),
    .B(\sa10_sr[5] ),
    .C(\sa00_sr[5] ),
    .X(_10515_));
 sky130_fd_sc_hd__xor2_1 _19735_ (.A(\sa20_sr[4] ),
    .B(\sa30_sr[5] ),
    .X(_10516_));
 sky130_fd_sc_hd__xnor2_1 _19736_ (.A(_10515_),
    .B(_10516_),
    .Y(_10517_));
 sky130_fd_sc_hd__mux2i_4 _19737_ (.A0(\text_in_r[109] ),
    .A1(_10517_),
    .S(_05879_),
    .Y(_10518_));
 sky130_fd_sc_hd__xnor2_4 _19738_ (.A(net4175),
    .B(_10518_),
    .Y(_10519_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_484 ();
 sky130_fd_sc_hd__xnor3_1 _19742_ (.A(\sa30_sr[5] ),
    .B(\sa10_sr[6] ),
    .C(\sa00_sr[6] ),
    .X(_10523_));
 sky130_fd_sc_hd__xnor2_1 _19743_ (.A(net4208),
    .B(\sa30_sr[6] ),
    .Y(_10524_));
 sky130_fd_sc_hd__xnor2_1 _19744_ (.A(_10523_),
    .B(_10524_),
    .Y(_10525_));
 sky130_fd_sc_hd__nor2_2 _19745_ (.A(net398),
    .B(_10525_),
    .Y(_10526_));
 sky130_fd_sc_hd__a21oi_4 _19746_ (.A1(net398),
    .A2(\text_in_r[110] ),
    .B1(_10526_),
    .Y(_10527_));
 sky130_fd_sc_hd__xor2_4 _19747_ (.A(\u0.w[0][14] ),
    .B(_10527_),
    .X(_10528_));
 sky130_fd_sc_hd__xor2_1 _19748_ (.A(net4229),
    .B(\sa30_sr[6] ),
    .X(_10529_));
 sky130_fd_sc_hd__xor2_1 _19749_ (.A(\sa20_sr[6] ),
    .B(net4189),
    .X(_10530_));
 sky130_fd_sc_hd__xnor2_1 _19750_ (.A(_10529_),
    .B(_10530_),
    .Y(_10531_));
 sky130_fd_sc_hd__xnor2_2 _19751_ (.A(net4216),
    .B(_10531_),
    .Y(_10532_));
 sky130_fd_sc_hd__mux2i_4 _19752_ (.A0(\text_in_r[111] ),
    .A1(_10532_),
    .S(net4118),
    .Y(_10533_));
 sky130_fd_sc_hd__xor2_4 _19753_ (.A(\u0.w[0][15] ),
    .B(_10533_),
    .X(_10534_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_483 ();
 sky130_fd_sc_hd__nand2_8 _19755_ (.A(_10528_),
    .B(_10534_),
    .Y(_10536_));
 sky130_fd_sc_hd__xnor2_1 _19756_ (.A(\sa00_sr[4] ),
    .B(net4189),
    .Y(_10537_));
 sky130_fd_sc_hd__xnor2_1 _19757_ (.A(\sa30_sr[3] ),
    .B(\sa10_sr[4] ),
    .Y(_10538_));
 sky130_fd_sc_hd__xnor3_1 _19758_ (.A(_08280_),
    .B(_10537_),
    .C(_10538_),
    .X(_10539_));
 sky130_fd_sc_hd__mux2i_4 _19759_ (.A0(\text_in_r[108] ),
    .A1(_10539_),
    .S(_05879_),
    .Y(_10540_));
 sky130_fd_sc_hd__xnor2_4 _19760_ (.A(net4176),
    .B(_10540_),
    .Y(_10541_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_480 ();
 sky130_fd_sc_hd__xnor2_1 _19764_ (.A(\sa00_sr[3] ),
    .B(net4189),
    .Y(_10545_));
 sky130_fd_sc_hd__xnor2_1 _19765_ (.A(\sa30_sr[2] ),
    .B(net4218),
    .Y(_10546_));
 sky130_fd_sc_hd__xnor3_1 _19766_ (.A(\sa20_sr[2] ),
    .B(\sa30_sr[3] ),
    .C(net4207),
    .X(_10547_));
 sky130_fd_sc_hd__xnor3_1 _19767_ (.A(_10545_),
    .B(_10546_),
    .C(_10547_),
    .X(_10548_));
 sky130_fd_sc_hd__mux2i_4 _19768_ (.A0(\text_in_r[107] ),
    .A1(_10548_),
    .S(net4117),
    .Y(_10549_));
 sky130_fd_sc_hd__xnor2_4 _19769_ (.A(_10549_),
    .B(\u0.w[0][11] ),
    .Y(_10550_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_479 ();
 sky130_fd_sc_hd__nor2_4 _19771_ (.A(net3883),
    .B(net390),
    .Y(_10552_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_478 ();
 sky130_fd_sc_hd__nand2_8 _19773_ (.A(_10509_),
    .B(net3879),
    .Y(_10554_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_477 ();
 sky130_fd_sc_hd__xor2_1 _19775_ (.A(net4177),
    .B(_10549_),
    .X(_10556_));
 sky130_fd_sc_hd__nand2_8 _19776_ (.A(net3883),
    .B(net3872),
    .Y(_10557_));
 sky130_fd_sc_hd__nand2_1 _19777_ (.A(_10554_),
    .B(_10557_),
    .Y(_10558_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_474 ();
 sky130_fd_sc_hd__nand2_8 _19781_ (.A(net3883),
    .B(net3879),
    .Y(_10562_));
 sky130_fd_sc_hd__nor2_4 _19782_ (.A(_12221_[0]),
    .B(_10562_),
    .Y(_10563_));
 sky130_fd_sc_hd__a221oi_2 _19783_ (.A1(_12230_[0]),
    .A2(_10552_),
    .B1(_10558_),
    .B2(_12220_[0]),
    .C1(_10563_),
    .Y(_10564_));
 sky130_fd_sc_hd__nor2_1 _19784_ (.A(_10495_),
    .B(net3883),
    .Y(_10565_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_473 ();
 sky130_fd_sc_hd__nand2_8 _19786_ (.A(_12221_[0]),
    .B(net3876),
    .Y(_10567_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_472 ();
 sky130_fd_sc_hd__nor2_2 _19788_ (.A(_10495_),
    .B(net3878),
    .Y(_10569_));
 sky130_fd_sc_hd__nand2b_4 _19789_ (.A_N(_12221_[0]),
    .B(_10509_),
    .Y(_10570_));
 sky130_fd_sc_hd__o221ai_1 _19790_ (.A1(net3611),
    .A2(_10567_),
    .B1(_10569_),
    .B2(_10570_),
    .C1(net3881),
    .Y(_10571_));
 sky130_fd_sc_hd__o21ai_0 _19791_ (.A1(net3881),
    .A2(_10564_),
    .B1(_10571_),
    .Y(_10572_));
 sky130_fd_sc_hd__nor3b_1 _19792_ (.A(net3882),
    .B(_10536_),
    .C_N(_10572_),
    .Y(_10573_));
 sky130_fd_sc_hd__xor2_4 _19793_ (.A(net4175),
    .B(_10518_),
    .X(_10574_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_468 ();
 sky130_fd_sc_hd__nor2_1 _19798_ (.A(_12220_[0]),
    .B(net3873),
    .Y(_10579_));
 sky130_fd_sc_hd__nor2_4 _19799_ (.A(_12234_[0]),
    .B(net3878),
    .Y(_10580_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_466 ();
 sky130_fd_sc_hd__a21oi_4 _19802_ (.A1(_12221_[0]),
    .A2(net3873),
    .B1(_10509_),
    .Y(_10583_));
 sky130_fd_sc_hd__o21ai_0 _19803_ (.A1(_12230_[0]),
    .A2(net3873),
    .B1(_10583_),
    .Y(_10584_));
 sky130_fd_sc_hd__xor2_4 _19804_ (.A(net4176),
    .B(_10540_),
    .X(_10585_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_463 ();
 sky130_fd_sc_hd__o311ai_0 _19808_ (.A1(net3884),
    .A2(_10579_),
    .A3(_10580_),
    .B1(_10584_),
    .C1(net3869),
    .Y(_10589_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_462 ();
 sky130_fd_sc_hd__nand2_2 _19810_ (.A(net3888),
    .B(net3886),
    .Y(_10590_));
 sky130_fd_sc_hd__nand2_8 _19811_ (.A(_10500_),
    .B(net3883),
    .Y(_10591_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_461 ();
 sky130_fd_sc_hd__nand2_1 _19813_ (.A(net3881),
    .B(net3878),
    .Y(_10593_));
 sky130_fd_sc_hd__a21o_1 _19814_ (.A1(_10590_),
    .A2(_10591_),
    .B1(_10593_),
    .X(_10594_));
 sky130_fd_sc_hd__nor2_4 _19815_ (.A(net3869),
    .B(net3878),
    .Y(_10595_));
 sky130_fd_sc_hd__nand3_1 _19816_ (.A(_10590_),
    .B(_10591_),
    .C(_10595_),
    .Y(_10596_));
 sky130_fd_sc_hd__nand3_1 _19817_ (.A(_10589_),
    .B(_10594_),
    .C(_10596_),
    .Y(_10597_));
 sky130_fd_sc_hd__nor3_1 _19818_ (.A(net3870),
    .B(_10536_),
    .C(_10597_),
    .Y(_10598_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_458 ();
 sky130_fd_sc_hd__nand2_4 _19822_ (.A(_10509_),
    .B(net3873),
    .Y(_10602_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_456 ();
 sky130_fd_sc_hd__nor3_1 _19825_ (.A(_12225_[0]),
    .B(_10509_),
    .C(net390),
    .Y(_10605_));
 sky130_fd_sc_hd__a311oi_1 _19826_ (.A1(_12222_[0]),
    .A2(net3883),
    .A3(net3879),
    .B1(_10605_),
    .C1(_10585_),
    .Y(_10606_));
 sky130_fd_sc_hd__o21ai_2 _19827_ (.A1(_12230_[0]),
    .A2(_10602_),
    .B1(_10606_),
    .Y(_10607_));
 sky130_fd_sc_hd__nor2_2 _19828_ (.A(net3595),
    .B(net3872),
    .Y(_10608_));
 sky130_fd_sc_hd__a21oi_1 _19829_ (.A1(_12222_[0]),
    .A2(net3874),
    .B1(_10608_),
    .Y(_10609_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_455 ();
 sky130_fd_sc_hd__nand3_2 _19831_ (.A(_12232_[0]),
    .B(_10509_),
    .C(net3877),
    .Y(_10611_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_453 ();
 sky130_fd_sc_hd__o211ai_1 _19834_ (.A1(net3675),
    .A2(_10609_),
    .B1(_10611_),
    .C1(net3869),
    .Y(_10614_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_451 ();
 sky130_fd_sc_hd__a221oi_1 _19837_ (.A1(_12243_[0]),
    .A2(net3878),
    .B1(_10552_),
    .B2(_12221_[0]),
    .C1(net3869),
    .Y(_10617_));
 sky130_fd_sc_hd__a21oi_4 _19838_ (.A1(_10504_),
    .A2(_10506_),
    .B1(_12227_[0]),
    .Y(_10618_));
 sky130_fd_sc_hd__a21oi_2 _19839_ (.A1(_12225_[0]),
    .A2(net3883),
    .B1(_10618_),
    .Y(_10619_));
 sky130_fd_sc_hd__a21o_4 _19840_ (.A1(net3873),
    .A2(_10619_),
    .B1(net3881),
    .X(_10620_));
 sky130_fd_sc_hd__nand2_4 _19841_ (.A(_12222_[0]),
    .B(net3874),
    .Y(_10621_));
 sky130_fd_sc_hd__nand2_4 _19842_ (.A(_10500_),
    .B(net3879),
    .Y(_10622_));
 sky130_fd_sc_hd__a21oi_1 _19843_ (.A1(_10621_),
    .A2(_10622_),
    .B1(net3883),
    .Y(_10623_));
 sky130_fd_sc_hd__nor2_2 _19844_ (.A(_12220_[0]),
    .B(_10562_),
    .Y(_10624_));
 sky130_fd_sc_hd__nor3_1 _19845_ (.A(_10620_),
    .B(_10623_),
    .C(_10624_),
    .Y(_10625_));
 sky130_fd_sc_hd__xnor2_4 _19846_ (.A(net4174),
    .B(_10527_),
    .Y(_10626_));
 sky130_fd_sc_hd__nor2_1 _19847_ (.A(_10626_),
    .B(_10534_),
    .Y(_10627_));
 sky130_fd_sc_hd__o31ai_1 _19848_ (.A1(net3882),
    .A2(_10617_),
    .A3(_10625_),
    .B1(_10627_),
    .Y(_10628_));
 sky130_fd_sc_hd__a31oi_1 _19849_ (.A1(net3882),
    .A2(_10607_),
    .A3(_10614_),
    .B1(_10628_),
    .Y(_10629_));
 sky130_fd_sc_hd__nor2_4 _19850_ (.A(net3886),
    .B(net3883),
    .Y(_10630_));
 sky130_fd_sc_hd__nor2_1 _19851_ (.A(_12234_[0]),
    .B(_10509_),
    .Y(_10631_));
 sky130_fd_sc_hd__o21ai_4 _19852_ (.A1(_10630_),
    .A2(_10631_),
    .B1(net3878),
    .Y(_10632_));
 sky130_fd_sc_hd__nor2_2 _19853_ (.A(_10509_),
    .B(net3878),
    .Y(_10633_));
 sky130_fd_sc_hd__and2_4 _19854_ (.A(_12221_[0]),
    .B(net3878),
    .X(_10634_));
 sky130_fd_sc_hd__a211oi_1 _19855_ (.A1(_12232_[0]),
    .A2(_10633_),
    .B1(_10634_),
    .C1(net3869),
    .Y(_10635_));
 sky130_fd_sc_hd__a21oi_1 _19856_ (.A1(net3869),
    .A2(_10632_),
    .B1(_10635_),
    .Y(_10636_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_450 ();
 sky130_fd_sc_hd__nand2_8 _19858_ (.A(net401),
    .B(net3872),
    .Y(_10638_));
 sky130_fd_sc_hd__a21oi_1 _19859_ (.A1(_10593_),
    .A2(_10638_),
    .B1(net3883),
    .Y(_10639_));
 sky130_fd_sc_hd__nor3_1 _19860_ (.A(net3882),
    .B(_10636_),
    .C(_10639_),
    .Y(_10640_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_449 ();
 sky130_fd_sc_hd__nand2_1 _19862_ (.A(_12220_[0]),
    .B(_10552_),
    .Y(_10642_));
 sky130_fd_sc_hd__nor2_4 _19863_ (.A(_12227_[0]),
    .B(net3873),
    .Y(_10643_));
 sky130_fd_sc_hd__nor2_4 _19864_ (.A(_12222_[0]),
    .B(net3879),
    .Y(_10644_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_448 ();
 sky130_fd_sc_hd__o21ai_0 _19866_ (.A1(_10643_),
    .A2(_10644_),
    .B1(net3884),
    .Y(_10646_));
 sky130_fd_sc_hd__nor2_4 _19867_ (.A(net3886),
    .B(net3872),
    .Y(_10647_));
 sky130_fd_sc_hd__o21ai_1 _19868_ (.A1(_10495_),
    .A2(net3879),
    .B1(net3883),
    .Y(_10648_));
 sky130_fd_sc_hd__o21ai_1 _19869_ (.A1(_12221_[0]),
    .A2(net3879),
    .B1(_10509_),
    .Y(_10649_));
 sky130_fd_sc_hd__nor2_2 _19870_ (.A(_12230_[0]),
    .B(net3873),
    .Y(_10650_));
 sky130_fd_sc_hd__o22ai_1 _19871_ (.A1(_10647_),
    .A2(_10648_),
    .B1(_10649_),
    .B2(_10650_),
    .Y(_10651_));
 sky130_fd_sc_hd__nor2_1 _19872_ (.A(net3881),
    .B(_10651_),
    .Y(_10652_));
 sky130_fd_sc_hd__a311oi_2 _19873_ (.A1(net3881),
    .A2(_10642_),
    .A3(_10646_),
    .B1(_10652_),
    .C1(net3870),
    .Y(_10653_));
 sky130_fd_sc_hd__nor2_1 _19874_ (.A(net3883),
    .B(_10585_),
    .Y(_10654_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_447 ();
 sky130_fd_sc_hd__nor2_1 _19876_ (.A(_12225_[0]),
    .B(net3877),
    .Y(_10656_));
 sky130_fd_sc_hd__nor2_1 _19877_ (.A(_10647_),
    .B(_10656_),
    .Y(_10657_));
 sky130_fd_sc_hd__nand2_1 _19878_ (.A(_10654_),
    .B(_10657_),
    .Y(_10658_));
 sky130_fd_sc_hd__nor2_1 _19879_ (.A(_12222_[0]),
    .B(_10509_),
    .Y(_10659_));
 sky130_fd_sc_hd__nand2_4 _19880_ (.A(_10495_),
    .B(_10509_),
    .Y(_10660_));
 sky130_fd_sc_hd__nand3b_1 _19881_ (.A_N(_10659_),
    .B(_10660_),
    .C(net3873),
    .Y(_10661_));
 sky130_fd_sc_hd__nor2_4 _19882_ (.A(net3888),
    .B(net3879),
    .Y(_10662_));
 sky130_fd_sc_hd__nand2_1 _19883_ (.A(_12236_[0]),
    .B(net3878),
    .Y(_10663_));
 sky130_fd_sc_hd__nor2_4 _19884_ (.A(_10509_),
    .B(_10585_),
    .Y(_10664_));
 sky130_fd_sc_hd__and3b_1 _19885_ (.A_N(_10662_),
    .B(_10663_),
    .C(_10664_),
    .X(_10665_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_446 ();
 sky130_fd_sc_hd__nand2_1 _19887_ (.A(net3870),
    .B(_10534_),
    .Y(_10667_));
 sky130_fd_sc_hd__a311oi_1 _19888_ (.A1(net3869),
    .A2(_10632_),
    .A3(_10661_),
    .B1(_10665_),
    .C1(_10667_),
    .Y(_10668_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_445 ();
 sky130_fd_sc_hd__a21oi_2 _19890_ (.A1(_10658_),
    .A2(_10668_),
    .B1(net3674),
    .Y(_10670_));
 sky130_fd_sc_hd__nor2_4 _19891_ (.A(net3886),
    .B(net3878),
    .Y(_10671_));
 sky130_fd_sc_hd__o32ai_1 _19892_ (.A1(net3883),
    .A2(_10608_),
    .A3(_10671_),
    .B1(_10562_),
    .B2(net402),
    .Y(_10672_));
 sky130_fd_sc_hd__nor2_1 _19893_ (.A(net3881),
    .B(_10672_),
    .Y(_10673_));
 sky130_fd_sc_hd__o21ai_1 _19894_ (.A1(_10634_),
    .A2(_10671_),
    .B1(net3883),
    .Y(_10674_));
 sky130_fd_sc_hd__nor2_1 _19895_ (.A(_12225_[0]),
    .B(net3883),
    .Y(_10675_));
 sky130_fd_sc_hd__nand2_2 _19896_ (.A(net3875),
    .B(_10675_),
    .Y(_10676_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_444 ();
 sky130_fd_sc_hd__nor2_4 _19898_ (.A(net3883),
    .B(net3871),
    .Y(_10678_));
 sky130_fd_sc_hd__nand2_4 _19899_ (.A(_12236_[0]),
    .B(_10678_),
    .Y(_10679_));
 sky130_fd_sc_hd__a31oi_1 _19900_ (.A1(_10674_),
    .A2(_10676_),
    .A3(_10679_),
    .B1(net3869),
    .Y(_10680_));
 sky130_fd_sc_hd__o211ai_1 _19901_ (.A1(_10673_),
    .A2(_10680_),
    .B1(net3882),
    .C1(_10534_),
    .Y(_10681_));
 sky130_fd_sc_hd__o311a_1 _19902_ (.A1(_10534_),
    .A2(_10640_),
    .A3(_10653_),
    .B1(_10670_),
    .C1(_10681_),
    .X(_10682_));
 sky130_fd_sc_hd__nor4_4 _19903_ (.A(_10573_),
    .B(_10598_),
    .C(_10629_),
    .D(_10682_),
    .Y(_00096_));
 sky130_fd_sc_hd__xnor2_4 _19904_ (.A(\u0.w[0][15] ),
    .B(_10533_),
    .Y(_10683_));
 sky130_fd_sc_hd__nand2_4 _19905_ (.A(net3674),
    .B(_10683_),
    .Y(_10684_));
 sky130_fd_sc_hd__nor2_2 _19906_ (.A(net3888),
    .B(_10509_),
    .Y(_10685_));
 sky130_fd_sc_hd__nor3_1 _19907_ (.A(_10550_),
    .B(_10618_),
    .C(_10685_),
    .Y(_10686_));
 sky130_fd_sc_hd__o21ai_1 _19908_ (.A1(_12250_[0]),
    .A2(net3875),
    .B1(net3881),
    .Y(_10687_));
 sky130_fd_sc_hd__nand2_1 _19909_ (.A(_12221_[0]),
    .B(_10509_),
    .Y(_10688_));
 sky130_fd_sc_hd__nand2_1 _19910_ (.A(_12236_[0]),
    .B(net3883),
    .Y(_10689_));
 sky130_fd_sc_hd__a21oi_1 _19911_ (.A1(_10688_),
    .A2(_10689_),
    .B1(net3873),
    .Y(_10690_));
 sky130_fd_sc_hd__o22ai_1 _19912_ (.A1(_10686_),
    .A2(_10687_),
    .B1(_10690_),
    .B2(_10620_),
    .Y(_10691_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_443 ();
 sky130_fd_sc_hd__o21ai_0 _19914_ (.A1(_10608_),
    .A2(_10662_),
    .B1(net3675),
    .Y(_10693_));
 sky130_fd_sc_hd__nand2_8 _19915_ (.A(_10519_),
    .B(_10585_),
    .Y(_10694_));
 sky130_fd_sc_hd__a21oi_1 _19916_ (.A1(net3888),
    .A2(_10671_),
    .B1(_10694_),
    .Y(_10695_));
 sky130_fd_sc_hd__nand2_4 _19917_ (.A(_12221_[0]),
    .B(net3877),
    .Y(_10696_));
 sky130_fd_sc_hd__a32oi_1 _19918_ (.A1(net3883),
    .A2(_10696_),
    .A3(_10638_),
    .B1(_10630_),
    .B2(net3872),
    .Y(_10697_));
 sky130_fd_sc_hd__o21ai_0 _19919_ (.A1(_10500_),
    .A2(_10554_),
    .B1(_10697_),
    .Y(_10698_));
 sky130_fd_sc_hd__nor2_4 _19920_ (.A(net3870),
    .B(net3869),
    .Y(_10699_));
 sky130_fd_sc_hd__a222oi_1 _19921_ (.A1(net3870),
    .A2(_10691_),
    .B1(_10693_),
    .B2(_10695_),
    .C1(_10698_),
    .C2(_10699_),
    .Y(_10700_));
 sky130_fd_sc_hd__nand2_8 _19922_ (.A(_10500_),
    .B(net3871),
    .Y(_10701_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_442 ();
 sky130_fd_sc_hd__a21oi_1 _19924_ (.A1(_10696_),
    .A2(_10701_),
    .B1(net3883),
    .Y(_10703_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_441 ();
 sky130_fd_sc_hd__a211oi_1 _19926_ (.A1(_12220_[0]),
    .A2(net3877),
    .B1(_10644_),
    .C1(_10509_),
    .Y(_10705_));
 sky130_fd_sc_hd__o21ai_0 _19927_ (.A1(_10703_),
    .A2(_10705_),
    .B1(_10699_),
    .Y(_10706_));
 sky130_fd_sc_hd__nor2_4 _19928_ (.A(net3882),
    .B(net3869),
    .Y(_10707_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_440 ();
 sky130_fd_sc_hd__nand2_2 _19930_ (.A(_12234_[0]),
    .B(net3879),
    .Y(_10709_));
 sky130_fd_sc_hd__o22a_4 _19931_ (.A1(_12222_[0]),
    .A2(_10602_),
    .B1(_10709_),
    .B2(net3884),
    .X(_10710_));
 sky130_fd_sc_hd__nand2b_4 _19932_ (.A_N(_12221_[0]),
    .B(net3878),
    .Y(_10711_));
 sky130_fd_sc_hd__nand2_4 _19933_ (.A(_12236_[0]),
    .B(net3872),
    .Y(_10712_));
 sky130_fd_sc_hd__nand3_1 _19934_ (.A(net3883),
    .B(_10711_),
    .C(_10712_),
    .Y(_10713_));
 sky130_fd_sc_hd__nand3_1 _19935_ (.A(_10707_),
    .B(_10710_),
    .C(_10713_),
    .Y(_10714_));
 sky130_fd_sc_hd__nor2_1 _19936_ (.A(_10519_),
    .B(net3881),
    .Y(_10715_));
 sky130_fd_sc_hd__and2_4 _19937_ (.A(_12234_[0]),
    .B(net3873),
    .X(_10716_));
 sky130_fd_sc_hd__nor2_4 _19938_ (.A(_12221_[0]),
    .B(net3873),
    .Y(_10717_));
 sky130_fd_sc_hd__o21ai_0 _19939_ (.A1(_10716_),
    .A2(_10717_),
    .B1(net3884),
    .Y(_10718_));
 sky130_fd_sc_hd__nand2_2 _19940_ (.A(net3885),
    .B(_10552_),
    .Y(_10719_));
 sky130_fd_sc_hd__nand2_8 _19941_ (.A(_10626_),
    .B(_10534_),
    .Y(_10720_));
 sky130_fd_sc_hd__a31oi_1 _19942_ (.A1(_10715_),
    .A2(_10718_),
    .A3(_10719_),
    .B1(_10720_),
    .Y(_10721_));
 sky130_fd_sc_hd__nor2_4 _19943_ (.A(net3888),
    .B(net3872),
    .Y(_10722_));
 sky130_fd_sc_hd__nor2_4 _19944_ (.A(_12220_[0]),
    .B(net3878),
    .Y(_10723_));
 sky130_fd_sc_hd__nor2_4 _19945_ (.A(_10574_),
    .B(net3881),
    .Y(_10724_));
 sky130_fd_sc_hd__o21ai_0 _19946_ (.A1(_10643_),
    .A2(_10671_),
    .B1(net3883),
    .Y(_10725_));
 sky130_fd_sc_hd__o311ai_0 _19947_ (.A1(net3883),
    .A2(_10722_),
    .A3(_10723_),
    .B1(_10724_),
    .C1(_10725_),
    .Y(_10726_));
 sky130_fd_sc_hd__nand4_1 _19948_ (.A(_10706_),
    .B(_10714_),
    .C(_10721_),
    .D(_10726_),
    .Y(_10727_));
 sky130_fd_sc_hd__o21ai_0 _19949_ (.A1(_10684_),
    .A2(_10700_),
    .B1(_10727_),
    .Y(_10728_));
 sky130_fd_sc_hd__nor2_1 _19950_ (.A(_12234_[0]),
    .B(_10554_),
    .Y(_10729_));
 sky130_fd_sc_hd__a21oi_1 _19951_ (.A1(_10638_),
    .A2(_10711_),
    .B1(net3675),
    .Y(_10730_));
 sky130_fd_sc_hd__o21ai_0 _19952_ (.A1(_10729_),
    .A2(_10730_),
    .B1(net3882),
    .Y(_10731_));
 sky130_fd_sc_hd__nor2_4 _19953_ (.A(_10678_),
    .B(_10633_),
    .Y(_10732_));
 sky130_fd_sc_hd__a22oi_1 _19954_ (.A1(_12221_[0]),
    .A2(_10552_),
    .B1(_10647_),
    .B2(net3888),
    .Y(_10733_));
 sky130_fd_sc_hd__o211ai_1 _19955_ (.A1(_10500_),
    .A2(_10732_),
    .B1(_10733_),
    .C1(net3870),
    .Y(_10734_));
 sky130_fd_sc_hd__nand3_1 _19956_ (.A(net3869),
    .B(_10731_),
    .C(_10734_),
    .Y(_10735_));
 sky130_fd_sc_hd__o21ai_0 _19957_ (.A1(_10580_),
    .A2(_10722_),
    .B1(net3884),
    .Y(_10736_));
 sky130_fd_sc_hd__and3_1 _19958_ (.A(net3882),
    .B(_10679_),
    .C(_10736_),
    .X(_10737_));
 sky130_fd_sc_hd__nor2_1 _19959_ (.A(_10500_),
    .B(net3878),
    .Y(_10738_));
 sky130_fd_sc_hd__o21ai_0 _19960_ (.A1(_10717_),
    .A2(_10723_),
    .B1(net3884),
    .Y(_10739_));
 sky130_fd_sc_hd__o311a_1 _19961_ (.A1(net3884),
    .A2(_10643_),
    .A3(_10738_),
    .B1(_10739_),
    .C1(net3870),
    .X(_10740_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_439 ();
 sky130_fd_sc_hd__o21ai_2 _19963_ (.A1(_10737_),
    .A2(_10740_),
    .B1(net3881),
    .Y(_10742_));
 sky130_fd_sc_hd__nand2_8 _19964_ (.A(_10626_),
    .B(_10683_),
    .Y(_10743_));
 sky130_fd_sc_hd__a21oi_2 _19965_ (.A1(_10735_),
    .A2(_10742_),
    .B1(_10743_),
    .Y(_10744_));
 sky130_fd_sc_hd__nor2_1 _19966_ (.A(_12234_[0]),
    .B(net3874),
    .Y(_10745_));
 sky130_fd_sc_hd__nor3_1 _19967_ (.A(net3675),
    .B(_10671_),
    .C(_10745_),
    .Y(_10746_));
 sky130_fd_sc_hd__nor3_1 _19968_ (.A(net3883),
    .B(_10608_),
    .C(_10723_),
    .Y(_10747_));
 sky130_fd_sc_hd__o21ai_0 _19969_ (.A1(_10746_),
    .A2(_10747_),
    .B1(_10699_),
    .Y(_10748_));
 sky130_fd_sc_hd__nor2_4 _19970_ (.A(_10495_),
    .B(net3871),
    .Y(_10749_));
 sky130_fd_sc_hd__o21ai_2 _19971_ (.A1(_10662_),
    .A2(_10749_),
    .B1(net3675),
    .Y(_10750_));
 sky130_fd_sc_hd__nand2_1 _19972_ (.A(_10725_),
    .B(_10750_),
    .Y(_10751_));
 sky130_fd_sc_hd__nand2_1 _19973_ (.A(_10707_),
    .B(_10751_),
    .Y(_10752_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_438 ();
 sky130_fd_sc_hd__mux2i_1 _19975_ (.A0(_12230_[0]),
    .A1(_12234_[0]),
    .S(net3883),
    .Y(_10754_));
 sky130_fd_sc_hd__nand2_2 _19976_ (.A(net3873),
    .B(_10754_),
    .Y(_10755_));
 sky130_fd_sc_hd__o311ai_0 _19977_ (.A1(_12246_[0]),
    .A2(net3882),
    .A3(net3874),
    .B1(_10755_),
    .C1(net3869),
    .Y(_10756_));
 sky130_fd_sc_hd__a31oi_1 _19978_ (.A1(_10748_),
    .A2(_10752_),
    .A3(_10756_),
    .B1(_10536_),
    .Y(_10757_));
 sky130_fd_sc_hd__nor3_2 _19979_ (.A(_10728_),
    .B(_10744_),
    .C(_10757_),
    .Y(_00097_));
 sky130_fd_sc_hd__nor3_2 _19980_ (.A(_12222_[0]),
    .B(_12227_[0]),
    .C(net3873),
    .Y(_10758_));
 sky130_fd_sc_hd__a222oi_1 _19981_ (.A1(_12230_[0]),
    .A2(_10552_),
    .B1(_10558_),
    .B2(_12234_[0]),
    .C1(_10758_),
    .C2(net3884),
    .Y(_10759_));
 sky130_fd_sc_hd__nor2_2 _19982_ (.A(net3870),
    .B(_10759_),
    .Y(_10760_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_437 ();
 sky130_fd_sc_hd__nand2_4 _19984_ (.A(_10495_),
    .B(net3883),
    .Y(_10762_));
 sky130_fd_sc_hd__a21oi_1 _19985_ (.A1(net3595),
    .A2(net3675),
    .B1(net3874),
    .Y(_10763_));
 sky130_fd_sc_hd__a221oi_1 _19986_ (.A1(_12252_[0]),
    .A2(net3874),
    .B1(_10762_),
    .B2(_10763_),
    .C1(net3882),
    .Y(_10764_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_436 ();
 sky130_fd_sc_hd__a22oi_1 _19988_ (.A1(_12241_[0]),
    .A2(net3878),
    .B1(_10552_),
    .B2(net3595),
    .Y(_10766_));
 sky130_fd_sc_hd__and2_4 _19989_ (.A(_12220_[0]),
    .B(net3872),
    .X(_10767_));
 sky130_fd_sc_hd__nand2_1 _19990_ (.A(net402),
    .B(_10678_),
    .Y(_10768_));
 sky130_fd_sc_hd__o311ai_0 _19991_ (.A1(net3675),
    .A2(_10717_),
    .A3(_10767_),
    .B1(_10768_),
    .C1(net3882),
    .Y(_10769_));
 sky130_fd_sc_hd__o2111ai_1 _19992_ (.A1(net3882),
    .A2(_10766_),
    .B1(_10769_),
    .C1(_10528_),
    .D1(net3869),
    .Y(_10770_));
 sky130_fd_sc_hd__o41ai_1 _19993_ (.A1(_10626_),
    .A2(net3869),
    .A3(_10760_),
    .A4(_10764_),
    .B1(_10770_),
    .Y(_10771_));
 sky130_fd_sc_hd__o21ai_0 _19994_ (.A1(net3611),
    .A2(_10662_),
    .B1(_12221_[0]),
    .Y(_10772_));
 sky130_fd_sc_hd__a22oi_1 _19995_ (.A1(_10622_),
    .A2(_10685_),
    .B1(_10749_),
    .B2(_10591_),
    .Y(_10773_));
 sky130_fd_sc_hd__nand2_4 _19996_ (.A(_10519_),
    .B(net3881),
    .Y(_10774_));
 sky130_fd_sc_hd__a21oi_2 _19997_ (.A1(_10772_),
    .A2(_10773_),
    .B1(_10774_),
    .Y(_10775_));
 sky130_fd_sc_hd__a211oi_1 _19998_ (.A1(_10590_),
    .A2(_10762_),
    .B1(net3882),
    .C1(net3874),
    .Y(_10776_));
 sky130_fd_sc_hd__a31oi_1 _19999_ (.A1(_12246_[0]),
    .A2(net3870),
    .A3(net3874),
    .B1(_10776_),
    .Y(_10777_));
 sky130_fd_sc_hd__nand2_1 _20000_ (.A(_12243_[0]),
    .B(net3874),
    .Y(_10778_));
 sky130_fd_sc_hd__nand2_1 _20001_ (.A(net3595),
    .B(net3883),
    .Y(_10779_));
 sky130_fd_sc_hd__nand3_1 _20002_ (.A(net3878),
    .B(_10570_),
    .C(_10779_),
    .Y(_10780_));
 sky130_fd_sc_hd__nand3_1 _20003_ (.A(net3882),
    .B(_10778_),
    .C(_10780_),
    .Y(_10781_));
 sky130_fd_sc_hd__a21oi_1 _20004_ (.A1(_10777_),
    .A2(_10781_),
    .B1(net3881),
    .Y(_10782_));
 sky130_fd_sc_hd__and2_4 _20005_ (.A(_12230_[0]),
    .B(net3878),
    .X(_10783_));
 sky130_fd_sc_hd__o21ai_0 _20006_ (.A1(_10634_),
    .A2(_10723_),
    .B1(net3675),
    .Y(_10784_));
 sky130_fd_sc_hd__o311a_1 _20007_ (.A1(net3675),
    .A2(_10569_),
    .A3(_10783_),
    .B1(_10784_),
    .C1(_10707_),
    .X(_10785_));
 sky130_fd_sc_hd__nor4_1 _20008_ (.A(_10528_),
    .B(_10775_),
    .C(_10782_),
    .D(_10785_),
    .Y(_10786_));
 sky130_fd_sc_hd__nand2_1 _20009_ (.A(_12225_[0]),
    .B(net3873),
    .Y(_10787_));
 sky130_fd_sc_hd__a21oi_1 _20010_ (.A1(_10787_),
    .A2(_10709_),
    .B1(net3884),
    .Y(_10788_));
 sky130_fd_sc_hd__nor2_1 _20011_ (.A(_12236_[0]),
    .B(_10562_),
    .Y(_10789_));
 sky130_fd_sc_hd__nor3_1 _20012_ (.A(_10694_),
    .B(_10788_),
    .C(_10789_),
    .Y(_10790_));
 sky130_fd_sc_hd__nor2_1 _20013_ (.A(_10536_),
    .B(_10790_),
    .Y(_10791_));
 sky130_fd_sc_hd__nor2_1 _20014_ (.A(_12222_[0]),
    .B(net3873),
    .Y(_10792_));
 sky130_fd_sc_hd__and2_4 _20015_ (.A(_12221_[0]),
    .B(net3873),
    .X(_10793_));
 sky130_fd_sc_hd__o21ai_2 _20016_ (.A1(_10793_),
    .A2(_10647_),
    .B1(net3883),
    .Y(_10794_));
 sky130_fd_sc_hd__o31ai_1 _20017_ (.A1(net3884),
    .A2(_10792_),
    .A3(_10662_),
    .B1(_10794_),
    .Y(_10795_));
 sky130_fd_sc_hd__nand2_1 _20018_ (.A(_10699_),
    .B(_10795_),
    .Y(_10796_));
 sky130_fd_sc_hd__nand2b_4 _20019_ (.A_N(net3595),
    .B(net3878),
    .Y(_10797_));
 sky130_fd_sc_hd__a211oi_1 _20020_ (.A1(net402),
    .A2(net3872),
    .B1(_10749_),
    .C1(_10509_),
    .Y(_10798_));
 sky130_fd_sc_hd__a31oi_1 _20021_ (.A1(_10509_),
    .A2(_10797_),
    .A3(_10712_),
    .B1(_10798_),
    .Y(_10799_));
 sky130_fd_sc_hd__o21ai_2 _20022_ (.A1(net3873),
    .A2(_10619_),
    .B1(net3869),
    .Y(_10800_));
 sky130_fd_sc_hd__a311oi_1 _20023_ (.A1(net3873),
    .A2(_10762_),
    .A3(_10688_),
    .B1(_10800_),
    .C1(net3882),
    .Y(_10801_));
 sky130_fd_sc_hd__a21oi_1 _20024_ (.A1(_10707_),
    .A2(_10799_),
    .B1(_10801_),
    .Y(_10802_));
 sky130_fd_sc_hd__nand3_1 _20025_ (.A(_10791_),
    .B(_10796_),
    .C(_10802_),
    .Y(_10803_));
 sky130_fd_sc_hd__a21oi_1 _20026_ (.A1(_12232_[0]),
    .A2(net3872),
    .B1(_10717_),
    .Y(_10804_));
 sky130_fd_sc_hd__o21ai_0 _20027_ (.A1(net3883),
    .A2(_10804_),
    .B1(_10674_),
    .Y(_10805_));
 sky130_fd_sc_hd__nand2_2 _20028_ (.A(_10495_),
    .B(net3877),
    .Y(_10806_));
 sky130_fd_sc_hd__nand2_2 _20029_ (.A(_12232_[0]),
    .B(net3872),
    .Y(_10807_));
 sky130_fd_sc_hd__a311oi_1 _20030_ (.A1(net3883),
    .A2(_10806_),
    .A3(_10807_),
    .B1(net3882),
    .C1(_10618_),
    .Y(_10808_));
 sky130_fd_sc_hd__a211oi_1 _20031_ (.A1(net3882),
    .A2(_10805_),
    .B1(_10808_),
    .C1(net3881),
    .Y(_10809_));
 sky130_fd_sc_hd__nand2_4 _20032_ (.A(_12232_[0]),
    .B(net3878),
    .Y(_10810_));
 sky130_fd_sc_hd__a21oi_1 _20033_ (.A1(_10701_),
    .A2(_10810_),
    .B1(_10509_),
    .Y(_10811_));
 sky130_fd_sc_hd__o21ai_4 _20034_ (.A1(_12236_[0]),
    .A2(net3878),
    .B1(_10509_),
    .Y(_10812_));
 sky130_fd_sc_hd__o21ai_0 _20035_ (.A1(_10722_),
    .A2(_10812_),
    .B1(_10699_),
    .Y(_10813_));
 sky130_fd_sc_hd__a21oi_1 _20036_ (.A1(_10622_),
    .A2(_10807_),
    .B1(_10509_),
    .Y(_10814_));
 sky130_fd_sc_hd__o21ai_0 _20037_ (.A1(_10643_),
    .A2(_10812_),
    .B1(_10707_),
    .Y(_10815_));
 sky130_fd_sc_hd__o22ai_1 _20038_ (.A1(_10811_),
    .A2(_10813_),
    .B1(_10814_),
    .B2(_10815_),
    .Y(_10816_));
 sky130_fd_sc_hd__o21bai_1 _20039_ (.A1(_10809_),
    .A2(_10816_),
    .B1_N(_10720_),
    .Y(_10817_));
 sky130_fd_sc_hd__o311a_4 _20040_ (.A1(net3673),
    .A2(_10771_),
    .A3(_10786_),
    .B1(_10803_),
    .C1(_10817_),
    .X(_00098_));
 sky130_fd_sc_hd__a21oi_1 _20041_ (.A1(_12221_[0]),
    .A2(net3882),
    .B1(_10509_),
    .Y(_10818_));
 sky130_fd_sc_hd__o21ai_0 _20042_ (.A1(net3888),
    .A2(net3882),
    .B1(_10818_),
    .Y(_10819_));
 sky130_fd_sc_hd__o311ai_0 _20043_ (.A1(_12230_[0]),
    .A2(net3883),
    .A3(net3882),
    .B1(_10595_),
    .C1(_10819_),
    .Y(_10820_));
 sky130_fd_sc_hd__nand2_2 _20044_ (.A(net3870),
    .B(_10585_),
    .Y(_10821_));
 sky130_fd_sc_hd__nor2_2 _20045_ (.A(net3883),
    .B(_10701_),
    .Y(_10822_));
 sky130_fd_sc_hd__nor2_1 _20046_ (.A(_10821_),
    .B(_10822_),
    .Y(_10823_));
 sky130_fd_sc_hd__nor2_1 _20047_ (.A(_12222_[0]),
    .B(_12227_[0]),
    .Y(_10824_));
 sky130_fd_sc_hd__nor2_1 _20048_ (.A(net3873),
    .B(_10824_),
    .Y(_10825_));
 sky130_fd_sc_hd__o21ai_0 _20049_ (.A1(_10793_),
    .A2(_10825_),
    .B1(net3883),
    .Y(_10826_));
 sky130_fd_sc_hd__nand3_1 _20050_ (.A(_10679_),
    .B(_10823_),
    .C(_10826_),
    .Y(_10827_));
 sky130_fd_sc_hd__nor2_1 _20051_ (.A(_10585_),
    .B(net3875),
    .Y(_10828_));
 sky130_fd_sc_hd__o21ai_0 _20052_ (.A1(_12221_[0]),
    .A2(net3882),
    .B1(_10509_),
    .Y(_10829_));
 sky130_fd_sc_hd__o21ai_0 _20053_ (.A1(_12222_[0]),
    .A2(_10509_),
    .B1(_10829_),
    .Y(_10830_));
 sky130_fd_sc_hd__nor2_2 _20054_ (.A(net3885),
    .B(_10509_),
    .Y(_10831_));
 sky130_fd_sc_hd__a221oi_1 _20055_ (.A1(_12232_[0]),
    .A2(_10732_),
    .B1(_10831_),
    .B2(net3876),
    .C1(_10694_),
    .Y(_10832_));
 sky130_fd_sc_hd__a21oi_1 _20056_ (.A1(_10828_),
    .A2(_10830_),
    .B1(_10832_),
    .Y(_10833_));
 sky130_fd_sc_hd__nand4_1 _20057_ (.A(_10528_),
    .B(_10820_),
    .C(_10827_),
    .D(_10833_),
    .Y(_10834_));
 sky130_fd_sc_hd__nand2_1 _20058_ (.A(_10583_),
    .B(_10810_),
    .Y(_10835_));
 sky130_fd_sc_hd__nor2_1 _20059_ (.A(_12236_[0]),
    .B(net3879),
    .Y(_10836_));
 sky130_fd_sc_hd__o21ai_0 _20060_ (.A1(_10647_),
    .A2(_10836_),
    .B1(_10509_),
    .Y(_10837_));
 sky130_fd_sc_hd__nand2_1 _20061_ (.A(_10835_),
    .B(_10837_),
    .Y(_10838_));
 sky130_fd_sc_hd__nand2_1 _20062_ (.A(_10699_),
    .B(_10838_),
    .Y(_10839_));
 sky130_fd_sc_hd__nand2_2 _20063_ (.A(_12236_[0]),
    .B(_10509_),
    .Y(_10840_));
 sky130_fd_sc_hd__a41oi_1 _20064_ (.A1(net3870),
    .A2(_10591_),
    .A3(_10595_),
    .A4(_10840_),
    .B1(_10528_),
    .Y(_10841_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_435 ();
 sky130_fd_sc_hd__nand2_2 _20066_ (.A(_12232_[0]),
    .B(_10509_),
    .Y(_10843_));
 sky130_fd_sc_hd__o21ai_0 _20067_ (.A1(_10509_),
    .A2(_10824_),
    .B1(_10843_),
    .Y(_10844_));
 sky130_fd_sc_hd__a21oi_1 _20068_ (.A1(net3879),
    .A2(_10844_),
    .B1(_10821_),
    .Y(_10845_));
 sky130_fd_sc_hd__nor2_1 _20069_ (.A(net3888),
    .B(_10602_),
    .Y(_10846_));
 sky130_fd_sc_hd__a2111oi_0 _20070_ (.A1(_10500_),
    .A2(_10648_),
    .B1(_10694_),
    .C1(_10846_),
    .D1(_10624_),
    .Y(_10847_));
 sky130_fd_sc_hd__a21oi_1 _20071_ (.A1(_10755_),
    .A2(_10845_),
    .B1(_10847_),
    .Y(_10848_));
 sky130_fd_sc_hd__a31oi_2 _20072_ (.A1(_10839_),
    .A2(_10841_),
    .A3(_10848_),
    .B1(_10683_),
    .Y(_10849_));
 sky130_fd_sc_hd__nor2_1 _20073_ (.A(_10500_),
    .B(_10541_),
    .Y(_10850_));
 sky130_fd_sc_hd__o32ai_1 _20074_ (.A1(_10495_),
    .A2(_10541_),
    .A3(_10831_),
    .B1(_10660_),
    .B2(_10850_),
    .Y(_10851_));
 sky130_fd_sc_hd__nor3_1 _20075_ (.A(_12221_[0]),
    .B(_10509_),
    .C(_10541_),
    .Y(_10852_));
 sky130_fd_sc_hd__nor3_1 _20076_ (.A(_12221_[0]),
    .B(net3883),
    .C(_10585_),
    .Y(_10853_));
 sky130_fd_sc_hd__a2111oi_0 _20077_ (.A1(_10585_),
    .A2(_10565_),
    .B1(_10852_),
    .C1(_10853_),
    .D1(net3876),
    .Y(_10854_));
 sky130_fd_sc_hd__a221oi_1 _20078_ (.A1(_10500_),
    .A2(_10664_),
    .B1(_10851_),
    .B2(net3876),
    .C1(_10854_),
    .Y(_10855_));
 sky130_fd_sc_hd__nand2_1 _20079_ (.A(_12225_[0]),
    .B(_10678_),
    .Y(_10856_));
 sky130_fd_sc_hd__nor2_1 _20080_ (.A(net3888),
    .B(_10500_),
    .Y(_10857_));
 sky130_fd_sc_hd__o21ai_0 _20081_ (.A1(_10831_),
    .A2(_10857_),
    .B1(net3876),
    .Y(_10858_));
 sky130_fd_sc_hd__a211oi_1 _20082_ (.A1(_10856_),
    .A2(_10858_),
    .B1(_10528_),
    .C1(net3881),
    .Y(_10859_));
 sky130_fd_sc_hd__nand2b_1 _20083_ (.A_N(_12221_[0]),
    .B(net3872),
    .Y(_10860_));
 sky130_fd_sc_hd__a21oi_2 _20084_ (.A1(_10860_),
    .A2(_10806_),
    .B1(net3675),
    .Y(_10861_));
 sky130_fd_sc_hd__a21oi_1 _20085_ (.A1(_10663_),
    .A2(_10807_),
    .B1(net3883),
    .Y(_10862_));
 sky130_fd_sc_hd__nor4_1 _20086_ (.A(_10528_),
    .B(net3869),
    .C(_10861_),
    .D(_10862_),
    .Y(_10863_));
 sky130_fd_sc_hd__a211oi_1 _20087_ (.A1(_10528_),
    .A2(_10855_),
    .B1(_10859_),
    .C1(_10863_),
    .Y(_10864_));
 sky130_fd_sc_hd__nor2_1 _20088_ (.A(net3870),
    .B(_10743_),
    .Y(_10865_));
 sky130_fd_sc_hd__nand3_1 _20089_ (.A(net3675),
    .B(_10567_),
    .C(_10797_),
    .Y(_10866_));
 sky130_fd_sc_hd__o311ai_1 _20090_ (.A1(net3675),
    .A2(_10580_),
    .A3(_10650_),
    .B1(_10866_),
    .C1(net3869),
    .Y(_10867_));
 sky130_fd_sc_hd__nand2_1 _20091_ (.A(_12230_[0]),
    .B(_10552_),
    .Y(_10868_));
 sky130_fd_sc_hd__nand3_2 _20092_ (.A(net3888),
    .B(net3886),
    .C(_10550_),
    .Y(_10869_));
 sky130_fd_sc_hd__nand4_1 _20093_ (.A(net3881),
    .B(_10868_),
    .C(_10794_),
    .D(_10869_),
    .Y(_10870_));
 sky130_fd_sc_hd__nand3_1 _20094_ (.A(_10865_),
    .B(_10867_),
    .C(_10870_),
    .Y(_10871_));
 sky130_fd_sc_hd__o21a_1 _20095_ (.A1(_12236_[0]),
    .A2(net3874),
    .B1(_10583_),
    .X(_10872_));
 sky130_fd_sc_hd__nor3_1 _20096_ (.A(net3883),
    .B(_10569_),
    .C(_10643_),
    .Y(_10873_));
 sky130_fd_sc_hd__o21ai_0 _20097_ (.A1(_10872_),
    .A2(_10873_),
    .B1(net3869),
    .Y(_10874_));
 sky130_fd_sc_hd__nand2_1 _20098_ (.A(_12220_[0]),
    .B(net3878),
    .Y(_10875_));
 sky130_fd_sc_hd__nand2_1 _20099_ (.A(_12230_[0]),
    .B(net3874),
    .Y(_10876_));
 sky130_fd_sc_hd__nor4_1 _20100_ (.A(net3883),
    .B(net3869),
    .C(_10634_),
    .D(_10738_),
    .Y(_10877_));
 sky130_fd_sc_hd__a31oi_1 _20101_ (.A1(_10875_),
    .A2(_10664_),
    .A3(_10876_),
    .B1(_10877_),
    .Y(_10878_));
 sky130_fd_sc_hd__nand4_1 _20102_ (.A(net3882),
    .B(_10627_),
    .C(_10874_),
    .D(_10878_),
    .Y(_10879_));
 sky130_fd_sc_hd__o311ai_2 _20103_ (.A1(net3882),
    .A2(net3673),
    .A3(_10864_),
    .B1(_10871_),
    .C1(_10879_),
    .Y(_10880_));
 sky130_fd_sc_hd__a21oi_4 _20104_ (.A1(_10834_),
    .A2(_10849_),
    .B1(_10880_),
    .Y(_00099_));
 sky130_fd_sc_hd__nand2_1 _20105_ (.A(net401),
    .B(net3883),
    .Y(_10881_));
 sky130_fd_sc_hd__a21oi_1 _20106_ (.A1(_10570_),
    .A2(_10881_),
    .B1(net3877),
    .Y(_10882_));
 sky130_fd_sc_hd__nand2_1 _20107_ (.A(net3869),
    .B(_10632_),
    .Y(_10883_));
 sky130_fd_sc_hd__o221ai_1 _20108_ (.A1(net3869),
    .A2(_10710_),
    .B1(_10882_),
    .B2(_10883_),
    .C1(_10626_),
    .Y(_10884_));
 sky130_fd_sc_hd__o21ai_0 _20109_ (.A1(_10656_),
    .A2(_10722_),
    .B1(net3883),
    .Y(_10885_));
 sky130_fd_sc_hd__a31oi_1 _20110_ (.A1(_12221_[0]),
    .A2(_10509_),
    .A3(net3877),
    .B1(_10716_),
    .Y(_10886_));
 sky130_fd_sc_hd__o21ai_0 _20111_ (.A1(net3881),
    .A2(_10886_),
    .B1(_10528_),
    .Y(_10887_));
 sky130_fd_sc_hd__a31oi_1 _20112_ (.A1(net3881),
    .A2(_10611_),
    .A3(_10885_),
    .B1(_10887_),
    .Y(_10888_));
 sky130_fd_sc_hd__nor3_1 _20113_ (.A(net3870),
    .B(_10683_),
    .C(_10888_),
    .Y(_10889_));
 sky130_fd_sc_hd__nand3_1 _20114_ (.A(_10509_),
    .B(_10567_),
    .C(_10810_),
    .Y(_10890_));
 sky130_fd_sc_hd__nand3_1 _20115_ (.A(net3674),
    .B(net3869),
    .C(_10890_),
    .Y(_10891_));
 sky130_fd_sc_hd__a31oi_1 _20116_ (.A1(net3883),
    .A2(_10797_),
    .A3(_10712_),
    .B1(_10891_),
    .Y(_10892_));
 sky130_fd_sc_hd__o21ai_0 _20117_ (.A1(_10509_),
    .A2(_10644_),
    .B1(_10810_),
    .Y(_10893_));
 sky130_fd_sc_hd__o311ai_0 _20118_ (.A1(net3883),
    .A2(_10722_),
    .A3(_10767_),
    .B1(net3869),
    .C1(_10591_),
    .Y(_10894_));
 sky130_fd_sc_hd__o21ai_0 _20119_ (.A1(net3869),
    .A2(_10893_),
    .B1(_10894_),
    .Y(_10895_));
 sky130_fd_sc_hd__nand3_1 _20120_ (.A(_10509_),
    .B(_10696_),
    .C(_10638_),
    .Y(_10896_));
 sky130_fd_sc_hd__o2111ai_1 _20121_ (.A1(_12232_[0]),
    .A2(_10509_),
    .B1(net3674),
    .C1(net3881),
    .D1(_10896_),
    .Y(_10897_));
 sky130_fd_sc_hd__o21ai_0 _20122_ (.A1(net3674),
    .A2(_10895_),
    .B1(_10897_),
    .Y(_10898_));
 sky130_fd_sc_hd__nor4_1 _20123_ (.A(net3870),
    .B(_10534_),
    .C(_10892_),
    .D(_10898_),
    .Y(_10899_));
 sky130_fd_sc_hd__nand2_2 _20124_ (.A(net3886),
    .B(net3877),
    .Y(_10900_));
 sky130_fd_sc_hd__o21bai_1 _20125_ (.A1(net3881),
    .A2(_10900_),
    .B1_N(_10664_),
    .Y(_10901_));
 sky130_fd_sc_hd__a221o_1 _20126_ (.A1(_12220_[0]),
    .A2(_10654_),
    .B1(_10685_),
    .B2(net3869),
    .C1(net3872),
    .X(_10902_));
 sky130_fd_sc_hd__a21oi_1 _20127_ (.A1(_10509_),
    .A2(net3869),
    .B1(_10500_),
    .Y(_10903_));
 sky130_fd_sc_hd__o211ai_1 _20128_ (.A1(net3888),
    .A2(_10903_),
    .B1(_10591_),
    .C1(net3873),
    .Y(_10904_));
 sky130_fd_sc_hd__a221oi_1 _20129_ (.A1(net3888),
    .A2(_10901_),
    .B1(_10902_),
    .B2(_10904_),
    .C1(_10743_),
    .Y(_10905_));
 sky130_fd_sc_hd__o211ai_1 _20130_ (.A1(_10500_),
    .A2(_10557_),
    .B1(_10812_),
    .C1(net3869),
    .Y(_10906_));
 sky130_fd_sc_hd__o21ai_0 _20131_ (.A1(_10643_),
    .A2(_10767_),
    .B1(_10664_),
    .Y(_10907_));
 sky130_fd_sc_hd__o211ai_1 _20132_ (.A1(net3869),
    .A2(_10750_),
    .B1(_10906_),
    .C1(_10907_),
    .Y(_10908_));
 sky130_fd_sc_hd__o21ai_0 _20133_ (.A1(_10720_),
    .A2(_10908_),
    .B1(net3870),
    .Y(_10909_));
 sky130_fd_sc_hd__o21ai_0 _20134_ (.A1(net3888),
    .A2(_10701_),
    .B1(_10611_),
    .Y(_10910_));
 sky130_fd_sc_hd__nand2_1 _20135_ (.A(net3888),
    .B(net3873),
    .Y(_10911_));
 sky130_fd_sc_hd__a21oi_1 _20136_ (.A1(_10911_),
    .A2(_10900_),
    .B1(_10509_),
    .Y(_10912_));
 sky130_fd_sc_hd__o21ai_0 _20137_ (.A1(_10910_),
    .A2(_10912_),
    .B1(net3881),
    .Y(_10913_));
 sky130_fd_sc_hd__a21oi_1 _20138_ (.A1(_10621_),
    .A2(_10622_),
    .B1(_10509_),
    .Y(_10914_));
 sky130_fd_sc_hd__o21ai_0 _20139_ (.A1(_12220_[0]),
    .A2(_10602_),
    .B1(_10869_),
    .Y(_10915_));
 sky130_fd_sc_hd__o21ai_0 _20140_ (.A1(_10914_),
    .A2(_10915_),
    .B1(net3869),
    .Y(_10916_));
 sky130_fd_sc_hd__a21oi_1 _20141_ (.A1(_10913_),
    .A2(_10916_),
    .B1(_10536_),
    .Y(_10917_));
 sky130_fd_sc_hd__nand3_1 _20142_ (.A(net3883),
    .B(_10797_),
    .C(_10638_),
    .Y(_10918_));
 sky130_fd_sc_hd__nand3_1 _20143_ (.A(_10509_),
    .B(_10712_),
    .C(_10806_),
    .Y(_10919_));
 sky130_fd_sc_hd__a21oi_1 _20144_ (.A1(_10918_),
    .A2(_10919_),
    .B1(net3869),
    .Y(_10920_));
 sky130_fd_sc_hd__o21ai_0 _20145_ (.A1(_12220_[0]),
    .A2(_10509_),
    .B1(_10660_),
    .Y(_10921_));
 sky130_fd_sc_hd__a21oi_1 _20146_ (.A1(net3877),
    .A2(_10921_),
    .B1(_10620_),
    .Y(_10922_));
 sky130_fd_sc_hd__nor3_1 _20147_ (.A(_10684_),
    .B(_10920_),
    .C(_10922_),
    .Y(_10923_));
 sky130_fd_sc_hd__nor4_1 _20148_ (.A(_10905_),
    .B(_10909_),
    .C(_10917_),
    .D(_10923_),
    .Y(_10924_));
 sky130_fd_sc_hd__a211oi_1 _20149_ (.A1(_10884_),
    .A2(_10889_),
    .B1(_10899_),
    .C1(_10924_),
    .Y(_00100_));
 sky130_fd_sc_hd__nand2_2 _20150_ (.A(net3884),
    .B(_10711_),
    .Y(_10925_));
 sky130_fd_sc_hd__nand2_2 _20151_ (.A(_12225_[0]),
    .B(net3879),
    .Y(_10926_));
 sky130_fd_sc_hd__nand2_2 _20152_ (.A(_10509_),
    .B(_10926_),
    .Y(_10927_));
 sky130_fd_sc_hd__nor2_1 _20153_ (.A(_12232_[0]),
    .B(net3878),
    .Y(_10928_));
 sky130_fd_sc_hd__o221ai_1 _20154_ (.A1(_10569_),
    .A2(_10925_),
    .B1(_10927_),
    .B2(_10928_),
    .C1(net3882),
    .Y(_10929_));
 sky130_fd_sc_hd__o221ai_1 _20155_ (.A1(_12234_[0]),
    .A2(_10557_),
    .B1(_10783_),
    .B2(_10812_),
    .C1(net3870),
    .Y(_10930_));
 sky130_fd_sc_hd__nand3_1 _20156_ (.A(net3885),
    .B(net3882),
    .C(_10662_),
    .Y(_10931_));
 sky130_fd_sc_hd__a21oi_1 _20157_ (.A1(_10574_),
    .A2(net3875),
    .B1(_10509_),
    .Y(_10932_));
 sky130_fd_sc_hd__nor3_1 _20158_ (.A(net3883),
    .B(_10519_),
    .C(_10550_),
    .Y(_10933_));
 sky130_fd_sc_hd__o22ai_1 _20159_ (.A1(_10574_),
    .A2(net3875),
    .B1(_10932_),
    .B2(_10933_),
    .Y(_10934_));
 sky130_fd_sc_hd__o2bb2ai_1 _20160_ (.A1_N(_12227_[0]),
    .A2_N(_10552_),
    .B1(_10562_),
    .B2(_12234_[0]),
    .Y(_10935_));
 sky130_fd_sc_hd__a22oi_1 _20161_ (.A1(_10500_),
    .A2(_10934_),
    .B1(_10935_),
    .B2(net3870),
    .Y(_10936_));
 sky130_fd_sc_hd__a21oi_2 _20162_ (.A1(_10931_),
    .A2(_10936_),
    .B1(net3881),
    .Y(_10937_));
 sky130_fd_sc_hd__a311oi_1 _20163_ (.A1(net3881),
    .A2(_10929_),
    .A3(_10930_),
    .B1(_10937_),
    .C1(_10683_),
    .Y(_10938_));
 sky130_fd_sc_hd__nand2_1 _20164_ (.A(_12227_[0]),
    .B(net3879),
    .Y(_10939_));
 sky130_fd_sc_hd__o211ai_1 _20165_ (.A1(net3879),
    .A2(_10843_),
    .B1(_10939_),
    .C1(_10606_),
    .Y(_10940_));
 sky130_fd_sc_hd__a21oi_1 _20166_ (.A1(_10840_),
    .A2(_10881_),
    .B1(net3872),
    .Y(_10941_));
 sky130_fd_sc_hd__nor2_1 _20167_ (.A(net3881),
    .B(_10941_),
    .Y(_10942_));
 sky130_fd_sc_hd__a21oi_1 _20168_ (.A1(_10661_),
    .A2(_10942_),
    .B1(net3870),
    .Y(_10943_));
 sky130_fd_sc_hd__nand2_2 _20169_ (.A(net3870),
    .B(net3881),
    .Y(_10944_));
 sky130_fd_sc_hd__a21oi_1 _20170_ (.A1(_10638_),
    .A2(_10927_),
    .B1(_10944_),
    .Y(_10945_));
 sky130_fd_sc_hd__a221oi_1 _20171_ (.A1(_10500_),
    .A2(_10678_),
    .B1(_10583_),
    .B2(_10810_),
    .C1(_10821_),
    .Y(_10946_));
 sky130_fd_sc_hd__a2111oi_1 _20172_ (.A1(_10940_),
    .A2(_10943_),
    .B1(_10945_),
    .C1(_10946_),
    .D1(net3673),
    .Y(_10947_));
 sky130_fd_sc_hd__nand2_1 _20173_ (.A(_12227_[0]),
    .B(_10552_),
    .Y(_10948_));
 sky130_fd_sc_hd__o21ai_0 _20174_ (.A1(_12236_[0]),
    .A2(net3884),
    .B1(net3878),
    .Y(_10949_));
 sky130_fd_sc_hd__o21ai_0 _20175_ (.A1(_10783_),
    .A2(_10812_),
    .B1(net3870),
    .Y(_10950_));
 sky130_fd_sc_hd__a21oi_1 _20176_ (.A1(_10583_),
    .A2(_10711_),
    .B1(_10950_),
    .Y(_10951_));
 sky130_fd_sc_hd__a31oi_1 _20177_ (.A1(net3882),
    .A2(_10948_),
    .A3(_10949_),
    .B1(_10951_),
    .Y(_10952_));
 sky130_fd_sc_hd__nand2_4 _20178_ (.A(_12225_[0]),
    .B(_10552_),
    .Y(_10953_));
 sky130_fd_sc_hd__o21ai_0 _20179_ (.A1(_10716_),
    .A2(_10758_),
    .B1(net3883),
    .Y(_10954_));
 sky130_fd_sc_hd__nand3_1 _20180_ (.A(net3882),
    .B(_10953_),
    .C(_10954_),
    .Y(_10955_));
 sky130_fd_sc_hd__a211o_1 _20181_ (.A1(_12234_[0]),
    .A2(_10633_),
    .B1(_10783_),
    .C1(net3882),
    .X(_10956_));
 sky130_fd_sc_hd__a31oi_1 _20182_ (.A1(net3869),
    .A2(_10955_),
    .A3(_10956_),
    .B1(_10536_),
    .Y(_10957_));
 sky130_fd_sc_hd__o21ai_1 _20183_ (.A1(net3869),
    .A2(_10952_),
    .B1(_10957_),
    .Y(_10958_));
 sky130_fd_sc_hd__a21oi_1 _20184_ (.A1(_10696_),
    .A2(_10621_),
    .B1(net3883),
    .Y(_10959_));
 sky130_fd_sc_hd__nor2_1 _20185_ (.A(_10495_),
    .B(_10557_),
    .Y(_10960_));
 sky130_fd_sc_hd__o21ai_2 _20186_ (.A1(_10959_),
    .A2(_10960_),
    .B1(net3881),
    .Y(_10961_));
 sky130_fd_sc_hd__nand2b_1 _20187_ (.A_N(_12220_[0]),
    .B(net3877),
    .Y(_10962_));
 sky130_fd_sc_hd__a21oi_2 _20188_ (.A1(_10962_),
    .A2(_10712_),
    .B1(net3883),
    .Y(_10963_));
 sky130_fd_sc_hd__o21ai_0 _20189_ (.A1(_10563_),
    .A2(_10963_),
    .B1(net3869),
    .Y(_10964_));
 sky130_fd_sc_hd__nand2_1 _20190_ (.A(net3881),
    .B(_10754_),
    .Y(_10965_));
 sky130_fd_sc_hd__o21ai_0 _20191_ (.A1(net3888),
    .A2(net3881),
    .B1(_10965_),
    .Y(_10966_));
 sky130_fd_sc_hd__a21oi_1 _20192_ (.A1(_10500_),
    .A2(_10595_),
    .B1(_10850_),
    .Y(_10967_));
 sky130_fd_sc_hd__nand3_1 _20193_ (.A(_10585_),
    .B(net3876),
    .C(net3611),
    .Y(_10968_));
 sky130_fd_sc_hd__o2111ai_1 _20194_ (.A1(net3888),
    .A2(_10967_),
    .B1(_10968_),
    .C1(_10719_),
    .D1(net3882),
    .Y(_10969_));
 sky130_fd_sc_hd__a21oi_2 _20195_ (.A1(net3880),
    .A2(_10966_),
    .B1(_10969_),
    .Y(_10970_));
 sky130_fd_sc_hd__a311o_1 _20196_ (.A1(net3870),
    .A2(_10961_),
    .A3(_10964_),
    .B1(_10684_),
    .C1(_10970_),
    .X(_10971_));
 sky130_fd_sc_hd__o311ai_2 _20197_ (.A1(_10528_),
    .A2(_10938_),
    .A3(_10947_),
    .B1(_10958_),
    .C1(_10971_),
    .Y(_00101_));
 sky130_fd_sc_hd__nor2_2 _20198_ (.A(_12232_[0]),
    .B(net3873),
    .Y(_10972_));
 sky130_fd_sc_hd__a21oi_1 _20199_ (.A1(_12230_[0]),
    .A2(net3873),
    .B1(_10972_),
    .Y(_10973_));
 sky130_fd_sc_hd__o221ai_1 _20200_ (.A1(_10495_),
    .A2(_10562_),
    .B1(_10973_),
    .B2(net3883),
    .C1(net3881),
    .Y(_10974_));
 sky130_fd_sc_hd__nand2_1 _20201_ (.A(_12240_[0]),
    .B(net3880),
    .Y(_10975_));
 sky130_fd_sc_hd__nand3_1 _20202_ (.A(net3873),
    .B(_10762_),
    .C(_10843_),
    .Y(_10976_));
 sky130_fd_sc_hd__a21oi_1 _20203_ (.A1(_10975_),
    .A2(_10976_),
    .B1(_10694_),
    .Y(_10977_));
 sky130_fd_sc_hd__nor4b_1 _20204_ (.A(_10563_),
    .B(_10774_),
    .C(_10822_),
    .D_N(_10679_),
    .Y(_10978_));
 sky130_fd_sc_hd__a311oi_1 _20205_ (.A1(net3870),
    .A2(_10800_),
    .A3(_10974_),
    .B1(_10977_),
    .C1(_10978_),
    .Y(_10979_));
 sky130_fd_sc_hd__nand2_1 _20206_ (.A(net3673),
    .B(_10979_),
    .Y(_10980_));
 sky130_fd_sc_hd__o21ai_0 _20207_ (.A1(_10644_),
    .A2(_10927_),
    .B1(_10724_),
    .Y(_10981_));
 sky130_fd_sc_hd__nor2_1 _20208_ (.A(_12221_[0]),
    .B(net3675),
    .Y(_10982_));
 sky130_fd_sc_hd__a211oi_1 _20209_ (.A1(net3595),
    .A2(net3675),
    .B1(net3878),
    .C1(_10982_),
    .Y(_10983_));
 sky130_fd_sc_hd__o21ai_0 _20210_ (.A1(_12241_[0]),
    .A2(net3874),
    .B1(_10699_),
    .Y(_10984_));
 sky130_fd_sc_hd__o22a_1 _20211_ (.A1(_10861_),
    .A2(_10981_),
    .B1(_10983_),
    .B2(_10984_),
    .X(_10985_));
 sky130_fd_sc_hd__a21oi_1 _20212_ (.A1(net3873),
    .A2(_10824_),
    .B1(_10509_),
    .Y(_10986_));
 sky130_fd_sc_hd__a32oi_1 _20213_ (.A1(_10509_),
    .A2(_10567_),
    .A3(_10622_),
    .B1(_10926_),
    .B2(_10986_),
    .Y(_10987_));
 sky130_fd_sc_hd__nand2_1 _20214_ (.A(_10715_),
    .B(_10987_),
    .Y(_10988_));
 sky130_fd_sc_hd__nor2_1 _20215_ (.A(_12230_[0]),
    .B(net3878),
    .Y(_10989_));
 sky130_fd_sc_hd__o21ai_0 _20216_ (.A1(_10749_),
    .A2(_10989_),
    .B1(net3675),
    .Y(_10990_));
 sky130_fd_sc_hd__o211ai_1 _20217_ (.A1(net3595),
    .A2(_10562_),
    .B1(_10707_),
    .C1(_10990_),
    .Y(_10991_));
 sky130_fd_sc_hd__nand4_1 _20218_ (.A(_10683_),
    .B(_10985_),
    .C(_10988_),
    .D(_10991_),
    .Y(_10992_));
 sky130_fd_sc_hd__nand2_1 _20219_ (.A(_12232_[0]),
    .B(net3883),
    .Y(_10993_));
 sky130_fd_sc_hd__nor2_1 _20220_ (.A(net3875),
    .B(_10993_),
    .Y(_10994_));
 sky130_fd_sc_hd__o22ai_1 _20221_ (.A1(_10509_),
    .A2(_10567_),
    .B1(_10554_),
    .B2(_10500_),
    .Y(_10995_));
 sky130_fd_sc_hd__nor3_1 _20222_ (.A(net3881),
    .B(_10994_),
    .C(_10995_),
    .Y(_10996_));
 sky130_fd_sc_hd__nor4_1 _20223_ (.A(_10585_),
    .B(_10550_),
    .C(_10831_),
    .D(_10675_),
    .Y(_10997_));
 sky130_fd_sc_hd__a2111oi_0 _20224_ (.A1(_12250_[0]),
    .A2(_10828_),
    .B1(_10996_),
    .C1(_10997_),
    .D1(_10519_),
    .Y(_10998_));
 sky130_fd_sc_hd__a21oi_1 _20225_ (.A1(_10509_),
    .A2(_10900_),
    .B1(net3888),
    .Y(_10999_));
 sky130_fd_sc_hd__o211ai_1 _20226_ (.A1(net3875),
    .A2(_10591_),
    .B1(_10724_),
    .C1(_10953_),
    .Y(_11000_));
 sky130_fd_sc_hd__nor2_1 _20227_ (.A(_10630_),
    .B(_10774_),
    .Y(_11001_));
 sky130_fd_sc_hd__o211ai_1 _20228_ (.A1(_12236_[0]),
    .A2(_10557_),
    .B1(_10869_),
    .C1(_11001_),
    .Y(_11002_));
 sky130_fd_sc_hd__o21ai_0 _20229_ (.A1(_10999_),
    .A2(_11000_),
    .B1(_11002_),
    .Y(_11003_));
 sky130_fd_sc_hd__mux2i_1 _20230_ (.A0(_12236_[0]),
    .A1(_12232_[0]),
    .S(_10509_),
    .Y(_11004_));
 sky130_fd_sc_hd__o21ai_0 _20231_ (.A1(net3880),
    .A2(_11004_),
    .B1(_10585_),
    .Y(_11005_));
 sky130_fd_sc_hd__a211oi_1 _20232_ (.A1(_12234_[0]),
    .A2(_10509_),
    .B1(net3873),
    .C1(_10659_),
    .Y(_11006_));
 sky130_fd_sc_hd__or4_1 _20233_ (.A(_12239_[0]),
    .B(_12248_[0]),
    .C(net3880),
    .D(_10694_),
    .X(_11007_));
 sky130_fd_sc_hd__o31ai_1 _20234_ (.A1(net3882),
    .A2(_11005_),
    .A3(_11006_),
    .B1(_11007_),
    .Y(_11008_));
 sky130_fd_sc_hd__or2_4 _20235_ (.A(_10649_),
    .B(_10825_),
    .X(_11009_));
 sky130_fd_sc_hd__o21ai_0 _20236_ (.A1(_10671_),
    .A2(_10972_),
    .B1(net3883),
    .Y(_11010_));
 sky130_fd_sc_hd__a21oi_2 _20237_ (.A1(_11009_),
    .A2(_11010_),
    .B1(_10944_),
    .Y(_11011_));
 sky130_fd_sc_hd__o21ai_2 _20238_ (.A1(net3611),
    .A2(_10857_),
    .B1(net3880),
    .Y(_11012_));
 sky130_fd_sc_hd__nor2_1 _20239_ (.A(_10694_),
    .B(_11012_),
    .Y(_11013_));
 sky130_fd_sc_hd__nor3_1 _20240_ (.A(_12220_[0]),
    .B(_10509_),
    .C(net390),
    .Y(_11014_));
 sky130_fd_sc_hd__a2111oi_0 _20241_ (.A1(_12222_[0]),
    .A2(_10678_),
    .B1(_10774_),
    .C1(_11014_),
    .D1(_10994_),
    .Y(_11015_));
 sky130_fd_sc_hd__nor4_1 _20242_ (.A(_11008_),
    .B(_11011_),
    .C(_11013_),
    .D(_11015_),
    .Y(_11016_));
 sky130_fd_sc_hd__o32ai_1 _20243_ (.A1(_10720_),
    .A2(_10998_),
    .A3(_11003_),
    .B1(_11016_),
    .B2(_10743_),
    .Y(_11017_));
 sky130_fd_sc_hd__a31oi_1 _20244_ (.A1(_10528_),
    .A2(_10980_),
    .A3(_10992_),
    .B1(_11017_),
    .Y(_00102_));
 sky130_fd_sc_hd__o22a_1 _20245_ (.A1(net402),
    .A2(_10562_),
    .B1(_10779_),
    .B2(net3878),
    .X(_11018_));
 sky130_fd_sc_hd__o21ai_0 _20246_ (.A1(_10662_),
    .A2(_10925_),
    .B1(net3870),
    .Y(_11019_));
 sky130_fd_sc_hd__a31oi_1 _20247_ (.A1(net3675),
    .A2(_10696_),
    .A3(_10701_),
    .B1(_11019_),
    .Y(_11020_));
 sky130_fd_sc_hd__a311oi_1 _20248_ (.A1(net3882),
    .A2(_10750_),
    .A3(_11018_),
    .B1(_11020_),
    .C1(net3869),
    .Y(_11021_));
 sky130_fd_sc_hd__nor2_1 _20249_ (.A(_12248_[0]),
    .B(net3875),
    .Y(_11022_));
 sky130_fd_sc_hd__a311oi_2 _20250_ (.A1(net3875),
    .A2(_10570_),
    .A3(_10993_),
    .B1(_11022_),
    .C1(net3882),
    .Y(_11023_));
 sky130_fd_sc_hd__a21oi_1 _20251_ (.A1(_12222_[0]),
    .A2(_10552_),
    .B1(_10745_),
    .Y(_11024_));
 sky130_fd_sc_hd__nor2_1 _20252_ (.A(net3870),
    .B(_11024_),
    .Y(_11025_));
 sky130_fd_sc_hd__nor3_2 _20253_ (.A(net3881),
    .B(_11023_),
    .C(_11025_),
    .Y(_11026_));
 sky130_fd_sc_hd__nor2_1 _20254_ (.A(net3885),
    .B(_10541_),
    .Y(_11027_));
 sky130_fd_sc_hd__o32ai_1 _20255_ (.A1(_10541_),
    .A2(_10550_),
    .A3(_10762_),
    .B1(_10554_),
    .B2(net3888),
    .Y(_11028_));
 sky130_fd_sc_hd__nor4_1 _20256_ (.A(_12234_[0]),
    .B(net3883),
    .C(_10541_),
    .D(_10550_),
    .Y(_11029_));
 sky130_fd_sc_hd__a2111oi_1 _20257_ (.A1(_10749_),
    .A2(_11027_),
    .B1(_11028_),
    .C1(_10574_),
    .D1(_11029_),
    .Y(_11030_));
 sky130_fd_sc_hd__o21ai_0 _20258_ (.A1(_10500_),
    .A2(_10562_),
    .B1(_10701_),
    .Y(_11031_));
 sky130_fd_sc_hd__nand2_1 _20259_ (.A(_10541_),
    .B(_11031_),
    .Y(_11032_));
 sky130_fd_sc_hd__a21oi_1 _20260_ (.A1(_12234_[0]),
    .A2(net3876),
    .B1(net3883),
    .Y(_11033_));
 sky130_fd_sc_hd__a31oi_1 _20261_ (.A1(net3883),
    .A2(_10567_),
    .A3(_10926_),
    .B1(_11033_),
    .Y(_11034_));
 sky130_fd_sc_hd__a31oi_1 _20262_ (.A1(_10585_),
    .A2(_10583_),
    .A3(_10709_),
    .B1(net3882),
    .Y(_11035_));
 sky130_fd_sc_hd__o21a_1 _20263_ (.A1(_10585_),
    .A2(_11034_),
    .B1(_11035_),
    .X(_11036_));
 sky130_fd_sc_hd__a211oi_1 _20264_ (.A1(_11030_),
    .A2(_11032_),
    .B1(_10536_),
    .C1(_11036_),
    .Y(_11037_));
 sky130_fd_sc_hd__o221ai_1 _20265_ (.A1(_12236_[0]),
    .A2(_10562_),
    .B1(_10732_),
    .B2(_12221_[0]),
    .C1(_10719_),
    .Y(_11038_));
 sky130_fd_sc_hd__nand2_1 _20266_ (.A(net3876),
    .B(_11004_),
    .Y(_11039_));
 sky130_fd_sc_hd__nand3_1 _20267_ (.A(net3880),
    .B(_10591_),
    .C(_10660_),
    .Y(_11040_));
 sky130_fd_sc_hd__a21oi_1 _20268_ (.A1(_11039_),
    .A2(_11040_),
    .B1(_10541_),
    .Y(_11041_));
 sky130_fd_sc_hd__a2111oi_0 _20269_ (.A1(_10541_),
    .A2(_11038_),
    .B1(_11041_),
    .C1(_10720_),
    .D1(net3882),
    .Y(_11042_));
 sky130_fd_sc_hd__nand3_1 _20270_ (.A(net3879),
    .B(_10762_),
    .C(_10843_),
    .Y(_11043_));
 sky130_fd_sc_hd__o211ai_1 _20271_ (.A1(_12236_[0]),
    .A2(_10557_),
    .B1(_11043_),
    .C1(_10585_),
    .Y(_11044_));
 sky130_fd_sc_hd__o41ai_1 _20272_ (.A1(_10624_),
    .A2(_10605_),
    .A3(_10822_),
    .A4(_10729_),
    .B1(net3881),
    .Y(_11045_));
 sky130_fd_sc_hd__a211oi_1 _20273_ (.A1(_11044_),
    .A2(_11045_),
    .B1(net3870),
    .C1(_10720_),
    .Y(_11046_));
 sky130_fd_sc_hd__nor3_2 _20274_ (.A(_11037_),
    .B(_11042_),
    .C(_11046_),
    .Y(_11047_));
 sky130_fd_sc_hd__o21ai_0 _20275_ (.A1(_12227_[0]),
    .A2(net3879),
    .B1(_11012_),
    .Y(_11048_));
 sky130_fd_sc_hd__nor3_1 _20276_ (.A(_10509_),
    .B(_10662_),
    .C(_10758_),
    .Y(_11049_));
 sky130_fd_sc_hd__nor3_1 _20277_ (.A(net3883),
    .B(_10716_),
    .C(_10972_),
    .Y(_11050_));
 sky130_fd_sc_hd__nor3_1 _20278_ (.A(net3870),
    .B(_11049_),
    .C(_11050_),
    .Y(_11051_));
 sky130_fd_sc_hd__a21oi_1 _20279_ (.A1(net3870),
    .A2(_11048_),
    .B1(_11051_),
    .Y(_11052_));
 sky130_fd_sc_hd__o32ai_1 _20280_ (.A1(net3883),
    .A2(_10580_),
    .A3(_10650_),
    .B1(_10925_),
    .B2(_10723_),
    .Y(_11053_));
 sky130_fd_sc_hd__nor2_1 _20281_ (.A(_12220_[0]),
    .B(_10509_),
    .Y(_11054_));
 sky130_fd_sc_hd__nor3_1 _20282_ (.A(net3883),
    .B(_10644_),
    .C(_10722_),
    .Y(_11055_));
 sky130_fd_sc_hd__nor3_1 _20283_ (.A(_10821_),
    .B(_11054_),
    .C(_11055_),
    .Y(_11056_));
 sky130_fd_sc_hd__a211oi_1 _20284_ (.A1(_10724_),
    .A2(_11053_),
    .B1(_11056_),
    .C1(_10743_),
    .Y(_11057_));
 sky130_fd_sc_hd__o21ai_2 _20285_ (.A1(net3869),
    .A2(_11052_),
    .B1(_11057_),
    .Y(_11058_));
 sky130_fd_sc_hd__o311ai_4 _20286_ (.A1(_10684_),
    .A2(_11021_),
    .A3(_11026_),
    .B1(_11047_),
    .C1(_11058_),
    .Y(_00103_));
 sky130_fd_sc_hd__xnor2_1 _20287_ (.A(net4227),
    .B(\sa30_sub[7] ),
    .Y(_11059_));
 sky130_fd_sc_hd__xnor2_1 _20288_ (.A(\sa11_sr[1] ),
    .B(\sa30_sub[0] ),
    .Y(_11060_));
 sky130_fd_sc_hd__xnor3_1 _20289_ (.A(\sa30_sub[1] ),
    .B(net4206),
    .C(net4202),
    .X(_11061_));
 sky130_fd_sc_hd__xnor3_1 _20290_ (.A(_11059_),
    .B(_11060_),
    .C(_11061_),
    .X(_11062_));
 sky130_fd_sc_hd__mux2i_1 _20291_ (.A0(\text_in_r[73] ),
    .A1(_11062_),
    .S(net4117),
    .Y(_11063_));
 sky130_fd_sc_hd__xor2_1 _20292_ (.A(\u0.w[1][9] ),
    .B(_11063_),
    .X(_11064_));
 sky130_fd_sc_hd__clkinv_8 _20293_ (.A(net3867),
    .Y(_11065_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_433 ();
 sky130_fd_sc_hd__xnor3_1 _20296_ (.A(net4215),
    .B(\sa21_sr[7] ),
    .C(\sa30_sub[7] ),
    .X(_11067_));
 sky130_fd_sc_hd__xnor2_1 _20297_ (.A(_08808_),
    .B(_11067_),
    .Y(_11068_));
 sky130_fd_sc_hd__mux2i_1 _20298_ (.A0(\text_in_r[72] ),
    .A1(_11068_),
    .S(net4119),
    .Y(_11069_));
 sky130_fd_sc_hd__xor2_1 _20299_ (.A(\u0.w[1][8] ),
    .B(_11069_),
    .X(_11070_));
 sky130_fd_sc_hd__clkinv_16 _20300_ (.A(net3865),
    .Y(_11071_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_432 ();
 sky130_fd_sc_hd__xnor3_1 _20302_ (.A(\sa11_sr[2] ),
    .B(\sa30_sub[2] ),
    .C(net4226),
    .X(_11072_));
 sky130_fd_sc_hd__xor2_1 _20303_ (.A(_06479_),
    .B(_11072_),
    .X(_11073_));
 sky130_fd_sc_hd__mux2i_4 _20304_ (.A0(\text_in_r[74] ),
    .A1(_11073_),
    .S(net4119),
    .Y(_11074_));
 sky130_fd_sc_hd__xnor2_4 _20305_ (.A(\u0.w[1][10] ),
    .B(_11074_),
    .Y(_11075_));
 sky130_fd_sc_hd__clkinv_16 _20306_ (.A(_11075_),
    .Y(_11076_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_424 ();
 sky130_fd_sc_hd__xnor2_1 _20315_ (.A(net4203),
    .B(\sa30_sub[6] ),
    .Y(_11082_));
 sky130_fd_sc_hd__xnor3_1 _20316_ (.A(\sa30_sub[5] ),
    .B(\sa11_sr[6] ),
    .C(\sa01_sr[6] ),
    .X(_11083_));
 sky130_fd_sc_hd__xnor2_2 _20317_ (.A(_11082_),
    .B(_11083_),
    .Y(_11084_));
 sky130_fd_sc_hd__nor2_2 _20318_ (.A(net398),
    .B(_11084_),
    .Y(_11085_));
 sky130_fd_sc_hd__a21oi_4 _20319_ (.A1(net398),
    .A2(\text_in_r[78] ),
    .B1(_11085_),
    .Y(_11086_));
 sky130_fd_sc_hd__xor2_4 _20320_ (.A(\u0.w[1][14] ),
    .B(_11086_),
    .X(_11087_));
 sky130_fd_sc_hd__xnor2_1 _20321_ (.A(\sa01_sr[7] ),
    .B(\sa30_sub[6] ),
    .Y(_11088_));
 sky130_fd_sc_hd__xnor2_1 _20322_ (.A(_08888_),
    .B(_11088_),
    .Y(_11089_));
 sky130_fd_sc_hd__xnor2_2 _20323_ (.A(net4214),
    .B(_11089_),
    .Y(_11090_));
 sky130_fd_sc_hd__mux2i_2 _20324_ (.A0(\text_in_r[79] ),
    .A1(_11090_),
    .S(_05879_),
    .Y(_11091_));
 sky130_fd_sc_hd__xnor2_4 _20325_ (.A(\u0.w[1][15] ),
    .B(_11091_),
    .Y(_11092_));
 sky130_fd_sc_hd__nor2_4 _20326_ (.A(_11087_),
    .B(_11092_),
    .Y(_11093_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_422 ();
 sky130_fd_sc_hd__xnor2_1 _20329_ (.A(net4225),
    .B(\sa30_sub[7] ),
    .Y(_11096_));
 sky130_fd_sc_hd__xnor2_1 _20330_ (.A(\sa30_sub[2] ),
    .B(\sa11_sr[3] ),
    .Y(_11097_));
 sky130_fd_sc_hd__xnor3_1 _20331_ (.A(_08831_),
    .B(_11096_),
    .C(_11097_),
    .X(_11098_));
 sky130_fd_sc_hd__nand2b_2 _20332_ (.A_N(\text_in_r[75] ),
    .B(net398),
    .Y(_11099_));
 sky130_fd_sc_hd__o211a_4 _20333_ (.A1(net398),
    .A2(_11098_),
    .B1(_11099_),
    .C1(\u0.w[1][11] ),
    .X(_11100_));
 sky130_fd_sc_hd__and2_4 _20334_ (.A(net398),
    .B(\text_in_r[75] ),
    .X(_11101_));
 sky130_fd_sc_hd__a211oi_2 _20335_ (.A1(net4121),
    .A2(_11098_),
    .B1(_11101_),
    .C1(\u0.w[1][11] ),
    .Y(_11102_));
 sky130_fd_sc_hd__nor2_4 _20336_ (.A(_11100_),
    .B(_11102_),
    .Y(_11103_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_421 ();
 sky130_fd_sc_hd__nor2_4 _20338_ (.A(net3672),
    .B(net3862),
    .Y(_11105_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_420 ();
 sky130_fd_sc_hd__o211ai_1 _20340_ (.A1(net398),
    .A2(_11098_),
    .B1(_11099_),
    .C1(\u0.w[1][11] ),
    .Y(_11107_));
 sky130_fd_sc_hd__a211o_4 _20341_ (.A1(net4121),
    .A2(_11098_),
    .B1(_11101_),
    .C1(\u0.w[1][11] ),
    .X(_11108_));
 sky130_fd_sc_hd__nand2_4 _20342_ (.A(_11107_),
    .B(_11108_),
    .Y(_11109_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_418 ();
 sky130_fd_sc_hd__nor2_4 _20345_ (.A(_12272_[0]),
    .B(net3860),
    .Y(_11112_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_417 ();
 sky130_fd_sc_hd__nand2_4 _20347_ (.A(_12261_[0]),
    .B(net3858),
    .Y(_11114_));
 sky130_fd_sc_hd__nand2_8 _20348_ (.A(net3866),
    .B(net3862),
    .Y(_11115_));
 sky130_fd_sc_hd__nand3_1 _20349_ (.A(net3670),
    .B(_11114_),
    .C(_11115_),
    .Y(_11116_));
 sky130_fd_sc_hd__xor2_1 _20350_ (.A(\sa01_sr[4] ),
    .B(\sa30_sub[7] ),
    .X(_11117_));
 sky130_fd_sc_hd__xnor2_1 _20351_ (.A(net4188),
    .B(\sa11_sr[4] ),
    .Y(_11118_));
 sky130_fd_sc_hd__xor3_1 _20352_ (.A(\sa21_sr[3] ),
    .B(\sa30_sub[4] ),
    .C(net4202),
    .X(_11119_));
 sky130_fd_sc_hd__xnor3_1 _20353_ (.A(_11117_),
    .B(_11118_),
    .C(_11119_),
    .X(_11120_));
 sky130_fd_sc_hd__mux2i_4 _20354_ (.A0(\text_in_r[76] ),
    .A1(_11120_),
    .S(net4121),
    .Y(_11121_));
 sky130_fd_sc_hd__xnor2_4 _20355_ (.A(\u0.w[1][12] ),
    .B(_11121_),
    .Y(_11122_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_416 ();
 sky130_fd_sc_hd__o311ai_1 _20357_ (.A1(net3670),
    .A2(_11105_),
    .A3(_11112_),
    .B1(_11116_),
    .C1(net3857),
    .Y(_11124_));
 sky130_fd_sc_hd__xor2_1 _20358_ (.A(\u0.w[1][12] ),
    .B(_11121_),
    .X(_11125_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_415 ();
 sky130_fd_sc_hd__nor2_1 _20360_ (.A(_12270_[0]),
    .B(_11076_),
    .Y(_11127_));
 sky130_fd_sc_hd__nor2_1 _20361_ (.A(net3866),
    .B(net3863),
    .Y(_11128_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_414 ();
 sky130_fd_sc_hd__o21ai_0 _20363_ (.A1(_11127_),
    .A2(_11128_),
    .B1(net3862),
    .Y(_11130_));
 sky130_fd_sc_hd__and2_0 _20364_ (.A(net3855),
    .B(_11130_),
    .X(_11131_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_411 ();
 sky130_fd_sc_hd__nand2_2 _20368_ (.A(net3672),
    .B(_11076_),
    .Y(_11135_));
 sky130_fd_sc_hd__o211ai_1 _20369_ (.A1(_12258_[0]),
    .A2(_11076_),
    .B1(net3858),
    .C1(_11135_),
    .Y(_11136_));
 sky130_fd_sc_hd__xor2_1 _20370_ (.A(\sa30_sub[4] ),
    .B(\sa11_sr[5] ),
    .X(_11137_));
 sky130_fd_sc_hd__xnor2_2 _20371_ (.A(_08823_),
    .B(_11137_),
    .Y(_11138_));
 sky130_fd_sc_hd__mux2i_4 _20372_ (.A0(\text_in_r[77] ),
    .A1(_11138_),
    .S(_05879_),
    .Y(_11139_));
 sky130_fd_sc_hd__xnor2_4 _20373_ (.A(net4156),
    .B(_11139_),
    .Y(_11140_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_408 ();
 sky130_fd_sc_hd__a21oi_1 _20377_ (.A1(_11131_),
    .A2(_11136_),
    .B1(net3854),
    .Y(_11144_));
 sky130_fd_sc_hd__nand2_1 _20378_ (.A(_11124_),
    .B(_11144_),
    .Y(_11145_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_407 ();
 sky130_fd_sc_hd__or3_4 _20380_ (.A(_12272_[0]),
    .B(_11100_),
    .C(_11102_),
    .X(_11147_));
 sky130_fd_sc_hd__nand3_4 _20381_ (.A(_12257_[0]),
    .B(_11107_),
    .C(_11108_),
    .Y(_11148_));
 sky130_fd_sc_hd__nand2_1 _20382_ (.A(net3671),
    .B(net3859),
    .Y(_11149_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_405 ();
 sky130_fd_sc_hd__a21oi_1 _20385_ (.A1(_11148_),
    .A2(net3610),
    .B1(net3670),
    .Y(_11152_));
 sky130_fd_sc_hd__a31oi_1 _20386_ (.A1(net3670),
    .A2(_11114_),
    .A3(_11147_),
    .B1(_11152_),
    .Y(_11153_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_403 ();
 sky130_fd_sc_hd__nand2_8 _20389_ (.A(net3863),
    .B(net3862),
    .Y(_11156_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_401 ();
 sky130_fd_sc_hd__nor2_4 _20392_ (.A(net3671),
    .B(net3862),
    .Y(_11159_));
 sky130_fd_sc_hd__a21oi_1 _20393_ (.A1(_12261_[0]),
    .A2(net3862),
    .B1(_11159_),
    .Y(_11160_));
 sky130_fd_sc_hd__o221ai_1 _20394_ (.A1(_12263_[0]),
    .A2(_11156_),
    .B1(_11160_),
    .B2(net3864),
    .C1(net3855),
    .Y(_11161_));
 sky130_fd_sc_hd__o21ai_1 _20395_ (.A1(net3855),
    .A2(_11153_),
    .B1(_11161_),
    .Y(_11162_));
 sky130_fd_sc_hd__nand2_1 _20396_ (.A(_11140_),
    .B(_11162_),
    .Y(_11163_));
 sky130_fd_sc_hd__nand2_8 _20397_ (.A(_11087_),
    .B(_11092_),
    .Y(_11164_));
 sky130_fd_sc_hd__clkinvlp_2 _20398_ (.A(_12261_[0]),
    .Y(_11165_));
 sky130_fd_sc_hd__mux2i_1 _20399_ (.A0(_12263_[0]),
    .A1(_11165_),
    .S(net3863),
    .Y(_11166_));
 sky130_fd_sc_hd__o21ai_4 _20400_ (.A1(net3861),
    .A2(_11166_),
    .B1(net3855),
    .Y(_11167_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_400 ();
 sky130_fd_sc_hd__nor2_2 _20402_ (.A(_12256_[0]),
    .B(_11156_),
    .Y(_11169_));
 sky130_fd_sc_hd__nand2_4 _20403_ (.A(_11071_),
    .B(net3861),
    .Y(_11170_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_399 ();
 sky130_fd_sc_hd__nand2_2 _20405_ (.A(_12258_[0]),
    .B(net3858),
    .Y(_11172_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_398 ();
 sky130_fd_sc_hd__a21oi_1 _20407_ (.A1(_11170_),
    .A2(_11172_),
    .B1(net3863),
    .Y(_11174_));
 sky130_fd_sc_hd__nor3_1 _20408_ (.A(_11167_),
    .B(_11169_),
    .C(_11174_),
    .Y(_11175_));
 sky130_fd_sc_hd__nor2_4 _20409_ (.A(net3863),
    .B(net3861),
    .Y(_11176_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_395 ();
 sky130_fd_sc_hd__a221oi_1 _20413_ (.A1(_12279_[0]),
    .A2(net3861),
    .B1(_11176_),
    .B2(_12257_[0]),
    .C1(net3855),
    .Y(_11180_));
 sky130_fd_sc_hd__nor3_1 _20414_ (.A(_11140_),
    .B(_11175_),
    .C(_11180_),
    .Y(_11181_));
 sky130_fd_sc_hd__nor2_4 _20415_ (.A(_12266_[0]),
    .B(net3861),
    .Y(_11182_));
 sky130_fd_sc_hd__nand2_1 _20416_ (.A(_11076_),
    .B(_11182_),
    .Y(_11183_));
 sky130_fd_sc_hd__nor2_2 _20417_ (.A(_12258_[0]),
    .B(net3858),
    .Y(_11184_));
 sky130_fd_sc_hd__nor2_1 _20418_ (.A(_11076_),
    .B(_11184_),
    .Y(_11185_));
 sky130_fd_sc_hd__nand2_4 _20419_ (.A(_11114_),
    .B(_11185_),
    .Y(_11186_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_394 ();
 sky130_fd_sc_hd__nor2_4 _20421_ (.A(net3863),
    .B(net3858),
    .Y(_11188_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_393 ();
 sky130_fd_sc_hd__nor2_4 _20423_ (.A(_12258_[0]),
    .B(net3862),
    .Y(_11190_));
 sky130_fd_sc_hd__a21oi_1 _20424_ (.A1(_12261_[0]),
    .A2(net3861),
    .B1(_11190_),
    .Y(_11191_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_392 ();
 sky130_fd_sc_hd__a221oi_1 _20426_ (.A1(_12268_[0]),
    .A2(_11188_),
    .B1(_11191_),
    .B2(net3863),
    .C1(net3856),
    .Y(_11193_));
 sky130_fd_sc_hd__xor2_4 _20427_ (.A(net4156),
    .B(_11139_),
    .X(_11194_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_390 ();
 sky130_fd_sc_hd__a311oi_1 _20430_ (.A1(net3856),
    .A2(_11183_),
    .A3(_11186_),
    .B1(_11193_),
    .C1(_11194_),
    .Y(_11197_));
 sky130_fd_sc_hd__nor3_1 _20431_ (.A(_11164_),
    .B(_11181_),
    .C(_11197_),
    .Y(_11198_));
 sky130_fd_sc_hd__nand2_8 _20432_ (.A(_11071_),
    .B(net3863),
    .Y(_11199_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_389 ();
 sky130_fd_sc_hd__nand2_1 _20434_ (.A(net3868),
    .B(net3866),
    .Y(_11201_));
 sky130_fd_sc_hd__a21oi_1 _20435_ (.A1(_11199_),
    .A2(_11201_),
    .B1(_11194_),
    .Y(_11202_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_388 ();
 sky130_fd_sc_hd__nor3_1 _20437_ (.A(_12257_[0]),
    .B(net3863),
    .C(_11140_),
    .Y(_11204_));
 sky130_fd_sc_hd__a21oi_1 _20438_ (.A1(net3866),
    .A2(_11140_),
    .B1(_11076_),
    .Y(_11205_));
 sky130_fd_sc_hd__nand3_1 _20439_ (.A(_12257_[0]),
    .B(net3863),
    .C(_11194_),
    .Y(_11206_));
 sky130_fd_sc_hd__nand3_1 _20440_ (.A(_11071_),
    .B(_11076_),
    .C(_11140_),
    .Y(_11207_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_387 ();
 sky130_fd_sc_hd__o2111ai_1 _20442_ (.A1(net3868),
    .A2(_11205_),
    .B1(_11206_),
    .C1(_11207_),
    .D1(net3858),
    .Y(_11209_));
 sky130_fd_sc_hd__o311a_1 _20443_ (.A1(net3858),
    .A2(_11202_),
    .A3(_11204_),
    .B1(_11209_),
    .C1(net3856),
    .X(_11210_));
 sky130_fd_sc_hd__nand2_4 _20444_ (.A(net3669),
    .B(net3862),
    .Y(_11211_));
 sky130_fd_sc_hd__nand2_4 _20445_ (.A(net3863),
    .B(net3859),
    .Y(_11212_));
 sky130_fd_sc_hd__nand2_1 _20446_ (.A(_11211_),
    .B(_11212_),
    .Y(_11213_));
 sky130_fd_sc_hd__nor2_2 _20447_ (.A(_11140_),
    .B(_11122_),
    .Y(_11214_));
 sky130_fd_sc_hd__nor2_2 _20448_ (.A(_12257_[0]),
    .B(_11076_),
    .Y(_11215_));
 sky130_fd_sc_hd__nand2_2 _20449_ (.A(net3861),
    .B(_11215_),
    .Y(_11216_));
 sky130_fd_sc_hd__nand2_1 _20450_ (.A(net3667),
    .B(_11216_),
    .Y(_11217_));
 sky130_fd_sc_hd__a221oi_1 _20451_ (.A1(_12266_[0]),
    .A2(_11176_),
    .B1(_11213_),
    .B2(_12256_[0]),
    .C1(_11217_),
    .Y(_11218_));
 sky130_fd_sc_hd__nand2_8 _20452_ (.A(_11140_),
    .B(net3855),
    .Y(_11219_));
 sky130_fd_sc_hd__inv_4 _20453_ (.A(_12257_[0]),
    .Y(_11220_));
 sky130_fd_sc_hd__nand2_8 _20454_ (.A(_11220_),
    .B(net3858),
    .Y(_11221_));
 sky130_fd_sc_hd__nand2_4 _20455_ (.A(_12266_[0]),
    .B(net3862),
    .Y(_11222_));
 sky130_fd_sc_hd__a21oi_1 _20456_ (.A1(_11221_),
    .A2(_11222_),
    .B1(net3668),
    .Y(_11223_));
 sky130_fd_sc_hd__nand2_1 _20457_ (.A(_12256_[0]),
    .B(net3862),
    .Y(_11224_));
 sky130_fd_sc_hd__nand2_4 _20458_ (.A(_12270_[0]),
    .B(net3860),
    .Y(_11225_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_386 ();
 sky130_fd_sc_hd__a21oi_1 _20460_ (.A1(_11224_),
    .A2(_11225_),
    .B1(net3863),
    .Y(_11227_));
 sky130_fd_sc_hd__xnor2_4 _20461_ (.A(\u0.w[1][14] ),
    .B(_11086_),
    .Y(_11228_));
 sky130_fd_sc_hd__nor2_4 _20462_ (.A(_11228_),
    .B(_11092_),
    .Y(_11229_));
 sky130_fd_sc_hd__o31ai_1 _20463_ (.A1(_11219_),
    .A2(_11223_),
    .A3(_11227_),
    .B1(_11229_),
    .Y(_11230_));
 sky130_fd_sc_hd__nor2_4 _20464_ (.A(net3866),
    .B(net3858),
    .Y(_11231_));
 sky130_fd_sc_hd__o211ai_1 _20465_ (.A1(_12266_[0]),
    .A2(net3858),
    .B1(_11221_),
    .C1(net3670),
    .Y(_11232_));
 sky130_fd_sc_hd__o311ai_0 _20466_ (.A1(net3670),
    .A2(_11231_),
    .A3(_11105_),
    .B1(_11232_),
    .C1(net3855),
    .Y(_11233_));
 sky130_fd_sc_hd__nor2_1 _20467_ (.A(_12263_[0]),
    .B(net3859),
    .Y(_11234_));
 sky130_fd_sc_hd__o21ai_0 _20468_ (.A1(net3581),
    .A2(_11190_),
    .B1(net3864),
    .Y(_11235_));
 sky130_fd_sc_hd__a21oi_1 _20469_ (.A1(_12256_[0]),
    .A2(_11176_),
    .B1(net3855),
    .Y(_11236_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_385 ();
 sky130_fd_sc_hd__a21oi_1 _20471_ (.A1(_11235_),
    .A2(_11236_),
    .B1(net3852),
    .Y(_11238_));
 sky130_fd_sc_hd__nand2_2 _20472_ (.A(_12268_[0]),
    .B(net3859),
    .Y(_11239_));
 sky130_fd_sc_hd__a21oi_1 _20473_ (.A1(_11148_),
    .A2(_11239_),
    .B1(net3855),
    .Y(_11240_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_384 ();
 sky130_fd_sc_hd__nor2_4 _20475_ (.A(net3857),
    .B(net3859),
    .Y(_11241_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_383 ();
 sky130_fd_sc_hd__nor3_1 _20477_ (.A(_12263_[0]),
    .B(net3863),
    .C(net3862),
    .Y(_11243_));
 sky130_fd_sc_hd__a21oi_1 _20478_ (.A1(net3866),
    .A2(_11241_),
    .B1(_11243_),
    .Y(_11244_));
 sky130_fd_sc_hd__o21ai_0 _20479_ (.A1(net3670),
    .A2(_11240_),
    .B1(_11244_),
    .Y(_11245_));
 sky130_fd_sc_hd__a21oi_1 _20480_ (.A1(_11241_),
    .A2(_11127_),
    .B1(net3854),
    .Y(_11246_));
 sky130_fd_sc_hd__a22oi_1 _20481_ (.A1(_11233_),
    .A2(_11238_),
    .B1(_11245_),
    .B2(_11246_),
    .Y(_11247_));
 sky130_fd_sc_hd__nand2_8 _20482_ (.A(_11228_),
    .B(_11092_),
    .Y(_11248_));
 sky130_fd_sc_hd__o32ai_1 _20483_ (.A1(_11210_),
    .A2(_11218_),
    .A3(_11230_),
    .B1(_11247_),
    .B2(_11248_),
    .Y(_11249_));
 sky130_fd_sc_hd__a311oi_2 _20484_ (.A1(_11093_),
    .A2(_11145_),
    .A3(_11163_),
    .B1(_11198_),
    .C1(_11249_),
    .Y(_00104_));
 sky130_fd_sc_hd__nor2_4 _20485_ (.A(_12261_[0]),
    .B(net3858),
    .Y(_11250_));
 sky130_fd_sc_hd__nor2_4 _20486_ (.A(net3868),
    .B(net3862),
    .Y(_11251_));
 sky130_fd_sc_hd__o21ai_0 _20487_ (.A1(_11250_),
    .A2(_11251_),
    .B1(net3668),
    .Y(_11252_));
 sky130_fd_sc_hd__nor2_2 _20488_ (.A(net3866),
    .B(net3862),
    .Y(_11253_));
 sky130_fd_sc_hd__a21oi_1 _20489_ (.A1(net3868),
    .A2(_11253_),
    .B1(_11219_),
    .Y(_11254_));
 sky130_fd_sc_hd__a21oi_1 _20490_ (.A1(_11252_),
    .A2(_11254_),
    .B1(_11164_),
    .Y(_11255_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_382 ();
 sky130_fd_sc_hd__nor2_1 _20492_ (.A(_12263_[0]),
    .B(net3863),
    .Y(_11257_));
 sky130_fd_sc_hd__nor2_1 _20493_ (.A(net3868),
    .B(net3668),
    .Y(_11258_));
 sky130_fd_sc_hd__nor3_1 _20494_ (.A(net3862),
    .B(net3580),
    .C(_11258_),
    .Y(_11259_));
 sky130_fd_sc_hd__o21ai_0 _20495_ (.A1(_12286_[0]),
    .A2(net3858),
    .B1(_11122_),
    .Y(_11260_));
 sky130_fd_sc_hd__nand2_2 _20496_ (.A(net3631),
    .B(_11076_),
    .Y(_11261_));
 sky130_fd_sc_hd__nand2_1 _20497_ (.A(net3594),
    .B(net3863),
    .Y(_11262_));
 sky130_fd_sc_hd__a21oi_1 _20498_ (.A1(_11261_),
    .A2(_11262_),
    .B1(net3858),
    .Y(_11263_));
 sky130_fd_sc_hd__o22ai_1 _20499_ (.A1(_11259_),
    .A2(_11260_),
    .B1(_11263_),
    .B2(_11167_),
    .Y(_11264_));
 sky130_fd_sc_hd__nor2_4 _20500_ (.A(_12257_[0]),
    .B(net3859),
    .Y(_11265_));
 sky130_fd_sc_hd__nor2_2 _20501_ (.A(_12263_[0]),
    .B(net3862),
    .Y(_11266_));
 sky130_fd_sc_hd__nor3_1 _20502_ (.A(net3669),
    .B(_11265_),
    .C(_11266_),
    .Y(_11267_));
 sky130_fd_sc_hd__nand2_8 _20503_ (.A(net3853),
    .B(_11122_),
    .Y(_11268_));
 sky130_fd_sc_hd__a311oi_1 _20504_ (.A1(net3669),
    .A2(net3610),
    .A3(_11115_),
    .B1(_11267_),
    .C1(_11268_),
    .Y(_11269_));
 sky130_fd_sc_hd__a21oi_1 _20505_ (.A1(net3852),
    .A2(_11264_),
    .B1(_11269_),
    .Y(_11270_));
 sky130_fd_sc_hd__nand2_1 _20506_ (.A(_11255_),
    .B(_11270_),
    .Y(_11271_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_381 ();
 sky130_fd_sc_hd__nor2_4 _20508_ (.A(net3670),
    .B(net3861),
    .Y(_11273_));
 sky130_fd_sc_hd__nor2_4 _20509_ (.A(_11188_),
    .B(_11273_),
    .Y(_11274_));
 sky130_fd_sc_hd__a22oi_1 _20510_ (.A1(net3868),
    .A2(_11231_),
    .B1(_11176_),
    .B2(_12257_[0]),
    .Y(_11275_));
 sky130_fd_sc_hd__o21ai_0 _20511_ (.A1(net3671),
    .A2(_11274_),
    .B1(_11275_),
    .Y(_11276_));
 sky130_fd_sc_hd__nand2_4 _20512_ (.A(_12256_[0]),
    .B(net3858),
    .Y(_11277_));
 sky130_fd_sc_hd__nand3_2 _20513_ (.A(net3863),
    .B(_11148_),
    .C(_11277_),
    .Y(_11278_));
 sky130_fd_sc_hd__nand2_8 _20514_ (.A(net3852),
    .B(_11122_),
    .Y(_11279_));
 sky130_fd_sc_hd__nand2_2 _20515_ (.A(_12263_[0]),
    .B(net3862),
    .Y(_11280_));
 sky130_fd_sc_hd__a21oi_1 _20516_ (.A1(_11280_),
    .A2(net3610),
    .B1(net3863),
    .Y(_11281_));
 sky130_fd_sc_hd__nor2_1 _20517_ (.A(_11279_),
    .B(_11281_),
    .Y(_11282_));
 sky130_fd_sc_hd__a22oi_1 _20518_ (.A1(net3667),
    .A2(_11276_),
    .B1(_11278_),
    .B2(_11282_),
    .Y(_11283_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_380 ();
 sky130_fd_sc_hd__nor2_4 _20520_ (.A(_11194_),
    .B(net3856),
    .Y(_11285_));
 sky130_fd_sc_hd__and2_4 _20521_ (.A(_12263_[0]),
    .B(net3858),
    .X(_11286_));
 sky130_fd_sc_hd__o21ai_0 _20522_ (.A1(_11265_),
    .A2(_11286_),
    .B1(net3863),
    .Y(_11287_));
 sky130_fd_sc_hd__o211ai_1 _20523_ (.A1(_12270_[0]),
    .A2(_11211_),
    .B1(_11285_),
    .C1(_11287_),
    .Y(_11288_));
 sky130_fd_sc_hd__nor2_4 _20524_ (.A(_11194_),
    .B(net3855),
    .Y(_11289_));
 sky130_fd_sc_hd__nor2_1 _20525_ (.A(_12270_[0]),
    .B(net3862),
    .Y(_11290_));
 sky130_fd_sc_hd__nor2_1 _20526_ (.A(net3868),
    .B(net3858),
    .Y(_11291_));
 sky130_fd_sc_hd__o21ai_0 _20527_ (.A1(_11290_),
    .A2(net3666),
    .B1(net3863),
    .Y(_11292_));
 sky130_fd_sc_hd__nand2_1 _20528_ (.A(net3594),
    .B(_11188_),
    .Y(_11293_));
 sky130_fd_sc_hd__a31oi_1 _20529_ (.A1(_11289_),
    .A2(_11292_),
    .A3(_11293_),
    .B1(_11248_),
    .Y(_11294_));
 sky130_fd_sc_hd__nand3_1 _20530_ (.A(_11283_),
    .B(_11288_),
    .C(_11294_),
    .Y(_11295_));
 sky130_fd_sc_hd__and2_0 _20531_ (.A(_12270_[0]),
    .B(net3859),
    .X(_11296_));
 sky130_fd_sc_hd__o21ai_0 _20532_ (.A1(_11296_),
    .A2(_11265_),
    .B1(net3863),
    .Y(_11297_));
 sky130_fd_sc_hd__nand2_1 _20533_ (.A(net3866),
    .B(_11176_),
    .Y(_11298_));
 sky130_fd_sc_hd__nor2_4 _20534_ (.A(net3854),
    .B(net3855),
    .Y(_11299_));
 sky130_fd_sc_hd__nand2_2 _20535_ (.A(_12270_[0]),
    .B(net3862),
    .Y(_11300_));
 sky130_fd_sc_hd__o21ai_1 _20536_ (.A1(_12258_[0]),
    .A2(net3862),
    .B1(_11300_),
    .Y(_11301_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_379 ();
 sky130_fd_sc_hd__and2_4 _20538_ (.A(_12272_[0]),
    .B(net3858),
    .X(_11303_));
 sky130_fd_sc_hd__nor3_1 _20539_ (.A(net3669),
    .B(_11265_),
    .C(_11303_),
    .Y(_11304_));
 sky130_fd_sc_hd__a21oi_1 _20540_ (.A1(net3669),
    .A2(_11301_),
    .B1(_11304_),
    .Y(_11305_));
 sky130_fd_sc_hd__a32o_1 _20541_ (.A1(net3667),
    .A2(_11297_),
    .A3(_11298_),
    .B1(_11299_),
    .B2(_11305_),
    .X(_11306_));
 sky130_fd_sc_hd__and3_4 _20542_ (.A(net3669),
    .B(_11148_),
    .C(net3610),
    .X(_11307_));
 sky130_fd_sc_hd__a21oi_1 _20543_ (.A1(_12256_[0]),
    .A2(net3862),
    .B1(_11190_),
    .Y(_11308_));
 sky130_fd_sc_hd__o21ai_0 _20544_ (.A1(net3669),
    .A2(_11308_),
    .B1(_11289_),
    .Y(_11309_));
 sky130_fd_sc_hd__nor2_1 _20545_ (.A(net3581),
    .B(_11253_),
    .Y(_11310_));
 sky130_fd_sc_hd__nor2_1 _20546_ (.A(net3670),
    .B(_11310_),
    .Y(_11311_));
 sky130_fd_sc_hd__nor2_1 _20547_ (.A(_12256_[0]),
    .B(net3862),
    .Y(_11312_));
 sky130_fd_sc_hd__o31ai_1 _20548_ (.A1(net3863),
    .A2(_11312_),
    .A3(net3666),
    .B1(_11285_),
    .Y(_11313_));
 sky130_fd_sc_hd__o22ai_1 _20549_ (.A1(_11307_),
    .A2(_11309_),
    .B1(_11311_),
    .B2(_11313_),
    .Y(_11314_));
 sky130_fd_sc_hd__o21ai_0 _20550_ (.A1(_11306_),
    .A2(_11314_),
    .B1(_11093_),
    .Y(_11315_));
 sky130_fd_sc_hd__nand2_4 _20551_ (.A(net3672),
    .B(net3860),
    .Y(_11316_));
 sky130_fd_sc_hd__nand2_1 _20552_ (.A(net3868),
    .B(net3862),
    .Y(_11317_));
 sky130_fd_sc_hd__a21oi_1 _20553_ (.A1(_11316_),
    .A2(_11317_),
    .B1(net3863),
    .Y(_11318_));
 sky130_fd_sc_hd__nor3_1 _20554_ (.A(_11279_),
    .B(_11311_),
    .C(_11318_),
    .Y(_11319_));
 sky130_fd_sc_hd__nand2_2 _20555_ (.A(_12261_[0]),
    .B(net3862),
    .Y(_11320_));
 sky130_fd_sc_hd__a21oi_1 _20556_ (.A1(_11320_),
    .A2(_11277_),
    .B1(net3863),
    .Y(_11321_));
 sky130_fd_sc_hd__nand2_4 _20557_ (.A(net3866),
    .B(net3858),
    .Y(_11322_));
 sky130_fd_sc_hd__a21oi_1 _20558_ (.A1(_11322_),
    .A2(_11300_),
    .B1(net3669),
    .Y(_11323_));
 sky130_fd_sc_hd__mux2i_1 _20559_ (.A0(_12266_[0]),
    .A1(_12270_[0]),
    .S(net3864),
    .Y(_11324_));
 sky130_fd_sc_hd__nor3_1 _20560_ (.A(_12282_[0]),
    .B(net3853),
    .C(net3858),
    .Y(_11325_));
 sky130_fd_sc_hd__a21oi_1 _20561_ (.A1(net3858),
    .A2(_11324_),
    .B1(_11325_),
    .Y(_11326_));
 sky130_fd_sc_hd__o32ai_1 _20562_ (.A1(_11268_),
    .A2(_11321_),
    .A3(_11323_),
    .B1(_11326_),
    .B2(net3857),
    .Y(_11327_));
 sky130_fd_sc_hd__o21ai_0 _20563_ (.A1(_11319_),
    .A2(_11327_),
    .B1(_11229_),
    .Y(_11328_));
 sky130_fd_sc_hd__nand4_1 _20564_ (.A(_11271_),
    .B(_11295_),
    .C(_11315_),
    .D(_11328_),
    .Y(_00105_));
 sky130_fd_sc_hd__o21ai_0 _20565_ (.A1(net3672),
    .A2(net3862),
    .B1(_11222_),
    .Y(_11329_));
 sky130_fd_sc_hd__o21ai_0 _20566_ (.A1(_12256_[0]),
    .A2(net3862),
    .B1(_11148_),
    .Y(_11330_));
 sky130_fd_sc_hd__nand2_1 _20567_ (.A(_11076_),
    .B(_11330_),
    .Y(_11331_));
 sky130_fd_sc_hd__o21ai_0 _20568_ (.A1(net3668),
    .A2(_11329_),
    .B1(_11331_),
    .Y(_11332_));
 sky130_fd_sc_hd__nor2_4 _20569_ (.A(net3672),
    .B(net3858),
    .Y(_11333_));
 sky130_fd_sc_hd__o21ai_1 _20570_ (.A1(net3672),
    .A2(net3863),
    .B1(_11316_),
    .Y(_11334_));
 sky130_fd_sc_hd__a222oi_1 _20571_ (.A1(_11170_),
    .A2(_11258_),
    .B1(_11333_),
    .B2(_11199_),
    .C1(_11334_),
    .C2(net3631),
    .Y(_11335_));
 sky130_fd_sc_hd__o22ai_1 _20572_ (.A1(_11279_),
    .A2(_11332_),
    .B1(_11335_),
    .B2(_11268_),
    .Y(_11336_));
 sky130_fd_sc_hd__nor2_1 _20573_ (.A(net3868),
    .B(_11140_),
    .Y(_11337_));
 sky130_fd_sc_hd__a21oi_1 _20574_ (.A1(_12257_[0]),
    .A2(_11140_),
    .B1(_11337_),
    .Y(_11338_));
 sky130_fd_sc_hd__nor3_1 _20575_ (.A(net3672),
    .B(net3866),
    .C(_11140_),
    .Y(_11339_));
 sky130_fd_sc_hd__a31oi_1 _20576_ (.A1(_11165_),
    .A2(net3863),
    .A3(_11140_),
    .B1(_11339_),
    .Y(_11340_));
 sky130_fd_sc_hd__o21ai_0 _20577_ (.A1(net3863),
    .A2(_11338_),
    .B1(_11340_),
    .Y(_11341_));
 sky130_fd_sc_hd__nor2_1 _20578_ (.A(_12279_[0]),
    .B(_11194_),
    .Y(_11342_));
 sky130_fd_sc_hd__a211oi_1 _20579_ (.A1(_12282_[0]),
    .A2(_11194_),
    .B1(net3862),
    .C1(_11342_),
    .Y(_11343_));
 sky130_fd_sc_hd__a211oi_1 _20580_ (.A1(net3862),
    .A2(_11341_),
    .B1(_11343_),
    .C1(net3856),
    .Y(_11344_));
 sky130_fd_sc_hd__nor3_1 _20581_ (.A(_11248_),
    .B(_11336_),
    .C(_11344_),
    .Y(_11345_));
 sky130_fd_sc_hd__a221oi_1 _20582_ (.A1(_12263_[0]),
    .A2(_11188_),
    .B1(_11330_),
    .B2(net3863),
    .C1(_11219_),
    .Y(_11346_));
 sky130_fd_sc_hd__nand2_1 _20583_ (.A(_12277_[0]),
    .B(net3861),
    .Y(_11347_));
 sky130_fd_sc_hd__nand2_2 _20584_ (.A(_12261_[0]),
    .B(_11176_),
    .Y(_11348_));
 sky130_fd_sc_hd__nand2_8 _20585_ (.A(_11194_),
    .B(net3855),
    .Y(_11349_));
 sky130_fd_sc_hd__a21oi_1 _20586_ (.A1(_11347_),
    .A2(_11348_),
    .B1(_11349_),
    .Y(_11350_));
 sky130_fd_sc_hd__nor2_4 _20587_ (.A(_12258_[0]),
    .B(_12263_[0]),
    .Y(_11351_));
 sky130_fd_sc_hd__o221ai_1 _20588_ (.A1(_12270_[0]),
    .A2(_11274_),
    .B1(_11351_),
    .B2(_11156_),
    .C1(_11183_),
    .Y(_11352_));
 sky130_fd_sc_hd__nand2_2 _20589_ (.A(_11065_),
    .B(net3863),
    .Y(_11353_));
 sky130_fd_sc_hd__a21oi_1 _20590_ (.A1(_12261_[0]),
    .A2(_11076_),
    .B1(net3858),
    .Y(_11354_));
 sky130_fd_sc_hd__a22oi_1 _20591_ (.A1(_12288_[0]),
    .A2(net3858),
    .B1(_11353_),
    .B2(_11354_),
    .Y(_11355_));
 sky130_fd_sc_hd__o21ai_0 _20592_ (.A1(_11140_),
    .A2(_11355_),
    .B1(net3856),
    .Y(_11356_));
 sky130_fd_sc_hd__a21oi_1 _20593_ (.A1(net3854),
    .A2(_11352_),
    .B1(_11356_),
    .Y(_11357_));
 sky130_fd_sc_hd__nor2_2 _20594_ (.A(_12272_[0]),
    .B(net3862),
    .Y(_11358_));
 sky130_fd_sc_hd__or3_1 _20595_ (.A(net3863),
    .B(_11234_),
    .C(_11358_),
    .X(_11359_));
 sky130_fd_sc_hd__o211ai_1 _20596_ (.A1(_12268_[0]),
    .A2(net3862),
    .B1(_11115_),
    .C1(net3864),
    .Y(_11360_));
 sky130_fd_sc_hd__a21oi_1 _20597_ (.A1(_11359_),
    .A2(_11360_),
    .B1(_11279_),
    .Y(_11361_));
 sky130_fd_sc_hd__or3_1 _20598_ (.A(net3863),
    .B(_11291_),
    .C(_11358_),
    .X(_11362_));
 sky130_fd_sc_hd__nor2_4 _20599_ (.A(_12268_[0]),
    .B(net3859),
    .Y(_11363_));
 sky130_fd_sc_hd__or3_1 _20600_ (.A(net3670),
    .B(_11159_),
    .C(_11363_),
    .X(_11364_));
 sky130_fd_sc_hd__a21oi_1 _20601_ (.A1(_11362_),
    .A2(_11364_),
    .B1(_11268_),
    .Y(_11365_));
 sky130_fd_sc_hd__and3_1 _20602_ (.A(net3863),
    .B(_11148_),
    .C(_11149_),
    .X(_11366_));
 sky130_fd_sc_hd__nor3b_1 _20603_ (.A(_11265_),
    .B(net3863),
    .C_N(_11239_),
    .Y(_11367_));
 sky130_fd_sc_hd__nand2_4 _20604_ (.A(_11065_),
    .B(net3861),
    .Y(_11368_));
 sky130_fd_sc_hd__a311o_1 _20605_ (.A1(net3863),
    .A2(_11239_),
    .A3(_11368_),
    .B1(_11257_),
    .C1(_11349_),
    .X(_11369_));
 sky130_fd_sc_hd__o31ai_1 _20606_ (.A1(_11219_),
    .A2(_11366_),
    .A3(_11367_),
    .B1(_11369_),
    .Y(_11370_));
 sky130_fd_sc_hd__o31ai_2 _20607_ (.A1(_11361_),
    .A2(_11365_),
    .A3(_11370_),
    .B1(_11093_),
    .Y(_11371_));
 sky130_fd_sc_hd__o41ai_1 _20608_ (.A1(_11164_),
    .A2(_11346_),
    .A3(_11350_),
    .A4(_11357_),
    .B1(_11371_),
    .Y(_11372_));
 sky130_fd_sc_hd__a21oi_1 _20609_ (.A1(net3861),
    .A2(_11166_),
    .B1(_11122_),
    .Y(_11373_));
 sky130_fd_sc_hd__nand3_1 _20610_ (.A(net3858),
    .B(_11261_),
    .C(_11353_),
    .Y(_11374_));
 sky130_fd_sc_hd__o21ai_0 _20611_ (.A1(_11250_),
    .A2(_11303_),
    .B1(_11076_),
    .Y(_11375_));
 sky130_fd_sc_hd__o311ai_1 _20612_ (.A1(net3669),
    .A2(_11266_),
    .A3(net3666),
    .B1(_11375_),
    .C1(net3852),
    .Y(_11376_));
 sky130_fd_sc_hd__nor2_1 _20613_ (.A(net3594),
    .B(_11156_),
    .Y(_11377_));
 sky130_fd_sc_hd__a21oi_1 _20614_ (.A1(_11114_),
    .A2(_11300_),
    .B1(net3863),
    .Y(_11378_));
 sky130_fd_sc_hd__o31ai_1 _20615_ (.A1(_11194_),
    .A2(_11377_),
    .A3(_11378_),
    .B1(net3855),
    .Y(_11379_));
 sky130_fd_sc_hd__a32oi_1 _20616_ (.A1(_11194_),
    .A2(_11373_),
    .A3(_11374_),
    .B1(_11376_),
    .B2(_11379_),
    .Y(_11380_));
 sky130_fd_sc_hd__nand3_1 _20617_ (.A(net3863),
    .B(_11221_),
    .C(_11115_),
    .Y(_11381_));
 sky130_fd_sc_hd__o311ai_0 _20618_ (.A1(net3863),
    .A2(_11184_),
    .A3(_11251_),
    .B1(_11381_),
    .C1(net3853),
    .Y(_11382_));
 sky130_fd_sc_hd__nor3_1 _20619_ (.A(_11122_),
    .B(_11377_),
    .C(_11378_),
    .Y(_11383_));
 sky130_fd_sc_hd__o21ai_0 _20620_ (.A1(_11382_),
    .A2(_11383_),
    .B1(_11229_),
    .Y(_11384_));
 sky130_fd_sc_hd__nor2_1 _20621_ (.A(_11380_),
    .B(_11384_),
    .Y(_11385_));
 sky130_fd_sc_hd__or3_4 _20622_ (.A(_11345_),
    .B(_11372_),
    .C(_11385_),
    .X(_00106_));
 sky130_fd_sc_hd__nor2_2 _20623_ (.A(_11071_),
    .B(net3858),
    .Y(_11386_));
 sky130_fd_sc_hd__nand2_2 _20624_ (.A(net3672),
    .B(_11386_),
    .Y(_11387_));
 sky130_fd_sc_hd__nand2_1 _20625_ (.A(net3858),
    .B(_11215_),
    .Y(_11388_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_378 ();
 sky130_fd_sc_hd__o21ai_0 _20627_ (.A1(_11231_),
    .A2(_11182_),
    .B1(_11076_),
    .Y(_11390_));
 sky130_fd_sc_hd__nand4_1 _20628_ (.A(_11289_),
    .B(_11387_),
    .C(_11388_),
    .D(_11390_),
    .Y(_11391_));
 sky130_fd_sc_hd__a21oi_1 _20629_ (.A1(_11221_),
    .A2(_11320_),
    .B1(net3864),
    .Y(_11392_));
 sky130_fd_sc_hd__a21oi_1 _20630_ (.A1(_11222_),
    .A2(_11225_),
    .B1(net3670),
    .Y(_11393_));
 sky130_fd_sc_hd__nor2_4 _20631_ (.A(_11220_),
    .B(net3861),
    .Y(_11394_));
 sky130_fd_sc_hd__o211ai_1 _20632_ (.A1(_12268_[0]),
    .A2(net3862),
    .B1(_11147_),
    .C1(net3670),
    .Y(_11395_));
 sky130_fd_sc_hd__o311a_1 _20633_ (.A1(net3670),
    .A2(_11394_),
    .A3(_11333_),
    .B1(_11395_),
    .C1(net3852),
    .X(_11396_));
 sky130_fd_sc_hd__o32ai_1 _20634_ (.A1(net3852),
    .A2(_11392_),
    .A3(_11393_),
    .B1(_11396_),
    .B2(net3855),
    .Y(_11397_));
 sky130_fd_sc_hd__o21ai_0 _20635_ (.A1(net3868),
    .A2(net3671),
    .B1(_11199_),
    .Y(_11398_));
 sky130_fd_sc_hd__a221oi_1 _20636_ (.A1(_12261_[0]),
    .A2(_11188_),
    .B1(_11398_),
    .B2(net3858),
    .C1(_11349_),
    .Y(_11399_));
 sky130_fd_sc_hd__a211oi_1 _20637_ (.A1(_11391_),
    .A2(_11397_),
    .B1(_11399_),
    .C1(_11087_),
    .Y(_11400_));
 sky130_fd_sc_hd__or3_1 _20638_ (.A(net3863),
    .B(_11105_),
    .C(net3581),
    .X(_11401_));
 sky130_fd_sc_hd__o31ai_1 _20639_ (.A1(net3670),
    .A2(_11394_),
    .A3(_11112_),
    .B1(_11401_),
    .Y(_11402_));
 sky130_fd_sc_hd__nor2_1 _20640_ (.A(_12256_[0]),
    .B(net3858),
    .Y(_11403_));
 sky130_fd_sc_hd__nor3_1 _20641_ (.A(_11076_),
    .B(_11182_),
    .C(_11403_),
    .Y(_11404_));
 sky130_fd_sc_hd__nor3_1 _20642_ (.A(net3863),
    .B(_11265_),
    .C(_11253_),
    .Y(_11405_));
 sky130_fd_sc_hd__o211ai_1 _20643_ (.A1(_11404_),
    .A2(_11405_),
    .B1(_11087_),
    .C1(_11289_),
    .Y(_11406_));
 sky130_fd_sc_hd__o311ai_0 _20644_ (.A1(_11228_),
    .A2(_11219_),
    .A3(_11402_),
    .B1(_11406_),
    .C1(_11092_),
    .Y(_11407_));
 sky130_fd_sc_hd__a211oi_1 _20645_ (.A1(net3866),
    .A2(net3855),
    .B1(net3863),
    .C1(net3868),
    .Y(_11408_));
 sky130_fd_sc_hd__a31oi_1 _20646_ (.A1(net3868),
    .A2(net3855),
    .A3(_11199_),
    .B1(_11408_),
    .Y(_11409_));
 sky130_fd_sc_hd__nand3_1 _20647_ (.A(net3672),
    .B(_11076_),
    .C(net3855),
    .Y(_11410_));
 sky130_fd_sc_hd__o21ai_0 _20648_ (.A1(_11076_),
    .A2(net3855),
    .B1(_11410_),
    .Y(_11411_));
 sky130_fd_sc_hd__a21oi_1 _20649_ (.A1(_11076_),
    .A2(net3855),
    .B1(_11220_),
    .Y(_11412_));
 sky130_fd_sc_hd__o21ai_0 _20650_ (.A1(_11411_),
    .A2(_11412_),
    .B1(net3861),
    .Y(_11413_));
 sky130_fd_sc_hd__o21ai_0 _20651_ (.A1(net3861),
    .A2(_11409_),
    .B1(_11413_),
    .Y(_11414_));
 sky130_fd_sc_hd__nor2_1 _20652_ (.A(net3855),
    .B(_11199_),
    .Y(_11415_));
 sky130_fd_sc_hd__nor4_1 _20653_ (.A(_11140_),
    .B(_11164_),
    .C(_11414_),
    .D(_11415_),
    .Y(_11416_));
 sky130_fd_sc_hd__nor3_1 _20654_ (.A(net3866),
    .B(net3852),
    .C(net3860),
    .Y(_11417_));
 sky130_fd_sc_hd__nor2_4 _20655_ (.A(net3631),
    .B(net3862),
    .Y(_11418_));
 sky130_fd_sc_hd__nor2_4 _20656_ (.A(_11418_),
    .B(_11363_),
    .Y(_11419_));
 sky130_fd_sc_hd__a21oi_1 _20657_ (.A1(net3852),
    .A2(_11159_),
    .B1(net3670),
    .Y(_11420_));
 sky130_fd_sc_hd__o21ai_0 _20658_ (.A1(net3852),
    .A2(_11419_),
    .B1(_11420_),
    .Y(_11421_));
 sky130_fd_sc_hd__o311ai_0 _20659_ (.A1(net3864),
    .A2(_11358_),
    .A3(_11417_),
    .B1(_11421_),
    .C1(net3857),
    .Y(_11422_));
 sky130_fd_sc_hd__o21ai_0 _20660_ (.A1(net3670),
    .A2(_11105_),
    .B1(_11071_),
    .Y(_11423_));
 sky130_fd_sc_hd__a21oi_1 _20661_ (.A1(net3672),
    .A2(_11176_),
    .B1(_11219_),
    .Y(_11424_));
 sky130_fd_sc_hd__nand3b_1 _20662_ (.A_N(_11169_),
    .B(_11423_),
    .C(_11424_),
    .Y(_11425_));
 sky130_fd_sc_hd__nand2_2 _20663_ (.A(_12268_[0]),
    .B(net3861),
    .Y(_11426_));
 sky130_fd_sc_hd__nor3b_4 _20664_ (.A(net3863),
    .B(_11182_),
    .C_N(_11426_),
    .Y(_11427_));
 sky130_fd_sc_hd__nand2_4 _20665_ (.A(net3862),
    .B(_11351_),
    .Y(_11428_));
 sky130_fd_sc_hd__a21oi_1 _20666_ (.A1(_11225_),
    .A2(_11428_),
    .B1(net3670),
    .Y(_11429_));
 sky130_fd_sc_hd__o21ai_0 _20667_ (.A1(_11427_),
    .A2(_11429_),
    .B1(net3667),
    .Y(_11430_));
 sky130_fd_sc_hd__a22oi_1 _20668_ (.A1(net3671),
    .A2(_11273_),
    .B1(_11274_),
    .B2(_12268_[0]),
    .Y(_11431_));
 sky130_fd_sc_hd__nor4_1 _20669_ (.A(_12257_[0]),
    .B(_11076_),
    .C(_11194_),
    .D(_11184_),
    .Y(_11432_));
 sky130_fd_sc_hd__nand3_1 _20670_ (.A(_11076_),
    .B(_11194_),
    .C(_11148_),
    .Y(_11433_));
 sky130_fd_sc_hd__a21oi_1 _20671_ (.A1(_12266_[0]),
    .A2(net3858),
    .B1(_11433_),
    .Y(_11434_));
 sky130_fd_sc_hd__nand2_1 _20672_ (.A(_12258_[0]),
    .B(net3861),
    .Y(_11435_));
 sky130_fd_sc_hd__nand3_1 _20673_ (.A(net3868),
    .B(_11194_),
    .C(net3858),
    .Y(_11436_));
 sky130_fd_sc_hd__a21oi_1 _20674_ (.A1(_11435_),
    .A2(_11436_),
    .B1(_11076_),
    .Y(_11437_));
 sky130_fd_sc_hd__nor4_1 _20675_ (.A(net3855),
    .B(_11432_),
    .C(_11434_),
    .D(_11437_),
    .Y(_11438_));
 sky130_fd_sc_hd__nor3_2 _20676_ (.A(net3864),
    .B(_11159_),
    .C(_11112_),
    .Y(_11439_));
 sky130_fd_sc_hd__a311oi_1 _20677_ (.A1(net3864),
    .A2(_11221_),
    .A3(_11428_),
    .B1(_11439_),
    .C1(_11349_),
    .Y(_11440_));
 sky130_fd_sc_hd__a2111oi_0 _20678_ (.A1(_11285_),
    .A2(_11431_),
    .B1(_11438_),
    .C1(_11440_),
    .D1(_11228_),
    .Y(_11441_));
 sky130_fd_sc_hd__a41oi_1 _20679_ (.A1(_11228_),
    .A2(_11422_),
    .A3(_11425_),
    .A4(_11430_),
    .B1(_11441_),
    .Y(_11442_));
 sky130_fd_sc_hd__o32ai_1 _20680_ (.A1(_11400_),
    .A2(_11407_),
    .A3(_11416_),
    .B1(_11442_),
    .B2(_11092_),
    .Y(_00107_));
 sky130_fd_sc_hd__nor2_1 _20681_ (.A(net3863),
    .B(net3855),
    .Y(_11443_));
 sky130_fd_sc_hd__nor2_1 _20682_ (.A(_12257_[0]),
    .B(net3863),
    .Y(_11444_));
 sky130_fd_sc_hd__and2_0 _20683_ (.A(_12263_[0]),
    .B(net3863),
    .X(_11445_));
 sky130_fd_sc_hd__o21ai_0 _20684_ (.A1(_11444_),
    .A2(_11445_),
    .B1(net3858),
    .Y(_11446_));
 sky130_fd_sc_hd__a221oi_1 _20685_ (.A1(_11301_),
    .A2(_11443_),
    .B1(_11446_),
    .B2(_11131_),
    .C1(net3852),
    .Y(_11447_));
 sky130_fd_sc_hd__nand3_1 _20686_ (.A(net3670),
    .B(_11316_),
    .C(_11317_),
    .Y(_11448_));
 sky130_fd_sc_hd__o211ai_1 _20687_ (.A1(_12263_[0]),
    .A2(net3859),
    .B1(_11277_),
    .C1(net3863),
    .Y(_11449_));
 sky130_fd_sc_hd__o22ai_1 _20688_ (.A1(net3671),
    .A2(_11212_),
    .B1(_11358_),
    .B2(net3863),
    .Y(_11450_));
 sky130_fd_sc_hd__o21ai_0 _20689_ (.A1(net3857),
    .A2(_11450_),
    .B1(net3852),
    .Y(_11451_));
 sky130_fd_sc_hd__a31oi_2 _20690_ (.A1(net3857),
    .A2(_11448_),
    .A3(_11449_),
    .B1(_11451_),
    .Y(_11452_));
 sky130_fd_sc_hd__a21oi_1 _20691_ (.A1(_11076_),
    .A2(_11426_),
    .B1(_11190_),
    .Y(_11453_));
 sky130_fd_sc_hd__and3_1 _20692_ (.A(_11076_),
    .B(_11277_),
    .C(_11368_),
    .X(_11454_));
 sky130_fd_sc_hd__nand2_1 _20693_ (.A(net3855),
    .B(_11199_),
    .Y(_11455_));
 sky130_fd_sc_hd__o221ai_1 _20694_ (.A1(net3855),
    .A2(_11453_),
    .B1(_11454_),
    .B2(_11455_),
    .C1(_11140_),
    .Y(_11456_));
 sky130_fd_sc_hd__o22ai_1 _20695_ (.A1(net3866),
    .A2(_11212_),
    .B1(_11115_),
    .B2(net3672),
    .Y(_11457_));
 sky130_fd_sc_hd__a211o_1 _20696_ (.A1(net3672),
    .A2(_11274_),
    .B1(_11457_),
    .C1(_11349_),
    .X(_11458_));
 sky130_fd_sc_hd__o21ai_2 _20697_ (.A1(net3868),
    .A2(net3610),
    .B1(_11299_),
    .Y(_11459_));
 sky130_fd_sc_hd__nor2_2 _20698_ (.A(net3672),
    .B(_11076_),
    .Y(_11460_));
 sky130_fd_sc_hd__a211o_1 _20699_ (.A1(_12256_[0]),
    .A2(_11188_),
    .B1(_11459_),
    .C1(_11460_),
    .X(_11461_));
 sky130_fd_sc_hd__nand4_1 _20700_ (.A(_11092_),
    .B(_11456_),
    .C(_11458_),
    .D(_11461_),
    .Y(_11462_));
 sky130_fd_sc_hd__o311ai_1 _20701_ (.A1(_11092_),
    .A2(_11447_),
    .A3(_11452_),
    .B1(_11462_),
    .C1(_11228_),
    .Y(_11463_));
 sky130_fd_sc_hd__nand2b_1 _20702_ (.A_N(_12256_[0]),
    .B(net3863),
    .Y(_11464_));
 sky130_fd_sc_hd__a21oi_1 _20703_ (.A1(_11135_),
    .A2(_11464_),
    .B1(net3858),
    .Y(_11465_));
 sky130_fd_sc_hd__nor3_1 _20704_ (.A(net3669),
    .B(_11250_),
    .C(_11286_),
    .Y(_11466_));
 sky130_fd_sc_hd__nor3_1 _20705_ (.A(net3863),
    .B(net3666),
    .C(_11303_),
    .Y(_11467_));
 sky130_fd_sc_hd__o21ai_0 _20706_ (.A1(_11466_),
    .A2(_11467_),
    .B1(_11122_),
    .Y(_11468_));
 sky130_fd_sc_hd__o21ai_0 _20707_ (.A1(_11167_),
    .A2(_11465_),
    .B1(_11468_),
    .Y(_11469_));
 sky130_fd_sc_hd__o21ai_0 _20708_ (.A1(_11418_),
    .A2(_11363_),
    .B1(net3855),
    .Y(_11470_));
 sky130_fd_sc_hd__o21ai_0 _20709_ (.A1(_11265_),
    .A2(_11266_),
    .B1(_11122_),
    .Y(_11471_));
 sky130_fd_sc_hd__nand2_1 _20710_ (.A(_12268_[0]),
    .B(_11122_),
    .Y(_11472_));
 sky130_fd_sc_hd__o21ai_0 _20711_ (.A1(_11250_),
    .A2(_11303_),
    .B1(net3855),
    .Y(_11473_));
 sky130_fd_sc_hd__a21oi_1 _20712_ (.A1(_11472_),
    .A2(_11473_),
    .B1(_11076_),
    .Y(_11474_));
 sky130_fd_sc_hd__a311oi_1 _20713_ (.A1(_11076_),
    .A2(_11470_),
    .A3(_11471_),
    .B1(_11474_),
    .C1(net3852),
    .Y(_11475_));
 sky130_fd_sc_hd__a211o_1 _20714_ (.A1(net3852),
    .A2(_11469_),
    .B1(_11475_),
    .C1(_11164_),
    .X(_11476_));
 sky130_fd_sc_hd__o21ai_0 _20715_ (.A1(_12258_[0]),
    .A2(_11212_),
    .B1(_11387_),
    .Y(_11477_));
 sky130_fd_sc_hd__a21oi_1 _20716_ (.A1(_11170_),
    .A2(_11277_),
    .B1(net3863),
    .Y(_11478_));
 sky130_fd_sc_hd__o211ai_1 _20717_ (.A1(net3858),
    .A2(_11261_),
    .B1(_11225_),
    .C1(_11140_),
    .Y(_11479_));
 sky130_fd_sc_hd__o311ai_0 _20718_ (.A1(_11140_),
    .A2(_11477_),
    .A3(_11478_),
    .B1(_11479_),
    .C1(net3855),
    .Y(_11480_));
 sky130_fd_sc_hd__nand2_1 _20719_ (.A(_12268_[0]),
    .B(_11076_),
    .Y(_11481_));
 sky130_fd_sc_hd__nand2_4 _20720_ (.A(_11165_),
    .B(net3858),
    .Y(_11482_));
 sky130_fd_sc_hd__a21oi_1 _20721_ (.A1(_11482_),
    .A2(_11368_),
    .B1(_11076_),
    .Y(_11483_));
 sky130_fd_sc_hd__o21a_1 _20722_ (.A1(_11105_),
    .A2(_11386_),
    .B1(net3863),
    .X(_11484_));
 sky130_fd_sc_hd__o22ai_1 _20723_ (.A1(_11268_),
    .A2(_11483_),
    .B1(_11484_),
    .B2(_11459_),
    .Y(_11485_));
 sky130_fd_sc_hd__o21ai_0 _20724_ (.A1(net3858),
    .A2(_11481_),
    .B1(_11485_),
    .Y(_11486_));
 sky130_fd_sc_hd__nand3_1 _20725_ (.A(_11229_),
    .B(_11480_),
    .C(_11486_),
    .Y(_11487_));
 sky130_fd_sc_hd__nand3_1 _20726_ (.A(_11463_),
    .B(_11476_),
    .C(_11487_),
    .Y(_00108_));
 sky130_fd_sc_hd__nand2_1 _20727_ (.A(net3854),
    .B(_11348_),
    .Y(_11488_));
 sky130_fd_sc_hd__o21ai_0 _20728_ (.A1(_11429_),
    .A2(_11488_),
    .B1(net3855),
    .Y(_11489_));
 sky130_fd_sc_hd__nand3b_1 _20729_ (.A_N(_11358_),
    .B(net3670),
    .C(_11222_),
    .Y(_11490_));
 sky130_fd_sc_hd__o31ai_1 _20730_ (.A1(net3670),
    .A2(_11394_),
    .A3(_11265_),
    .B1(_11490_),
    .Y(_11491_));
 sky130_fd_sc_hd__nand2_1 _20731_ (.A(_12263_[0]),
    .B(_11176_),
    .Y(_11492_));
 sky130_fd_sc_hd__o21ai_0 _20732_ (.A1(_12272_[0]),
    .A2(net3864),
    .B1(net3862),
    .Y(_11493_));
 sky130_fd_sc_hd__a31oi_1 _20733_ (.A1(net3857),
    .A2(_11492_),
    .A3(_11493_),
    .B1(net3852),
    .Y(_11494_));
 sky130_fd_sc_hd__a21o_1 _20734_ (.A1(net3852),
    .A2(_11491_),
    .B1(_11494_),
    .X(_11495_));
 sky130_fd_sc_hd__o211ai_1 _20735_ (.A1(net3670),
    .A2(_11225_),
    .B1(_11222_),
    .C1(net3667),
    .Y(_11496_));
 sky130_fd_sc_hd__nand2_1 _20736_ (.A(_11229_),
    .B(_11496_),
    .Y(_11497_));
 sky130_fd_sc_hd__a21oi_1 _20737_ (.A1(_11489_),
    .A2(_11495_),
    .B1(_11497_),
    .Y(_11498_));
 sky130_fd_sc_hd__o221ai_1 _20738_ (.A1(_12270_[0]),
    .A2(_11156_),
    .B1(_11274_),
    .B2(net3866),
    .C1(_11492_),
    .Y(_11499_));
 sky130_fd_sc_hd__o21ai_0 _20739_ (.A1(_12270_[0]),
    .A2(_11212_),
    .B1(_11490_),
    .Y(_11500_));
 sky130_fd_sc_hd__o21ai_0 _20740_ (.A1(_12261_[0]),
    .A2(net3859),
    .B1(_11239_),
    .Y(_11501_));
 sky130_fd_sc_hd__a21oi_1 _20741_ (.A1(_11148_),
    .A2(_11316_),
    .B1(net3670),
    .Y(_11502_));
 sky130_fd_sc_hd__a21oi_1 _20742_ (.A1(net3670),
    .A2(_11501_),
    .B1(_11502_),
    .Y(_11503_));
 sky130_fd_sc_hd__o2bb2ai_1 _20743_ (.A1_N(_11299_),
    .A2_N(_11500_),
    .B1(_11503_),
    .B2(_11268_),
    .Y(_11504_));
 sky130_fd_sc_hd__a22oi_1 _20744_ (.A1(net3671),
    .A2(_11212_),
    .B1(_11159_),
    .B2(net3672),
    .Y(_11505_));
 sky130_fd_sc_hd__o21ai_0 _20745_ (.A1(_11219_),
    .A2(_11505_),
    .B1(_11093_),
    .Y(_11506_));
 sky130_fd_sc_hd__a211oi_1 _20746_ (.A1(net3667),
    .A2(_11499_),
    .B1(_11504_),
    .C1(_11506_),
    .Y(_11507_));
 sky130_fd_sc_hd__o21ai_0 _20747_ (.A1(_11403_),
    .A2(_11303_),
    .B1(_11076_),
    .Y(_11508_));
 sky130_fd_sc_hd__a21oi_1 _20748_ (.A1(_11172_),
    .A2(_11148_),
    .B1(net3863),
    .Y(_11509_));
 sky130_fd_sc_hd__a211oi_1 _20749_ (.A1(net3868),
    .A2(_11273_),
    .B1(_11279_),
    .C1(_11509_),
    .Y(_11510_));
 sky130_fd_sc_hd__a31oi_1 _20750_ (.A1(net3667),
    .A2(_11216_),
    .A3(_11508_),
    .B1(_11510_),
    .Y(_11511_));
 sky130_fd_sc_hd__nor3_1 _20751_ (.A(net3866),
    .B(net3855),
    .C(net3862),
    .Y(_11512_));
 sky130_fd_sc_hd__o21ai_0 _20752_ (.A1(_11241_),
    .A2(_11512_),
    .B1(net3672),
    .Y(_11513_));
 sky130_fd_sc_hd__nor2_1 _20753_ (.A(net3868),
    .B(net3857),
    .Y(_11514_));
 sky130_fd_sc_hd__o21ai_0 _20754_ (.A1(_11176_),
    .A2(_11514_),
    .B1(net3866),
    .Y(_11515_));
 sky130_fd_sc_hd__nor2_1 _20755_ (.A(net3857),
    .B(net3862),
    .Y(_11516_));
 sky130_fd_sc_hd__nor2_1 _20756_ (.A(net3855),
    .B(net3858),
    .Y(_11517_));
 sky130_fd_sc_hd__a32oi_1 _20757_ (.A1(net3868),
    .A2(net3670),
    .A3(_11516_),
    .B1(_11517_),
    .B2(_11324_),
    .Y(_11518_));
 sky130_fd_sc_hd__nand4_1 _20758_ (.A(net3854),
    .B(_11513_),
    .C(_11515_),
    .D(_11518_),
    .Y(_11519_));
 sky130_fd_sc_hd__a21oi_1 _20759_ (.A1(_11511_),
    .A2(_11519_),
    .B1(_11164_),
    .Y(_11520_));
 sky130_fd_sc_hd__nand2_1 _20760_ (.A(net3854),
    .B(_11280_),
    .Y(_11521_));
 sky130_fd_sc_hd__a21oi_1 _20761_ (.A1(_12268_[0]),
    .A2(_11176_),
    .B1(_11521_),
    .Y(_11522_));
 sky130_fd_sc_hd__o21ai_0 _20762_ (.A1(net3670),
    .A2(_11286_),
    .B1(_11320_),
    .Y(_11523_));
 sky130_fd_sc_hd__a221oi_1 _20763_ (.A1(_11186_),
    .A2(_11522_),
    .B1(_11523_),
    .B2(net3852),
    .C1(net3855),
    .Y(_11524_));
 sky130_fd_sc_hd__o21ai_0 _20764_ (.A1(_11112_),
    .A2(_11251_),
    .B1(net3670),
    .Y(_11525_));
 sky130_fd_sc_hd__and3_1 _20765_ (.A(_11235_),
    .B(_11285_),
    .C(_11525_),
    .X(_11526_));
 sky130_fd_sc_hd__o221a_1 _20766_ (.A1(net3866),
    .A2(_11211_),
    .B1(_11419_),
    .B2(net3670),
    .C1(net3667),
    .X(_11527_));
 sky130_fd_sc_hd__nor4_1 _20767_ (.A(_11248_),
    .B(_11524_),
    .C(_11526_),
    .D(_11527_),
    .Y(_11528_));
 sky130_fd_sc_hd__nor4_1 _20768_ (.A(_11498_),
    .B(_11507_),
    .C(_11520_),
    .D(_11528_),
    .Y(_00109_));
 sky130_fd_sc_hd__o21ai_0 _20769_ (.A1(net3868),
    .A2(net3866),
    .B1(net3862),
    .Y(_11529_));
 sky130_fd_sc_hd__o32ai_1 _20770_ (.A1(_12275_[0]),
    .A2(_12284_[0]),
    .A3(net3862),
    .B1(_11460_),
    .B2(_11529_),
    .Y(_11530_));
 sky130_fd_sc_hd__nand3_1 _20771_ (.A(net3863),
    .B(_11322_),
    .C(_11426_),
    .Y(_11531_));
 sky130_fd_sc_hd__o211ai_1 _20772_ (.A1(net3858),
    .A2(_11351_),
    .B1(_11221_),
    .C1(_11076_),
    .Y(_11532_));
 sky130_fd_sc_hd__a21oi_1 _20773_ (.A1(_11531_),
    .A2(_11532_),
    .B1(_11279_),
    .Y(_11533_));
 sky130_fd_sc_hd__a21oi_1 _20774_ (.A1(_11285_),
    .A2(_11530_),
    .B1(_11533_),
    .Y(_11534_));
 sky130_fd_sc_hd__a21oi_1 _20775_ (.A1(_11076_),
    .A2(_11268_),
    .B1(_12258_[0]),
    .Y(_11535_));
 sky130_fd_sc_hd__o211ai_1 _20776_ (.A1(net3862),
    .A2(_11481_),
    .B1(_11214_),
    .C1(_11076_),
    .Y(_11536_));
 sky130_fd_sc_hd__a21boi_0 _20777_ (.A1(_12258_[0]),
    .A2(_11536_),
    .B1_N(_12270_[0]),
    .Y(_11537_));
 sky130_fd_sc_hd__a211oi_1 _20778_ (.A1(_12256_[0]),
    .A2(net3858),
    .B1(_11363_),
    .C1(_11076_),
    .Y(_11538_));
 sky130_fd_sc_hd__nor3_1 _20779_ (.A(_11076_),
    .B(_11268_),
    .C(_11538_),
    .Y(_11539_));
 sky130_fd_sc_hd__a21oi_1 _20780_ (.A1(_11481_),
    .A2(_11262_),
    .B1(net3862),
    .Y(_11540_));
 sky130_fd_sc_hd__o22ai_1 _20781_ (.A1(_11268_),
    .A2(_11538_),
    .B1(_11540_),
    .B2(_11349_),
    .Y(_11541_));
 sky130_fd_sc_hd__o41ai_1 _20782_ (.A1(net3858),
    .A2(_11535_),
    .A3(_11537_),
    .A4(_11539_),
    .B1(_11541_),
    .Y(_11542_));
 sky130_fd_sc_hd__a21oi_2 _20783_ (.A1(_11534_),
    .A2(_11542_),
    .B1(_11248_),
    .Y(_11543_));
 sky130_fd_sc_hd__o22ai_1 _20784_ (.A1(net3594),
    .A2(_11212_),
    .B1(_11115_),
    .B2(net3672),
    .Y(_11544_));
 sky130_fd_sc_hd__o211ai_1 _20785_ (.A1(_12261_[0]),
    .A2(net3863),
    .B1(net3858),
    .C1(_11199_),
    .Y(_11545_));
 sky130_fd_sc_hd__a21oi_1 _20786_ (.A1(_12286_[0]),
    .A2(net3862),
    .B1(net3853),
    .Y(_11546_));
 sky130_fd_sc_hd__nand2_1 _20787_ (.A(_11545_),
    .B(_11546_),
    .Y(_11547_));
 sky130_fd_sc_hd__o31ai_1 _20788_ (.A1(_11194_),
    .A2(_11128_),
    .A3(_11544_),
    .B1(_11547_),
    .Y(_11548_));
 sky130_fd_sc_hd__a21oi_1 _20789_ (.A1(_11076_),
    .A2(_11115_),
    .B1(net3868),
    .Y(_11549_));
 sky130_fd_sc_hd__o21ai_0 _20790_ (.A1(net3866),
    .A2(_11156_),
    .B1(_11348_),
    .Y(_11550_));
 sky130_fd_sc_hd__nand2_1 _20791_ (.A(_11076_),
    .B(_11115_),
    .Y(_11551_));
 sky130_fd_sc_hd__o211ai_1 _20792_ (.A1(_11076_),
    .A2(_11419_),
    .B1(_11551_),
    .C1(net3667),
    .Y(_11552_));
 sky130_fd_sc_hd__o311ai_0 _20793_ (.A1(_11219_),
    .A2(_11549_),
    .A3(_11550_),
    .B1(_11093_),
    .C1(_11552_),
    .Y(_11553_));
 sky130_fd_sc_hd__a21oi_1 _20794_ (.A1(net3856),
    .A2(_11548_),
    .B1(_11553_),
    .Y(_11554_));
 sky130_fd_sc_hd__o21ai_0 _20795_ (.A1(_11182_),
    .A2(_11333_),
    .B1(_11076_),
    .Y(_11555_));
 sky130_fd_sc_hd__o211ai_1 _20796_ (.A1(_12261_[0]),
    .A2(_11156_),
    .B1(_11299_),
    .C1(_11555_),
    .Y(_11556_));
 sky130_fd_sc_hd__nand4_1 _20797_ (.A(net3863),
    .B(_11221_),
    .C(_11285_),
    .D(_11368_),
    .Y(_11557_));
 sky130_fd_sc_hd__o311a_1 _20798_ (.A1(net3863),
    .A2(_11219_),
    .A3(_11191_),
    .B1(_11556_),
    .C1(_11557_),
    .X(_11558_));
 sky130_fd_sc_hd__o21ai_0 _20799_ (.A1(_11165_),
    .A2(net3863),
    .B1(net3858),
    .Y(_11559_));
 sky130_fd_sc_hd__o221ai_1 _20800_ (.A1(_12277_[0]),
    .A2(net3858),
    .B1(_11215_),
    .B2(_11559_),
    .C1(_11289_),
    .Y(_11560_));
 sky130_fd_sc_hd__nor3_1 _20801_ (.A(net3863),
    .B(_11418_),
    .C(_11386_),
    .Y(_11561_));
 sky130_fd_sc_hd__nor2_1 _20802_ (.A(net3861),
    .B(_11351_),
    .Y(_11562_));
 sky130_fd_sc_hd__nor3_1 _20803_ (.A(_11076_),
    .B(_11250_),
    .C(_11562_),
    .Y(_11563_));
 sky130_fd_sc_hd__o21ai_0 _20804_ (.A1(_11561_),
    .A2(_11563_),
    .B1(net3667),
    .Y(_11564_));
 sky130_fd_sc_hd__a31oi_1 _20805_ (.A1(_11558_),
    .A2(_11560_),
    .A3(_11564_),
    .B1(_11164_),
    .Y(_11565_));
 sky130_fd_sc_hd__nor2_1 _20806_ (.A(net3672),
    .B(_11156_),
    .Y(_11566_));
 sky130_fd_sc_hd__nor3_1 _20807_ (.A(net3855),
    .B(_11427_),
    .C(_11566_),
    .Y(_11567_));
 sky130_fd_sc_hd__nor3_1 _20808_ (.A(_11140_),
    .B(_11373_),
    .C(_11567_),
    .Y(_11568_));
 sky130_fd_sc_hd__nand2_1 _20809_ (.A(_11216_),
    .B(_11289_),
    .Y(_11569_));
 sky130_fd_sc_hd__a21oi_1 _20810_ (.A1(_12268_[0]),
    .A2(_11076_),
    .B1(net3861),
    .Y(_11570_));
 sky130_fd_sc_hd__a22oi_1 _20811_ (.A1(_12276_[0]),
    .A2(net3861),
    .B1(_11353_),
    .B2(_11570_),
    .Y(_11571_));
 sky130_fd_sc_hd__o22ai_1 _20812_ (.A1(_11439_),
    .A2(_11569_),
    .B1(_11571_),
    .B2(_11219_),
    .Y(_11572_));
 sky130_fd_sc_hd__o21ai_0 _20813_ (.A1(_11568_),
    .A2(_11572_),
    .B1(_11229_),
    .Y(_11573_));
 sky130_fd_sc_hd__nor4b_1 _20814_ (.A(_11543_),
    .B(_11554_),
    .C(_11565_),
    .D_N(_11573_),
    .Y(_00110_));
 sky130_fd_sc_hd__nand3_1 _20815_ (.A(net3863),
    .B(_11316_),
    .C(_11428_),
    .Y(_11574_));
 sky130_fd_sc_hd__o311ai_0 _20816_ (.A1(net3863),
    .A2(_11296_),
    .A3(_11363_),
    .B1(_11574_),
    .C1(net3857),
    .Y(_11575_));
 sky130_fd_sc_hd__nand3_1 _20817_ (.A(net3670),
    .B(_11222_),
    .C(_11225_),
    .Y(_11576_));
 sky130_fd_sc_hd__nand3_1 _20818_ (.A(net3855),
    .B(_11278_),
    .C(_11576_),
    .Y(_11577_));
 sky130_fd_sc_hd__a21oi_2 _20819_ (.A1(_11575_),
    .A2(_11577_),
    .B1(net3852),
    .Y(_11578_));
 sky130_fd_sc_hd__nor2_1 _20820_ (.A(_11460_),
    .B(_11529_),
    .Y(_11579_));
 sky130_fd_sc_hd__o31ai_1 _20821_ (.A1(net3863),
    .A2(_11190_),
    .A3(net3666),
    .B1(_11464_),
    .Y(_11580_));
 sky130_fd_sc_hd__nand2_1 _20822_ (.A(net3855),
    .B(_11580_),
    .Y(_11581_));
 sky130_fd_sc_hd__o311a_1 _20823_ (.A1(net3855),
    .A2(_11266_),
    .A3(_11579_),
    .B1(_11581_),
    .C1(net3852),
    .X(_11582_));
 sky130_fd_sc_hd__o21bai_1 _20824_ (.A1(_11578_),
    .A2(_11582_),
    .B1_N(_11248_),
    .Y(_11583_));
 sky130_fd_sc_hd__nor3_1 _20825_ (.A(net3669),
    .B(_11265_),
    .C(_11251_),
    .Y(_11584_));
 sky130_fd_sc_hd__a211o_1 _20826_ (.A1(_12268_[0]),
    .A2(net3863),
    .B1(net3862),
    .C1(_11444_),
    .X(_11585_));
 sky130_fd_sc_hd__o211ai_1 _20827_ (.A1(_12284_[0]),
    .A2(net3858),
    .B1(net3667),
    .C1(_11585_),
    .Y(_11586_));
 sky130_fd_sc_hd__nand2_1 _20828_ (.A(_12258_[0]),
    .B(_11176_),
    .Y(_11587_));
 sky130_fd_sc_hd__o21ai_0 _20829_ (.A1(_12270_[0]),
    .A2(net3858),
    .B1(_11587_),
    .Y(_11588_));
 sky130_fd_sc_hd__a31oi_1 _20830_ (.A1(net3863),
    .A2(_11280_),
    .A3(_11482_),
    .B1(_11318_),
    .Y(_11589_));
 sky130_fd_sc_hd__a221oi_1 _20831_ (.A1(_11285_),
    .A2(_11588_),
    .B1(_11589_),
    .B2(_11289_),
    .C1(_11164_),
    .Y(_11590_));
 sky130_fd_sc_hd__o311ai_0 _20832_ (.A1(_11279_),
    .A2(_11307_),
    .A3(_11584_),
    .B1(_11586_),
    .C1(_11590_),
    .Y(_11591_));
 sky130_fd_sc_hd__nand3_1 _20833_ (.A(net3863),
    .B(_11224_),
    .C(_11114_),
    .Y(_11592_));
 sky130_fd_sc_hd__nand3_1 _20834_ (.A(net3668),
    .B(_11322_),
    .C(_11300_),
    .Y(_11593_));
 sky130_fd_sc_hd__a21oi_1 _20835_ (.A1(_11199_),
    .A2(_11135_),
    .B1(net3858),
    .Y(_11594_));
 sky130_fd_sc_hd__nor3_1 _20836_ (.A(_11349_),
    .B(_11540_),
    .C(_11594_),
    .Y(_11595_));
 sky130_fd_sc_hd__a31o_1 _20837_ (.A1(_11289_),
    .A2(_11592_),
    .A3(_11593_),
    .B1(_11595_),
    .X(_11596_));
 sky130_fd_sc_hd__o32ai_1 _20838_ (.A1(net3669),
    .A2(net3666),
    .A3(_11303_),
    .B1(_11211_),
    .B2(_12268_[0]),
    .Y(_11597_));
 sky130_fd_sc_hd__o221ai_1 _20839_ (.A1(net3594),
    .A2(_11156_),
    .B1(_11274_),
    .B2(_12257_[0]),
    .C1(_11298_),
    .Y(_11598_));
 sky130_fd_sc_hd__a22o_1 _20840_ (.A1(_11285_),
    .A2(_11597_),
    .B1(_11598_),
    .B2(_11299_),
    .X(_11599_));
 sky130_fd_sc_hd__o21ai_0 _20841_ (.A1(_11596_),
    .A2(_11599_),
    .B1(_11093_),
    .Y(_11600_));
 sky130_fd_sc_hd__nor2_1 _20842_ (.A(net3855),
    .B(net3862),
    .Y(_11601_));
 sky130_fd_sc_hd__a21oi_1 _20843_ (.A1(net3868),
    .A2(_11241_),
    .B1(_11601_),
    .Y(_11602_));
 sky130_fd_sc_hd__a21oi_1 _20844_ (.A1(net3863),
    .A2(_11516_),
    .B1(_11188_),
    .Y(_11603_));
 sky130_fd_sc_hd__nor2_1 _20845_ (.A(_12270_[0]),
    .B(net3863),
    .Y(_11604_));
 sky130_fd_sc_hd__a32oi_1 _20846_ (.A1(net3866),
    .A2(net3863),
    .A3(_11517_),
    .B1(_11604_),
    .B2(_11516_),
    .Y(_11605_));
 sky130_fd_sc_hd__o221ai_1 _20847_ (.A1(net3866),
    .A2(_11602_),
    .B1(_11603_),
    .B2(net3868),
    .C1(_11605_),
    .Y(_11606_));
 sky130_fd_sc_hd__nand2_1 _20848_ (.A(net3854),
    .B(_11606_),
    .Y(_11607_));
 sky130_fd_sc_hd__a211oi_1 _20849_ (.A1(_12261_[0]),
    .A2(_11517_),
    .B1(_11394_),
    .C1(net3670),
    .Y(_11608_));
 sky130_fd_sc_hd__o21ai_0 _20850_ (.A1(_11176_),
    .A2(_11241_),
    .B1(_12270_[0]),
    .Y(_11609_));
 sky130_fd_sc_hd__o211ai_1 _20851_ (.A1(_11443_),
    .A2(_11608_),
    .B1(_11609_),
    .C1(net3852),
    .Y(_11610_));
 sky130_fd_sc_hd__nand3_1 _20852_ (.A(_11229_),
    .B(_11607_),
    .C(_11610_),
    .Y(_11611_));
 sky130_fd_sc_hd__and4_4 _20853_ (.A(_11583_),
    .B(_11591_),
    .C(_11600_),
    .D(_11611_),
    .X(_00111_));
 sky130_fd_sc_hd__xnor2_1 _20854_ (.A(\sa02_sr[1] ),
    .B(\sa31_sub[7] ),
    .Y(_11612_));
 sky130_fd_sc_hd__xnor2_1 _20855_ (.A(\sa12_sr[1] ),
    .B(\sa31_sub[0] ),
    .Y(_11613_));
 sky130_fd_sc_hd__xnor3_1 _20856_ (.A(\sa31_sub[1] ),
    .B(\sa20_sub[0] ),
    .C(net4196),
    .X(_11614_));
 sky130_fd_sc_hd__xnor3_1 _20857_ (.A(_11612_),
    .B(_11613_),
    .C(_11614_),
    .X(_11615_));
 sky130_fd_sc_hd__mux2i_2 _20858_ (.A0(\text_in_r[41] ),
    .A1(_11615_),
    .S(net4111),
    .Y(_11616_));
 sky130_fd_sc_hd__xor2_4 _20859_ (.A(net4135),
    .B(_11616_),
    .X(_11617_));
 sky130_fd_sc_hd__inv_8 _20860_ (.A(_11617_),
    .Y(_11618_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_377 ();
 sky130_fd_sc_hd__xnor3_1 _20862_ (.A(\sa12_sr[0] ),
    .B(net4196),
    .C(net4182),
    .X(_11619_));
 sky130_fd_sc_hd__xnor2_1 _20863_ (.A(_09366_),
    .B(_11619_),
    .Y(_11620_));
 sky130_fd_sc_hd__mux2i_2 _20864_ (.A0(\text_in_r[40] ),
    .A1(_11620_),
    .S(net4111),
    .Y(_11621_));
 sky130_fd_sc_hd__xor2_4 _20865_ (.A(net4136),
    .B(_11621_),
    .X(_11622_));
 sky130_fd_sc_hd__inv_16 _20866_ (.A(_11622_),
    .Y(_11623_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_376 ();
 sky130_fd_sc_hd__xnor3_1 _20868_ (.A(\sa12_sr[2] ),
    .B(\sa31_sub[2] ),
    .C(\sa02_sr[2] ),
    .X(_11624_));
 sky130_fd_sc_hd__xnor2_1 _20869_ (.A(_07075_),
    .B(_11624_),
    .Y(_11625_));
 sky130_fd_sc_hd__mux2i_2 _20870_ (.A0(\text_in_r[42] ),
    .A1(_11625_),
    .S(net4111),
    .Y(_11626_));
 sky130_fd_sc_hd__xnor2_4 _20871_ (.A(\u0.w[2][10] ),
    .B(_11626_),
    .Y(_11627_));
 sky130_fd_sc_hd__clkinv_16 _20872_ (.A(_11627_),
    .Y(_11628_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_367 ();
 sky130_fd_sc_hd__xnor3_1 _20882_ (.A(\sa31_sub[4] ),
    .B(\sa12_sr[5] ),
    .C(\sa02_sr[5] ),
    .X(_11635_));
 sky130_fd_sc_hd__xor2_1 _20883_ (.A(\sa20_sub[4] ),
    .B(\sa31_sub[5] ),
    .X(_11636_));
 sky130_fd_sc_hd__xnor2_2 _20884_ (.A(_11635_),
    .B(_11636_),
    .Y(_11637_));
 sky130_fd_sc_hd__mux2i_4 _20885_ (.A0(\text_in_r[45] ),
    .A1(_11637_),
    .S(net4113),
    .Y(_11638_));
 sky130_fd_sc_hd__xnor2_4 _20886_ (.A(\u0.w[2][13] ),
    .B(_11638_),
    .Y(_11639_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_363 ();
 sky130_fd_sc_hd__nor2b_2 _20891_ (.A(net4230),
    .B_N(\u0.w[2][11] ),
    .Y(_11644_));
 sky130_fd_sc_hd__nor2_1 _20892_ (.A(\u0.w[2][11] ),
    .B(net4230),
    .Y(_11645_));
 sky130_fd_sc_hd__xor2_1 _20893_ (.A(\sa02_sr[3] ),
    .B(\sa31_sub[7] ),
    .X(_11646_));
 sky130_fd_sc_hd__xnor2_1 _20894_ (.A(\sa31_sub[2] ),
    .B(\sa12_sr[3] ),
    .Y(_11647_));
 sky130_fd_sc_hd__xor3_1 _20895_ (.A(\sa20_sub[2] ),
    .B(\sa31_sub[3] ),
    .C(net4196),
    .X(_11648_));
 sky130_fd_sc_hd__xnor3_1 _20896_ (.A(_11646_),
    .B(_11647_),
    .C(_11648_),
    .X(_11649_));
 sky130_fd_sc_hd__mux2i_4 _20897_ (.A0(_11644_),
    .A1(_11645_),
    .S(_11649_),
    .Y(_11650_));
 sky130_fd_sc_hd__nor2_2 _20898_ (.A(\u0.w[2][11] ),
    .B(net4118),
    .Y(_11651_));
 sky130_fd_sc_hd__nand2_1 _20899_ (.A(\u0.w[2][11] ),
    .B(net398),
    .Y(_11652_));
 sky130_fd_sc_hd__nor2_2 _20900_ (.A(\text_in_r[43] ),
    .B(_11652_),
    .Y(_11653_));
 sky130_fd_sc_hd__a21oi_4 _20901_ (.A1(\text_in_r[43] ),
    .A2(_11651_),
    .B1(_11653_),
    .Y(_11654_));
 sky130_fd_sc_hd__and2_4 _20902_ (.A(_11650_),
    .B(_11654_),
    .X(_11655_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_358 ();
 sky130_fd_sc_hd__nor2_2 _20908_ (.A(_12297_[0]),
    .B(net3845),
    .Y(_11661_));
 sky130_fd_sc_hd__a21oi_1 _20909_ (.A1(_12294_[0]),
    .A2(net3845),
    .B1(_11661_),
    .Y(_11662_));
 sky130_fd_sc_hd__nor2_4 _20910_ (.A(net3848),
    .B(_11655_),
    .Y(_11663_));
 sky130_fd_sc_hd__nand2_4 _20911_ (.A(_12304_[0]),
    .B(_11663_),
    .Y(_11664_));
 sky130_fd_sc_hd__xor2_1 _20912_ (.A(\sa12_sr[4] ),
    .B(\sa02_sr[4] ),
    .X(_11665_));
 sky130_fd_sc_hd__xnor2_1 _20913_ (.A(net4183),
    .B(net4182),
    .Y(_11666_));
 sky130_fd_sc_hd__xor3_1 _20914_ (.A(\sa20_sub[3] ),
    .B(\sa31_sub[4] ),
    .C(net4196),
    .X(_11667_));
 sky130_fd_sc_hd__xnor3_1 _20915_ (.A(_11665_),
    .B(_11666_),
    .C(_11667_),
    .X(_11668_));
 sky130_fd_sc_hd__mux2i_4 _20916_ (.A0(\text_in_r[44] ),
    .A1(_11668_),
    .S(net4112),
    .Y(_11669_));
 sky130_fd_sc_hd__xor2_4 _20917_ (.A(\u0.w[2][12] ),
    .B(_11669_),
    .X(_11670_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_356 ();
 sky130_fd_sc_hd__o211ai_1 _20920_ (.A1(net3663),
    .A2(_11662_),
    .B1(_11664_),
    .C1(net3841),
    .Y(_11673_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_354 ();
 sky130_fd_sc_hd__nand2_8 _20923_ (.A(net3663),
    .B(net3845),
    .Y(_11676_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_352 ();
 sky130_fd_sc_hd__nor2_1 _20926_ (.A(_12294_[0]),
    .B(net3843),
    .Y(_11679_));
 sky130_fd_sc_hd__a211oi_2 _20927_ (.A1(_12297_[0]),
    .A2(net3843),
    .B1(_11679_),
    .C1(net3662),
    .Y(_11680_));
 sky130_fd_sc_hd__nor2_1 _20928_ (.A(net3840),
    .B(_11680_),
    .Y(_11681_));
 sky130_fd_sc_hd__o21ai_0 _20929_ (.A1(_12302_[0]),
    .A2(_11676_),
    .B1(_11681_),
    .Y(_11682_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_351 ();
 sky130_fd_sc_hd__nand2_8 _20931_ (.A(_11650_),
    .B(_11654_),
    .Y(_11684_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_350 ();
 sky130_fd_sc_hd__nand2_8 _20933_ (.A(net3848),
    .B(net3838),
    .Y(_11686_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_349 ();
 sky130_fd_sc_hd__mux2i_1 _20935_ (.A0(_12294_[0]),
    .A1(_11623_),
    .S(net3839),
    .Y(_11688_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_348 ();
 sky130_fd_sc_hd__nor2_2 _20937_ (.A(_12299_[0]),
    .B(net3848),
    .Y(_11690_));
 sky130_fd_sc_hd__a21o_1 _20938_ (.A1(_12297_[0]),
    .A2(net3848),
    .B1(_11684_),
    .X(_11691_));
 sky130_fd_sc_hd__o21a_4 _20939_ (.A1(_11690_),
    .A2(_11691_),
    .B1(net3841),
    .X(_11692_));
 sky130_fd_sc_hd__o221ai_2 _20940_ (.A1(_12292_[0]),
    .A2(_11686_),
    .B1(_11688_),
    .B2(net3848),
    .C1(_11692_),
    .Y(_11693_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_346 ();
 sky130_fd_sc_hd__nor2_2 _20943_ (.A(net3848),
    .B(_11684_),
    .Y(_11696_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_343 ();
 sky130_fd_sc_hd__a221oi_1 _20947_ (.A1(_12315_[0]),
    .A2(net3836),
    .B1(net3661),
    .B2(_12293_[0]),
    .C1(net3840),
    .Y(_11700_));
 sky130_fd_sc_hd__nor2_2 _20948_ (.A(_11639_),
    .B(_11700_),
    .Y(_11701_));
 sky130_fd_sc_hd__a32oi_2 _20949_ (.A1(net3847),
    .A2(_11673_),
    .A3(_11682_),
    .B1(_11693_),
    .B2(_11701_),
    .Y(_11702_));
 sky130_fd_sc_hd__xor2_1 _20950_ (.A(net4197),
    .B(\sa31_sub[5] ),
    .X(_11703_));
 sky130_fd_sc_hd__xnor2_1 _20951_ (.A(_11703_),
    .B(_09455_),
    .Y(_11704_));
 sky130_fd_sc_hd__xnor2_1 _20952_ (.A(\sa12_sr[6] ),
    .B(_11704_),
    .Y(_11705_));
 sky130_fd_sc_hd__mux2_8 _20953_ (.A0(\text_in_r[46] ),
    .A1(_11705_),
    .S(net4112),
    .X(_11706_));
 sky130_fd_sc_hd__xor2_4 _20954_ (.A(\u0.w[2][14] ),
    .B(_11706_),
    .X(_11707_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_342 ();
 sky130_fd_sc_hd__xnor2_1 _20956_ (.A(_07084_),
    .B(_09491_),
    .Y(_11709_));
 sky130_fd_sc_hd__xnor2_2 _20957_ (.A(\sa31_sub[6] ),
    .B(_11709_),
    .Y(_11710_));
 sky130_fd_sc_hd__mux2i_4 _20958_ (.A0(\text_in_r[47] ),
    .A1(_11710_),
    .S(net4113),
    .Y(_11711_));
 sky130_fd_sc_hd__xnor2_4 _20959_ (.A(\u0.w[2][15] ),
    .B(_11711_),
    .Y(_11712_));
 sky130_fd_sc_hd__nand2b_4 _20960_ (.A_N(_11707_),
    .B(_11712_),
    .Y(_11713_));
 sky130_fd_sc_hd__or2_4 _20961_ (.A(_11712_),
    .B(_11707_),
    .X(_11714_));
 sky130_fd_sc_hd__xnor2_4 _20962_ (.A(\u0.w[2][12] ),
    .B(_11669_),
    .Y(_11715_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_339 ();
 sky130_fd_sc_hd__xor2_4 _20966_ (.A(\u0.w[2][13] ),
    .B(_11638_),
    .X(_11719_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_336 ();
 sky130_fd_sc_hd__nand2_1 _20970_ (.A(_11623_),
    .B(net3664),
    .Y(_11723_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_333 ();
 sky130_fd_sc_hd__a21oi_1 _20974_ (.A1(net3849),
    .A2(net3847),
    .B1(net3664),
    .Y(_11726_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_328 ();
 sky130_fd_sc_hd__a31oi_1 _20980_ (.A1(_12293_[0]),
    .A2(net3848),
    .A3(net3833),
    .B1(_11684_),
    .Y(_11732_));
 sky130_fd_sc_hd__o221ai_2 _20981_ (.A1(net3833),
    .A2(_11723_),
    .B1(_11726_),
    .B2(net3851),
    .C1(_11732_),
    .Y(_11733_));
 sky130_fd_sc_hd__nor2_4 _20982_ (.A(_12293_[0]),
    .B(net3848),
    .Y(_11734_));
 sky130_fd_sc_hd__nand2_1 _20983_ (.A(_11623_),
    .B(net3848),
    .Y(_11735_));
 sky130_fd_sc_hd__nand2_1 _20984_ (.A(net3850),
    .B(net3849),
    .Y(_11736_));
 sky130_fd_sc_hd__a21oi_1 _20985_ (.A1(_11735_),
    .A2(_11736_),
    .B1(net3832),
    .Y(_11737_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_326 ();
 sky130_fd_sc_hd__a211o_4 _20988_ (.A1(net3832),
    .A2(_11734_),
    .B1(_11737_),
    .C1(net3842),
    .X(_11740_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_324 ();
 sky130_fd_sc_hd__nor2_4 _20991_ (.A(net3846),
    .B(net3834),
    .Y(_11743_));
 sky130_fd_sc_hd__nand2_1 _20992_ (.A(_12302_[0]),
    .B(_11628_),
    .Y(_11744_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_323 ();
 sky130_fd_sc_hd__nand2_4 _20994_ (.A(_11639_),
    .B(_11670_),
    .Y(_11746_));
 sky130_fd_sc_hd__a21oi_1 _20995_ (.A1(_12306_[0]),
    .A2(net3661),
    .B1(_11746_),
    .Y(_11747_));
 sky130_fd_sc_hd__o32ai_1 _20996_ (.A1(_12293_[0]),
    .A2(_11628_),
    .A3(_11743_),
    .B1(_11744_),
    .B2(_11747_),
    .Y(_11748_));
 sky130_fd_sc_hd__inv_1 _20997_ (.A(_12302_[0]),
    .Y(_11749_));
 sky130_fd_sc_hd__nand2_2 _20998_ (.A(_11719_),
    .B(_11670_),
    .Y(_11750_));
 sky130_fd_sc_hd__nand2_1 _20999_ (.A(_12302_[0]),
    .B(_11750_),
    .Y(_11751_));
 sky130_fd_sc_hd__a221oi_1 _21000_ (.A1(_11749_),
    .A2(_11747_),
    .B1(_11751_),
    .B2(_12293_[0]),
    .C1(_11686_),
    .Y(_11752_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_322 ();
 sky130_fd_sc_hd__a311oi_1 _21002_ (.A1(_12293_[0]),
    .A2(_11639_),
    .A3(net3840),
    .B1(_11684_),
    .C1(_11628_),
    .Y(_11754_));
 sky130_fd_sc_hd__o21ai_0 _21003_ (.A1(_11663_),
    .A2(_11754_),
    .B1(_12292_[0]),
    .Y(_11755_));
 sky130_fd_sc_hd__o21ai_0 _21004_ (.A1(_11747_),
    .A2(_11743_),
    .B1(_11755_),
    .Y(_11756_));
 sky130_fd_sc_hd__a211oi_1 _21005_ (.A1(_11655_),
    .A2(_11748_),
    .B1(_11752_),
    .C1(_11756_),
    .Y(_11757_));
 sky130_fd_sc_hd__a31oi_2 _21006_ (.A1(net3834),
    .A2(_11733_),
    .A3(_11740_),
    .B1(_11757_),
    .Y(_11758_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_320 ();
 sky130_fd_sc_hd__nor2_4 _21009_ (.A(_12299_[0]),
    .B(_11655_),
    .Y(_11761_));
 sky130_fd_sc_hd__nor2_4 _21010_ (.A(_12294_[0]),
    .B(_11684_),
    .Y(_11762_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_318 ();
 sky130_fd_sc_hd__o21ai_2 _21013_ (.A1(_11761_),
    .A2(_11762_),
    .B1(net3848),
    .Y(_11765_));
 sky130_fd_sc_hd__nand2_1 _21014_ (.A(_12292_[0]),
    .B(net3661),
    .Y(_11766_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_317 ();
 sky130_fd_sc_hd__nand2_4 _21016_ (.A(net3851),
    .B(net3843),
    .Y(_11768_));
 sky130_fd_sc_hd__nand2_8 _21017_ (.A(_11623_),
    .B(_11684_),
    .Y(_11769_));
 sky130_fd_sc_hd__nor2_2 _21018_ (.A(_12302_[0]),
    .B(net3843),
    .Y(_11770_));
 sky130_fd_sc_hd__nor2_2 _21019_ (.A(_12293_[0]),
    .B(_11684_),
    .Y(_11771_));
 sky130_fd_sc_hd__nor3_1 _21020_ (.A(net3848),
    .B(_11770_),
    .C(net3608),
    .Y(_11772_));
 sky130_fd_sc_hd__a311oi_1 _21021_ (.A1(net3848),
    .A2(_11768_),
    .A3(_11769_),
    .B1(_11772_),
    .C1(net3834),
    .Y(_11773_));
 sky130_fd_sc_hd__a311o_1 _21022_ (.A1(net3834),
    .A2(_11765_),
    .A3(_11766_),
    .B1(_11773_),
    .C1(_11719_),
    .X(_11774_));
 sky130_fd_sc_hd__nor2_1 _21023_ (.A(net3849),
    .B(net3848),
    .Y(_11775_));
 sky130_fd_sc_hd__nor2_1 _21024_ (.A(_12306_[0]),
    .B(_11628_),
    .Y(_11776_));
 sky130_fd_sc_hd__o21ai_2 _21025_ (.A1(_11775_),
    .A2(_11776_),
    .B1(net3836),
    .Y(_11777_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_315 ();
 sky130_fd_sc_hd__nand2_1 _21028_ (.A(_12304_[0]),
    .B(net3848),
    .Y(_11780_));
 sky130_fd_sc_hd__a2bb2oi_1 _21029_ (.A1_N(_12293_[0]),
    .A2_N(_11686_),
    .B1(_11780_),
    .B2(net3842),
    .Y(_11781_));
 sky130_fd_sc_hd__a221oi_1 _21030_ (.A1(_12299_[0]),
    .A2(net3661),
    .B1(_11781_),
    .B2(net3834),
    .C1(net3846),
    .Y(_11782_));
 sky130_fd_sc_hd__o21ai_1 _21031_ (.A1(net3834),
    .A2(_11777_),
    .B1(_11782_),
    .Y(_11783_));
 sky130_fd_sc_hd__and2_4 _21032_ (.A(_11712_),
    .B(_11707_),
    .X(_11784_));
 sky130_fd_sc_hd__nand2_2 _21033_ (.A(net3665),
    .B(_11628_),
    .Y(_11785_));
 sky130_fd_sc_hd__o211ai_1 _21034_ (.A1(_12294_[0]),
    .A2(_11628_),
    .B1(net3844),
    .C1(_11785_),
    .Y(_11786_));
 sky130_fd_sc_hd__xor2_4 _21035_ (.A(\u0.w[2][15] ),
    .B(_11711_),
    .X(_11787_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_314 ();
 sky130_fd_sc_hd__nand2_8 _21037_ (.A(_11787_),
    .B(_11707_),
    .Y(_11789_));
 sky130_fd_sc_hd__a41oi_1 _21038_ (.A1(_11719_),
    .A2(net3840),
    .A3(_11786_),
    .A4(_11777_),
    .B1(_11789_),
    .Y(_11790_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_313 ();
 sky130_fd_sc_hd__nand2b_2 _21040_ (.A_N(_12308_[0]),
    .B(net3837),
    .Y(_11792_));
 sky130_fd_sc_hd__nand3_1 _21041_ (.A(net3848),
    .B(_11792_),
    .C(_11768_),
    .Y(_11793_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_312 ();
 sky130_fd_sc_hd__nand2_2 _21043_ (.A(_12297_[0]),
    .B(net3843),
    .Y(_11795_));
 sky130_fd_sc_hd__nand2_8 _21044_ (.A(net3849),
    .B(net3838),
    .Y(_11796_));
 sky130_fd_sc_hd__nand3_1 _21045_ (.A(net3662),
    .B(_11795_),
    .C(_11796_),
    .Y(_11797_));
 sky130_fd_sc_hd__nor2_4 _21046_ (.A(net3846),
    .B(net3840),
    .Y(_11798_));
 sky130_fd_sc_hd__nand3_1 _21047_ (.A(_11793_),
    .B(_11797_),
    .C(_11798_),
    .Y(_11799_));
 sky130_fd_sc_hd__a21oi_4 _21048_ (.A1(net4072),
    .A2(_11654_),
    .B1(_12293_[0]),
    .Y(_11800_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_311 ();
 sky130_fd_sc_hd__a211oi_2 _21050_ (.A1(net3849),
    .A2(_11655_),
    .B1(_11800_),
    .C1(net3664),
    .Y(_11802_));
 sky130_fd_sc_hd__a31oi_1 _21051_ (.A1(net3662),
    .A2(_11792_),
    .A3(_11795_),
    .B1(_11802_),
    .Y(_11803_));
 sky130_fd_sc_hd__mux2i_1 _21052_ (.A0(_12297_[0]),
    .A1(net3849),
    .S(net3843),
    .Y(_11804_));
 sky130_fd_sc_hd__o221ai_1 _21053_ (.A1(_12299_[0]),
    .A2(_11686_),
    .B1(_11804_),
    .B2(net3848),
    .C1(net3840),
    .Y(_11805_));
 sky130_fd_sc_hd__o211ai_1 _21054_ (.A1(net3840),
    .A2(_11803_),
    .B1(_11805_),
    .C1(net3846),
    .Y(_11806_));
 sky130_fd_sc_hd__and3_4 _21055_ (.A(_11790_),
    .B(_11799_),
    .C(_11806_),
    .X(_11807_));
 sky130_fd_sc_hd__a31oi_2 _21056_ (.A1(_11774_),
    .A2(_11783_),
    .A3(_11784_),
    .B1(_11807_),
    .Y(_11808_));
 sky130_fd_sc_hd__o221ai_4 _21057_ (.A1(_11702_),
    .A2(_11713_),
    .B1(_11714_),
    .B2(_11758_),
    .C1(_11808_),
    .Y(_00112_));
 sky130_fd_sc_hd__nand2_4 _21058_ (.A(_12293_[0]),
    .B(net3839),
    .Y(_11809_));
 sky130_fd_sc_hd__nand2_2 _21059_ (.A(_12292_[0]),
    .B(net3845),
    .Y(_11810_));
 sky130_fd_sc_hd__nand3_2 _21060_ (.A(net3848),
    .B(_11809_),
    .C(_11810_),
    .Y(_11811_));
 sky130_fd_sc_hd__a22oi_1 _21061_ (.A1(_11623_),
    .A2(net3661),
    .B1(_11663_),
    .B2(net3593),
    .Y(_11812_));
 sky130_fd_sc_hd__nand2_8 _21062_ (.A(net3665),
    .B(net3839),
    .Y(_11813_));
 sky130_fd_sc_hd__nor2_1 _21063_ (.A(net3663),
    .B(_11813_),
    .Y(_11814_));
 sky130_fd_sc_hd__nand2_8 _21064_ (.A(net3848),
    .B(_11655_),
    .Y(_11815_));
 sky130_fd_sc_hd__nor2_2 _21065_ (.A(_12306_[0]),
    .B(_11815_),
    .Y(_11816_));
 sky130_fd_sc_hd__a2111oi_0 _21066_ (.A1(_12308_[0]),
    .A2(_11663_),
    .B1(_11814_),
    .C1(_11816_),
    .D1(_11719_),
    .Y(_11817_));
 sky130_fd_sc_hd__a311o_1 _21067_ (.A1(_11719_),
    .A2(_11811_),
    .A3(_11812_),
    .B1(net3841),
    .C1(_11817_),
    .X(_11818_));
 sky130_fd_sc_hd__xnor2_2 _21068_ (.A(_11628_),
    .B(_11655_),
    .Y(_11819_));
 sky130_fd_sc_hd__o22ai_1 _21069_ (.A1(net3665),
    .A2(_11769_),
    .B1(_11819_),
    .B2(_11623_),
    .Y(_11820_));
 sky130_fd_sc_hd__a21oi_1 _21070_ (.A1(_12293_[0]),
    .A2(net3661),
    .B1(_11820_),
    .Y(_11821_));
 sky130_fd_sc_hd__nand2_4 _21071_ (.A(_11628_),
    .B(_11684_),
    .Y(_11822_));
 sky130_fd_sc_hd__a21oi_1 _21072_ (.A1(net3593),
    .A2(net3845),
    .B1(_11800_),
    .Y(_11823_));
 sky130_fd_sc_hd__o221ai_1 _21073_ (.A1(_12306_[0]),
    .A2(_11822_),
    .B1(_11823_),
    .B2(net3662),
    .C1(net3847),
    .Y(_11824_));
 sky130_fd_sc_hd__o211ai_1 _21074_ (.A1(net3847),
    .A2(_11821_),
    .B1(_11824_),
    .C1(net3841),
    .Y(_11825_));
 sky130_fd_sc_hd__nor2_4 _21075_ (.A(_11670_),
    .B(_11655_),
    .Y(_00421_));
 sky130_fd_sc_hd__mux2i_1 _21076_ (.A0(_12293_[0]),
    .A1(_12308_[0]),
    .S(net3848),
    .Y(_00422_));
 sky130_fd_sc_hd__nand2_1 _21077_ (.A(_12297_[0]),
    .B(_11670_),
    .Y(_00423_));
 sky130_fd_sc_hd__a21oi_1 _21078_ (.A1(net3665),
    .A2(_11715_),
    .B1(_11628_),
    .Y(_00424_));
 sky130_fd_sc_hd__and2_0 _21079_ (.A(_12299_[0]),
    .B(_11628_),
    .X(_00425_));
 sky130_fd_sc_hd__a211oi_1 _21080_ (.A1(_00423_),
    .A2(_00424_),
    .B1(_11684_),
    .C1(_00425_),
    .Y(_00426_));
 sky130_fd_sc_hd__a221oi_2 _21081_ (.A1(_12322_[0]),
    .A2(_00421_),
    .B1(_00422_),
    .B2(_11692_),
    .C1(_00426_),
    .Y(_00427_));
 sky130_fd_sc_hd__nor3_1 _21082_ (.A(_11707_),
    .B(net3847),
    .C(_00427_),
    .Y(_00428_));
 sky130_fd_sc_hd__nor2_2 _21083_ (.A(net3593),
    .B(_11684_),
    .Y(_00429_));
 sky130_fd_sc_hd__nand2_2 _21084_ (.A(_11623_),
    .B(_11655_),
    .Y(_00430_));
 sky130_fd_sc_hd__nand3_1 _21085_ (.A(net3662),
    .B(_00430_),
    .C(_11796_),
    .Y(_00431_));
 sky130_fd_sc_hd__o311ai_0 _21086_ (.A1(net3662),
    .A2(_11800_),
    .A3(_00429_),
    .B1(_00431_),
    .C1(net3835),
    .Y(_00432_));
 sky130_fd_sc_hd__nor2_4 _21087_ (.A(net3849),
    .B(net3839),
    .Y(_00433_));
 sky130_fd_sc_hd__nand2b_4 _21088_ (.A_N(_12297_[0]),
    .B(net3838),
    .Y(_00434_));
 sky130_fd_sc_hd__nand2_2 _21089_ (.A(net3665),
    .B(_11655_),
    .Y(_00435_));
 sky130_fd_sc_hd__nand2_1 _21090_ (.A(_00434_),
    .B(_00435_),
    .Y(_00436_));
 sky130_fd_sc_hd__a221o_1 _21091_ (.A1(net3851),
    .A2(_00433_),
    .B1(_00436_),
    .B2(net3663),
    .C1(net3835),
    .X(_00437_));
 sky130_fd_sc_hd__a211oi_1 _21092_ (.A1(_00432_),
    .A2(_00437_),
    .B1(_11707_),
    .C1(_11719_),
    .Y(_00438_));
 sky130_fd_sc_hd__a311o_1 _21093_ (.A1(_11707_),
    .A2(_11818_),
    .A3(_11825_),
    .B1(_00428_),
    .C1(_00438_),
    .X(_00439_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_310 ();
 sky130_fd_sc_hd__a21oi_1 _21095_ (.A1(_12292_[0]),
    .A2(_11684_),
    .B1(_11762_),
    .Y(_00441_));
 sky130_fd_sc_hd__nand3_2 _21096_ (.A(net3662),
    .B(_11809_),
    .C(_00430_),
    .Y(_00442_));
 sky130_fd_sc_hd__o21ai_0 _21097_ (.A1(net3662),
    .A2(_00441_),
    .B1(_00442_),
    .Y(_00443_));
 sky130_fd_sc_hd__and3_4 _21098_ (.A(_12308_[0]),
    .B(net4072),
    .C(_11654_),
    .X(_00444_));
 sky130_fd_sc_hd__a21oi_4 _21099_ (.A1(net4072),
    .A2(_11654_),
    .B1(_12306_[0]),
    .Y(_00445_));
 sky130_fd_sc_hd__a21oi_1 _21100_ (.A1(_12294_[0]),
    .A2(_11655_),
    .B1(_00445_),
    .Y(_00446_));
 sky130_fd_sc_hd__nand2_1 _21101_ (.A(net3662),
    .B(_00446_),
    .Y(_00447_));
 sky130_fd_sc_hd__o311ai_0 _21102_ (.A1(net3662),
    .A2(_11800_),
    .A3(_00444_),
    .B1(_00447_),
    .C1(_11719_),
    .Y(_00448_));
 sky130_fd_sc_hd__o21ai_0 _21103_ (.A1(_11719_),
    .A2(_00443_),
    .B1(_00448_),
    .Y(_00449_));
 sky130_fd_sc_hd__o21ai_2 _21104_ (.A1(_00433_),
    .A2(_11761_),
    .B1(net3848),
    .Y(_00450_));
 sky130_fd_sc_hd__o211ai_1 _21105_ (.A1(_12292_[0]),
    .A2(_11684_),
    .B1(_11813_),
    .C1(net3662),
    .Y(_00451_));
 sky130_fd_sc_hd__nand3_1 _21106_ (.A(net3847),
    .B(_00450_),
    .C(_00451_),
    .Y(_00452_));
 sky130_fd_sc_hd__clkinv_2 _21107_ (.A(_12306_[0]),
    .Y(_00453_));
 sky130_fd_sc_hd__nor2_4 _21108_ (.A(_00453_),
    .B(net3837),
    .Y(_00454_));
 sky130_fd_sc_hd__o21ai_0 _21109_ (.A1(_11800_),
    .A2(_00454_),
    .B1(net3848),
    .Y(_00455_));
 sky130_fd_sc_hd__o211ai_1 _21110_ (.A1(_11623_),
    .A2(_11676_),
    .B1(_00455_),
    .C1(_11719_),
    .Y(_00456_));
 sky130_fd_sc_hd__a31oi_1 _21111_ (.A1(net3841),
    .A2(_00452_),
    .A3(_00456_),
    .B1(_11789_),
    .Y(_00457_));
 sky130_fd_sc_hd__o21ai_0 _21112_ (.A1(net3841),
    .A2(_00449_),
    .B1(_00457_),
    .Y(_00458_));
 sky130_fd_sc_hd__nor2_4 _21113_ (.A(_11712_),
    .B(_11707_),
    .Y(_00459_));
 sky130_fd_sc_hd__nand2_1 _21114_ (.A(_12306_[0]),
    .B(net3848),
    .Y(_00460_));
 sky130_fd_sc_hd__nand3_1 _21115_ (.A(net3843),
    .B(_11744_),
    .C(_00460_),
    .Y(_00461_));
 sky130_fd_sc_hd__o311ai_2 _21116_ (.A1(_12318_[0]),
    .A2(_11639_),
    .A3(net3843),
    .B1(_00461_),
    .C1(net3840),
    .Y(_00462_));
 sky130_fd_sc_hd__o211ai_1 _21117_ (.A1(_12292_[0]),
    .A2(_11684_),
    .B1(_00434_),
    .C1(net3662),
    .Y(_00463_));
 sky130_fd_sc_hd__o31ai_1 _21118_ (.A1(net3662),
    .A2(_00433_),
    .A3(_00445_),
    .B1(_00463_),
    .Y(_00464_));
 sky130_fd_sc_hd__nor2_4 _21119_ (.A(net3850),
    .B(_11684_),
    .Y(_00465_));
 sky130_fd_sc_hd__nor2_2 _21120_ (.A(net3665),
    .B(_11655_),
    .Y(_00466_));
 sky130_fd_sc_hd__o21ai_2 _21121_ (.A1(_00465_),
    .A2(_00466_),
    .B1(_11628_),
    .Y(_00467_));
 sky130_fd_sc_hd__nand2_2 _21122_ (.A(_11719_),
    .B(_11715_),
    .Y(_00468_));
 sky130_fd_sc_hd__a21oi_1 _21123_ (.A1(_00450_),
    .A2(_00467_),
    .B1(_00468_),
    .Y(_00469_));
 sky130_fd_sc_hd__a31oi_1 _21124_ (.A1(net3847),
    .A2(net3835),
    .A3(_00464_),
    .B1(_00469_),
    .Y(_00470_));
 sky130_fd_sc_hd__nand3_2 _21125_ (.A(_00459_),
    .B(_00462_),
    .C(_00470_),
    .Y(_00471_));
 sky130_fd_sc_hd__o211ai_1 _21126_ (.A1(_11787_),
    .A2(_00439_),
    .B1(_00458_),
    .C1(_00471_),
    .Y(_00113_));
 sky130_fd_sc_hd__o21ai_2 _21127_ (.A1(_11770_),
    .A2(_00465_),
    .B1(net3848),
    .Y(_00472_));
 sky130_fd_sc_hd__a21oi_1 _21128_ (.A1(_12292_[0]),
    .A2(net3842),
    .B1(_11800_),
    .Y(_00473_));
 sky130_fd_sc_hd__nand2_1 _21129_ (.A(_11628_),
    .B(_00473_),
    .Y(_00474_));
 sky130_fd_sc_hd__nor2_1 _21130_ (.A(_11618_),
    .B(net3848),
    .Y(_00475_));
 sky130_fd_sc_hd__o21ai_0 _21131_ (.A1(_00465_),
    .A2(_00475_),
    .B1(_12293_[0]),
    .Y(_00476_));
 sky130_fd_sc_hd__nor2_1 _21132_ (.A(net3850),
    .B(_11628_),
    .Y(_00477_));
 sky130_fd_sc_hd__a22oi_1 _21133_ (.A1(_11735_),
    .A2(_00466_),
    .B1(_00477_),
    .B2(_11769_),
    .Y(_00478_));
 sky130_fd_sc_hd__a21oi_1 _21134_ (.A1(_00476_),
    .A2(_00478_),
    .B1(net3832),
    .Y(_00479_));
 sky130_fd_sc_hd__a311oi_1 _21135_ (.A1(net3832),
    .A2(_00472_),
    .A3(_00474_),
    .B1(_00479_),
    .C1(net3840),
    .Y(_00480_));
 sky130_fd_sc_hd__a211oi_1 _21136_ (.A1(_12297_[0]),
    .A2(net3848),
    .B1(net3842),
    .C1(_11734_),
    .Y(_00481_));
 sky130_fd_sc_hd__a211oi_1 _21137_ (.A1(_12315_[0]),
    .A2(net3842),
    .B1(_00481_),
    .C1(net3832),
    .Y(_00482_));
 sky130_fd_sc_hd__nand2_1 _21138_ (.A(_11618_),
    .B(net3848),
    .Y(_00483_));
 sky130_fd_sc_hd__o21ai_0 _21139_ (.A1(_12318_[0]),
    .A2(net3836),
    .B1(net3832),
    .Y(_00484_));
 sky130_fd_sc_hd__a31oi_1 _21140_ (.A1(net3836),
    .A2(_11736_),
    .A3(_00483_),
    .B1(_00484_),
    .Y(_00485_));
 sky130_fd_sc_hd__nor3_1 _21141_ (.A(net3834),
    .B(_00482_),
    .C(_00485_),
    .Y(_00486_));
 sky130_fd_sc_hd__o21ai_1 _21142_ (.A1(_00480_),
    .A2(_00486_),
    .B1(_11784_),
    .Y(_00487_));
 sky130_fd_sc_hd__nor2_2 _21143_ (.A(_12294_[0]),
    .B(_12299_[0]),
    .Y(_00488_));
 sky130_fd_sc_hd__inv_1 _21144_ (.A(_00488_),
    .Y(_00489_));
 sky130_fd_sc_hd__nand3_1 _21145_ (.A(net3848),
    .B(_11684_),
    .C(_00489_),
    .Y(_00490_));
 sky130_fd_sc_hd__o221ai_1 _21146_ (.A1(_12302_[0]),
    .A2(_11676_),
    .B1(_11819_),
    .B2(_12306_[0]),
    .C1(_00490_),
    .Y(_00491_));
 sky130_fd_sc_hd__nor2_1 _21147_ (.A(net3840),
    .B(_00491_),
    .Y(_00492_));
 sky130_fd_sc_hd__a221oi_1 _21148_ (.A1(_12299_[0]),
    .A2(_11663_),
    .B1(_00473_),
    .B2(net3848),
    .C1(net3834),
    .Y(_00493_));
 sky130_fd_sc_hd__nor3_1 _21149_ (.A(net3833),
    .B(_00492_),
    .C(_00493_),
    .Y(_00494_));
 sky130_fd_sc_hd__nand2_1 _21150_ (.A(_12297_[0]),
    .B(_11628_),
    .Y(_00495_));
 sky130_fd_sc_hd__nand3_1 _21151_ (.A(_00421_),
    .B(_00483_),
    .C(_00495_),
    .Y(_00496_));
 sky130_fd_sc_hd__nor2_2 _21152_ (.A(net3834),
    .B(net3836),
    .Y(_00497_));
 sky130_fd_sc_hd__nand2_4 _21153_ (.A(net3840),
    .B(net3836),
    .Y(_00498_));
 sky130_fd_sc_hd__nor2_1 _21154_ (.A(_12313_[0]),
    .B(_00498_),
    .Y(_00499_));
 sky130_fd_sc_hd__a21oi_1 _21155_ (.A1(_00495_),
    .A2(_00497_),
    .B1(_00499_),
    .Y(_00500_));
 sky130_fd_sc_hd__nand3_1 _21156_ (.A(_12324_[0]),
    .B(net3834),
    .C(net3842),
    .Y(_00501_));
 sky130_fd_sc_hd__a31oi_1 _21157_ (.A1(_00496_),
    .A2(_00500_),
    .A3(_00501_),
    .B1(net3846),
    .Y(_00502_));
 sky130_fd_sc_hd__nor2_4 _21158_ (.A(_11787_),
    .B(net3660),
    .Y(_00503_));
 sky130_fd_sc_hd__o21ai_0 _21159_ (.A1(_00494_),
    .A2(_00502_),
    .B1(_00503_),
    .Y(_00504_));
 sky130_fd_sc_hd__nand2_1 _21160_ (.A(_12306_[0]),
    .B(_11684_),
    .Y(_00505_));
 sky130_fd_sc_hd__a21oi_1 _21161_ (.A1(_11795_),
    .A2(_00505_),
    .B1(net3848),
    .Y(_00506_));
 sky130_fd_sc_hd__nor2_1 _21162_ (.A(_12308_[0]),
    .B(_11686_),
    .Y(_00507_));
 sky130_fd_sc_hd__nor2_1 _21163_ (.A(_11623_),
    .B(net3843),
    .Y(_00508_));
 sky130_fd_sc_hd__nor2_1 _21164_ (.A(_00508_),
    .B(net3609),
    .Y(_00509_));
 sky130_fd_sc_hd__o21ai_0 _21165_ (.A1(_11679_),
    .A2(_00465_),
    .B1(net3662),
    .Y(_00510_));
 sky130_fd_sc_hd__o211ai_1 _21166_ (.A1(net3662),
    .A2(_00509_),
    .B1(_00510_),
    .C1(net3834),
    .Y(_00511_));
 sky130_fd_sc_hd__o311ai_0 _21167_ (.A1(net3834),
    .A2(_00506_),
    .A3(_00507_),
    .B1(_00511_),
    .C1(_11639_),
    .Y(_00512_));
 sky130_fd_sc_hd__nand2_1 _21168_ (.A(net3848),
    .B(_00436_),
    .Y(_00513_));
 sky130_fd_sc_hd__o311ai_0 _21169_ (.A1(net3848),
    .A2(net3608),
    .A3(_11761_),
    .B1(_11743_),
    .C1(_00513_),
    .Y(_00514_));
 sky130_fd_sc_hd__nor2_4 _21170_ (.A(net3851),
    .B(net3845),
    .Y(_00515_));
 sky130_fd_sc_hd__o21ai_0 _21171_ (.A1(_11661_),
    .A2(_00444_),
    .B1(net3662),
    .Y(_00516_));
 sky130_fd_sc_hd__o311ai_1 _21172_ (.A1(net3662),
    .A2(_00515_),
    .A3(_00429_),
    .B1(_00516_),
    .C1(_11798_),
    .Y(_00517_));
 sky130_fd_sc_hd__nand4_1 _21173_ (.A(_00459_),
    .B(_00512_),
    .C(_00514_),
    .D(_00517_),
    .Y(_00518_));
 sky130_fd_sc_hd__o21ai_0 _21174_ (.A1(_12304_[0]),
    .A2(net3839),
    .B1(_11796_),
    .Y(_00519_));
 sky130_fd_sc_hd__nor2_1 _21175_ (.A(_12308_[0]),
    .B(net3839),
    .Y(_00520_));
 sky130_fd_sc_hd__or3_1 _21176_ (.A(net3848),
    .B(_11761_),
    .C(_00520_),
    .X(_00521_));
 sky130_fd_sc_hd__o21ai_0 _21177_ (.A1(net3664),
    .A2(_00519_),
    .B1(_00521_),
    .Y(_00522_));
 sky130_fd_sc_hd__nand2_4 _21178_ (.A(_12304_[0]),
    .B(_11655_),
    .Y(_00523_));
 sky130_fd_sc_hd__a311oi_1 _21179_ (.A1(net3848),
    .A2(_11813_),
    .A3(_00523_),
    .B1(net3835),
    .C1(_11690_),
    .Y(_00524_));
 sky130_fd_sc_hd__a21oi_1 _21180_ (.A1(net3835),
    .A2(_00522_),
    .B1(_00524_),
    .Y(_00525_));
 sky130_fd_sc_hd__clkinv_1 _21181_ (.A(_12293_[0]),
    .Y(_00526_));
 sky130_fd_sc_hd__nand2_2 _21182_ (.A(_00526_),
    .B(_11684_),
    .Y(_00527_));
 sky130_fd_sc_hd__a21oi_1 _21183_ (.A1(_00527_),
    .A2(_00523_),
    .B1(net3848),
    .Y(_00528_));
 sky130_fd_sc_hd__o21ai_2 _21184_ (.A1(_11802_),
    .A2(_00528_),
    .B1(net3841),
    .Y(_00529_));
 sky130_fd_sc_hd__o21ai_0 _21185_ (.A1(_12304_[0]),
    .A2(_11628_),
    .B1(_11785_),
    .Y(_00530_));
 sky130_fd_sc_hd__nor2_4 _21186_ (.A(net3849),
    .B(_11628_),
    .Y(_00531_));
 sky130_fd_sc_hd__and2_0 _21187_ (.A(_12308_[0]),
    .B(_11628_),
    .X(_00532_));
 sky130_fd_sc_hd__o31ai_1 _21188_ (.A1(_11684_),
    .A2(_00531_),
    .A3(_00532_),
    .B1(_11715_),
    .Y(_00533_));
 sky130_fd_sc_hd__a21oi_1 _21189_ (.A1(_11684_),
    .A2(_00530_),
    .B1(_00533_),
    .Y(_00534_));
 sky130_fd_sc_hd__nor2_1 _21190_ (.A(net3833),
    .B(_00534_),
    .Y(_00535_));
 sky130_fd_sc_hd__a221o_4 _21191_ (.A1(net3833),
    .A2(_00525_),
    .B1(_00529_),
    .B2(_00535_),
    .C1(_11789_),
    .X(_00536_));
 sky130_fd_sc_hd__nand4_1 _21192_ (.A(_00487_),
    .B(_00504_),
    .C(_00518_),
    .D(_00536_),
    .Y(_00114_));
 sky130_fd_sc_hd__o22ai_1 _21193_ (.A1(_12292_[0]),
    .A2(_11686_),
    .B1(_11676_),
    .B2(net3851),
    .Y(_00537_));
 sky130_fd_sc_hd__a21oi_1 _21194_ (.A1(net3848),
    .A2(_11768_),
    .B1(net3849),
    .Y(_00538_));
 sky130_fd_sc_hd__o21a_1 _21195_ (.A1(_00537_),
    .A2(_00538_),
    .B1(net3841),
    .X(_00539_));
 sky130_fd_sc_hd__nand2_4 _21196_ (.A(_12308_[0]),
    .B(_11655_),
    .Y(_00540_));
 sky130_fd_sc_hd__nand2_4 _21197_ (.A(_12293_[0]),
    .B(net3843),
    .Y(_00541_));
 sky130_fd_sc_hd__nand2_2 _21198_ (.A(_12304_[0]),
    .B(_11684_),
    .Y(_00542_));
 sky130_fd_sc_hd__and3_4 _21199_ (.A(net3848),
    .B(_00541_),
    .C(_00542_),
    .X(_00543_));
 sky130_fd_sc_hd__a311oi_1 _21200_ (.A1(_11628_),
    .A2(_11796_),
    .A3(_00540_),
    .B1(_00543_),
    .C1(net3841),
    .Y(_00544_));
 sky130_fd_sc_hd__nor2_1 _21201_ (.A(_12304_[0]),
    .B(net3843),
    .Y(_00545_));
 sky130_fd_sc_hd__a21oi_1 _21202_ (.A1(_12302_[0]),
    .A2(net3843),
    .B1(_00545_),
    .Y(_00546_));
 sky130_fd_sc_hd__nor2_2 _21203_ (.A(net3843),
    .B(_00489_),
    .Y(_00547_));
 sky130_fd_sc_hd__o21ai_1 _21204_ (.A1(_00454_),
    .A2(_00547_),
    .B1(net3848),
    .Y(_00548_));
 sky130_fd_sc_hd__o211ai_1 _21205_ (.A1(net3848),
    .A2(_00546_),
    .B1(_00548_),
    .C1(_11670_),
    .Y(_00549_));
 sky130_fd_sc_hd__nand3_1 _21206_ (.A(net3833),
    .B(_00533_),
    .C(_00549_),
    .Y(_00550_));
 sky130_fd_sc_hd__o311ai_2 _21207_ (.A1(net3833),
    .A2(_00539_),
    .A3(_00544_),
    .B1(_00550_),
    .C1(net3660),
    .Y(_00551_));
 sky130_fd_sc_hd__nand2_2 _21208_ (.A(_12308_[0]),
    .B(_11684_),
    .Y(_00552_));
 sky130_fd_sc_hd__a21oi_1 _21209_ (.A1(_00430_),
    .A2(_00552_),
    .B1(net3848),
    .Y(_00553_));
 sky130_fd_sc_hd__nor2_1 _21210_ (.A(_11623_),
    .B(net3848),
    .Y(_00554_));
 sky130_fd_sc_hd__o211ai_1 _21211_ (.A1(_00554_),
    .A2(_00541_),
    .B1(_00490_),
    .C1(_11743_),
    .Y(_00555_));
 sky130_fd_sc_hd__a22oi_1 _21212_ (.A1(_12294_[0]),
    .A2(net3848),
    .B1(_11719_),
    .B2(_11734_),
    .Y(_00556_));
 sky130_fd_sc_hd__nand2_1 _21213_ (.A(_11715_),
    .B(_11655_),
    .Y(_00557_));
 sky130_fd_sc_hd__nor2_1 _21214_ (.A(_11617_),
    .B(_11639_),
    .Y(_00558_));
 sky130_fd_sc_hd__a211oi_1 _21215_ (.A1(_12293_[0]),
    .A2(_11639_),
    .B1(_00558_),
    .C1(_11628_),
    .Y(_00559_));
 sky130_fd_sc_hd__a311oi_1 _21216_ (.A1(_11749_),
    .A2(_11628_),
    .A3(_11719_),
    .B1(_00557_),
    .C1(_00559_),
    .Y(_00560_));
 sky130_fd_sc_hd__nor2_4 _21217_ (.A(net3849),
    .B(_11815_),
    .Y(_00561_));
 sky130_fd_sc_hd__a211oi_1 _21218_ (.A1(_12304_[0]),
    .A2(_11819_),
    .B1(_00561_),
    .C1(_11746_),
    .Y(_00562_));
 sky130_fd_sc_hd__a2111oi_0 _21219_ (.A1(_00421_),
    .A2(_00556_),
    .B1(_00560_),
    .C1(_00562_),
    .D1(_11707_),
    .Y(_00563_));
 sky130_fd_sc_hd__o21ai_1 _21220_ (.A1(_00553_),
    .A2(_00555_),
    .B1(net3570),
    .Y(_00564_));
 sky130_fd_sc_hd__nand2_4 _21221_ (.A(_12299_[0]),
    .B(_11684_),
    .Y(_00565_));
 sky130_fd_sc_hd__a21oi_1 _21222_ (.A1(_11792_),
    .A2(_00541_),
    .B1(net3662),
    .Y(_00566_));
 sky130_fd_sc_hd__a311oi_1 _21223_ (.A1(net3664),
    .A2(_00435_),
    .A3(_00565_),
    .B1(_00566_),
    .C1(net3835),
    .Y(_00567_));
 sky130_fd_sc_hd__nor2_1 _21224_ (.A(_12302_[0]),
    .B(_11684_),
    .Y(_00568_));
 sky130_fd_sc_hd__nor2_2 _21225_ (.A(_12292_[0]),
    .B(_11655_),
    .Y(_00569_));
 sky130_fd_sc_hd__nor3_1 _21226_ (.A(net3662),
    .B(_00568_),
    .C(_00569_),
    .Y(_00570_));
 sky130_fd_sc_hd__a311oi_1 _21227_ (.A1(net3664),
    .A2(_00527_),
    .A3(_00430_),
    .B1(_00570_),
    .C1(net3841),
    .Y(_00571_));
 sky130_fd_sc_hd__nor3_1 _21228_ (.A(_11707_),
    .B(_00567_),
    .C(_00571_),
    .Y(_00572_));
 sky130_fd_sc_hd__o21ai_0 _21229_ (.A1(_12302_[0]),
    .A2(_11684_),
    .B1(_11769_),
    .Y(_00573_));
 sky130_fd_sc_hd__o32ai_1 _21230_ (.A1(_12293_[0]),
    .A2(net3663),
    .A3(net3839),
    .B1(_11796_),
    .B2(net3851),
    .Y(_00574_));
 sky130_fd_sc_hd__nand2_1 _21231_ (.A(_11707_),
    .B(net3835),
    .Y(_00575_));
 sky130_fd_sc_hd__a211oi_1 _21232_ (.A1(net3663),
    .A2(_00573_),
    .B1(_00574_),
    .C1(_00575_),
    .Y(_00576_));
 sky130_fd_sc_hd__a21oi_2 _21233_ (.A1(_12302_[0]),
    .A2(_11684_),
    .B1(_00454_),
    .Y(_00577_));
 sky130_fd_sc_hd__a211oi_1 _21234_ (.A1(_12297_[0]),
    .A2(_11684_),
    .B1(net3609),
    .C1(net3848),
    .Y(_00578_));
 sky130_fd_sc_hd__nand2_2 _21235_ (.A(_11707_),
    .B(net3841),
    .Y(_00579_));
 sky130_fd_sc_hd__a211oi_1 _21236_ (.A1(net3848),
    .A2(_00577_),
    .B1(_00578_),
    .C1(_00579_),
    .Y(_00580_));
 sky130_fd_sc_hd__o311a_1 _21237_ (.A1(_00572_),
    .A2(_00576_),
    .A3(_00580_),
    .B1(net3847),
    .C1(_11712_),
    .X(_00581_));
 sky130_fd_sc_hd__o21ai_1 _21238_ (.A1(net3609),
    .A2(_00515_),
    .B1(net3848),
    .Y(_00582_));
 sky130_fd_sc_hd__a21o_1 _21239_ (.A1(_00523_),
    .A2(_00552_),
    .B1(net3848),
    .X(_00583_));
 sky130_fd_sc_hd__nand2_1 _21240_ (.A(_12297_[0]),
    .B(_11663_),
    .Y(_00584_));
 sky130_fd_sc_hd__nor2_1 _21241_ (.A(net3851),
    .B(_11623_),
    .Y(_00585_));
 sky130_fd_sc_hd__o21ai_0 _21242_ (.A1(_00531_),
    .A2(_00585_),
    .B1(net3845),
    .Y(_00586_));
 sky130_fd_sc_hd__a21oi_1 _21243_ (.A1(_00584_),
    .A2(_00586_),
    .B1(net3835),
    .Y(_00587_));
 sky130_fd_sc_hd__a31oi_1 _21244_ (.A1(net3835),
    .A2(_00582_),
    .A3(_00583_),
    .B1(_00587_),
    .Y(_00588_));
 sky130_fd_sc_hd__nand2_1 _21245_ (.A(net3833),
    .B(_11784_),
    .Y(_00589_));
 sky130_fd_sc_hd__nand2_2 _21246_ (.A(net3663),
    .B(net3841),
    .Y(_00590_));
 sky130_fd_sc_hd__nand2_1 _21247_ (.A(net3848),
    .B(net3835),
    .Y(_00591_));
 sky130_fd_sc_hd__o21ai_0 _21248_ (.A1(net3851),
    .A2(_00590_),
    .B1(_00591_),
    .Y(_00592_));
 sky130_fd_sc_hd__o211ai_1 _21249_ (.A1(_11623_),
    .A2(net3835),
    .B1(net3663),
    .C1(net3665),
    .Y(_00593_));
 sky130_fd_sc_hd__o311ai_0 _21250_ (.A1(net3665),
    .A2(net3835),
    .A3(_00531_),
    .B1(_00593_),
    .C1(net3845),
    .Y(_00594_));
 sky130_fd_sc_hd__o21ai_0 _21251_ (.A1(net3845),
    .A2(_00592_),
    .B1(_00594_),
    .Y(_00595_));
 sky130_fd_sc_hd__a32oi_1 _21252_ (.A1(_12293_[0]),
    .A2(net3839),
    .A3(_00590_),
    .B1(_00531_),
    .B2(net3835),
    .Y(_00596_));
 sky130_fd_sc_hd__nand4_1 _21253_ (.A(net3833),
    .B(_00503_),
    .C(_00595_),
    .D(_00596_),
    .Y(_00597_));
 sky130_fd_sc_hd__o21ai_0 _21254_ (.A1(_00588_),
    .A2(_00589_),
    .B1(_00597_),
    .Y(_00598_));
 sky130_fd_sc_hd__a311oi_1 _21255_ (.A1(_11787_),
    .A2(_00551_),
    .A3(_00564_),
    .B1(_00581_),
    .C1(_00598_),
    .Y(_00115_));
 sky130_fd_sc_hd__a211oi_1 _21256_ (.A1(net3593),
    .A2(net3845),
    .B1(_11661_),
    .C1(net3662),
    .Y(_00599_));
 sky130_fd_sc_hd__a31oi_1 _21257_ (.A1(net3663),
    .A2(_11813_),
    .A3(_00540_),
    .B1(_00599_),
    .Y(_00600_));
 sky130_fd_sc_hd__nor2_1 _21258_ (.A(net3841),
    .B(_00600_),
    .Y(_00601_));
 sky130_fd_sc_hd__o21ai_0 _21259_ (.A1(_12292_[0]),
    .A2(_11628_),
    .B1(_11785_),
    .Y(_00602_));
 sky130_fd_sc_hd__a21boi_2 _21260_ (.A1(net3839),
    .A2(_00602_),
    .B1_N(_11692_),
    .Y(_00603_));
 sky130_fd_sc_hd__nand2_1 _21261_ (.A(_12292_[0]),
    .B(_11663_),
    .Y(_00604_));
 sky130_fd_sc_hd__nand2_2 _21262_ (.A(net3665),
    .B(_00433_),
    .Y(_00605_));
 sky130_fd_sc_hd__a21oi_1 _21263_ (.A1(net3851),
    .A2(net3848),
    .B1(_00575_),
    .Y(_00606_));
 sky130_fd_sc_hd__a311oi_1 _21264_ (.A1(_00604_),
    .A2(_00605_),
    .A3(_00606_),
    .B1(net3847),
    .C1(_11787_),
    .Y(_00607_));
 sky130_fd_sc_hd__nand3_2 _21265_ (.A(net3851),
    .B(net3849),
    .C(net3839),
    .Y(_00608_));
 sky130_fd_sc_hd__a21oi_1 _21266_ (.A1(net3665),
    .A2(_11819_),
    .B1(_00579_),
    .Y(_00609_));
 sky130_fd_sc_hd__nand3b_1 _21267_ (.A_N(_00561_),
    .B(_00608_),
    .C(_00609_),
    .Y(_00610_));
 sky130_fd_sc_hd__o311a_1 _21268_ (.A1(_11707_),
    .A2(_00601_),
    .A3(_00603_),
    .B1(_00607_),
    .C1(_00610_),
    .X(_00611_));
 sky130_fd_sc_hd__a21oi_1 _21269_ (.A1(_12299_[0]),
    .A2(net3848),
    .B1(_11734_),
    .Y(_00612_));
 sky130_fd_sc_hd__o211ai_1 _21270_ (.A1(net3836),
    .A2(_00612_),
    .B1(_11777_),
    .C1(net3840),
    .Y(_00613_));
 sky130_fd_sc_hd__nand3_1 _21271_ (.A(net3662),
    .B(_11715_),
    .C(_00446_),
    .Y(_00614_));
 sky130_fd_sc_hd__nor2_1 _21272_ (.A(_12297_[0]),
    .B(_11684_),
    .Y(_00615_));
 sky130_fd_sc_hd__o21ai_0 _21273_ (.A1(_00515_),
    .A2(_00615_),
    .B1(net3848),
    .Y(_00616_));
 sky130_fd_sc_hd__nand3_1 _21274_ (.A(_12306_[0]),
    .B(net4072),
    .C(_11654_),
    .Y(_00617_));
 sky130_fd_sc_hd__nand3_1 _21275_ (.A(_12293_[0]),
    .B(net3662),
    .C(_11684_),
    .Y(_00618_));
 sky130_fd_sc_hd__a21oi_1 _21276_ (.A1(_00617_),
    .A2(_00618_),
    .B1(net3835),
    .Y(_00619_));
 sky130_fd_sc_hd__a311oi_1 _21277_ (.A1(net3835),
    .A2(_11664_),
    .A3(_00616_),
    .B1(_00619_),
    .C1(_11707_),
    .Y(_00620_));
 sky130_fd_sc_hd__a31oi_1 _21278_ (.A1(_11707_),
    .A2(_00613_),
    .A3(_00614_),
    .B1(_00620_),
    .Y(_00621_));
 sky130_fd_sc_hd__and3_4 _21279_ (.A(_11787_),
    .B(net3847),
    .C(_00621_),
    .X(_00622_));
 sky130_fd_sc_hd__nand2_1 _21280_ (.A(_11768_),
    .B(_11796_),
    .Y(_00623_));
 sky130_fd_sc_hd__nand2_1 _21281_ (.A(net3848),
    .B(_00623_),
    .Y(_00624_));
 sky130_fd_sc_hd__o221ai_1 _21282_ (.A1(_12292_[0]),
    .A2(_11676_),
    .B1(_11688_),
    .B2(net3664),
    .C1(_00608_),
    .Y(_00625_));
 sky130_fd_sc_hd__nor2_1 _21283_ (.A(net3835),
    .B(_00625_),
    .Y(_00626_));
 sky130_fd_sc_hd__a41o_1 _21284_ (.A1(net3835),
    .A2(_11664_),
    .A3(_00605_),
    .A4(_00624_),
    .B1(_00626_),
    .X(_00627_));
 sky130_fd_sc_hd__o21ai_0 _21285_ (.A1(_12292_[0]),
    .A2(_11684_),
    .B1(_00565_),
    .Y(_00628_));
 sky130_fd_sc_hd__o21a_1 _21286_ (.A1(net3664),
    .A2(_00628_),
    .B1(_00467_),
    .X(_00629_));
 sky130_fd_sc_hd__o221ai_1 _21287_ (.A1(_11623_),
    .A2(_11815_),
    .B1(_00520_),
    .B2(net3848),
    .C1(net3841),
    .Y(_00630_));
 sky130_fd_sc_hd__o211ai_1 _21288_ (.A1(net3841),
    .A2(_00629_),
    .B1(_00630_),
    .C1(net3660),
    .Y(_00631_));
 sky130_fd_sc_hd__o2111a_1 _21289_ (.A1(net3660),
    .A2(_00627_),
    .B1(_00631_),
    .C1(net3833),
    .D1(_11787_),
    .X(_00632_));
 sky130_fd_sc_hd__nand2_2 _21290_ (.A(_11707_),
    .B(_11762_),
    .Y(_00633_));
 sky130_fd_sc_hd__o211ai_1 _21291_ (.A1(_12304_[0]),
    .A2(_11707_),
    .B1(_00633_),
    .C1(net3848),
    .Y(_00634_));
 sky130_fd_sc_hd__nor4_1 _21292_ (.A(net3848),
    .B(_11707_),
    .C(_11800_),
    .D(_00429_),
    .Y(_00635_));
 sky130_fd_sc_hd__a31oi_1 _21293_ (.A1(_12304_[0]),
    .A2(_11707_),
    .A3(net3839),
    .B1(_00635_),
    .Y(_00636_));
 sky130_fd_sc_hd__nand3_1 _21294_ (.A(net3848),
    .B(_00434_),
    .C(_00540_),
    .Y(_00637_));
 sky130_fd_sc_hd__nand3_1 _21295_ (.A(_11628_),
    .B(_00541_),
    .C(_00542_),
    .Y(_00638_));
 sky130_fd_sc_hd__a211oi_1 _21296_ (.A1(_00637_),
    .A2(_00638_),
    .B1(net3660),
    .C1(net3835),
    .Y(_00639_));
 sky130_fd_sc_hd__a311oi_1 _21297_ (.A1(net3663),
    .A2(_11813_),
    .A3(_11810_),
    .B1(_00579_),
    .C1(_00531_),
    .Y(_00640_));
 sky130_fd_sc_hd__a311oi_1 _21298_ (.A1(net3835),
    .A2(_00634_),
    .A3(_00636_),
    .B1(_00639_),
    .C1(_00640_),
    .Y(_00641_));
 sky130_fd_sc_hd__nor3_1 _21299_ (.A(_11787_),
    .B(_11719_),
    .C(_00641_),
    .Y(_00642_));
 sky130_fd_sc_hd__nor4_1 _21300_ (.A(_00611_),
    .B(_00622_),
    .C(_00632_),
    .D(_00642_),
    .Y(_00116_));
 sky130_fd_sc_hd__o21a_4 _21301_ (.A1(_11770_),
    .A2(_00444_),
    .B1(net3662),
    .X(_00643_));
 sky130_fd_sc_hd__a31oi_1 _21302_ (.A1(net3848),
    .A2(_00527_),
    .A3(_00541_),
    .B1(_00643_),
    .Y(_00644_));
 sky130_fd_sc_hd__o221ai_1 _21303_ (.A1(_11684_),
    .A2(_00425_),
    .B1(_11822_),
    .B2(_12308_[0]),
    .C1(net3847),
    .Y(_00645_));
 sky130_fd_sc_hd__o211ai_1 _21304_ (.A1(net3847),
    .A2(_00644_),
    .B1(_00645_),
    .C1(_11715_),
    .Y(_00646_));
 sky130_fd_sc_hd__nand2_2 _21305_ (.A(_12297_[0]),
    .B(_11696_),
    .Y(_00647_));
 sky130_fd_sc_hd__a221oi_1 _21306_ (.A1(_12302_[0]),
    .A2(_11684_),
    .B1(_00454_),
    .B2(net3848),
    .C1(_11639_),
    .Y(_00648_));
 sky130_fd_sc_hd__a311o_1 _21307_ (.A1(_11639_),
    .A2(_00548_),
    .A3(_00647_),
    .B1(_00648_),
    .C1(_11715_),
    .X(_00649_));
 sky130_fd_sc_hd__and3_1 _21308_ (.A(_00459_),
    .B(_00646_),
    .C(_00649_),
    .X(_00650_));
 sky130_fd_sc_hd__nand2_1 _21309_ (.A(_12304_[0]),
    .B(_11696_),
    .Y(_00651_));
 sky130_fd_sc_hd__nand2_1 _21310_ (.A(_00565_),
    .B(_00651_),
    .Y(_00652_));
 sky130_fd_sc_hd__a21oi_1 _21311_ (.A1(_12299_[0]),
    .A2(net3848),
    .B1(_00532_),
    .Y(_00653_));
 sky130_fd_sc_hd__o211ai_1 _21312_ (.A1(net3844),
    .A2(_00653_),
    .B1(_11786_),
    .C1(_11670_),
    .Y(_00654_));
 sky130_fd_sc_hd__o311a_1 _21313_ (.A1(_11670_),
    .A2(_11680_),
    .A3(_00652_),
    .B1(_00654_),
    .C1(_11639_),
    .X(_00655_));
 sky130_fd_sc_hd__nor2_1 _21314_ (.A(net3849),
    .B(_11822_),
    .Y(_00656_));
 sky130_fd_sc_hd__o21ai_0 _21315_ (.A1(_00543_),
    .A2(_00656_),
    .B1(_11670_),
    .Y(_00657_));
 sky130_fd_sc_hd__a21oi_1 _21316_ (.A1(_12297_[0]),
    .A2(net3838),
    .B1(net3848),
    .Y(_00658_));
 sky130_fd_sc_hd__a21oi_1 _21317_ (.A1(_12299_[0]),
    .A2(net3844),
    .B1(_00658_),
    .Y(_00659_));
 sky130_fd_sc_hd__nand2_1 _21318_ (.A(_11715_),
    .B(_00659_),
    .Y(_00660_));
 sky130_fd_sc_hd__and3_1 _21319_ (.A(net3833),
    .B(_00657_),
    .C(_00660_),
    .X(_00661_));
 sky130_fd_sc_hd__o21a_1 _21320_ (.A1(_00655_),
    .A2(_00661_),
    .B1(_11784_),
    .X(_00662_));
 sky130_fd_sc_hd__nor2_1 _21321_ (.A(net3849),
    .B(_11819_),
    .Y(_00663_));
 sky130_fd_sc_hd__nand2_1 _21322_ (.A(_12299_[0]),
    .B(net3661),
    .Y(_00664_));
 sky130_fd_sc_hd__o21ai_0 _21323_ (.A1(_12306_[0]),
    .A2(_11686_),
    .B1(_00664_),
    .Y(_00665_));
 sky130_fd_sc_hd__o21ai_0 _21324_ (.A1(_00663_),
    .A2(_00665_),
    .B1(net3841),
    .Y(_00666_));
 sky130_fd_sc_hd__o21ai_0 _21325_ (.A1(_11816_),
    .A2(_00643_),
    .B1(_11715_),
    .Y(_00667_));
 sky130_fd_sc_hd__nand3_1 _21326_ (.A(net3848),
    .B(_11809_),
    .C(_00435_),
    .Y(_00668_));
 sky130_fd_sc_hd__nand3_1 _21327_ (.A(net3664),
    .B(_00434_),
    .C(_00523_),
    .Y(_00669_));
 sky130_fd_sc_hd__a211oi_1 _21328_ (.A1(net3849),
    .A2(_00435_),
    .B1(_00561_),
    .C1(net3835),
    .Y(_00670_));
 sky130_fd_sc_hd__a311oi_1 _21329_ (.A1(net3835),
    .A2(_00668_),
    .A3(_00669_),
    .B1(_00670_),
    .C1(net3833),
    .Y(_00671_));
 sky130_fd_sc_hd__a311oi_1 _21330_ (.A1(net3833),
    .A2(_00666_),
    .A3(_00667_),
    .B1(_00671_),
    .C1(_11789_),
    .Y(_00672_));
 sky130_fd_sc_hd__nand3_1 _21331_ (.A(_11744_),
    .B(_00421_),
    .C(_00460_),
    .Y(_00673_));
 sky130_fd_sc_hd__nand3_1 _21332_ (.A(net3850),
    .B(_11628_),
    .C(_00497_),
    .Y(_00674_));
 sky130_fd_sc_hd__o21ai_0 _21333_ (.A1(net3849),
    .A2(_00557_),
    .B1(_00498_),
    .Y(_00675_));
 sky130_fd_sc_hd__o21ai_0 _21334_ (.A1(net3850),
    .A2(net3834),
    .B1(_11676_),
    .Y(_00676_));
 sky130_fd_sc_hd__a221oi_1 _21335_ (.A1(net3665),
    .A2(_00675_),
    .B1(_00676_),
    .B2(net3849),
    .C1(net3832),
    .Y(_00677_));
 sky130_fd_sc_hd__nand2_1 _21336_ (.A(_12294_[0]),
    .B(_11655_),
    .Y(_00678_));
 sky130_fd_sc_hd__a21oi_1 _21337_ (.A1(_11809_),
    .A2(_00678_),
    .B1(net3848),
    .Y(_00679_));
 sky130_fd_sc_hd__nor2_1 _21338_ (.A(net3665),
    .B(_11815_),
    .Y(_00680_));
 sky130_fd_sc_hd__o21ai_0 _21339_ (.A1(_00444_),
    .A2(_00569_),
    .B1(net3662),
    .Y(_00681_));
 sky130_fd_sc_hd__o211ai_1 _21340_ (.A1(_12293_[0]),
    .A2(_11686_),
    .B1(_11743_),
    .C1(_00681_),
    .Y(_00682_));
 sky130_fd_sc_hd__o311ai_0 _21341_ (.A1(_00468_),
    .A2(_00679_),
    .A3(_00680_),
    .B1(_00682_),
    .C1(_00503_),
    .Y(_00683_));
 sky130_fd_sc_hd__a31oi_1 _21342_ (.A1(_00673_),
    .A2(_00674_),
    .A3(_00677_),
    .B1(_00683_),
    .Y(_00684_));
 sky130_fd_sc_hd__or4_1 _21343_ (.A(_00650_),
    .B(_00662_),
    .C(_00672_),
    .D(_00684_),
    .X(_00117_));
 sky130_fd_sc_hd__nor2_1 _21344_ (.A(net3848),
    .B(_00508_),
    .Y(_00685_));
 sky130_fd_sc_hd__o221ai_1 _21345_ (.A1(net3849),
    .A2(_11686_),
    .B1(_00685_),
    .B2(net3851),
    .C1(_00647_),
    .Y(_00686_));
 sky130_fd_sc_hd__nand2_1 _21346_ (.A(_11639_),
    .B(_00686_),
    .Y(_00687_));
 sky130_fd_sc_hd__o21ai_0 _21347_ (.A1(_00543_),
    .A2(_00685_),
    .B1(net3833),
    .Y(_00688_));
 sky130_fd_sc_hd__nor2_1 _21348_ (.A(_12297_[0]),
    .B(net3848),
    .Y(_00689_));
 sky130_fd_sc_hd__nand2_1 _21349_ (.A(_12322_[0]),
    .B(net3839),
    .Y(_00690_));
 sky130_fd_sc_hd__o311ai_0 _21350_ (.A1(net3839),
    .A2(_00531_),
    .A3(_00689_),
    .B1(_00690_),
    .C1(_11719_),
    .Y(_00691_));
 sky130_fd_sc_hd__o2111ai_1 _21351_ (.A1(_12308_[0]),
    .A2(_11815_),
    .B1(_00608_),
    .C1(net3847),
    .D1(_11723_),
    .Y(_00692_));
 sky130_fd_sc_hd__a21oi_1 _21352_ (.A1(_00691_),
    .A2(_00692_),
    .B1(net3841),
    .Y(_00693_));
 sky130_fd_sc_hd__a311oi_2 _21353_ (.A1(net3841),
    .A2(_00687_),
    .A3(_00688_),
    .B1(_00693_),
    .C1(_11789_),
    .Y(_00694_));
 sky130_fd_sc_hd__o21ai_0 _21354_ (.A1(_00568_),
    .A2(_00466_),
    .B1(_11628_),
    .Y(_00695_));
 sky130_fd_sc_hd__o21ai_0 _21355_ (.A1(_12297_[0]),
    .A2(_11686_),
    .B1(_00695_),
    .Y(_00696_));
 sky130_fd_sc_hd__o211ai_1 _21356_ (.A1(_12293_[0]),
    .A2(_11628_),
    .B1(net3842),
    .C1(_00495_),
    .Y(_00697_));
 sky130_fd_sc_hd__o211ai_1 _21357_ (.A1(_12313_[0]),
    .A2(net3842),
    .B1(_00697_),
    .C1(net3846),
    .Y(_00698_));
 sky130_fd_sc_hd__o211ai_1 _21358_ (.A1(net3846),
    .A2(_00696_),
    .B1(_00698_),
    .C1(net3834),
    .Y(_00699_));
 sky130_fd_sc_hd__nand2_1 _21359_ (.A(net3662),
    .B(_00509_),
    .Y(_00700_));
 sky130_fd_sc_hd__o211ai_1 _21360_ (.A1(_11684_),
    .A2(_00488_),
    .B1(_00434_),
    .C1(net3848),
    .Y(_00701_));
 sky130_fd_sc_hd__nor3_1 _21361_ (.A(net3663),
    .B(_11771_),
    .C(_00515_),
    .Y(_00702_));
 sky130_fd_sc_hd__a211oi_1 _21362_ (.A1(net3663),
    .A2(_11662_),
    .B1(_00702_),
    .C1(_11746_),
    .Y(_00703_));
 sky130_fd_sc_hd__a31oi_1 _21363_ (.A1(_11743_),
    .A2(_00700_),
    .A3(_00701_),
    .B1(_00703_),
    .Y(_00704_));
 sky130_fd_sc_hd__and3_1 _21364_ (.A(_00503_),
    .B(_00699_),
    .C(_00704_),
    .X(_00705_));
 sky130_fd_sc_hd__a211oi_1 _21365_ (.A1(_12304_[0]),
    .A2(_11628_),
    .B1(net3836),
    .C1(_00477_),
    .Y(_00706_));
 sky130_fd_sc_hd__a21oi_2 _21366_ (.A1(_12312_[0]),
    .A2(net3836),
    .B1(_00706_),
    .Y(_00707_));
 sky130_fd_sc_hd__o21ai_0 _21367_ (.A1(_12293_[0]),
    .A2(_11686_),
    .B1(_11715_),
    .Y(_00708_));
 sky130_fd_sc_hd__o221ai_2 _21368_ (.A1(_11715_),
    .A2(_00707_),
    .B1(_00708_),
    .B2(_00553_),
    .C1(net3847),
    .Y(_00709_));
 sky130_fd_sc_hd__nor2_1 _21369_ (.A(_12299_[0]),
    .B(_00590_),
    .Y(_00710_));
 sky130_fd_sc_hd__nand2_1 _21370_ (.A(net3851),
    .B(_11715_),
    .Y(_00711_));
 sky130_fd_sc_hd__a21oi_1 _21371_ (.A1(_00423_),
    .A2(_00711_),
    .B1(_11628_),
    .Y(_00712_));
 sky130_fd_sc_hd__o21ai_0 _21372_ (.A1(_00710_),
    .A2(_00712_),
    .B1(_11684_),
    .Y(_00713_));
 sky130_fd_sc_hd__o311ai_0 _21373_ (.A1(net3848),
    .A2(_11670_),
    .A3(_00546_),
    .B1(_00713_),
    .C1(net3833),
    .Y(_00714_));
 sky130_fd_sc_hd__and3_1 _21374_ (.A(_00459_),
    .B(_00709_),
    .C(_00714_),
    .X(_00715_));
 sky130_fd_sc_hd__nor2_1 _21375_ (.A(net3843),
    .B(_00488_),
    .Y(_00716_));
 sky130_fd_sc_hd__o211ai_1 _21376_ (.A1(_11623_),
    .A2(net3838),
    .B1(_00542_),
    .C1(net3848),
    .Y(_00717_));
 sky130_fd_sc_hd__o31ai_1 _21377_ (.A1(net3848),
    .A2(net3609),
    .A3(_00716_),
    .B1(_00717_),
    .Y(_00718_));
 sky130_fd_sc_hd__o21ai_0 _21378_ (.A1(_12292_[0]),
    .A2(net3838),
    .B1(_00542_),
    .Y(_00719_));
 sky130_fd_sc_hd__a221oi_1 _21379_ (.A1(_12294_[0]),
    .A2(_11663_),
    .B1(_00719_),
    .B2(net3848),
    .C1(net3833),
    .Y(_00720_));
 sky130_fd_sc_hd__a21oi_1 _21380_ (.A1(net3833),
    .A2(_00718_),
    .B1(_00720_),
    .Y(_00721_));
 sky130_fd_sc_hd__a211oi_1 _21381_ (.A1(_12304_[0]),
    .A2(_11655_),
    .B1(_00445_),
    .C1(net3848),
    .Y(_00722_));
 sky130_fd_sc_hd__a211oi_1 _21382_ (.A1(_12294_[0]),
    .A2(_11684_),
    .B1(_00444_),
    .C1(_11628_),
    .Y(_00723_));
 sky130_fd_sc_hd__nand2_1 _21383_ (.A(net3851),
    .B(net3848),
    .Y(_00724_));
 sky130_fd_sc_hd__nand2_1 _21384_ (.A(net3665),
    .B(_11623_),
    .Y(_00725_));
 sky130_fd_sc_hd__nor3_1 _21385_ (.A(_12311_[0]),
    .B(_12320_[0]),
    .C(net3836),
    .Y(_00726_));
 sky130_fd_sc_hd__a311o_1 _21386_ (.A1(_11684_),
    .A2(_00724_),
    .A3(_00725_),
    .B1(_00726_),
    .C1(_11746_),
    .X(_00727_));
 sky130_fd_sc_hd__o311ai_4 _21387_ (.A1(_11750_),
    .A2(_00722_),
    .A3(_00723_),
    .B1(_00727_),
    .C1(_11784_),
    .Y(_00728_));
 sky130_fd_sc_hd__a21oi_1 _21388_ (.A1(net3834),
    .A2(_00721_),
    .B1(_00728_),
    .Y(_00729_));
 sky130_fd_sc_hd__nor4_1 _21389_ (.A(_00694_),
    .B(_00705_),
    .C(_00715_),
    .D(_00729_),
    .Y(_00118_));
 sky130_fd_sc_hd__nor2_1 _21390_ (.A(_12304_[0]),
    .B(_11822_),
    .Y(_00730_));
 sky130_fd_sc_hd__a311oi_1 _21391_ (.A1(net3848),
    .A2(_11813_),
    .A3(_00540_),
    .B1(_00730_),
    .C1(_11746_),
    .Y(_00731_));
 sky130_fd_sc_hd__nand2_1 _21392_ (.A(_11815_),
    .B(_11822_),
    .Y(_00732_));
 sky130_fd_sc_hd__a221o_1 _21393_ (.A1(net3849),
    .A2(net3661),
    .B1(_00732_),
    .B2(_00526_),
    .C1(_00507_),
    .X(_00733_));
 sky130_fd_sc_hd__nand2_1 _21394_ (.A(_11769_),
    .B(_00540_),
    .Y(_00734_));
 sky130_fd_sc_hd__nand3_1 _21395_ (.A(net3664),
    .B(_11813_),
    .C(_00523_),
    .Y(_00735_));
 sky130_fd_sc_hd__o211ai_1 _21396_ (.A1(net3664),
    .A2(_00734_),
    .B1(_00735_),
    .C1(_11743_),
    .Y(_00736_));
 sky130_fd_sc_hd__o21ai_0 _21397_ (.A1(_00468_),
    .A2(_00733_),
    .B1(_00736_),
    .Y(_00737_));
 sky130_fd_sc_hd__o21ai_0 _21398_ (.A1(_00433_),
    .A2(_00445_),
    .B1(net3662),
    .Y(_00738_));
 sky130_fd_sc_hd__o21ai_0 _21399_ (.A1(_00569_),
    .A2(_00615_),
    .B1(net3848),
    .Y(_00739_));
 sky130_fd_sc_hd__a211oi_1 _21400_ (.A1(_00738_),
    .A2(_00739_),
    .B1(_11719_),
    .C1(net3841),
    .Y(_00740_));
 sky130_fd_sc_hd__nor3_1 _21401_ (.A(_00731_),
    .B(_00737_),
    .C(_00740_),
    .Y(_00741_));
 sky130_fd_sc_hd__a21oi_1 _21402_ (.A1(_12294_[0]),
    .A2(net3661),
    .B1(_00445_),
    .Y(_00742_));
 sky130_fd_sc_hd__o211ai_1 _21403_ (.A1(_12297_[0]),
    .A2(_11684_),
    .B1(_00565_),
    .C1(net3848),
    .Y(_00743_));
 sky130_fd_sc_hd__nand3_1 _21404_ (.A(_11715_),
    .B(_00467_),
    .C(_00743_),
    .Y(_00744_));
 sky130_fd_sc_hd__o21ai_0 _21405_ (.A1(_11715_),
    .A2(_00742_),
    .B1(_00744_),
    .Y(_00745_));
 sky130_fd_sc_hd__nor3b_1 _21406_ (.A(_11734_),
    .B(net3836),
    .C_N(_11780_),
    .Y(_00746_));
 sky130_fd_sc_hd__o21ai_0 _21407_ (.A1(_12320_[0]),
    .A2(_11655_),
    .B1(_11743_),
    .Y(_00747_));
 sky130_fd_sc_hd__o311ai_0 _21408_ (.A1(net3662),
    .A2(_11800_),
    .A3(_00465_),
    .B1(_00442_),
    .C1(_11798_),
    .Y(_00748_));
 sky130_fd_sc_hd__o21ai_0 _21409_ (.A1(_00746_),
    .A2(_00747_),
    .B1(_00748_),
    .Y(_00749_));
 sky130_fd_sc_hd__a21oi_1 _21410_ (.A1(net3847),
    .A2(_00745_),
    .B1(_00749_),
    .Y(_00750_));
 sky130_fd_sc_hd__a21oi_1 _21411_ (.A1(net3848),
    .A2(_00497_),
    .B1(_11663_),
    .Y(_00751_));
 sky130_fd_sc_hd__o21ai_0 _21412_ (.A1(net3665),
    .A2(_00498_),
    .B1(_00557_),
    .Y(_00752_));
 sky130_fd_sc_hd__nor4_1 _21413_ (.A(_12306_[0]),
    .B(net3848),
    .C(net3834),
    .D(net3836),
    .Y(_00753_));
 sky130_fd_sc_hd__a311o_1 _21414_ (.A1(net3849),
    .A2(net3848),
    .A3(_00421_),
    .B1(_00753_),
    .C1(net3832),
    .X(_00754_));
 sky130_fd_sc_hd__a21oi_1 _21415_ (.A1(_11623_),
    .A2(_00752_),
    .B1(_00754_),
    .Y(_00755_));
 sky130_fd_sc_hd__o21ai_1 _21416_ (.A1(net3850),
    .A2(_00751_),
    .B1(_00755_),
    .Y(_00756_));
 sky130_fd_sc_hd__a21boi_0 _21417_ (.A1(_12297_[0]),
    .A2(_00421_),
    .B1_N(_00541_),
    .Y(_00757_));
 sky130_fd_sc_hd__a21o_4 _21418_ (.A1(_11676_),
    .A2(_00498_),
    .B1(_00453_),
    .X(_00758_));
 sky130_fd_sc_hd__o211ai_1 _21419_ (.A1(net3662),
    .A2(_00757_),
    .B1(_00758_),
    .C1(_00590_),
    .Y(_00759_));
 sky130_fd_sc_hd__a21oi_1 _21420_ (.A1(_11719_),
    .A2(_00759_),
    .B1(_11714_),
    .Y(_00760_));
 sky130_fd_sc_hd__a21oi_1 _21421_ (.A1(net3662),
    .A2(_00577_),
    .B1(_11746_),
    .Y(_00761_));
 sky130_fd_sc_hd__o211ai_1 _21422_ (.A1(_12304_[0]),
    .A2(_11655_),
    .B1(_00617_),
    .C1(net3662),
    .Y(_00762_));
 sky130_fd_sc_hd__o31ai_1 _21423_ (.A1(net3662),
    .A2(_00465_),
    .A3(_00547_),
    .B1(_00762_),
    .Y(_00763_));
 sky130_fd_sc_hd__a311oi_1 _21424_ (.A1(_11684_),
    .A2(_00724_),
    .A3(_00725_),
    .B1(_00429_),
    .C1(net3847),
    .Y(_00764_));
 sky130_fd_sc_hd__a21oi_1 _21425_ (.A1(net3847),
    .A2(_00763_),
    .B1(_00764_),
    .Y(_00765_));
 sky130_fd_sc_hd__o21ai_0 _21426_ (.A1(_12292_[0]),
    .A2(net3662),
    .B1(_11743_),
    .Y(_00766_));
 sky130_fd_sc_hd__nor3_1 _21427_ (.A(net3848),
    .B(_11762_),
    .C(_00515_),
    .Y(_00767_));
 sky130_fd_sc_hd__o21ai_0 _21428_ (.A1(_00766_),
    .A2(_00767_),
    .B1(_11784_),
    .Y(_00768_));
 sky130_fd_sc_hd__a221oi_1 _21429_ (.A1(_11811_),
    .A2(_00761_),
    .B1(_00765_),
    .B2(net3835),
    .C1(_00768_),
    .Y(_00769_));
 sky130_fd_sc_hd__a21oi_1 _21430_ (.A1(_00756_),
    .A2(_00760_),
    .B1(_00769_),
    .Y(_00770_));
 sky130_fd_sc_hd__o221ai_2 _21431_ (.A1(_11789_),
    .A2(_00741_),
    .B1(_00750_),
    .B2(_11713_),
    .C1(_00770_),
    .Y(_00119_));
 sky130_fd_sc_hd__xnor2_1 _21432_ (.A(\sa03_sr[1] ),
    .B(\sa32_sub[7] ),
    .Y(_00771_));
 sky130_fd_sc_hd__xnor2_1 _21433_ (.A(\sa10_sub[1] ),
    .B(\sa32_sub[0] ),
    .Y(_00772_));
 sky130_fd_sc_hd__xnor3_1 _21434_ (.A(\sa32_sub[1] ),
    .B(\sa21_sub[0] ),
    .C(\sa21_sub[7] ),
    .X(_00773_));
 sky130_fd_sc_hd__xnor3_1 _21435_ (.A(_00771_),
    .B(_00772_),
    .C(_00773_),
    .X(_00774_));
 sky130_fd_sc_hd__mux2i_2 _21436_ (.A0(\text_in_r[9] ),
    .A1(_00774_),
    .S(_05879_),
    .Y(_00775_));
 sky130_fd_sc_hd__xor2_4 _21437_ (.A(\u0.tmp_w[9] ),
    .B(_00775_),
    .X(_00776_));
 sky130_fd_sc_hd__clkinv_16 _21438_ (.A(_00776_),
    .Y(_00777_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_308 ();
 sky130_fd_sc_hd__xnor3_1 _21441_ (.A(net4211),
    .B(\sa21_sub[7] ),
    .C(net4179),
    .X(_00779_));
 sky130_fd_sc_hd__xor2_1 _21442_ (.A(_09925_),
    .B(_00779_),
    .X(_00780_));
 sky130_fd_sc_hd__nand2_1 _21443_ (.A(net4230),
    .B(\text_in_r[8] ),
    .Y(_00781_));
 sky130_fd_sc_hd__o21a_4 _21444_ (.A1(net4230),
    .A2(_00780_),
    .B1(_00781_),
    .X(_00782_));
 sky130_fd_sc_hd__xor2_4 _21445_ (.A(net4126),
    .B(_00782_),
    .X(_00783_));
 sky130_fd_sc_hd__clkinv_16 _21446_ (.A(_00783_),
    .Y(_00784_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_307 ();
 sky130_fd_sc_hd__xnor3_1 _21448_ (.A(\sa10_sub[2] ),
    .B(\sa32_sub[2] ),
    .C(net4222),
    .X(_00785_));
 sky130_fd_sc_hd__xor2_1 _21449_ (.A(net4194),
    .B(net4181),
    .X(_00786_));
 sky130_fd_sc_hd__nor2_1 _21450_ (.A(\u0.tmp_w[10] ),
    .B(net4230),
    .Y(_00787_));
 sky130_fd_sc_hd__nand2_1 _21451_ (.A(_00786_),
    .B(_00787_),
    .Y(_00788_));
 sky130_fd_sc_hd__nor2b_1 _21452_ (.A(net4230),
    .B_N(\u0.tmp_w[10] ),
    .Y(_00789_));
 sky130_fd_sc_hd__or3b_1 _21453_ (.A(_00786_),
    .B(_00785_),
    .C_N(_00789_),
    .X(_00790_));
 sky130_fd_sc_hd__nand3_1 _21454_ (.A(_00786_),
    .B(_00785_),
    .C(_00789_),
    .Y(_00791_));
 sky130_fd_sc_hd__nand3_1 _21455_ (.A(_07660_),
    .B(_00785_),
    .C(_00787_),
    .Y(_00792_));
 sky130_fd_sc_hd__o2111ai_2 _21456_ (.A1(_00785_),
    .A2(_00788_),
    .B1(_00790_),
    .C1(_00791_),
    .D1(_00792_),
    .Y(_00793_));
 sky130_fd_sc_hd__nand2b_1 _21457_ (.A_N(\u0.tmp_w[10] ),
    .B(net398),
    .Y(_00794_));
 sky130_fd_sc_hd__nand3_1 _21458_ (.A(\u0.tmp_w[10] ),
    .B(net398),
    .C(\text_in_r[10] ),
    .Y(_00795_));
 sky130_fd_sc_hd__o21ai_2 _21459_ (.A1(\text_in_r[10] ),
    .A2(_00794_),
    .B1(_00795_),
    .Y(_00796_));
 sky130_fd_sc_hd__nor2_4 _21460_ (.A(_00793_),
    .B(_00796_),
    .Y(_00797_));
 sky130_fd_sc_hd__clkinv_16 _21461_ (.A(_00797_),
    .Y(_00798_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_300 ();
 sky130_fd_sc_hd__xnor3_1 _21469_ (.A(\sa21_sub[5] ),
    .B(\sa32_sub[5] ),
    .C(\sa10_sub[6] ),
    .X(_00803_));
 sky130_fd_sc_hd__xor2_1 _21470_ (.A(_09941_),
    .B(_00803_),
    .X(_00804_));
 sky130_fd_sc_hd__mux2i_4 _21471_ (.A0(\text_in_r[14] ),
    .A1(_00804_),
    .S(net4116),
    .Y(_00805_));
 sky130_fd_sc_hd__xnor2_4 _21472_ (.A(\u0.tmp_w[14] ),
    .B(_00805_),
    .Y(_00806_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_298 ();
 sky130_fd_sc_hd__xor3_1 _21475_ (.A(\sa32_sub[6] ),
    .B(_07670_),
    .C(_09946_),
    .X(_00809_));
 sky130_fd_sc_hd__mux2i_4 _21476_ (.A0(\text_in_r[15] ),
    .A1(_00809_),
    .S(net4121),
    .Y(_00810_));
 sky130_fd_sc_hd__xnor2_4 _21477_ (.A(\u0.tmp_w[15] ),
    .B(_00810_),
    .Y(_00811_));
 sky130_fd_sc_hd__nand2_4 _21478_ (.A(net3826),
    .B(_00811_),
    .Y(_00812_));
 sky130_fd_sc_hd__xor2_1 _21479_ (.A(\sa32_sub[4] ),
    .B(\sa10_sub[5] ),
    .X(_00813_));
 sky130_fd_sc_hd__xnor2_2 _21480_ (.A(_09953_),
    .B(_00813_),
    .Y(_00814_));
 sky130_fd_sc_hd__mux2i_4 _21481_ (.A0(\text_in_r[13] ),
    .A1(_00814_),
    .S(net4121),
    .Y(_00815_));
 sky130_fd_sc_hd__xnor2_4 _21482_ (.A(\u0.tmp_w[13] ),
    .B(_00815_),
    .Y(_00816_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_297 ();
 sky130_fd_sc_hd__xnor2_1 _21484_ (.A(net4180),
    .B(net4179),
    .Y(_00818_));
 sky130_fd_sc_hd__xor3_1 _21485_ (.A(net4192),
    .B(\sa32_sub[4] ),
    .C(net4191),
    .X(_00819_));
 sky130_fd_sc_hd__xnor3_1 _21486_ (.A(_07701_),
    .B(_00818_),
    .C(_00819_),
    .X(_00820_));
 sky130_fd_sc_hd__mux2i_4 _21487_ (.A0(\text_in_r[12] ),
    .A1(_00820_),
    .S(net4116),
    .Y(_00821_));
 sky130_fd_sc_hd__xnor2_4 _21488_ (.A(\u0.tmp_w[12] ),
    .B(_00821_),
    .Y(_00822_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_295 ();
 sky130_fd_sc_hd__xnor2_1 _21491_ (.A(\sa03_sr[3] ),
    .B(net4179),
    .Y(_00825_));
 sky130_fd_sc_hd__xnor2_1 _21492_ (.A(\sa32_sub[2] ),
    .B(\sa10_sub[3] ),
    .Y(_00826_));
 sky130_fd_sc_hd__xnor3_1 _21493_ (.A(_09964_),
    .B(_00825_),
    .C(_00826_),
    .X(_00827_));
 sky130_fd_sc_hd__nand2b_1 _21494_ (.A_N(\text_in_r[11] ),
    .B(net4230),
    .Y(_00828_));
 sky130_fd_sc_hd__o21a_4 _21495_ (.A1(net398),
    .A2(_00827_),
    .B1(_00828_),
    .X(_00829_));
 sky130_fd_sc_hd__xor2_4 _21496_ (.A(\u0.tmp_w[11] ),
    .B(_00829_),
    .X(_00830_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_294 ();
 sky130_fd_sc_hd__nand2_8 _21498_ (.A(net3827),
    .B(net3811),
    .Y(_00832_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_293 ();
 sky130_fd_sc_hd__clkinvlp_4 _21500_ (.A(_12330_[0]),
    .Y(_00834_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_292 ();
 sky130_fd_sc_hd__mux2i_2 _21502_ (.A0(_00834_),
    .A1(_12328_[0]),
    .S(_00798_),
    .Y(_00836_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_291 ();
 sky130_fd_sc_hd__o22ai_2 _21504_ (.A1(_12335_[0]),
    .A2(_00832_),
    .B1(_00836_),
    .B2(net3816),
    .Y(_00838_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_290 ();
 sky130_fd_sc_hd__nor2_2 _21506_ (.A(_12338_[0]),
    .B(net3827),
    .Y(_00840_));
 sky130_fd_sc_hd__nor2_4 _21507_ (.A(net3830),
    .B(_00798_),
    .Y(_00841_));
 sky130_fd_sc_hd__o21ai_2 _21508_ (.A1(_00840_),
    .A2(_00841_),
    .B1(net3818),
    .Y(_00842_));
 sky130_fd_sc_hd__xnor2_4 _21509_ (.A(\u0.tmp_w[11] ),
    .B(_00829_),
    .Y(_00843_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_289 ();
 sky130_fd_sc_hd__nand2_4 _21511_ (.A(net3659),
    .B(net3827),
    .Y(_00845_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_288 ();
 sky130_fd_sc_hd__nand2_1 _21513_ (.A(_12329_[0]),
    .B(_00798_),
    .Y(_00847_));
 sky130_fd_sc_hd__a31oi_1 _21514_ (.A1(net3807),
    .A2(_00845_),
    .A3(_00847_),
    .B1(net3821),
    .Y(_00848_));
 sky130_fd_sc_hd__a22o_1 _21515_ (.A1(net3821),
    .A2(_00838_),
    .B1(_00842_),
    .B2(_00848_),
    .X(_00849_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_285 ();
 sky130_fd_sc_hd__inv_8 _21519_ (.A(_12329_[0]),
    .Y(_00853_));
 sky130_fd_sc_hd__nand2_1 _21520_ (.A(_00853_),
    .B(_00822_),
    .Y(_00854_));
 sky130_fd_sc_hd__xor2_4 _21521_ (.A(\u0.tmp_w[12] ),
    .B(_00821_),
    .X(_00855_));
 sky130_fd_sc_hd__nand2_1 _21522_ (.A(_12342_[0]),
    .B(_00855_),
    .Y(_00856_));
 sky130_fd_sc_hd__nor2_4 _21523_ (.A(_00855_),
    .B(net3819),
    .Y(_00857_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_284 ();
 sky130_fd_sc_hd__a32o_1 _21525_ (.A1(net3819),
    .A2(_00854_),
    .A3(_00856_),
    .B1(_00857_),
    .B2(_12340_[0]),
    .X(_00859_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_282 ();
 sky130_fd_sc_hd__nor2_4 _21528_ (.A(_00784_),
    .B(_00843_),
    .Y(_00862_));
 sky130_fd_sc_hd__nand2_1 _21529_ (.A(net3806),
    .B(_00862_),
    .Y(_00863_));
 sky130_fd_sc_hd__nor2_4 _21530_ (.A(_12335_[0]),
    .B(net3817),
    .Y(_00864_));
 sky130_fd_sc_hd__nor2_1 _21531_ (.A(net3827),
    .B(_00864_),
    .Y(_00865_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_281 ();
 sky130_fd_sc_hd__a221oi_2 _21533_ (.A1(net3827),
    .A2(_00859_),
    .B1(_00863_),
    .B2(_00865_),
    .C1(_00816_),
    .Y(_00867_));
 sky130_fd_sc_hd__a21oi_1 _21534_ (.A1(net3824),
    .A2(_00849_),
    .B1(_00867_),
    .Y(_00868_));
 sky130_fd_sc_hd__nor2_1 _21535_ (.A(_00812_),
    .B(_00868_),
    .Y(_00869_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_280 ();
 sky130_fd_sc_hd__nand2_8 _21537_ (.A(net3657),
    .B(net3819),
    .Y(_00871_));
 sky130_fd_sc_hd__nand2_2 _21538_ (.A(_12330_[0]),
    .B(net3807),
    .Y(_00872_));
 sky130_fd_sc_hd__a21oi_1 _21539_ (.A1(_00871_),
    .A2(_00872_),
    .B1(net3828),
    .Y(_00873_));
 sky130_fd_sc_hd__nor2_2 _21540_ (.A(_12328_[0]),
    .B(_00832_),
    .Y(_00874_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_279 ();
 sky130_fd_sc_hd__nand2b_4 _21542_ (.A_N(_12335_[0]),
    .B(_00798_),
    .Y(_00876_));
 sky130_fd_sc_hd__nand2_2 _21543_ (.A(_12333_[0]),
    .B(net3827),
    .Y(_00877_));
 sky130_fd_sc_hd__a31oi_4 _21544_ (.A1(net3807),
    .A2(_00876_),
    .A3(_00877_),
    .B1(net3821),
    .Y(_00878_));
 sky130_fd_sc_hd__nor3b_1 _21545_ (.A(_00873_),
    .B(_00874_),
    .C_N(_00878_),
    .Y(_00879_));
 sky130_fd_sc_hd__nor2_4 _21546_ (.A(net3827),
    .B(net3811),
    .Y(_00880_));
 sky130_fd_sc_hd__a221oi_1 _21547_ (.A1(_12351_[0]),
    .A2(net3811),
    .B1(_00880_),
    .B2(_12329_[0]),
    .C1(net3805),
    .Y(_00881_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_277 ();
 sky130_fd_sc_hd__nand2_8 _21550_ (.A(_12340_[0]),
    .B(net3810),
    .Y(_00884_));
 sky130_fd_sc_hd__nor2_1 _21551_ (.A(net3827),
    .B(_00884_),
    .Y(_00885_));
 sky130_fd_sc_hd__and2_0 _21552_ (.A(net398),
    .B(\text_in_r[11] ),
    .X(_00886_));
 sky130_fd_sc_hd__a211oi_1 _21553_ (.A1(net4121),
    .A2(_00827_),
    .B1(_00886_),
    .C1(\u0.tmp_w[11] ),
    .Y(_00887_));
 sky130_fd_sc_hd__o211ai_1 _21554_ (.A1(net398),
    .A2(_00827_),
    .B1(_00828_),
    .C1(\u0.tmp_w[11] ),
    .Y(_00888_));
 sky130_fd_sc_hd__nand3b_1 _21555_ (.A_N(_00887_),
    .B(_12333_[0]),
    .C(_00888_),
    .Y(_00889_));
 sky130_fd_sc_hd__o21ai_1 _21556_ (.A1(_12330_[0]),
    .A2(net3811),
    .B1(net3579),
    .Y(_00890_));
 sky130_fd_sc_hd__nor2_1 _21557_ (.A(_00798_),
    .B(_00890_),
    .Y(_00891_));
 sky130_fd_sc_hd__nand2_8 _21558_ (.A(_00798_),
    .B(net3809),
    .Y(_00892_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_276 ();
 sky130_fd_sc_hd__nand2_4 _21560_ (.A(_12333_[0]),
    .B(net3807),
    .Y(_00894_));
 sky130_fd_sc_hd__nand2_2 _21561_ (.A(_00834_),
    .B(net3815),
    .Y(_00895_));
 sky130_fd_sc_hd__a31oi_2 _21562_ (.A1(net3827),
    .A2(_00894_),
    .A3(_00895_),
    .B1(_00855_),
    .Y(_00896_));
 sky130_fd_sc_hd__o21ai_2 _21563_ (.A1(_12338_[0]),
    .A2(_00892_),
    .B1(_00896_),
    .Y(_00897_));
 sky130_fd_sc_hd__o311ai_0 _21564_ (.A1(net3821),
    .A2(_00885_),
    .A3(_00891_),
    .B1(_00897_),
    .C1(net3824),
    .Y(_00898_));
 sky130_fd_sc_hd__xor2_4 _21565_ (.A(\u0.tmp_w[15] ),
    .B(_00810_),
    .X(_00899_));
 sky130_fd_sc_hd__nor2_4 _21566_ (.A(_00806_),
    .B(_00899_),
    .Y(_00900_));
 sky130_fd_sc_hd__o311a_1 _21567_ (.A1(net3824),
    .A2(_00879_),
    .A3(_00881_),
    .B1(_00898_),
    .C1(_00900_),
    .X(_00901_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_275 ();
 sky130_fd_sc_hd__xor2_4 _21569_ (.A(\u0.tmp_w[13] ),
    .B(_00815_),
    .X(_00903_));
 sky130_fd_sc_hd__o21ai_0 _21570_ (.A1(net3657),
    .A2(_00903_),
    .B1(net3827),
    .Y(_00904_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_274 ();
 sky130_fd_sc_hd__nor2_2 _21572_ (.A(net3830),
    .B(net3827),
    .Y(_00905_));
 sky130_fd_sc_hd__nor3_1 _21573_ (.A(_00853_),
    .B(_00798_),
    .C(_00816_),
    .Y(_00906_));
 sky130_fd_sc_hd__a221oi_1 _21574_ (.A1(_00777_),
    .A2(_00904_),
    .B1(_00905_),
    .B2(_00816_),
    .C1(_00906_),
    .Y(_00907_));
 sky130_fd_sc_hd__nor3_1 _21575_ (.A(_12329_[0]),
    .B(net3827),
    .C(_00816_),
    .Y(_00908_));
 sky130_fd_sc_hd__nand2_1 _21576_ (.A(net3814),
    .B(_00908_),
    .Y(_00909_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_273 ();
 sky130_fd_sc_hd__nand2_8 _21578_ (.A(net3658),
    .B(net3827),
    .Y(_00911_));
 sky130_fd_sc_hd__nand2_1 _21579_ (.A(net3831),
    .B(net3830),
    .Y(_00912_));
 sky130_fd_sc_hd__nand2_1 _21580_ (.A(_00911_),
    .B(_00912_),
    .Y(_00913_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_272 ();
 sky130_fd_sc_hd__a31oi_1 _21582_ (.A1(_00816_),
    .A2(net3818),
    .A3(_00913_),
    .B1(_00855_),
    .Y(_00915_));
 sky130_fd_sc_hd__o211ai_1 _21583_ (.A1(net3814),
    .A2(_00907_),
    .B1(_00909_),
    .C1(_00915_),
    .Y(_00916_));
 sky130_fd_sc_hd__nor2_4 _21584_ (.A(_00798_),
    .B(_00830_),
    .Y(_00917_));
 sky130_fd_sc_hd__nor2_4 _21585_ (.A(net3827),
    .B(net3807),
    .Y(_00918_));
 sky130_fd_sc_hd__nor2_4 _21586_ (.A(_00917_),
    .B(_00918_),
    .Y(_00919_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_270 ();
 sky130_fd_sc_hd__nor2_1 _21589_ (.A(_00853_),
    .B(net3807),
    .Y(_00922_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_269 ();
 sky130_fd_sc_hd__nand2_4 _21591_ (.A(_00903_),
    .B(net3806),
    .Y(_00924_));
 sky130_fd_sc_hd__a21oi_1 _21592_ (.A1(net3827),
    .A2(_00922_),
    .B1(_00924_),
    .Y(_00925_));
 sky130_fd_sc_hd__o221ai_1 _21593_ (.A1(_12338_[0]),
    .A2(_00892_),
    .B1(_00919_),
    .B2(_12328_[0]),
    .C1(_00925_),
    .Y(_00926_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_267 ();
 sky130_fd_sc_hd__nor2_2 _21596_ (.A(_12338_[0]),
    .B(net3807),
    .Y(_00929_));
 sky130_fd_sc_hd__nor2_1 _21597_ (.A(_00853_),
    .B(net3813),
    .Y(_00930_));
 sky130_fd_sc_hd__nor3_1 _21598_ (.A(_00798_),
    .B(_00929_),
    .C(_00930_),
    .Y(_00931_));
 sky130_fd_sc_hd__nor2_1 _21599_ (.A(_12328_[0]),
    .B(net3807),
    .Y(_00932_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_266 ();
 sky130_fd_sc_hd__nor2_2 _21601_ (.A(_12342_[0]),
    .B(net3816),
    .Y(_00934_));
 sky130_fd_sc_hd__nor3_1 _21602_ (.A(net3827),
    .B(_00932_),
    .C(_00934_),
    .Y(_00935_));
 sky130_fd_sc_hd__nor2_4 _21603_ (.A(_00903_),
    .B(net3823),
    .Y(_00936_));
 sky130_fd_sc_hd__o21ai_0 _21604_ (.A1(_00931_),
    .A2(_00935_),
    .B1(_00936_),
    .Y(_00937_));
 sky130_fd_sc_hd__xor2_4 _21605_ (.A(\u0.tmp_w[14] ),
    .B(_00805_),
    .X(_00938_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_265 ();
 sky130_fd_sc_hd__nand2_8 _21607_ (.A(net3803),
    .B(_00899_),
    .Y(_00940_));
 sky130_fd_sc_hd__a31oi_2 _21608_ (.A1(_00916_),
    .A2(_00926_),
    .A3(_00937_),
    .B1(_00940_),
    .Y(_00941_));
 sky130_fd_sc_hd__nand2_4 _21609_ (.A(_00777_),
    .B(net3809),
    .Y(_00942_));
 sky130_fd_sc_hd__nor2_4 _21610_ (.A(net3825),
    .B(net3806),
    .Y(_00943_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_264 ();
 sky130_fd_sc_hd__nand2_2 _21612_ (.A(_12344_[0]),
    .B(net3811),
    .Y(_00945_));
 sky130_fd_sc_hd__nand4_1 _21613_ (.A(net3828),
    .B(_00942_),
    .C(_00943_),
    .D(_00945_),
    .Y(_00946_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_263 ();
 sky130_fd_sc_hd__nor2_1 _21615_ (.A(_00816_),
    .B(net3822),
    .Y(_00948_));
 sky130_fd_sc_hd__nor2_1 _21616_ (.A(_12330_[0]),
    .B(_00798_),
    .Y(_00949_));
 sky130_fd_sc_hd__nand2_4 _21617_ (.A(net3659),
    .B(_00798_),
    .Y(_00950_));
 sky130_fd_sc_hd__inv_4 _21618_ (.A(_00950_),
    .Y(_00951_));
 sky130_fd_sc_hd__or3_4 _21619_ (.A(net3813),
    .B(_00949_),
    .C(_00951_),
    .X(_00952_));
 sky130_fd_sc_hd__nor2_2 _21620_ (.A(_12342_[0]),
    .B(_00798_),
    .Y(_00953_));
 sky130_fd_sc_hd__o21ai_2 _21621_ (.A1(_00905_),
    .A2(_00953_),
    .B1(net3813),
    .Y(_00954_));
 sky130_fd_sc_hd__nand3_1 _21622_ (.A(_00948_),
    .B(_00952_),
    .C(_00954_),
    .Y(_00955_));
 sky130_fd_sc_hd__nor2_4 _21623_ (.A(net3657),
    .B(_00892_),
    .Y(_00956_));
 sky130_fd_sc_hd__o22ai_1 _21624_ (.A1(_12335_[0]),
    .A2(_00832_),
    .B1(net3579),
    .B2(net3828),
    .Y(_00957_));
 sky130_fd_sc_hd__o21ai_0 _21625_ (.A1(_00956_),
    .A2(_00957_),
    .B1(_00936_),
    .Y(_00958_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_262 ();
 sky130_fd_sc_hd__nand2b_1 _21627_ (.A_N(_12333_[0]),
    .B(net3807),
    .Y(_00960_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_261 ();
 sky130_fd_sc_hd__nor2_2 _21629_ (.A(net3830),
    .B(net3807),
    .Y(_00962_));
 sky130_fd_sc_hd__nand2_4 _21630_ (.A(_00903_),
    .B(net3821),
    .Y(_00963_));
 sky130_fd_sc_hd__nand2_8 _21631_ (.A(_12329_[0]),
    .B(net3811),
    .Y(_00964_));
 sky130_fd_sc_hd__nand2_8 _21632_ (.A(_00784_),
    .B(net3807),
    .Y(_00965_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_260 ();
 sky130_fd_sc_hd__a21oi_1 _21634_ (.A1(_00964_),
    .A2(_00965_),
    .B1(_00798_),
    .Y(_00967_));
 sky130_fd_sc_hd__nand2_2 _21635_ (.A(_12344_[0]),
    .B(_00798_),
    .Y(_00968_));
 sky130_fd_sc_hd__nor2_4 _21636_ (.A(_00903_),
    .B(net3805),
    .Y(_00969_));
 sky130_fd_sc_hd__o21ai_0 _21637_ (.A1(_00843_),
    .A2(_00968_),
    .B1(_00969_),
    .Y(_00970_));
 sky130_fd_sc_hd__o32ai_1 _21638_ (.A1(net3828),
    .A2(_00962_),
    .A3(_00963_),
    .B1(_00967_),
    .B2(_00970_),
    .Y(_00971_));
 sky130_fd_sc_hd__o21ai_0 _21639_ (.A1(net3828),
    .A2(_00960_),
    .B1(_00971_),
    .Y(_00972_));
 sky130_fd_sc_hd__nand2_2 _21640_ (.A(_00806_),
    .B(_00899_),
    .Y(_00973_));
 sky130_fd_sc_hd__a41oi_1 _21641_ (.A1(_00946_),
    .A2(_00955_),
    .A3(_00958_),
    .A4(_00972_),
    .B1(_00973_),
    .Y(_00974_));
 sky130_fd_sc_hd__nor4_2 _21642_ (.A(_00869_),
    .B(_00901_),
    .C(_00941_),
    .D(_00974_),
    .Y(_00120_));
 sky130_fd_sc_hd__nor2_4 _21643_ (.A(net3830),
    .B(net3818),
    .Y(_00975_));
 sky130_fd_sc_hd__nor2_2 _21644_ (.A(_12342_[0]),
    .B(net3809),
    .Y(_00976_));
 sky130_fd_sc_hd__o21ai_0 _21645_ (.A1(_00975_),
    .A2(_00976_),
    .B1(net3827),
    .Y(_00977_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_259 ();
 sky130_fd_sc_hd__nand2_4 _21647_ (.A(_12328_[0]),
    .B(net3809),
    .Y(_00979_));
 sky130_fd_sc_hd__nand3_1 _21648_ (.A(_00798_),
    .B(_00979_),
    .C(net3579),
    .Y(_00980_));
 sky130_fd_sc_hd__nand2_8 _21649_ (.A(_00816_),
    .B(net3823),
    .Y(_00981_));
 sky130_fd_sc_hd__a21oi_1 _21650_ (.A1(_00977_),
    .A2(_00980_),
    .B1(_00981_),
    .Y(_00982_));
 sky130_fd_sc_hd__nand2b_2 _21651_ (.A_N(_12335_[0]),
    .B(net3817),
    .Y(_00983_));
 sky130_fd_sc_hd__a21oi_1 _21652_ (.A1(_00983_),
    .A2(_00965_),
    .B1(_00798_),
    .Y(_00984_));
 sky130_fd_sc_hd__nand2_1 _21653_ (.A(net3831),
    .B(net3813),
    .Y(_00985_));
 sky130_fd_sc_hd__a21oi_2 _21654_ (.A1(_00942_),
    .A2(_00985_),
    .B1(net3827),
    .Y(_00986_));
 sky130_fd_sc_hd__nor3_1 _21655_ (.A(_00963_),
    .B(_00984_),
    .C(_00986_),
    .Y(_00987_));
 sky130_fd_sc_hd__o21ai_0 _21656_ (.A1(_00840_),
    .A2(_00953_),
    .B1(net3809),
    .Y(_00988_));
 sky130_fd_sc_hd__o31ai_1 _21657_ (.A1(_12354_[0]),
    .A2(_00816_),
    .A3(net3809),
    .B1(_00988_),
    .Y(_00989_));
 sky130_fd_sc_hd__a21o_1 _21658_ (.A1(_00855_),
    .A2(_00989_),
    .B1(_00940_),
    .X(_00990_));
 sky130_fd_sc_hd__nand3_1 _21659_ (.A(_00806_),
    .B(_00899_),
    .C(_00903_),
    .Y(_00991_));
 sky130_fd_sc_hd__nand2_8 _21660_ (.A(_00853_),
    .B(net3817),
    .Y(_00992_));
 sky130_fd_sc_hd__nand2_8 _21661_ (.A(_12344_[0]),
    .B(_00843_),
    .Y(_00993_));
 sky130_fd_sc_hd__nand2_2 _21662_ (.A(_00834_),
    .B(net3809),
    .Y(_00994_));
 sky130_fd_sc_hd__nand2_4 _21663_ (.A(_12342_[0]),
    .B(net3819),
    .Y(_00995_));
 sky130_fd_sc_hd__a21oi_1 _21664_ (.A1(_00994_),
    .A2(_00995_),
    .B1(net3827),
    .Y(_00996_));
 sky130_fd_sc_hd__a311oi_1 _21665_ (.A1(net3827),
    .A2(_00992_),
    .A3(_00993_),
    .B1(_00996_),
    .C1(_00855_),
    .Y(_00997_));
 sky130_fd_sc_hd__nand2_4 _21666_ (.A(_12342_[0]),
    .B(net3808),
    .Y(_00998_));
 sky130_fd_sc_hd__a21oi_1 _21667_ (.A1(_00992_),
    .A2(_00998_),
    .B1(_00798_),
    .Y(_00999_));
 sky130_fd_sc_hd__nor3_1 _21668_ (.A(net3823),
    .B(_00956_),
    .C(_00999_),
    .Y(_01000_));
 sky130_fd_sc_hd__or3_4 _21669_ (.A(_00991_),
    .B(_00997_),
    .C(_01000_),
    .X(_01001_));
 sky130_fd_sc_hd__o31ai_1 _21670_ (.A1(_00982_),
    .A2(_00987_),
    .A3(_00990_),
    .B1(_01001_),
    .Y(_01002_));
 sky130_fd_sc_hd__nor2_1 _21671_ (.A(net3657),
    .B(_00919_),
    .Y(_01003_));
 sky130_fd_sc_hd__o22ai_1 _21672_ (.A1(_00853_),
    .A2(_00892_),
    .B1(_00871_),
    .B2(_00777_),
    .Y(_01004_));
 sky130_fd_sc_hd__o21ai_0 _21673_ (.A1(_01003_),
    .A2(_01004_),
    .B1(_00855_),
    .Y(_01005_));
 sky130_fd_sc_hd__nand3_1 _21674_ (.A(net3827),
    .B(_00979_),
    .C(_00964_),
    .Y(_01006_));
 sky130_fd_sc_hd__nand2_4 _21675_ (.A(_12335_[0]),
    .B(net3813),
    .Y(_01007_));
 sky130_fd_sc_hd__a21oi_1 _21676_ (.A1(_00965_),
    .A2(_01007_),
    .B1(net3827),
    .Y(_01008_));
 sky130_fd_sc_hd__nor2_1 _21677_ (.A(net3806),
    .B(_01008_),
    .Y(_01009_));
 sky130_fd_sc_hd__a21oi_1 _21678_ (.A1(_01006_),
    .A2(_01009_),
    .B1(net3825),
    .Y(_01010_));
 sky130_fd_sc_hd__nand2_2 _21679_ (.A(_12344_[0]),
    .B(_00918_),
    .Y(_01011_));
 sky130_fd_sc_hd__nor2_4 _21680_ (.A(net3831),
    .B(net3807),
    .Y(_01012_));
 sky130_fd_sc_hd__o21ai_0 _21681_ (.A1(_00934_),
    .A2(_01012_),
    .B1(net3827),
    .Y(_01013_));
 sky130_fd_sc_hd__nor3_2 _21682_ (.A(_12329_[0]),
    .B(_00798_),
    .C(net3808),
    .Y(_01014_));
 sky130_fd_sc_hd__nand2_1 _21683_ (.A(_00798_),
    .B(net3813),
    .Y(_01015_));
 sky130_fd_sc_hd__nand2_1 _21684_ (.A(_12335_[0]),
    .B(net3827),
    .Y(_01016_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_258 ();
 sky130_fd_sc_hd__o22ai_1 _21686_ (.A1(_12342_[0]),
    .A2(_01015_),
    .B1(_01016_),
    .B2(net3811),
    .Y(_01018_));
 sky130_fd_sc_hd__nor3_1 _21687_ (.A(net3821),
    .B(_01014_),
    .C(_01018_),
    .Y(_01019_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_257 ();
 sky130_fd_sc_hd__a311oi_2 _21689_ (.A1(net3822),
    .A2(_01011_),
    .A3(_01013_),
    .B1(_01019_),
    .C1(net3804),
    .Y(_01021_));
 sky130_fd_sc_hd__a211oi_1 _21690_ (.A1(_01005_),
    .A2(_01010_),
    .B1(_01021_),
    .C1(_00812_),
    .Y(_01022_));
 sky130_fd_sc_hd__nand2_2 _21691_ (.A(_12344_[0]),
    .B(net3827),
    .Y(_01023_));
 sky130_fd_sc_hd__a21o_1 _21692_ (.A1(_00847_),
    .A2(_01023_),
    .B1(net3807),
    .X(_01024_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_256 ();
 sky130_fd_sc_hd__o21ai_0 _21694_ (.A1(_12358_[0]),
    .A2(net3807),
    .B1(net3821),
    .Y(_01026_));
 sky130_fd_sc_hd__a31oi_1 _21695_ (.A1(net3807),
    .A2(_00845_),
    .A3(_00876_),
    .B1(_01026_),
    .Y(_01027_));
 sky130_fd_sc_hd__a21oi_1 _21696_ (.A1(_00878_),
    .A2(_01024_),
    .B1(_01027_),
    .Y(_01028_));
 sky130_fd_sc_hd__nor2_4 _21697_ (.A(net3831),
    .B(net3816),
    .Y(_01029_));
 sky130_fd_sc_hd__nor2_1 _21698_ (.A(_12333_[0]),
    .B(net3807),
    .Y(_01030_));
 sky130_fd_sc_hd__o21ai_0 _21699_ (.A1(_01029_),
    .A2(_01030_),
    .B1(_00798_),
    .Y(_01031_));
 sky130_fd_sc_hd__o211ai_1 _21700_ (.A1(_00777_),
    .A2(_00965_),
    .B1(_01031_),
    .C1(_00936_),
    .Y(_01032_));
 sky130_fd_sc_hd__nand2_4 _21701_ (.A(_12335_[0]),
    .B(net3807),
    .Y(_01033_));
 sky130_fd_sc_hd__nand3_1 _21702_ (.A(net3827),
    .B(_00964_),
    .C(_01033_),
    .Y(_01034_));
 sky130_fd_sc_hd__o21ai_0 _21703_ (.A1(_00862_),
    .A2(_00975_),
    .B1(_00798_),
    .Y(_01035_));
 sky130_fd_sc_hd__a21o_1 _21704_ (.A1(_01034_),
    .A2(_01035_),
    .B1(_00981_),
    .X(_01036_));
 sky130_fd_sc_hd__o211ai_1 _21705_ (.A1(net3825),
    .A2(_01028_),
    .B1(_01032_),
    .C1(_01036_),
    .Y(_01037_));
 sky130_fd_sc_hd__nor2_4 _21706_ (.A(_00938_),
    .B(_00811_),
    .Y(_01038_));
 sky130_fd_sc_hd__nand2_4 _21707_ (.A(net3824),
    .B(_01038_),
    .Y(_01039_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_255 ();
 sky130_fd_sc_hd__a21oi_1 _21709_ (.A1(_00979_),
    .A2(_00985_),
    .B1(net3827),
    .Y(_01041_));
 sky130_fd_sc_hd__nor2_1 _21710_ (.A(_12330_[0]),
    .B(net3811),
    .Y(_01042_));
 sky130_fd_sc_hd__a21oi_1 _21711_ (.A1(_12328_[0]),
    .A2(net3817),
    .B1(_01042_),
    .Y(_01043_));
 sky130_fd_sc_hd__nand3_1 _21712_ (.A(_00798_),
    .B(_00964_),
    .C(_00965_),
    .Y(_01044_));
 sky130_fd_sc_hd__o211ai_1 _21713_ (.A1(_00798_),
    .A2(_01043_),
    .B1(_01044_),
    .C1(net3822),
    .Y(_01045_));
 sky130_fd_sc_hd__o31ai_1 _21714_ (.A1(net3822),
    .A2(_00984_),
    .A3(_01041_),
    .B1(_01045_),
    .Y(_01046_));
 sky130_fd_sc_hd__o2bb2ai_1 _21715_ (.A1_N(_00900_),
    .A2_N(_01037_),
    .B1(_01039_),
    .B2(_01046_),
    .Y(_01047_));
 sky130_fd_sc_hd__nor3_1 _21716_ (.A(_01002_),
    .B(_01022_),
    .C(_01047_),
    .Y(_00121_));
 sky130_fd_sc_hd__nand2_8 _21717_ (.A(_00777_),
    .B(net3811),
    .Y(_01048_));
 sky130_fd_sc_hd__nand2_4 _21718_ (.A(_12340_[0]),
    .B(net3807),
    .Y(_01049_));
 sky130_fd_sc_hd__nand3_1 _21719_ (.A(net3828),
    .B(_01048_),
    .C(_01049_),
    .Y(_01050_));
 sky130_fd_sc_hd__nand2_1 _21720_ (.A(_00876_),
    .B(_01050_),
    .Y(_01051_));
 sky130_fd_sc_hd__a21oi_1 _21721_ (.A1(_00992_),
    .A2(_01049_),
    .B1(net3828),
    .Y(_01052_));
 sky130_fd_sc_hd__o21ai_0 _21722_ (.A1(_00967_),
    .A2(_01052_),
    .B1(net3824),
    .Y(_01053_));
 sky130_fd_sc_hd__o21ai_0 _21723_ (.A1(net3824),
    .A2(_01051_),
    .B1(_01053_),
    .Y(_01054_));
 sky130_fd_sc_hd__a21oi_1 _21724_ (.A1(_00871_),
    .A2(_01049_),
    .B1(_00798_),
    .Y(_01055_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_254 ();
 sky130_fd_sc_hd__nor2_1 _21726_ (.A(_12335_[0]),
    .B(_00843_),
    .Y(_01057_));
 sky130_fd_sc_hd__o21ai_4 _21727_ (.A1(_12344_[0]),
    .A2(_00830_),
    .B1(_00798_),
    .Y(_01058_));
 sky130_fd_sc_hd__o21ai_0 _21728_ (.A1(_01057_),
    .A2(_01058_),
    .B1(_00943_),
    .Y(_01059_));
 sky130_fd_sc_hd__nor2_1 _21729_ (.A(_01055_),
    .B(_01059_),
    .Y(_01060_));
 sky130_fd_sc_hd__a21oi_1 _21730_ (.A1(_00884_),
    .A2(_00965_),
    .B1(_00798_),
    .Y(_01061_));
 sky130_fd_sc_hd__o21ai_0 _21731_ (.A1(_01012_),
    .A2(_01058_),
    .B1(_00969_),
    .Y(_01062_));
 sky130_fd_sc_hd__o21ai_0 _21732_ (.A1(_01061_),
    .A2(_01062_),
    .B1(_01038_),
    .Y(_01063_));
 sky130_fd_sc_hd__nor2_1 _21733_ (.A(_01060_),
    .B(_01063_),
    .Y(_01064_));
 sky130_fd_sc_hd__o21ai_0 _21734_ (.A1(net3821),
    .A2(_01054_),
    .B1(_01064_),
    .Y(_01065_));
 sky130_fd_sc_hd__a32oi_1 _21735_ (.A1(net3827),
    .A2(_00979_),
    .A3(_00992_),
    .B1(_00918_),
    .B2(_12335_[0]),
    .Y(_01066_));
 sky130_fd_sc_hd__nor3_1 _21736_ (.A(_12330_[0]),
    .B(_12335_[0]),
    .C(_00843_),
    .Y(_01067_));
 sky130_fd_sc_hd__a22oi_1 _21737_ (.A1(_12338_[0]),
    .A2(_00880_),
    .B1(net3578),
    .B2(net3827),
    .Y(_01068_));
 sky130_fd_sc_hd__o21ai_0 _21738_ (.A1(_00917_),
    .A2(_00918_),
    .B1(_12342_[0]),
    .Y(_01069_));
 sky130_fd_sc_hd__nand3_1 _21739_ (.A(net3822),
    .B(_01068_),
    .C(_01069_),
    .Y(_01070_));
 sky130_fd_sc_hd__o211ai_1 _21740_ (.A1(net3821),
    .A2(_01066_),
    .B1(_01070_),
    .C1(net3824),
    .Y(_01071_));
 sky130_fd_sc_hd__a21oi_1 _21741_ (.A1(_12333_[0]),
    .A2(_00798_),
    .B1(net3807),
    .Y(_01072_));
 sky130_fd_sc_hd__a221oi_1 _21742_ (.A1(_12360_[0]),
    .A2(net3807),
    .B1(_00845_),
    .B2(_01072_),
    .C1(net3805),
    .Y(_01073_));
 sky130_fd_sc_hd__nand2_1 _21743_ (.A(_12349_[0]),
    .B(net3811),
    .Y(_01074_));
 sky130_fd_sc_hd__nand2_4 _21744_ (.A(_12333_[0]),
    .B(_00880_),
    .Y(_01075_));
 sky130_fd_sc_hd__a21oi_1 _21745_ (.A1(_01074_),
    .A2(_01075_),
    .B1(net3821),
    .Y(_01076_));
 sky130_fd_sc_hd__o21ai_0 _21746_ (.A1(_01073_),
    .A2(_01076_),
    .B1(net3804),
    .Y(_01077_));
 sky130_fd_sc_hd__nand3_1 _21747_ (.A(_00900_),
    .B(_01071_),
    .C(_01077_),
    .Y(_01078_));
 sky130_fd_sc_hd__nand3_1 _21748_ (.A(_00798_),
    .B(_00979_),
    .C(_00992_),
    .Y(_01079_));
 sky130_fd_sc_hd__o21ai_0 _21749_ (.A1(_00929_),
    .A2(_01029_),
    .B1(net3827),
    .Y(_01080_));
 sky130_fd_sc_hd__a31oi_1 _21750_ (.A1(_00943_),
    .A2(_01079_),
    .A3(_01080_),
    .B1(_00812_),
    .Y(_01081_));
 sky130_fd_sc_hd__nor2_1 _21751_ (.A(_12329_[0]),
    .B(net3827),
    .Y(_01082_));
 sky130_fd_sc_hd__nor3b_1 _21752_ (.A(_01082_),
    .B(net3807),
    .C_N(_00877_),
    .Y(_01083_));
 sky130_fd_sc_hd__a21oi_1 _21753_ (.A1(_12351_[0]),
    .A2(net3807),
    .B1(_01083_),
    .Y(_01084_));
 sky130_fd_sc_hd__nor2_1 _21754_ (.A(_12354_[0]),
    .B(net3818),
    .Y(_01085_));
 sky130_fd_sc_hd__a31oi_1 _21755_ (.A1(net3818),
    .A2(_00845_),
    .A3(_00912_),
    .B1(_01085_),
    .Y(_01086_));
 sky130_fd_sc_hd__nand3_1 _21756_ (.A(_00777_),
    .B(net3827),
    .C(_00871_),
    .Y(_01087_));
 sky130_fd_sc_hd__nand3_1 _21757_ (.A(net3831),
    .B(net3815),
    .C(_00911_),
    .Y(_01088_));
 sky130_fd_sc_hd__nand2_1 _21758_ (.A(net3831),
    .B(_00798_),
    .Y(_01089_));
 sky130_fd_sc_hd__a21o_1 _21759_ (.A1(_00942_),
    .A2(_01089_),
    .B1(_00853_),
    .X(_01090_));
 sky130_fd_sc_hd__a31oi_1 _21760_ (.A1(_01087_),
    .A2(_01088_),
    .A3(_01090_),
    .B1(_00981_),
    .Y(_01091_));
 sky130_fd_sc_hd__a221oi_1 _21761_ (.A1(_00936_),
    .A2(_01084_),
    .B1(_01086_),
    .B2(_00948_),
    .C1(_01091_),
    .Y(_01092_));
 sky130_fd_sc_hd__nand2_1 _21762_ (.A(_01081_),
    .B(_01092_),
    .Y(_01093_));
 sky130_fd_sc_hd__o21ai_1 _21763_ (.A1(_12344_[0]),
    .A2(net3817),
    .B1(net3579),
    .Y(_01094_));
 sky130_fd_sc_hd__or3_1 _21764_ (.A(_00798_),
    .B(_00864_),
    .C(_01012_),
    .X(_01095_));
 sky130_fd_sc_hd__o21ai_0 _21765_ (.A1(net3827),
    .A2(_01094_),
    .B1(_01095_),
    .Y(_01096_));
 sky130_fd_sc_hd__nand2_2 _21766_ (.A(_00876_),
    .B(_00877_),
    .Y(_01097_));
 sky130_fd_sc_hd__nand2_4 _21767_ (.A(net3817),
    .B(_01097_),
    .Y(_01098_));
 sky130_fd_sc_hd__a22o_1 _21768_ (.A1(net3821),
    .A2(_01096_),
    .B1(_01098_),
    .B2(_00848_),
    .X(_01099_));
 sky130_fd_sc_hd__o221ai_1 _21769_ (.A1(_12344_[0]),
    .A2(_00832_),
    .B1(_00995_),
    .B2(net3827),
    .C1(_01075_),
    .Y(_01100_));
 sky130_fd_sc_hd__nand2_8 _21770_ (.A(_12329_[0]),
    .B(_00843_),
    .Y(_01101_));
 sky130_fd_sc_hd__a21oi_1 _21771_ (.A1(_00871_),
    .A2(_01101_),
    .B1(_00798_),
    .Y(_01102_));
 sky130_fd_sc_hd__a311oi_1 _21772_ (.A1(_00798_),
    .A2(_00895_),
    .A3(_00942_),
    .B1(_00981_),
    .C1(_01102_),
    .Y(_01103_));
 sky130_fd_sc_hd__a211oi_1 _21773_ (.A1(_00936_),
    .A2(_01100_),
    .B1(_01103_),
    .C1(_00940_),
    .Y(_01104_));
 sky130_fd_sc_hd__o21ai_0 _21774_ (.A1(net3824),
    .A2(_01099_),
    .B1(_01104_),
    .Y(_01105_));
 sky130_fd_sc_hd__nand4_1 _21775_ (.A(_01065_),
    .B(_01078_),
    .C(_01093_),
    .D(_01105_),
    .Y(_00122_));
 sky130_fd_sc_hd__nor2_1 _21776_ (.A(_12329_[0]),
    .B(_00798_),
    .Y(_01106_));
 sky130_fd_sc_hd__nand2_8 _21777_ (.A(_00806_),
    .B(_00822_),
    .Y(_01107_));
 sky130_fd_sc_hd__a221oi_1 _21778_ (.A1(_00777_),
    .A2(_00862_),
    .B1(_01106_),
    .B2(_00843_),
    .C1(_01107_),
    .Y(_01108_));
 sky130_fd_sc_hd__nor2_1 _21779_ (.A(_12338_[0]),
    .B(net3811),
    .Y(_01109_));
 sky130_fd_sc_hd__o21ai_0 _21780_ (.A1(_00962_),
    .A2(_01109_),
    .B1(_00798_),
    .Y(_01110_));
 sky130_fd_sc_hd__nand2_1 _21781_ (.A(_01108_),
    .B(_01110_),
    .Y(_01111_));
 sky130_fd_sc_hd__nor3_1 _21782_ (.A(_00798_),
    .B(_00932_),
    .C(_01109_),
    .Y(_01112_));
 sky130_fd_sc_hd__a31oi_1 _21783_ (.A1(_00798_),
    .A2(_00992_),
    .A3(_00965_),
    .B1(_01112_),
    .Y(_01113_));
 sky130_fd_sc_hd__or3_1 _21784_ (.A(_00806_),
    .B(net3805),
    .C(_01113_),
    .X(_01114_));
 sky130_fd_sc_hd__nor2_2 _21785_ (.A(_00806_),
    .B(_00822_),
    .Y(_01115_));
 sky130_fd_sc_hd__o21ai_0 _21786_ (.A1(_12329_[0]),
    .A2(net3812),
    .B1(_00945_),
    .Y(_01116_));
 sky130_fd_sc_hd__nand3_1 _21787_ (.A(_00798_),
    .B(_00942_),
    .C(_01007_),
    .Y(_01117_));
 sky130_fd_sc_hd__o21ai_0 _21788_ (.A1(_00798_),
    .A2(_01116_),
    .B1(_01117_),
    .Y(_01118_));
 sky130_fd_sc_hd__nor2_4 _21789_ (.A(_00938_),
    .B(_00822_),
    .Y(_01119_));
 sky130_fd_sc_hd__nand2_2 _21790_ (.A(_00798_),
    .B(_01101_),
    .Y(_01120_));
 sky130_fd_sc_hd__o32ai_1 _21791_ (.A1(_00798_),
    .A2(_00929_),
    .A3(_00934_),
    .B1(_01030_),
    .B2(_01120_),
    .Y(_01121_));
 sky130_fd_sc_hd__a22oi_1 _21792_ (.A1(_01115_),
    .A2(_01118_),
    .B1(_01119_),
    .B2(_01121_),
    .Y(_01122_));
 sky130_fd_sc_hd__nand2_2 _21793_ (.A(_00811_),
    .B(net3824),
    .Y(_01123_));
 sky130_fd_sc_hd__a31oi_1 _21794_ (.A1(_01111_),
    .A2(_01114_),
    .A3(_01122_),
    .B1(_01123_),
    .Y(_01124_));
 sky130_fd_sc_hd__nor2_2 _21795_ (.A(net3827),
    .B(_00862_),
    .Y(_01125_));
 sky130_fd_sc_hd__a32o_1 _21796_ (.A1(net3827),
    .A2(_00884_),
    .A3(_01101_),
    .B1(_00993_),
    .B2(_01125_),
    .X(_01126_));
 sky130_fd_sc_hd__nor2_2 _21797_ (.A(_00777_),
    .B(net3811),
    .Y(_01127_));
 sky130_fd_sc_hd__o21ai_0 _21798_ (.A1(_00798_),
    .A2(_01127_),
    .B1(_00784_),
    .Y(_01128_));
 sky130_fd_sc_hd__a211oi_1 _21799_ (.A1(_00798_),
    .A2(_01029_),
    .B1(_00874_),
    .C1(net3821),
    .Y(_01129_));
 sky130_fd_sc_hd__a221oi_1 _21800_ (.A1(net3821),
    .A2(_01126_),
    .B1(_01128_),
    .B2(_01129_),
    .C1(net3804),
    .Y(_01130_));
 sky130_fd_sc_hd__a22oi_1 _21801_ (.A1(_12342_[0]),
    .A2(_00917_),
    .B1(_01067_),
    .B2(net3827),
    .Y(_01131_));
 sky130_fd_sc_hd__a2bb2oi_1 _21802_ (.A1_N(_12340_[0]),
    .A2_N(_01015_),
    .B1(_00880_),
    .B2(_12338_[0]),
    .Y(_01132_));
 sky130_fd_sc_hd__a21oi_1 _21803_ (.A1(_01131_),
    .A2(_01132_),
    .B1(net3821),
    .Y(_01133_));
 sky130_fd_sc_hd__a311oi_1 _21804_ (.A1(_00911_),
    .A2(_00857_),
    .A3(_00968_),
    .B1(_01133_),
    .C1(net3824),
    .Y(_01134_));
 sky130_fd_sc_hd__nor3_1 _21805_ (.A(_00973_),
    .B(_01130_),
    .C(_01134_),
    .Y(_01135_));
 sky130_fd_sc_hd__nand2_2 _21806_ (.A(_00811_),
    .B(_00903_),
    .Y(_01136_));
 sky130_fd_sc_hd__a21oi_2 _21807_ (.A1(_00853_),
    .A2(net3807),
    .B1(_00798_),
    .Y(_01137_));
 sky130_fd_sc_hd__a32oi_2 _21808_ (.A1(_00798_),
    .A2(_00945_),
    .A3(_01049_),
    .B1(_01137_),
    .B2(_01048_),
    .Y(_01138_));
 sky130_fd_sc_hd__nand2_2 _21809_ (.A(net3808),
    .B(_00841_),
    .Y(_01139_));
 sky130_fd_sc_hd__nand3_1 _21810_ (.A(net3659),
    .B(net3830),
    .C(net3808),
    .Y(_01140_));
 sky130_fd_sc_hd__o211ai_1 _21811_ (.A1(net3827),
    .A2(net3579),
    .B1(_01139_),
    .C1(_01140_),
    .Y(_01141_));
 sky130_fd_sc_hd__a2bb2oi_1 _21812_ (.A1_N(_01107_),
    .A2_N(_01138_),
    .B1(_01119_),
    .B2(_01141_),
    .Y(_01142_));
 sky130_fd_sc_hd__nand2_2 _21813_ (.A(net3831),
    .B(_00855_),
    .Y(_01143_));
 sky130_fd_sc_hd__nor2_1 _21814_ (.A(net3827),
    .B(_00855_),
    .Y(_01144_));
 sky130_fd_sc_hd__nor2_2 _21815_ (.A(_00798_),
    .B(_00822_),
    .Y(_01145_));
 sky130_fd_sc_hd__nor2_1 _21816_ (.A(_01144_),
    .B(_01145_),
    .Y(_01146_));
 sky130_fd_sc_hd__o221ai_1 _21817_ (.A1(net3827),
    .A2(_01143_),
    .B1(_01146_),
    .B2(_12329_[0]),
    .C1(net3818),
    .Y(_01147_));
 sky130_fd_sc_hd__nor2_1 _21818_ (.A(_00806_),
    .B(_01136_),
    .Y(_01148_));
 sky130_fd_sc_hd__nor2_1 _21819_ (.A(net3658),
    .B(_00822_),
    .Y(_01149_));
 sky130_fd_sc_hd__o22ai_1 _21820_ (.A1(_00841_),
    .A2(_01143_),
    .B1(_01149_),
    .B2(_00950_),
    .Y(_01150_));
 sky130_fd_sc_hd__a22oi_1 _21821_ (.A1(_00822_),
    .A2(_00841_),
    .B1(_01150_),
    .B2(net3808),
    .Y(_01151_));
 sky130_fd_sc_hd__nand3_1 _21822_ (.A(_01147_),
    .B(_01148_),
    .C(_01151_),
    .Y(_01152_));
 sky130_fd_sc_hd__o21ai_2 _21823_ (.A1(_01136_),
    .A2(_01142_),
    .B1(_01152_),
    .Y(_01153_));
 sky130_fd_sc_hd__a21oi_1 _21824_ (.A1(_12330_[0]),
    .A2(net3827),
    .B1(_00908_),
    .Y(_01154_));
 sky130_fd_sc_hd__nand2_1 _21825_ (.A(_00777_),
    .B(_00903_),
    .Y(_01155_));
 sky130_fd_sc_hd__o211ai_1 _21826_ (.A1(_00853_),
    .A2(_00903_),
    .B1(_01155_),
    .C1(net3827),
    .Y(_01156_));
 sky130_fd_sc_hd__a21oi_1 _21827_ (.A1(_00903_),
    .A2(_00840_),
    .B1(net3815),
    .Y(_01157_));
 sky130_fd_sc_hd__a221oi_1 _21828_ (.A1(net3813),
    .A2(_01154_),
    .B1(_01156_),
    .B2(_01157_),
    .C1(_00855_),
    .Y(_01158_));
 sky130_fd_sc_hd__nand2_1 _21829_ (.A(_12340_[0]),
    .B(_00919_),
    .Y(_01159_));
 sky130_fd_sc_hd__nand2_4 _21830_ (.A(net3825),
    .B(net3806),
    .Y(_01160_));
 sky130_fd_sc_hd__a21oi_1 _21831_ (.A1(_01139_),
    .A2(_01159_),
    .B1(_01160_),
    .Y(_01161_));
 sky130_fd_sc_hd__nand2_1 _21832_ (.A(net3808),
    .B(_00905_),
    .Y(_01162_));
 sky130_fd_sc_hd__nand2b_1 _21833_ (.A_N(net3578),
    .B(_01137_),
    .Y(_01163_));
 sky130_fd_sc_hd__a31oi_1 _21834_ (.A1(_01011_),
    .A2(_01162_),
    .A3(_01163_),
    .B1(_00924_),
    .Y(_01164_));
 sky130_fd_sc_hd__nor4_1 _21835_ (.A(_00940_),
    .B(_01158_),
    .C(_01161_),
    .D(_01164_),
    .Y(_01165_));
 sky130_fd_sc_hd__nor4_1 _21836_ (.A(_01124_),
    .B(_01135_),
    .C(_01153_),
    .D(_01165_),
    .Y(_00123_));
 sky130_fd_sc_hd__nand4_1 _21837_ (.A(_00798_),
    .B(net3803),
    .C(_00884_),
    .D(_01101_),
    .Y(_01166_));
 sky130_fd_sc_hd__nand3_1 _21838_ (.A(net3827),
    .B(net3803),
    .C(_01094_),
    .Y(_01167_));
 sky130_fd_sc_hd__nand3_1 _21839_ (.A(_00798_),
    .B(_00979_),
    .C(_01048_),
    .Y(_01168_));
 sky130_fd_sc_hd__a31oi_1 _21840_ (.A1(net3826),
    .A2(_00911_),
    .A3(_01168_),
    .B1(_01160_),
    .Y(_01169_));
 sky130_fd_sc_hd__nand2_1 _21841_ (.A(net3827),
    .B(net3823),
    .Y(_01170_));
 sky130_fd_sc_hd__a21oi_1 _21842_ (.A1(_00863_),
    .A2(_01170_),
    .B1(_00777_),
    .Y(_01171_));
 sky130_fd_sc_hd__o21ai_0 _21843_ (.A1(net3827),
    .A2(_00822_),
    .B1(net3830),
    .Y(_01172_));
 sky130_fd_sc_hd__a21oi_1 _21844_ (.A1(net3659),
    .A2(_01172_),
    .B1(_00841_),
    .Y(_01173_));
 sky130_fd_sc_hd__a221oi_1 _21845_ (.A1(_12328_[0]),
    .A2(_01144_),
    .B1(_01145_),
    .B2(net3659),
    .C1(net3808),
    .Y(_01174_));
 sky130_fd_sc_hd__a21oi_2 _21846_ (.A1(net3808),
    .A2(_01173_),
    .B1(_01174_),
    .Y(_01175_));
 sky130_fd_sc_hd__nor4_1 _21847_ (.A(net3803),
    .B(_00816_),
    .C(_01171_),
    .D(_01175_),
    .Y(_01176_));
 sky130_fd_sc_hd__a31oi_1 _21848_ (.A1(_01166_),
    .A2(_01167_),
    .A3(_01169_),
    .B1(_01176_),
    .Y(_01177_));
 sky130_fd_sc_hd__nor2_1 _21849_ (.A(_12328_[0]),
    .B(_00798_),
    .Y(_01178_));
 sky130_fd_sc_hd__o21ai_0 _21850_ (.A1(_01178_),
    .A2(_00951_),
    .B1(net3817),
    .Y(_01179_));
 sky130_fd_sc_hd__nor3b_1 _21851_ (.A(_00798_),
    .B(_00864_),
    .C_N(net3579),
    .Y(_01180_));
 sky130_fd_sc_hd__a21oi_1 _21852_ (.A1(_00993_),
    .A2(_01048_),
    .B1(net3827),
    .Y(_01181_));
 sky130_fd_sc_hd__nor3_1 _21853_ (.A(net3806),
    .B(_01180_),
    .C(_01181_),
    .Y(_01182_));
 sky130_fd_sc_hd__a21oi_1 _21854_ (.A1(_00878_),
    .A2(_01179_),
    .B1(_01182_),
    .Y(_01183_));
 sky130_fd_sc_hd__nand3_1 _21855_ (.A(net3803),
    .B(net3804),
    .C(_01183_),
    .Y(_01184_));
 sky130_fd_sc_hd__o21ai_0 _21856_ (.A1(_12329_[0]),
    .A2(net3826),
    .B1(net3817),
    .Y(_01185_));
 sky130_fd_sc_hd__o211ai_1 _21857_ (.A1(net3826),
    .A2(_01033_),
    .B1(_01185_),
    .C1(_00798_),
    .Y(_01186_));
 sky130_fd_sc_hd__nand2_1 _21858_ (.A(net3827),
    .B(net3803),
    .Y(_01187_));
 sky130_fd_sc_hd__nand2_1 _21859_ (.A(_00798_),
    .B(net3826),
    .Y(_01188_));
 sky130_fd_sc_hd__a21oi_1 _21860_ (.A1(_01187_),
    .A2(_01188_),
    .B1(_12340_[0]),
    .Y(_01189_));
 sky130_fd_sc_hd__a21oi_1 _21861_ (.A1(net3826),
    .A2(_01042_),
    .B1(_01189_),
    .Y(_01190_));
 sky130_fd_sc_hd__a31oi_1 _21862_ (.A1(_00969_),
    .A2(_01186_),
    .A3(_01190_),
    .B1(_00899_),
    .Y(_01191_));
 sky130_fd_sc_hd__nand2_1 _21863_ (.A(net3827),
    .B(_00995_),
    .Y(_01192_));
 sky130_fd_sc_hd__o22ai_1 _21864_ (.A1(_00862_),
    .A2(_01120_),
    .B1(_01192_),
    .B2(_00864_),
    .Y(_01193_));
 sky130_fd_sc_hd__a21oi_1 _21865_ (.A1(net3823),
    .A2(_00996_),
    .B1(net3803),
    .Y(_01194_));
 sky130_fd_sc_hd__o21ai_2 _21866_ (.A1(net3823),
    .A2(_01193_),
    .B1(_01194_),
    .Y(_01195_));
 sky130_fd_sc_hd__nand3_1 _21867_ (.A(_12329_[0]),
    .B(_00798_),
    .C(net3818),
    .Y(_01196_));
 sky130_fd_sc_hd__nand2_1 _21868_ (.A(_00899_),
    .B(net3824),
    .Y(_01197_));
 sky130_fd_sc_hd__a31oi_1 _21869_ (.A1(_00998_),
    .A2(_01115_),
    .A3(_01196_),
    .B1(_01197_),
    .Y(_01198_));
 sky130_fd_sc_hd__a21oi_1 _21870_ (.A1(_00960_),
    .A2(_01048_),
    .B1(_00798_),
    .Y(_01199_));
 sky130_fd_sc_hd__o211ai_1 _21871_ (.A1(_00885_),
    .A2(_01199_),
    .B1(_00938_),
    .C1(net3821),
    .Y(_01200_));
 sky130_fd_sc_hd__nand2_2 _21872_ (.A(net3827),
    .B(net3808),
    .Y(_01201_));
 sky130_fd_sc_hd__o21ai_0 _21873_ (.A1(net3658),
    .A2(_01201_),
    .B1(_01058_),
    .Y(_01202_));
 sky130_fd_sc_hd__a21oi_1 _21874_ (.A1(_00979_),
    .A2(_00983_),
    .B1(_00798_),
    .Y(_01203_));
 sky130_fd_sc_hd__nor3_2 _21875_ (.A(_00986_),
    .B(_01107_),
    .C(_01203_),
    .Y(_01204_));
 sky130_fd_sc_hd__nand2_1 _21876_ (.A(_00899_),
    .B(_00903_),
    .Y(_01205_));
 sky130_fd_sc_hd__a211oi_1 _21877_ (.A1(_01119_),
    .A2(_01202_),
    .B1(_01204_),
    .C1(_01205_),
    .Y(_01206_));
 sky130_fd_sc_hd__nand2_2 _21878_ (.A(_00822_),
    .B(net3818),
    .Y(_01207_));
 sky130_fd_sc_hd__nand3_1 _21879_ (.A(_00855_),
    .B(net3809),
    .C(_00836_),
    .Y(_01208_));
 sky130_fd_sc_hd__a31o_1 _21880_ (.A1(net3830),
    .A2(_00884_),
    .A3(_01144_),
    .B1(_00806_),
    .X(_01209_));
 sky130_fd_sc_hd__a41oi_1 _21881_ (.A1(net3659),
    .A2(net3830),
    .A3(_01207_),
    .A4(_01208_),
    .B1(_01209_),
    .Y(_01210_));
 sky130_fd_sc_hd__o22ai_1 _21882_ (.A1(net3659),
    .A2(_00892_),
    .B1(_00911_),
    .B2(net3808),
    .Y(_01211_));
 sky130_fd_sc_hd__a21oi_1 _21883_ (.A1(_00871_),
    .A2(_01089_),
    .B1(_12340_[0]),
    .Y(_01212_));
 sky130_fd_sc_hd__o221ai_1 _21884_ (.A1(net3818),
    .A2(_00836_),
    .B1(_00871_),
    .B2(net3827),
    .C1(_00855_),
    .Y(_01213_));
 sky130_fd_sc_hd__o31ai_1 _21885_ (.A1(_00855_),
    .A2(_01211_),
    .A3(_01212_),
    .B1(_01213_),
    .Y(_01214_));
 sky130_fd_sc_hd__nand2_1 _21886_ (.A(_01210_),
    .B(_01214_),
    .Y(_01215_));
 sky130_fd_sc_hd__a32o_4 _21887_ (.A1(_01195_),
    .A2(_01198_),
    .A3(_01200_),
    .B1(_01206_),
    .B2(_01215_),
    .X(_01216_));
 sky130_fd_sc_hd__a31oi_1 _21888_ (.A1(_01177_),
    .A2(_01184_),
    .A3(_01191_),
    .B1(_01216_),
    .Y(_00124_));
 sky130_fd_sc_hd__o21ai_0 _21889_ (.A1(net3830),
    .A2(_00917_),
    .B1(_01140_),
    .Y(_01217_));
 sky130_fd_sc_hd__nand2_2 _21890_ (.A(_12335_[0]),
    .B(_00880_),
    .Y(_01218_));
 sky130_fd_sc_hd__o21ai_0 _21891_ (.A1(_12344_[0]),
    .A2(net3827),
    .B1(_00830_),
    .Y(_01219_));
 sky130_fd_sc_hd__a21oi_1 _21892_ (.A1(_01075_),
    .A2(_01131_),
    .B1(net3821),
    .Y(_01220_));
 sky130_fd_sc_hd__a311oi_1 _21893_ (.A1(_00822_),
    .A2(_01218_),
    .A3(_01219_),
    .B1(_01220_),
    .C1(_00806_),
    .Y(_01221_));
 sky130_fd_sc_hd__o22ai_1 _21894_ (.A1(_12340_[0]),
    .A2(_00892_),
    .B1(net3579),
    .B2(net3827),
    .Y(_01222_));
 sky130_fd_sc_hd__a311oi_1 _21895_ (.A1(net3827),
    .A2(_00964_),
    .A3(_00942_),
    .B1(_01107_),
    .C1(_01222_),
    .Y(_01223_));
 sky130_fd_sc_hd__a2111oi_0 _21896_ (.A1(_01119_),
    .A2(_01217_),
    .B1(_01221_),
    .C1(_01197_),
    .D1(_01223_),
    .Y(_01224_));
 sky130_fd_sc_hd__nand2b_1 _21897_ (.A_N(_12328_[0]),
    .B(net3810),
    .Y(_01225_));
 sky130_fd_sc_hd__a21oi_1 _21898_ (.A1(_01225_),
    .A2(_00993_),
    .B1(net3827),
    .Y(_01226_));
 sky130_fd_sc_hd__a21oi_2 _21899_ (.A1(_00872_),
    .A2(_00964_),
    .B1(net3828),
    .Y(_01227_));
 sky130_fd_sc_hd__a211o_1 _21900_ (.A1(net3831),
    .A2(_00917_),
    .B1(_01227_),
    .C1(net3805),
    .X(_01228_));
 sky130_fd_sc_hd__o311a_1 _21901_ (.A1(net3821),
    .A2(_01014_),
    .A3(_01226_),
    .B1(_01228_),
    .C1(_00938_),
    .X(_01229_));
 sky130_fd_sc_hd__nor2_1 _21902_ (.A(net3827),
    .B(_00871_),
    .Y(_01230_));
 sky130_fd_sc_hd__nand2_1 _21903_ (.A(_00806_),
    .B(net3805),
    .Y(_01231_));
 sky130_fd_sc_hd__a311oi_1 _21904_ (.A1(net3827),
    .A2(_00884_),
    .A3(_01101_),
    .B1(_01230_),
    .C1(_01231_),
    .Y(_01232_));
 sky130_fd_sc_hd__a221oi_1 _21905_ (.A1(_12333_[0]),
    .A2(_00830_),
    .B1(_01033_),
    .B2(net3827),
    .C1(_01107_),
    .Y(_01233_));
 sky130_fd_sc_hd__nor4_1 _21906_ (.A(_01136_),
    .B(_01229_),
    .C(_01232_),
    .D(_01233_),
    .Y(_01234_));
 sky130_fd_sc_hd__a21oi_1 _21907_ (.A1(_00968_),
    .A2(_01016_),
    .B1(_00843_),
    .Y(_01235_));
 sky130_fd_sc_hd__nor2_1 _21908_ (.A(_01231_),
    .B(_01235_),
    .Y(_01236_));
 sky130_fd_sc_hd__nand2_1 _21909_ (.A(_00952_),
    .B(_01236_),
    .Y(_01237_));
 sky130_fd_sc_hd__nand2_2 _21910_ (.A(_12340_[0]),
    .B(_00798_),
    .Y(_01238_));
 sky130_fd_sc_hd__o2111ai_2 _21911_ (.A1(net3818),
    .A2(_01238_),
    .B1(_00896_),
    .C1(_00806_),
    .D1(_01007_),
    .Y(_01239_));
 sky130_fd_sc_hd__nor2_1 _21912_ (.A(net3823),
    .B(_00975_),
    .Y(_01240_));
 sky130_fd_sc_hd__a21oi_1 _21913_ (.A1(net3658),
    .A2(_00857_),
    .B1(_01240_),
    .Y(_01241_));
 sky130_fd_sc_hd__o22ai_1 _21914_ (.A1(_12338_[0]),
    .A2(_01207_),
    .B1(_01143_),
    .B2(net3814),
    .Y(_01242_));
 sky130_fd_sc_hd__nor3_1 _21915_ (.A(_12342_[0]),
    .B(_00798_),
    .C(_01207_),
    .Y(_01243_));
 sky130_fd_sc_hd__a2111oi_0 _21916_ (.A1(_00798_),
    .A2(_01242_),
    .B1(_01243_),
    .C1(_00806_),
    .D1(_00956_),
    .Y(_01244_));
 sky130_fd_sc_hd__o21ai_1 _21917_ (.A1(net3831),
    .A2(_01241_),
    .B1(_01244_),
    .Y(_01245_));
 sky130_fd_sc_hd__a31oi_1 _21918_ (.A1(_01237_),
    .A2(_01239_),
    .A3(_01245_),
    .B1(_01123_),
    .Y(_01246_));
 sky130_fd_sc_hd__a21oi_1 _21919_ (.A1(_12338_[0]),
    .A2(_00830_),
    .B1(_01058_),
    .Y(_01247_));
 sky130_fd_sc_hd__a31oi_1 _21920_ (.A1(net3827),
    .A2(_00992_),
    .A3(_01101_),
    .B1(_01247_),
    .Y(_01248_));
 sky130_fd_sc_hd__nand2_1 _21921_ (.A(_12342_[0]),
    .B(_00917_),
    .Y(_01249_));
 sky130_fd_sc_hd__nand2_2 _21922_ (.A(_12338_[0]),
    .B(net3814),
    .Y(_01250_));
 sky130_fd_sc_hd__a31oi_1 _21923_ (.A1(_00855_),
    .A2(_01249_),
    .A3(_01250_),
    .B1(_00806_),
    .Y(_01251_));
 sky130_fd_sc_hd__o21ai_0 _21924_ (.A1(net3805),
    .A2(_01248_),
    .B1(_01251_),
    .Y(_01252_));
 sky130_fd_sc_hd__nor2_1 _21925_ (.A(_12342_[0]),
    .B(_01201_),
    .Y(_01253_));
 sky130_fd_sc_hd__nor3_1 _21926_ (.A(_01107_),
    .B(_01247_),
    .C(_01253_),
    .Y(_01254_));
 sky130_fd_sc_hd__a41oi_1 _21927_ (.A1(_00954_),
    .A2(_01139_),
    .A3(_01119_),
    .A4(_01218_),
    .B1(_01254_),
    .Y(_01255_));
 sky130_fd_sc_hd__a21oi_1 _21928_ (.A1(_01252_),
    .A2(_01255_),
    .B1(_01205_),
    .Y(_01256_));
 sky130_fd_sc_hd__nor4_1 _21929_ (.A(net3568),
    .B(_01234_),
    .C(_01246_),
    .D(_01256_),
    .Y(_00125_));
 sky130_fd_sc_hd__o311a_1 _21930_ (.A1(_12330_[0]),
    .A2(_12335_[0]),
    .A3(net3812),
    .B1(net3579),
    .C1(net3828),
    .X(_01257_));
 sky130_fd_sc_hd__a31oi_1 _21931_ (.A1(_00798_),
    .A2(_00871_),
    .A3(_01101_),
    .B1(_01257_),
    .Y(_01258_));
 sky130_fd_sc_hd__nor2_1 _21932_ (.A(_12349_[0]),
    .B(net3807),
    .Y(_01259_));
 sky130_fd_sc_hd__a211oi_1 _21933_ (.A1(_12333_[0]),
    .A2(_00798_),
    .B1(net3812),
    .C1(_01106_),
    .Y(_01260_));
 sky130_fd_sc_hd__a221oi_1 _21934_ (.A1(_00798_),
    .A2(_00890_),
    .B1(_01048_),
    .B2(_01137_),
    .C1(net3804),
    .Y(_01261_));
 sky130_fd_sc_hd__o32ai_1 _21935_ (.A1(_00981_),
    .A2(_01259_),
    .A3(_01260_),
    .B1(_01261_),
    .B2(net3821),
    .Y(_01262_));
 sky130_fd_sc_hd__o21ai_0 _21936_ (.A1(net3824),
    .A2(_01258_),
    .B1(_01262_),
    .Y(_01263_));
 sky130_fd_sc_hd__a21oi_1 _21937_ (.A1(net3831),
    .A2(net3812),
    .B1(_01109_),
    .Y(_01264_));
 sky130_fd_sc_hd__o221ai_1 _21938_ (.A1(_12333_[0]),
    .A2(_00832_),
    .B1(_01264_),
    .B2(net3827),
    .C1(_00943_),
    .Y(_01265_));
 sky130_fd_sc_hd__nand3_1 _21939_ (.A(_00900_),
    .B(_01263_),
    .C(_01265_),
    .Y(_01266_));
 sky130_fd_sc_hd__a31oi_1 _21940_ (.A1(net3827),
    .A2(_00884_),
    .A3(_01101_),
    .B1(_01125_),
    .Y(_01267_));
 sky130_fd_sc_hd__nor2_4 _21941_ (.A(_12344_[0]),
    .B(_01201_),
    .Y(_01268_));
 sky130_fd_sc_hd__a2111oi_2 _21942_ (.A1(net3831),
    .A2(_00862_),
    .B1(_00905_),
    .C1(_00981_),
    .D1(_01268_),
    .Y(_01269_));
 sky130_fd_sc_hd__a21oi_1 _21943_ (.A1(_12333_[0]),
    .A2(_00880_),
    .B1(net3821),
    .Y(_01270_));
 sky130_fd_sc_hd__o221ai_1 _21944_ (.A1(_00843_),
    .A2(_00911_),
    .B1(_01125_),
    .B2(net3831),
    .C1(_01270_),
    .Y(_01271_));
 sky130_fd_sc_hd__nand2_1 _21945_ (.A(_12358_[0]),
    .B(net3812),
    .Y(_01272_));
 sky130_fd_sc_hd__o211ai_1 _21946_ (.A1(_12333_[0]),
    .A2(net3827),
    .B1(_00843_),
    .C1(_00911_),
    .Y(_01273_));
 sky130_fd_sc_hd__a21oi_1 _21947_ (.A1(_01272_),
    .A2(_01273_),
    .B1(net3805),
    .Y(_01274_));
 sky130_fd_sc_hd__a21oi_1 _21948_ (.A1(net3824),
    .A2(_01271_),
    .B1(_01274_),
    .Y(_01275_));
 sky130_fd_sc_hd__o221ai_1 _21949_ (.A1(_00924_),
    .A2(_01267_),
    .B1(_01269_),
    .B2(_01275_),
    .C1(_01038_),
    .Y(_01276_));
 sky130_fd_sc_hd__o21ai_0 _21950_ (.A1(_12328_[0]),
    .A2(net3812),
    .B1(_00884_),
    .Y(_01277_));
 sky130_fd_sc_hd__a221oi_1 _21951_ (.A1(_12330_[0]),
    .A2(_00918_),
    .B1(_01277_),
    .B2(net3827),
    .C1(_00981_),
    .Y(_01278_));
 sky130_fd_sc_hd__a21o_1 _21952_ (.A1(_01023_),
    .A2(_01238_),
    .B1(net3820),
    .X(_01279_));
 sky130_fd_sc_hd__nand2_2 _21953_ (.A(_00855_),
    .B(_01279_),
    .Y(_01280_));
 sky130_fd_sc_hd__a211oi_1 _21954_ (.A1(_12342_[0]),
    .A2(_00798_),
    .B1(net3808),
    .C1(_00949_),
    .Y(_01281_));
 sky130_fd_sc_hd__o211ai_1 _21955_ (.A1(_12340_[0]),
    .A2(net3807),
    .B1(_00965_),
    .C1(net3827),
    .Y(_01282_));
 sky130_fd_sc_hd__o311ai_0 _21956_ (.A1(net3827),
    .A2(_00930_),
    .A3(net3578),
    .B1(_01282_),
    .C1(_00943_),
    .Y(_01283_));
 sky130_fd_sc_hd__o31ai_1 _21957_ (.A1(_00816_),
    .A2(_01280_),
    .A3(_01281_),
    .B1(_01283_),
    .Y(_01284_));
 sky130_fd_sc_hd__o21ai_0 _21958_ (.A1(_00777_),
    .A2(_00798_),
    .B1(net3820),
    .Y(_01285_));
 sky130_fd_sc_hd__a21oi_1 _21959_ (.A1(_00777_),
    .A2(net3657),
    .B1(_01285_),
    .Y(_01286_));
 sky130_fd_sc_hd__nor3_1 _21960_ (.A(_12347_[0]),
    .B(_12356_[0]),
    .C(net3818),
    .Y(_01287_));
 sky130_fd_sc_hd__o21ai_0 _21961_ (.A1(_01286_),
    .A2(_01287_),
    .B1(_00936_),
    .Y(_01288_));
 sky130_fd_sc_hd__nand3_1 _21962_ (.A(net3826),
    .B(_00811_),
    .C(_01288_),
    .Y(_01289_));
 sky130_fd_sc_hd__nand3_1 _21963_ (.A(net3808),
    .B(_00845_),
    .C(_01238_),
    .Y(_01290_));
 sky130_fd_sc_hd__a21oi_1 _21964_ (.A1(_12348_[0]),
    .A2(net3818),
    .B1(_00903_),
    .Y(_01291_));
 sky130_fd_sc_hd__a221oi_2 _21965_ (.A1(_00903_),
    .A2(_01098_),
    .B1(_01290_),
    .B2(_01291_),
    .C1(_00822_),
    .Y(_01292_));
 sky130_fd_sc_hd__o21a_1 _21966_ (.A1(net3659),
    .A2(_00832_),
    .B1(_01132_),
    .X(_01293_));
 sky130_fd_sc_hd__nor2_1 _21967_ (.A(_01014_),
    .B(_00981_),
    .Y(_01294_));
 sky130_fd_sc_hd__a31oi_1 _21968_ (.A1(_01011_),
    .A2(_01162_),
    .A3(_01294_),
    .B1(_00940_),
    .Y(_01295_));
 sky130_fd_sc_hd__o21ai_0 _21969_ (.A1(_00963_),
    .A2(_01293_),
    .B1(_01295_),
    .Y(_01296_));
 sky130_fd_sc_hd__o32a_1 _21970_ (.A1(_01278_),
    .A2(_01284_),
    .A3(_01289_),
    .B1(_01292_),
    .B2(_01296_),
    .X(_01297_));
 sky130_fd_sc_hd__nand3_1 _21971_ (.A(_01266_),
    .B(_01276_),
    .C(_01297_),
    .Y(_00126_));
 sky130_fd_sc_hd__a21oi_1 _21972_ (.A1(_12340_[0]),
    .A2(net3827),
    .B1(_01082_),
    .Y(_01298_));
 sky130_fd_sc_hd__nor2_1 _21973_ (.A(_12356_[0]),
    .B(net3809),
    .Y(_01299_));
 sky130_fd_sc_hd__a21oi_1 _21974_ (.A1(net3807),
    .A2(_01298_),
    .B1(_01299_),
    .Y(_01300_));
 sky130_fd_sc_hd__nor2_1 _21975_ (.A(_01160_),
    .B(_00976_),
    .Y(_01301_));
 sky130_fd_sc_hd__o21ai_0 _21976_ (.A1(_00834_),
    .A2(_00892_),
    .B1(_01301_),
    .Y(_01302_));
 sky130_fd_sc_hd__a21oi_1 _21977_ (.A1(_00983_),
    .A2(_00894_),
    .B1(_00798_),
    .Y(_01303_));
 sky130_fd_sc_hd__o21ai_0 _21978_ (.A1(_00922_),
    .A2(_01127_),
    .B1(net3827),
    .Y(_01304_));
 sky130_fd_sc_hd__nand3_1 _21979_ (.A(net3804),
    .B(_01044_),
    .C(_01304_),
    .Y(_01305_));
 sky130_fd_sc_hd__o311ai_0 _21980_ (.A1(net3804),
    .A2(_00986_),
    .A3(_01303_),
    .B1(_01305_),
    .C1(net3822),
    .Y(_01306_));
 sky130_fd_sc_hd__o2111ai_1 _21981_ (.A1(_00924_),
    .A2(_01300_),
    .B1(_01302_),
    .C1(_01306_),
    .D1(_00900_),
    .Y(_01307_));
 sky130_fd_sc_hd__a21oi_1 _21982_ (.A1(_00911_),
    .A2(_00950_),
    .B1(net3808),
    .Y(_01308_));
 sky130_fd_sc_hd__nor2_1 _21983_ (.A(_01280_),
    .B(_01308_),
    .Y(_01309_));
 sky130_fd_sc_hd__nor2_1 _21984_ (.A(_12344_[0]),
    .B(_00832_),
    .Y(_01310_));
 sky130_fd_sc_hd__o21ai_0 _21985_ (.A1(_00956_),
    .A2(_01310_),
    .B1(net3823),
    .Y(_01311_));
 sky130_fd_sc_hd__o21ai_0 _21986_ (.A1(_00854_),
    .A2(_00919_),
    .B1(_01311_),
    .Y(_01312_));
 sky130_fd_sc_hd__a31oi_1 _21987_ (.A1(net3820),
    .A2(_00845_),
    .A3(_01238_),
    .B1(_01268_),
    .Y(_01313_));
 sky130_fd_sc_hd__nand2_1 _21988_ (.A(_12328_[0]),
    .B(net3819),
    .Y(_01314_));
 sky130_fd_sc_hd__a21oi_1 _21989_ (.A1(_00894_),
    .A2(_01314_),
    .B1(_01170_),
    .Y(_01315_));
 sky130_fd_sc_hd__nor4_1 _21990_ (.A(net3827),
    .B(net3806),
    .C(_00975_),
    .D(_00976_),
    .Y(_01316_));
 sky130_fd_sc_hd__nor3_1 _21991_ (.A(_01039_),
    .B(_01315_),
    .C(_01316_),
    .Y(_01317_));
 sky130_fd_sc_hd__o21ai_0 _21992_ (.A1(net3823),
    .A2(_01313_),
    .B1(_01317_),
    .Y(_01318_));
 sky130_fd_sc_hd__o31a_1 _21993_ (.A1(_00991_),
    .A2(_01309_),
    .A3(_01312_),
    .B1(_01318_),
    .X(_01319_));
 sky130_fd_sc_hd__o21ai_0 _21994_ (.A1(_00864_),
    .A2(_01286_),
    .B1(_00943_),
    .Y(_01320_));
 sky130_fd_sc_hd__o211ai_1 _21995_ (.A1(_12340_[0]),
    .A2(net3808),
    .B1(_00998_),
    .C1(_00798_),
    .Y(_01321_));
 sky130_fd_sc_hd__o311ai_1 _21996_ (.A1(_00798_),
    .A2(_01029_),
    .A3(net3578),
    .B1(_01321_),
    .C1(_00969_),
    .Y(_01322_));
 sky130_fd_sc_hd__nand3_2 _21997_ (.A(_00798_),
    .B(_00998_),
    .C(_01250_),
    .Y(_01323_));
 sky130_fd_sc_hd__a311oi_1 _21998_ (.A1(_00798_),
    .A2(_00994_),
    .A3(_01048_),
    .B1(_00924_),
    .C1(_01178_),
    .Y(_01324_));
 sky130_fd_sc_hd__a311oi_1 _21999_ (.A1(_00936_),
    .A2(_01006_),
    .A3(_01323_),
    .B1(_01324_),
    .C1(_00812_),
    .Y(_01325_));
 sky130_fd_sc_hd__a22oi_1 _22000_ (.A1(_00777_),
    .A2(_00918_),
    .B1(_01029_),
    .B2(_01145_),
    .Y(_01326_));
 sky130_fd_sc_hd__nand2_1 _22001_ (.A(net3830),
    .B(net3827),
    .Y(_01327_));
 sky130_fd_sc_hd__o32ai_1 _22002_ (.A1(_12342_[0]),
    .A2(net3823),
    .A3(_00892_),
    .B1(_01207_),
    .B2(_01327_),
    .Y(_01328_));
 sky130_fd_sc_hd__nor2_1 _22003_ (.A(_00903_),
    .B(_01328_),
    .Y(_01329_));
 sky130_fd_sc_hd__nor2_1 _22004_ (.A(net3808),
    .B(_01143_),
    .Y(_01330_));
 sky130_fd_sc_hd__o21ai_0 _22005_ (.A1(_00857_),
    .A2(_01330_),
    .B1(net3657),
    .Y(_01331_));
 sky130_fd_sc_hd__nand3_1 _22006_ (.A(_01326_),
    .B(_01329_),
    .C(_01331_),
    .Y(_01332_));
 sky130_fd_sc_hd__a21oi_1 _22007_ (.A1(net3579),
    .A2(_01101_),
    .B1(_00798_),
    .Y(_01333_));
 sky130_fd_sc_hd__a211o_1 _22008_ (.A1(_12342_[0]),
    .A2(_00880_),
    .B1(_01333_),
    .C1(_00855_),
    .X(_01334_));
 sky130_fd_sc_hd__a31oi_1 _22009_ (.A1(_01101_),
    .A2(_00995_),
    .A3(_01145_),
    .B1(_00816_),
    .Y(_01335_));
 sky130_fd_sc_hd__a21oi_1 _22010_ (.A1(_01334_),
    .A2(_01335_),
    .B1(_00940_),
    .Y(_01336_));
 sky130_fd_sc_hd__a32oi_2 _22011_ (.A1(_01320_),
    .A2(_01322_),
    .A3(_01325_),
    .B1(_01332_),
    .B2(_01336_),
    .Y(_01337_));
 sky130_fd_sc_hd__nand3_4 _22012_ (.A(_01307_),
    .B(_01319_),
    .C(_01337_),
    .Y(_00127_));
 sky130_fd_sc_hd__xor3_1 _22013_ (.A(\sa00_sr[7] ),
    .B(\sa00_sr[0] ),
    .C(\sa20_sr[1] ),
    .X(_01338_));
 sky130_fd_sc_hd__xnor3_1 _22014_ (.A(_10489_),
    .B(_10490_),
    .C(_01338_),
    .X(_01339_));
 sky130_fd_sc_hd__nand2_1 _22015_ (.A(net4230),
    .B(\text_in_r[97] ),
    .Y(_01340_));
 sky130_fd_sc_hd__o21a_4 _22016_ (.A1(net4230),
    .A2(_01339_),
    .B1(_01340_),
    .X(_01341_));
 sky130_fd_sc_hd__xor2_4 _22017_ (.A(net4173),
    .B(_01341_),
    .X(_01342_));
 sky130_fd_sc_hd__clkinv_16 _22018_ (.A(_01342_),
    .Y(_01343_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_251 ();
 sky130_fd_sc_hd__xnor3_1 _22022_ (.A(net4189),
    .B(_05874_),
    .C(net4110),
    .X(_01346_));
 sky130_fd_sc_hd__mux2i_1 _22023_ (.A0(\text_in_r[96] ),
    .A1(_01346_),
    .S(net4119),
    .Y(_01347_));
 sky130_fd_sc_hd__xor2_1 _22024_ (.A(net4178),
    .B(_01347_),
    .X(_01348_));
 sky130_fd_sc_hd__clkinv_16 _22025_ (.A(net3799),
    .Y(_01349_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_250 ();
 sky130_fd_sc_hd__xor2_1 _22027_ (.A(\sa30_sr[1] ),
    .B(\sa00_sr[2] ),
    .X(_01350_));
 sky130_fd_sc_hd__xnor2_2 _22028_ (.A(_05893_),
    .B(_01350_),
    .Y(_01351_));
 sky130_fd_sc_hd__mux2i_2 _22029_ (.A0(\text_in_r[98] ),
    .A1(_01351_),
    .S(net4111),
    .Y(_01352_));
 sky130_fd_sc_hd__xnor2_4 _22030_ (.A(\u0.w[0][2] ),
    .B(_01352_),
    .Y(_01353_));
 sky130_fd_sc_hd__clkinv_16 _22031_ (.A(_01353_),
    .Y(_01354_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_240 ();
 sky130_fd_sc_hd__xnor3_1 _22042_ (.A(_05927_),
    .B(_10545_),
    .C(_10546_),
    .X(_01362_));
 sky130_fd_sc_hd__nand2b_2 _22043_ (.A_N(\text_in_r[99] ),
    .B(net398),
    .Y(_01363_));
 sky130_fd_sc_hd__o211a_4 _22044_ (.A1(net398),
    .A2(_01362_),
    .B1(_01363_),
    .C1(net4163),
    .X(_01364_));
 sky130_fd_sc_hd__and2_4 _22045_ (.A(net398),
    .B(\text_in_r[99] ),
    .X(_01365_));
 sky130_fd_sc_hd__a211oi_4 _22046_ (.A1(net4118),
    .A2(_01362_),
    .B1(_01365_),
    .C1(net4163),
    .Y(_01366_));
 sky130_fd_sc_hd__nor2_4 _22047_ (.A(_01366_),
    .B(_01364_),
    .Y(_01367_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_239 ();
 sky130_fd_sc_hd__nand2_8 _22049_ (.A(net3797),
    .B(net3792),
    .Y(_01369_));
 sky130_fd_sc_hd__nand2_4 _22050_ (.A(net3800),
    .B(net3655),
    .Y(_01370_));
 sky130_fd_sc_hd__o211ai_1 _22051_ (.A1(net398),
    .A2(_01362_),
    .B1(_01363_),
    .C1(net4163),
    .Y(_01371_));
 sky130_fd_sc_hd__a211o_4 _22052_ (.A1(net4118),
    .A2(_01362_),
    .B1(_01365_),
    .C1(net4163),
    .X(_01372_));
 sky130_fd_sc_hd__nand2_8 _22053_ (.A(net4071),
    .B(_01372_),
    .Y(_01373_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_238 ();
 sky130_fd_sc_hd__nor2_4 _22055_ (.A(_01343_),
    .B(_01373_),
    .Y(_01375_));
 sky130_fd_sc_hd__o22ai_1 _22056_ (.A1(_12369_[0]),
    .A2(_01369_),
    .B1(_01370_),
    .B2(_01375_),
    .Y(_01376_));
 sky130_fd_sc_hd__xnor3_1 _22057_ (.A(_05949_),
    .B(_10537_),
    .C(_10538_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2i_4 _22058_ (.A0(\text_in_r[100] ),
    .A1(_01377_),
    .S(net4118),
    .Y(_01378_));
 sky130_fd_sc_hd__xnor2_4 _22059_ (.A(net4162),
    .B(_01378_),
    .Y(_01379_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_237 ();
 sky130_fd_sc_hd__xor2_1 _22061_ (.A(\sa00_sr[4] ),
    .B(net4208),
    .X(_01381_));
 sky130_fd_sc_hd__xnor2_2 _22062_ (.A(_10515_),
    .B(_01381_),
    .Y(_01382_));
 sky130_fd_sc_hd__mux2i_4 _22063_ (.A0(\text_in_r[101] ),
    .A1(_01382_),
    .S(net4118),
    .Y(_01383_));
 sky130_fd_sc_hd__xor2_4 _22064_ (.A(net4161),
    .B(_01383_),
    .X(_01384_));
 sky130_fd_sc_hd__nor2_4 _22065_ (.A(net3786),
    .B(_01384_),
    .Y(_01385_));
 sky130_fd_sc_hd__xnor2_4 _22066_ (.A(net4161),
    .B(_01383_),
    .Y(_01386_));
 sky130_fd_sc_hd__nand3_1 _22067_ (.A(_01343_),
    .B(_01349_),
    .C(net3797),
    .Y(_01387_));
 sky130_fd_sc_hd__a31o_4 _22068_ (.A1(net3792),
    .A2(_01370_),
    .A3(_01387_),
    .B1(net3786),
    .X(_01388_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_234 ();
 sky130_fd_sc_hd__nand2_2 _22072_ (.A(_01343_),
    .B(_01354_),
    .Y(_01392_));
 sky130_fd_sc_hd__o211a_1 _22073_ (.A1(_12366_[0]),
    .A2(_01354_),
    .B1(net3789),
    .C1(_01392_),
    .X(_01393_));
 sky130_fd_sc_hd__nor3_1 _22074_ (.A(_01386_),
    .B(_01388_),
    .C(_01393_),
    .Y(_01394_));
 sky130_fd_sc_hd__xor2_4 _22075_ (.A(net4162),
    .B(_01378_),
    .X(_01395_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_231 ();
 sky130_fd_sc_hd__nand2_8 _22079_ (.A(_12378_[0]),
    .B(net3795),
    .Y(_01399_));
 sky130_fd_sc_hd__nand2_8 _22080_ (.A(_01343_),
    .B(net3789),
    .Y(_01400_));
 sky130_fd_sc_hd__nor2_4 _22081_ (.A(_01343_),
    .B(net3792),
    .Y(_01401_));
 sky130_fd_sc_hd__o21ai_0 _22082_ (.A1(_01401_),
    .A2(_01370_),
    .B1(net3785),
    .Y(_01402_));
 sky130_fd_sc_hd__a31oi_1 _22083_ (.A1(net3797),
    .A2(_01399_),
    .A3(_01400_),
    .B1(_01402_),
    .Y(_01403_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_230 ();
 sky130_fd_sc_hd__nor2_2 _22085_ (.A(net3802),
    .B(net393),
    .Y(_01405_));
 sky130_fd_sc_hd__nor2_1 _22086_ (.A(_12378_[0]),
    .B(_01373_),
    .Y(_01406_));
 sky130_fd_sc_hd__or3_1 _22087_ (.A(net3796),
    .B(_01405_),
    .C(_01406_),
    .X(_01407_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_229 ();
 sky130_fd_sc_hd__nor2_4 _22089_ (.A(_01354_),
    .B(_01373_),
    .Y(_01409_));
 sky130_fd_sc_hd__nand2_1 _22090_ (.A(_12365_[0]),
    .B(_01409_),
    .Y(_01410_));
 sky130_fd_sc_hd__nand2_4 _22091_ (.A(_01349_),
    .B(_01373_),
    .Y(_01411_));
 sky130_fd_sc_hd__a31oi_1 _22092_ (.A1(_01407_),
    .A2(_01410_),
    .A3(_01411_),
    .B1(_01384_),
    .Y(_01412_));
 sky130_fd_sc_hd__xnor2_1 _22093_ (.A(\sa00_sr[5] ),
    .B(\sa20_sr[6] ),
    .Y(_01413_));
 sky130_fd_sc_hd__xnor2_2 _22094_ (.A(_10523_),
    .B(_01413_),
    .Y(_01414_));
 sky130_fd_sc_hd__nor2_2 _22095_ (.A(net398),
    .B(_01414_),
    .Y(_01415_));
 sky130_fd_sc_hd__a21oi_4 _22096_ (.A1(net398),
    .A2(\text_in_r[102] ),
    .B1(_01415_),
    .Y(_01416_));
 sky130_fd_sc_hd__xor2_4 _22097_ (.A(net4160),
    .B(_01416_),
    .X(_01417_));
 sky130_fd_sc_hd__xnor2_1 _22098_ (.A(_05971_),
    .B(_10529_),
    .Y(_01418_));
 sky130_fd_sc_hd__mux2i_4 _22099_ (.A0(\text_in_r[103] ),
    .A1(_01418_),
    .S(net4119),
    .Y(_01419_));
 sky130_fd_sc_hd__xnor2_4 _22100_ (.A(net4159),
    .B(_01419_),
    .Y(_01420_));
 sky130_fd_sc_hd__nor2_4 _22101_ (.A(_01417_),
    .B(_01420_),
    .Y(_01421_));
 sky130_fd_sc_hd__o31ai_1 _22102_ (.A1(net3780),
    .A2(_01403_),
    .A3(_01412_),
    .B1(_01421_),
    .Y(_01422_));
 sky130_fd_sc_hd__a211oi_1 _22103_ (.A1(_01376_),
    .A2(_01385_),
    .B1(_01394_),
    .C1(_01422_),
    .Y(_01423_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_226 ();
 sky130_fd_sc_hd__nor2_4 _22107_ (.A(_01354_),
    .B(net394),
    .Y(_01427_));
 sky130_fd_sc_hd__nand2_1 _22108_ (.A(_12374_[0]),
    .B(net3607),
    .Y(_01428_));
 sky130_fd_sc_hd__nand3_4 _22109_ (.A(net3630),
    .B(net4071),
    .C(_01372_),
    .Y(_01429_));
 sky130_fd_sc_hd__nand3_1 _22110_ (.A(net3786),
    .B(_01428_),
    .C(_01429_),
    .Y(_01430_));
 sky130_fd_sc_hd__nand2_1 _22111_ (.A(_01388_),
    .B(_01430_),
    .Y(_01431_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_225 ();
 sky130_fd_sc_hd__nor2_1 _22113_ (.A(_01349_),
    .B(_01373_),
    .Y(_01433_));
 sky130_fd_sc_hd__nand2_8 _22114_ (.A(net3780),
    .B(net3606),
    .Y(_01434_));
 sky130_fd_sc_hd__o211ai_1 _22115_ (.A1(_12369_[0]),
    .A2(net3792),
    .B1(_01434_),
    .C1(net3655),
    .Y(_01435_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_224 ();
 sky130_fd_sc_hd__nand2_1 _22117_ (.A(_12366_[0]),
    .B(_01373_),
    .Y(_01437_));
 sky130_fd_sc_hd__nand2_8 _22118_ (.A(_12369_[0]),
    .B(net3794),
    .Y(_01438_));
 sky130_fd_sc_hd__nor2_2 _22119_ (.A(net3797),
    .B(net3792),
    .Y(_01439_));
 sky130_fd_sc_hd__a32oi_1 _22120_ (.A1(net3797),
    .A2(_01437_),
    .A3(_01438_),
    .B1(net3651),
    .B2(_12364_[0]),
    .Y(_01440_));
 sky130_fd_sc_hd__nand2_8 _22121_ (.A(net3802),
    .B(net3788),
    .Y(_01441_));
 sky130_fd_sc_hd__nand2_8 _22122_ (.A(_01349_),
    .B(net3792),
    .Y(_01442_));
 sky130_fd_sc_hd__nor2_1 _22123_ (.A(_12372_[0]),
    .B(_01373_),
    .Y(_01443_));
 sky130_fd_sc_hd__nor2_2 _22124_ (.A(_12365_[0]),
    .B(_01367_),
    .Y(_01444_));
 sky130_fd_sc_hd__nor3_1 _22125_ (.A(net3798),
    .B(_01443_),
    .C(_01444_),
    .Y(_01445_));
 sky130_fd_sc_hd__a311oi_2 _22126_ (.A1(net3798),
    .A2(_01441_),
    .A3(_01442_),
    .B1(_01445_),
    .C1(net3786),
    .Y(_01446_));
 sky130_fd_sc_hd__a211oi_1 _22127_ (.A1(net3786),
    .A2(_01440_),
    .B1(_01446_),
    .C1(net3785),
    .Y(_01447_));
 sky130_fd_sc_hd__xnor2_4 _22128_ (.A(net4160),
    .B(_01416_),
    .Y(_01448_));
 sky130_fd_sc_hd__nand2_4 _22129_ (.A(_01448_),
    .B(_01420_),
    .Y(_01449_));
 sky130_fd_sc_hd__a311oi_1 _22130_ (.A1(net3785),
    .A2(_01431_),
    .A3(_01435_),
    .B1(_01447_),
    .C1(_01449_),
    .Y(_01450_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_223 ();
 sky130_fd_sc_hd__xor2_4 _22132_ (.A(\u0.w[0][7] ),
    .B(_01419_),
    .X(_01452_));
 sky130_fd_sc_hd__nor2_2 _22133_ (.A(_01448_),
    .B(_01452_),
    .Y(_01453_));
 sky130_fd_sc_hd__nand2_2 _22134_ (.A(net3783),
    .B(_01453_),
    .Y(_01454_));
 sky130_fd_sc_hd__nor2_2 _22135_ (.A(_12366_[0]),
    .B(_01373_),
    .Y(_01455_));
 sky130_fd_sc_hd__nor3_1 _22136_ (.A(net3802),
    .B(_01349_),
    .C(net3795),
    .Y(_01456_));
 sky130_fd_sc_hd__nor3_1 _22137_ (.A(_01354_),
    .B(_01455_),
    .C(_01456_),
    .Y(_01457_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_222 ();
 sky130_fd_sc_hd__nand2_8 _22139_ (.A(_01354_),
    .B(net3789),
    .Y(_01459_));
 sky130_fd_sc_hd__o21ai_2 _22140_ (.A1(_12372_[0]),
    .A2(_01459_),
    .B1(_01379_),
    .Y(_01460_));
 sky130_fd_sc_hd__nor2_4 _22141_ (.A(_12366_[0]),
    .B(net393),
    .Y(_01461_));
 sky130_fd_sc_hd__a21oi_2 _22142_ (.A1(net3656),
    .A2(_01433_),
    .B1(_01461_),
    .Y(_01462_));
 sky130_fd_sc_hd__nor2_4 _22143_ (.A(net3796),
    .B(_01373_),
    .Y(_01463_));
 sky130_fd_sc_hd__a221o_1 _22144_ (.A1(net3796),
    .A2(_01462_),
    .B1(_01463_),
    .B2(_12374_[0]),
    .C1(net3787),
    .X(_01464_));
 sky130_fd_sc_hd__o21ai_2 _22145_ (.A1(_01457_),
    .A2(_01460_),
    .B1(_01464_),
    .Y(_01465_));
 sky130_fd_sc_hd__nand3_2 _22146_ (.A(_01343_),
    .B(net3800),
    .C(_01353_),
    .Y(_01466_));
 sky130_fd_sc_hd__o21ai_2 _22147_ (.A1(_12369_[0]),
    .A2(net3797),
    .B1(_01466_),
    .Y(_01467_));
 sky130_fd_sc_hd__o21ai_2 _22148_ (.A1(net3792),
    .A2(_01467_),
    .B1(_01395_),
    .Y(_01468_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_221 ();
 sky130_fd_sc_hd__nor2_2 _22150_ (.A(_12364_[0]),
    .B(_01369_),
    .Y(_01470_));
 sky130_fd_sc_hd__a21oi_1 _22151_ (.A1(_01442_),
    .A2(_01437_),
    .B1(net3797),
    .Y(_01471_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_220 ();
 sky130_fd_sc_hd__a221o_1 _22153_ (.A1(_12385_[0]),
    .A2(net3792),
    .B1(_01439_),
    .B2(_12365_[0]),
    .C1(net3780),
    .X(_01473_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_219 ();
 sky130_fd_sc_hd__nor3_2 _22155_ (.A(_01386_),
    .B(_01448_),
    .C(_01452_),
    .Y(_01475_));
 sky130_fd_sc_hd__o311ai_0 _22156_ (.A1(_01468_),
    .A2(_01470_),
    .A3(_01471_),
    .B1(_01473_),
    .C1(_01475_),
    .Y(_01476_));
 sky130_fd_sc_hd__o21ai_0 _22157_ (.A1(_01454_),
    .A2(_01465_),
    .B1(_01476_),
    .Y(_01477_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_218 ();
 sky130_fd_sc_hd__nand2_4 _22159_ (.A(_01354_),
    .B(net3791),
    .Y(_01479_));
 sky130_fd_sc_hd__nand2b_4 _22160_ (.A_N(_01427_),
    .B(_01479_),
    .Y(_01480_));
 sky130_fd_sc_hd__nor2_2 _22161_ (.A(_12365_[0]),
    .B(_01369_),
    .Y(_01481_));
 sky130_fd_sc_hd__a221oi_1 _22162_ (.A1(_12372_[0]),
    .A2(net3651),
    .B1(_01480_),
    .B2(_12364_[0]),
    .C1(_01481_),
    .Y(_01482_));
 sky130_fd_sc_hd__nand2_1 _22163_ (.A(net3785),
    .B(_01482_),
    .Y(_01483_));
 sky130_fd_sc_hd__nor2_1 _22164_ (.A(net3802),
    .B(net3800),
    .Y(_01484_));
 sky130_fd_sc_hd__nor2_2 _22165_ (.A(net3792),
    .B(_01484_),
    .Y(_01485_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_217 ();
 sky130_fd_sc_hd__o21ai_0 _22167_ (.A1(_12364_[0]),
    .A2(_01373_),
    .B1(net3655),
    .Y(_01487_));
 sky130_fd_sc_hd__or3_4 _22168_ (.A(_12372_[0]),
    .B(_01364_),
    .C(_01366_),
    .X(_01488_));
 sky130_fd_sc_hd__nand2_8 _22169_ (.A(net3630),
    .B(net3788),
    .Y(_01489_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_216 ();
 sky130_fd_sc_hd__nand3_1 _22171_ (.A(net3797),
    .B(_01488_),
    .C(_01489_),
    .Y(_01491_));
 sky130_fd_sc_hd__o211ai_1 _22172_ (.A1(_01485_),
    .A2(_01487_),
    .B1(net3781),
    .C1(_01491_),
    .Y(_01492_));
 sky130_fd_sc_hd__nor2_4 _22173_ (.A(net3800),
    .B(_01354_),
    .Y(_01493_));
 sky130_fd_sc_hd__nor2_4 _22174_ (.A(_01343_),
    .B(_01349_),
    .Y(_01494_));
 sky130_fd_sc_hd__o21ai_0 _22175_ (.A1(_01493_),
    .A2(_01494_),
    .B1(net3793),
    .Y(_01495_));
 sky130_fd_sc_hd__or3_1 _22176_ (.A(net3793),
    .B(_01493_),
    .C(_01494_),
    .X(_01496_));
 sky130_fd_sc_hd__nand3_1 _22177_ (.A(net3781),
    .B(_01495_),
    .C(_01496_),
    .Y(_01497_));
 sky130_fd_sc_hd__nand2b_4 _22178_ (.A_N(_12365_[0]),
    .B(_01354_),
    .Y(_01498_));
 sky130_fd_sc_hd__nor2_1 _22179_ (.A(_01343_),
    .B(net3797),
    .Y(_01499_));
 sky130_fd_sc_hd__o221ai_1 _22180_ (.A1(_01401_),
    .A2(_01498_),
    .B1(_01489_),
    .B2(_01499_),
    .C1(_01384_),
    .Y(_01500_));
 sky130_fd_sc_hd__a21oi_1 _22181_ (.A1(_01497_),
    .A2(_01500_),
    .B1(net3780),
    .Y(_01501_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_215 ();
 sky130_fd_sc_hd__nand2_4 _22183_ (.A(_01417_),
    .B(_01452_),
    .Y(_01503_));
 sky130_fd_sc_hd__a311oi_1 _22184_ (.A1(net3780),
    .A2(_01483_),
    .A3(_01492_),
    .B1(_01501_),
    .C1(_01503_),
    .Y(_01504_));
 sky130_fd_sc_hd__or4_1 _22185_ (.A(_01423_),
    .B(_01450_),
    .C(_01477_),
    .D(_01504_),
    .X(_00128_));
 sky130_fd_sc_hd__nor2_4 _22186_ (.A(_01349_),
    .B(_01354_),
    .Y(_01505_));
 sky130_fd_sc_hd__nor2_4 _22187_ (.A(net3800),
    .B(net3796),
    .Y(_01506_));
 sky130_fd_sc_hd__nand2_8 _22188_ (.A(_01343_),
    .B(net394),
    .Y(_01507_));
 sky130_fd_sc_hd__a21oi_1 _22189_ (.A1(_12364_[0]),
    .A2(net3652),
    .B1(_01505_),
    .Y(_01508_));
 sky130_fd_sc_hd__o32a_1 _22190_ (.A1(_01505_),
    .A2(_01506_),
    .A3(_01507_),
    .B1(_01508_),
    .B2(net3791),
    .X(_01509_));
 sky130_fd_sc_hd__nand2_8 _22191_ (.A(net3800),
    .B(net3789),
    .Y(_01510_));
 sky130_fd_sc_hd__a21oi_1 _22192_ (.A1(_01438_),
    .A2(_01510_),
    .B1(net3654),
    .Y(_01511_));
 sky130_fd_sc_hd__o31ai_2 _22193_ (.A1(net3797),
    .A2(_01405_),
    .A3(_01375_),
    .B1(_01384_),
    .Y(_01512_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_214 ();
 sky130_fd_sc_hd__o221ai_1 _22195_ (.A1(net3784),
    .A2(_01509_),
    .B1(_01511_),
    .B2(_01512_),
    .C1(net3786),
    .Y(_01514_));
 sky130_fd_sc_hd__a221oi_1 _22196_ (.A1(_12372_[0]),
    .A2(_01354_),
    .B1(_01493_),
    .B2(_01343_),
    .C1(net3792),
    .Y(_01515_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_213 ();
 sky130_fd_sc_hd__nor3_1 _22198_ (.A(_12388_[0]),
    .B(net3783),
    .C(_01373_),
    .Y(_01517_));
 sky130_fd_sc_hd__o21ai_0 _22199_ (.A1(_01515_),
    .A2(_01517_),
    .B1(_01395_),
    .Y(_01518_));
 sky130_fd_sc_hd__a21oi_1 _22200_ (.A1(_01514_),
    .A2(_01518_),
    .B1(_01448_),
    .Y(_01519_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_212 ();
 sky130_fd_sc_hd__nor3_2 _22202_ (.A(net3802),
    .B(net3801),
    .C(_01373_),
    .Y(_01521_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_211 ();
 sky130_fd_sc_hd__o21ai_2 _22204_ (.A1(_01461_),
    .A2(_01521_),
    .B1(_01354_),
    .Y(_01523_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_210 ();
 sky130_fd_sc_hd__or3_4 _22206_ (.A(_12365_[0]),
    .B(_01364_),
    .C(_01366_),
    .X(_01525_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_209 ();
 sky130_fd_sc_hd__nand2_2 _22208_ (.A(_12378_[0]),
    .B(_01373_),
    .Y(_01527_));
 sky130_fd_sc_hd__a31oi_1 _22209_ (.A1(net3798),
    .A2(_01525_),
    .A3(_01527_),
    .B1(_01386_),
    .Y(_01528_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_208 ();
 sky130_fd_sc_hd__nand2_1 _22211_ (.A(_12364_[0]),
    .B(net3790),
    .Y(_01530_));
 sky130_fd_sc_hd__o21ai_0 _22212_ (.A1(_12366_[0]),
    .A2(net3790),
    .B1(_01530_),
    .Y(_01531_));
 sky130_fd_sc_hd__a21oi_2 _22213_ (.A1(_01510_),
    .A2(_01525_),
    .B1(net3798),
    .Y(_01532_));
 sky130_fd_sc_hd__a211oi_1 _22214_ (.A1(net3798),
    .A2(_01531_),
    .B1(_01532_),
    .C1(net3784),
    .Y(_01533_));
 sky130_fd_sc_hd__a21oi_1 _22215_ (.A1(_01523_),
    .A2(_01528_),
    .B1(_01533_),
    .Y(_01534_));
 sky130_fd_sc_hd__nor3_1 _22216_ (.A(_01395_),
    .B(_01417_),
    .C(_01534_),
    .Y(_01535_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_206 ();
 sky130_fd_sc_hd__nand2b_4 _22219_ (.A_N(_12364_[0]),
    .B(_01373_),
    .Y(_01538_));
 sky130_fd_sc_hd__a21oi_1 _22220_ (.A1(_01538_),
    .A2(_01507_),
    .B1(net3798),
    .Y(_01539_));
 sky130_fd_sc_hd__nand3_4 _22221_ (.A(net3656),
    .B(_01349_),
    .C(_01373_),
    .Y(_01540_));
 sky130_fd_sc_hd__a21oi_1 _22222_ (.A1(_01525_),
    .A2(_01540_),
    .B1(_01354_),
    .Y(_01541_));
 sky130_fd_sc_hd__nor2_2 _22223_ (.A(_01349_),
    .B(_01459_),
    .Y(_01542_));
 sky130_fd_sc_hd__o21ai_1 _22224_ (.A1(_01541_),
    .A2(_01542_),
    .B1(net3784),
    .Y(_01543_));
 sky130_fd_sc_hd__o31ai_1 _22225_ (.A1(net3784),
    .A2(_01511_),
    .A3(_01539_),
    .B1(_01543_),
    .Y(_01544_));
 sky130_fd_sc_hd__nor3_1 _22226_ (.A(net3786),
    .B(_01417_),
    .C(_01544_),
    .Y(_01545_));
 sky130_fd_sc_hd__nand2_4 _22227_ (.A(net3786),
    .B(net3784),
    .Y(_01546_));
 sky130_fd_sc_hd__nand2_2 _22228_ (.A(_12364_[0]),
    .B(_01373_),
    .Y(_01547_));
 sky130_fd_sc_hd__nor2_4 _22229_ (.A(_12369_[0]),
    .B(_01373_),
    .Y(_01548_));
 sky130_fd_sc_hd__nor2_4 _22230_ (.A(_01349_),
    .B(net3790),
    .Y(_01549_));
 sky130_fd_sc_hd__nor3_1 _22231_ (.A(net3798),
    .B(_01548_),
    .C(_01549_),
    .Y(_01550_));
 sky130_fd_sc_hd__a31oi_1 _22232_ (.A1(net3798),
    .A2(_01547_),
    .A3(_01429_),
    .B1(_01550_),
    .Y(_01551_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_205 ();
 sky130_fd_sc_hd__nand2_4 _22234_ (.A(_01379_),
    .B(_01386_),
    .Y(_01552_));
 sky130_fd_sc_hd__a21oi_1 _22235_ (.A1(net3802),
    .A2(_01409_),
    .B1(_01552_),
    .Y(_01553_));
 sky130_fd_sc_hd__nand2_1 _22236_ (.A(_01354_),
    .B(_01399_),
    .Y(_01554_));
 sky130_fd_sc_hd__a31oi_1 _22237_ (.A1(_01553_),
    .A2(_01540_),
    .A3(_01554_),
    .B1(_01449_),
    .Y(_01555_));
 sky130_fd_sc_hd__o21a_1 _22238_ (.A1(_01546_),
    .A2(_01551_),
    .B1(_01555_),
    .X(_01556_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_204 ();
 sky130_fd_sc_hd__nand2_2 _22240_ (.A(_12365_[0]),
    .B(_01354_),
    .Y(_01558_));
 sky130_fd_sc_hd__o22ai_1 _22241_ (.A1(_01343_),
    .A2(_01442_),
    .B1(_01558_),
    .B2(net3792),
    .Y(_01559_));
 sky130_fd_sc_hd__a211oi_1 _22242_ (.A1(net3800),
    .A2(_01480_),
    .B1(_01559_),
    .C1(net3783),
    .Y(_01560_));
 sky130_fd_sc_hd__nand2_4 _22243_ (.A(_12369_[0]),
    .B(net3789),
    .Y(_01561_));
 sky130_fd_sc_hd__a21oi_2 _22244_ (.A1(_01343_),
    .A2(_01349_),
    .B1(net3789),
    .Y(_01562_));
 sky130_fd_sc_hd__nor2_1 _22245_ (.A(net3798),
    .B(_01562_),
    .Y(_01563_));
 sky130_fd_sc_hd__a311oi_1 _22246_ (.A1(net3798),
    .A2(_01525_),
    .A3(_01561_),
    .B1(_01563_),
    .C1(net3784),
    .Y(_01564_));
 sky130_fd_sc_hd__o21ai_0 _22247_ (.A1(_01560_),
    .A2(_01564_),
    .B1(_01395_),
    .Y(_01565_));
 sky130_fd_sc_hd__a21oi_1 _22248_ (.A1(_01411_),
    .A2(_01479_),
    .B1(net3656),
    .Y(_01566_));
 sky130_fd_sc_hd__o21ai_2 _22249_ (.A1(_01506_),
    .A2(_01566_),
    .B1(net3780),
    .Y(_01567_));
 sky130_fd_sc_hd__nand2_2 _22250_ (.A(_01429_),
    .B(_01561_),
    .Y(_01568_));
 sky130_fd_sc_hd__o21ai_0 _22251_ (.A1(_01343_),
    .A2(net3786),
    .B1(_01549_),
    .Y(_01569_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_203 ();
 sky130_fd_sc_hd__a21oi_1 _22253_ (.A1(_01442_),
    .A2(_01569_),
    .B1(net3798),
    .Y(_01571_));
 sky130_fd_sc_hd__a311oi_1 _22254_ (.A1(net3798),
    .A2(net3786),
    .A3(_01568_),
    .B1(_01571_),
    .C1(_01454_),
    .Y(_01572_));
 sky130_fd_sc_hd__nand2_1 _22255_ (.A(_12378_[0]),
    .B(net3798),
    .Y(_01573_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_202 ();
 sky130_fd_sc_hd__a21oi_1 _22257_ (.A1(_01558_),
    .A2(_01573_),
    .B1(net3789),
    .Y(_01575_));
 sky130_fd_sc_hd__a2bb2oi_1 _22258_ (.A1_N(_12369_[0]),
    .A2_N(_01459_),
    .B1(_01480_),
    .B2(_01343_),
    .Y(_01576_));
 sky130_fd_sc_hd__o22ai_1 _22259_ (.A1(_01468_),
    .A2(_01575_),
    .B1(_01576_),
    .B2(net3780),
    .Y(_01577_));
 sky130_fd_sc_hd__a222oi_1 _22260_ (.A1(_01556_),
    .A2(_01565_),
    .B1(_01567_),
    .B2(_01572_),
    .C1(_01577_),
    .C2(_01475_),
    .Y(_01578_));
 sky130_fd_sc_hd__o41a_1 _22261_ (.A1(_01420_),
    .A2(_01519_),
    .A3(_01535_),
    .A4(_01545_),
    .B1(_01578_),
    .X(_00129_));
 sky130_fd_sc_hd__nand2_2 _22262_ (.A(_01448_),
    .B(_01452_),
    .Y(_01579_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_201 ();
 sky130_fd_sc_hd__a21boi_0 _22264_ (.A1(_12374_[0]),
    .A2(_01373_),
    .B1_N(_01507_),
    .Y(_01581_));
 sky130_fd_sc_hd__nand2_2 _22265_ (.A(net3780),
    .B(_01384_),
    .Y(_01582_));
 sky130_fd_sc_hd__nor2_1 _22266_ (.A(_12369_[0]),
    .B(net3797),
    .Y(_01583_));
 sky130_fd_sc_hd__a211oi_1 _22267_ (.A1(net3797),
    .A2(_01581_),
    .B1(_01582_),
    .C1(_01583_),
    .Y(_01584_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_200 ();
 sky130_fd_sc_hd__nand2b_2 _22269_ (.A_N(net3592),
    .B(_01373_),
    .Y(_01586_));
 sky130_fd_sc_hd__nor2_1 _22270_ (.A(_12374_[0]),
    .B(_01373_),
    .Y(_01587_));
 sky130_fd_sc_hd__nor3_1 _22271_ (.A(net3654),
    .B(_01549_),
    .C(_01587_),
    .Y(_01588_));
 sky130_fd_sc_hd__a31oi_1 _22272_ (.A1(net3654),
    .A2(_01507_),
    .A3(_01586_),
    .B1(_01588_),
    .Y(_01589_));
 sky130_fd_sc_hd__nor2_4 _22273_ (.A(_12374_[0]),
    .B(net3795),
    .Y(_01590_));
 sky130_fd_sc_hd__nor3_1 _22274_ (.A(net3655),
    .B(net3606),
    .C(_01590_),
    .Y(_01591_));
 sky130_fd_sc_hd__nor2_4 _22275_ (.A(_12378_[0]),
    .B(net3795),
    .Y(_01592_));
 sky130_fd_sc_hd__nor3_1 _22276_ (.A(net3797),
    .B(_01548_),
    .C(_01592_),
    .Y(_01593_));
 sky130_fd_sc_hd__nor2_1 _22277_ (.A(_01591_),
    .B(_01593_),
    .Y(_01594_));
 sky130_fd_sc_hd__o22ai_1 _22278_ (.A1(_01552_),
    .A2(_01589_),
    .B1(_01594_),
    .B2(_01546_),
    .Y(_01595_));
 sky130_fd_sc_hd__nand3_1 _22279_ (.A(net3797),
    .B(_01510_),
    .C(_01525_),
    .Y(_01596_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_199 ();
 sky130_fd_sc_hd__o211ai_1 _22281_ (.A1(_12374_[0]),
    .A2(net3790),
    .B1(_01429_),
    .C1(net3654),
    .Y(_01598_));
 sky130_fd_sc_hd__nand2_8 _22282_ (.A(_01395_),
    .B(net3782),
    .Y(_01599_));
 sky130_fd_sc_hd__a21oi_1 _22283_ (.A1(_01596_),
    .A2(_01598_),
    .B1(_01599_),
    .Y(_01600_));
 sky130_fd_sc_hd__a21oi_1 _22284_ (.A1(_01429_),
    .A2(_01538_),
    .B1(_01354_),
    .Y(_01601_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_198 ();
 sky130_fd_sc_hd__and3_1 _22286_ (.A(_12369_[0]),
    .B(_01354_),
    .C(net3792),
    .X(_01603_));
 sky130_fd_sc_hd__o21ai_2 _22287_ (.A1(_01601_),
    .A2(_01603_),
    .B1(_01385_),
    .Y(_01604_));
 sky130_fd_sc_hd__nand2_2 _22288_ (.A(_01379_),
    .B(net3788),
    .Y(_01605_));
 sky130_fd_sc_hd__nor2_1 _22289_ (.A(net3780),
    .B(net3788),
    .Y(_01606_));
 sky130_fd_sc_hd__nor3_1 _22290_ (.A(net3796),
    .B(_01379_),
    .C(net3791),
    .Y(_01607_));
 sky130_fd_sc_hd__o221ai_1 _22291_ (.A1(net3800),
    .A2(net3796),
    .B1(_01606_),
    .B2(_01607_),
    .C1(net3656),
    .Y(_01608_));
 sky130_fd_sc_hd__nor2_1 _22292_ (.A(_01379_),
    .B(net3788),
    .Y(_01609_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_197 ();
 sky130_fd_sc_hd__a21oi_1 _22294_ (.A1(_12383_[0]),
    .A2(_01609_),
    .B1(net3781),
    .Y(_01611_));
 sky130_fd_sc_hd__o211ai_1 _22295_ (.A1(_12392_[0]),
    .A2(_01605_),
    .B1(_01608_),
    .C1(_01611_),
    .Y(_01612_));
 sky130_fd_sc_hd__nor2_4 _22296_ (.A(_12366_[0]),
    .B(_12369_[0]),
    .Y(_01613_));
 sky130_fd_sc_hd__o21ai_1 _22297_ (.A1(net3789),
    .A2(_01613_),
    .B1(net3798),
    .Y(_01614_));
 sky130_fd_sc_hd__o21ai_0 _22298_ (.A1(_12372_[0]),
    .A2(net3794),
    .B1(_01354_),
    .Y(_01615_));
 sky130_fd_sc_hd__nor2_4 _22299_ (.A(net3780),
    .B(_01384_),
    .Y(_01616_));
 sky130_fd_sc_hd__o221ai_1 _22300_ (.A1(_01485_),
    .A2(_01614_),
    .B1(_01615_),
    .B2(_01562_),
    .C1(_01616_),
    .Y(_01617_));
 sky130_fd_sc_hd__nand4_1 _22301_ (.A(_01453_),
    .B(_01604_),
    .C(_01612_),
    .D(_01617_),
    .Y(_01618_));
 sky130_fd_sc_hd__o41ai_1 _22302_ (.A1(_01579_),
    .A2(_01584_),
    .A3(_01595_),
    .A4(_01600_),
    .B1(_01618_),
    .Y(_01619_));
 sky130_fd_sc_hd__o21ai_0 _22303_ (.A1(_01405_),
    .A2(_01499_),
    .B1(_12365_[0]),
    .Y(_01620_));
 sky130_fd_sc_hd__nand2_8 _22304_ (.A(_01349_),
    .B(net3796),
    .Y(_01621_));
 sky130_fd_sc_hd__nor2_4 _22305_ (.A(net3802),
    .B(_01354_),
    .Y(_01622_));
 sky130_fd_sc_hd__a22oi_1 _22306_ (.A1(_01375_),
    .A2(_01621_),
    .B1(_01442_),
    .B2(_01622_),
    .Y(_01623_));
 sky130_fd_sc_hd__o211a_1 _22307_ (.A1(_12364_[0]),
    .A2(net3793),
    .B1(_01429_),
    .C1(net3655),
    .X(_01624_));
 sky130_fd_sc_hd__a311oi_1 _22308_ (.A1(net3797),
    .A2(_01400_),
    .A3(_01488_),
    .B1(_01624_),
    .C1(net3781),
    .Y(_01625_));
 sky130_fd_sc_hd__a31oi_1 _22309_ (.A1(net3781),
    .A2(_01620_),
    .A3(_01623_),
    .B1(_01625_),
    .Y(_01626_));
 sky130_fd_sc_hd__nor2_1 _22310_ (.A(net3780),
    .B(_01626_),
    .Y(_01627_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_196 ();
 sky130_fd_sc_hd__nor3_1 _22312_ (.A(_01373_),
    .B(_01494_),
    .C(_01622_),
    .Y(_01629_));
 sky130_fd_sc_hd__nor2_1 _22313_ (.A(_12388_[0]),
    .B(net3792),
    .Y(_01630_));
 sky130_fd_sc_hd__nor2_1 _22314_ (.A(_01629_),
    .B(_01630_),
    .Y(_01631_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_195 ();
 sky130_fd_sc_hd__nand3_1 _22316_ (.A(net3792),
    .B(_01466_),
    .C(_01498_),
    .Y(_01633_));
 sky130_fd_sc_hd__a21oi_1 _22317_ (.A1(_12385_[0]),
    .A2(_01373_),
    .B1(net3785),
    .Y(_01634_));
 sky130_fd_sc_hd__a221oi_1 _22318_ (.A1(net3785),
    .A2(_01631_),
    .B1(_01633_),
    .B2(_01634_),
    .C1(net3786),
    .Y(_01635_));
 sky130_fd_sc_hd__nor3_1 _22319_ (.A(_01449_),
    .B(_01627_),
    .C(_01635_),
    .Y(_01636_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_194 ();
 sky130_fd_sc_hd__nor2_2 _22321_ (.A(_12378_[0]),
    .B(_01369_),
    .Y(_01638_));
 sky130_fd_sc_hd__a21oi_2 _22322_ (.A1(_01442_),
    .A2(_01510_),
    .B1(_01392_),
    .Y(_01639_));
 sky130_fd_sc_hd__a21oi_1 _22323_ (.A1(_01442_),
    .A2(_01489_),
    .B1(_01354_),
    .Y(_01640_));
 sky130_fd_sc_hd__nor3_1 _22324_ (.A(net3796),
    .B(_01405_),
    .C(_01455_),
    .Y(_01641_));
 sky130_fd_sc_hd__o21ai_0 _22325_ (.A1(_01640_),
    .A2(_01641_),
    .B1(net3787),
    .Y(_01642_));
 sky130_fd_sc_hd__o31ai_1 _22326_ (.A1(net3787),
    .A2(_01638_),
    .A3(_01639_),
    .B1(_01642_),
    .Y(_01643_));
 sky130_fd_sc_hd__nand3_4 _22327_ (.A(_01343_),
    .B(net3801),
    .C(net3792),
    .Y(_01644_));
 sky130_fd_sc_hd__a21oi_1 _22328_ (.A1(_01438_),
    .A2(_01489_),
    .B1(net3796),
    .Y(_01645_));
 sky130_fd_sc_hd__a311oi_2 _22329_ (.A1(net3796),
    .A2(_01441_),
    .A3(_01644_),
    .B1(_01645_),
    .C1(net3787),
    .Y(_01646_));
 sky130_fd_sc_hd__a21oi_1 _22330_ (.A1(_01442_),
    .A2(_01527_),
    .B1(net3797),
    .Y(_01647_));
 sky130_fd_sc_hd__a2111oi_0 _22331_ (.A1(_12369_[0]),
    .A2(net3607),
    .B1(_01647_),
    .C1(net3780),
    .D1(_01375_),
    .Y(_01648_));
 sky130_fd_sc_hd__nor3_1 _22332_ (.A(net3781),
    .B(_01646_),
    .C(_01648_),
    .Y(_01649_));
 sky130_fd_sc_hd__a211oi_1 _22333_ (.A1(net3781),
    .A2(_01643_),
    .B1(_01649_),
    .C1(_01503_),
    .Y(_01650_));
 sky130_fd_sc_hd__nor3_1 _22334_ (.A(_01619_),
    .B(_01636_),
    .C(_01650_),
    .Y(_00130_));
 sky130_fd_sc_hd__nand2_1 _22335_ (.A(_12372_[0]),
    .B(_01373_),
    .Y(_01651_));
 sky130_fd_sc_hd__nand3b_1 _22336_ (.A_N(_01587_),
    .B(_01651_),
    .C(net3654),
    .Y(_01652_));
 sky130_fd_sc_hd__nand2_2 _22337_ (.A(net3791),
    .B(_01613_),
    .Y(_01653_));
 sky130_fd_sc_hd__a31oi_1 _22338_ (.A1(net3796),
    .A2(_01540_),
    .A3(_01653_),
    .B1(_01379_),
    .Y(_01654_));
 sky130_fd_sc_hd__a211oi_1 _22339_ (.A1(net3592),
    .A2(net3652),
    .B1(net3604),
    .C1(_01605_),
    .Y(_01655_));
 sky130_fd_sc_hd__a21oi_1 _22340_ (.A1(_01652_),
    .A2(_01654_),
    .B1(_01655_),
    .Y(_01656_));
 sky130_fd_sc_hd__nor2_1 _22341_ (.A(net3782),
    .B(_01656_),
    .Y(_01657_));
 sky130_fd_sc_hd__a21oi_1 _22342_ (.A1(net3797),
    .A2(_01441_),
    .B1(net3801),
    .Y(_01658_));
 sky130_fd_sc_hd__a2111oi_4 _22343_ (.A1(_01343_),
    .A2(net3651),
    .B1(_01470_),
    .C1(_01658_),
    .D1(_01599_),
    .Y(_01659_));
 sky130_fd_sc_hd__nand2_4 _22344_ (.A(_12374_[0]),
    .B(net3790),
    .Y(_01660_));
 sky130_fd_sc_hd__a21oi_1 _22345_ (.A1(_01442_),
    .A2(_01586_),
    .B1(net3797),
    .Y(_01661_));
 sky130_fd_sc_hd__a31oi_1 _22346_ (.A1(net3797),
    .A2(_01489_),
    .A3(_01660_),
    .B1(_01661_),
    .Y(_01662_));
 sky130_fd_sc_hd__o21ai_0 _22347_ (.A1(_01552_),
    .A2(_01662_),
    .B1(_01421_),
    .Y(_01663_));
 sky130_fd_sc_hd__nor2_4 _22348_ (.A(_01417_),
    .B(_01452_),
    .Y(_01664_));
 sky130_fd_sc_hd__a221oi_1 _22349_ (.A1(_12372_[0]),
    .A2(net3651),
    .B1(net3606),
    .B2(net3802),
    .C1(_01640_),
    .Y(_01665_));
 sky130_fd_sc_hd__nand2_2 _22350_ (.A(_01373_),
    .B(_01493_),
    .Y(_01666_));
 sky130_fd_sc_hd__o21ai_0 _22351_ (.A1(_01373_),
    .A2(_01370_),
    .B1(_01666_),
    .Y(_01667_));
 sky130_fd_sc_hd__a2bb2oi_1 _22352_ (.A1_N(_12365_[0]),
    .A2_N(_01459_),
    .B1(_01409_),
    .B2(_12372_[0]),
    .Y(_01668_));
 sky130_fd_sc_hd__nand3_1 _22353_ (.A(_01385_),
    .B(_01664_),
    .C(_01668_),
    .Y(_01669_));
 sky130_fd_sc_hd__a21oi_1 _22354_ (.A1(_01343_),
    .A2(_01667_),
    .B1(_01669_),
    .Y(_01670_));
 sky130_fd_sc_hd__nand2_1 _22355_ (.A(net3802),
    .B(net3795),
    .Y(_01671_));
 sky130_fd_sc_hd__nor3_1 _22356_ (.A(net3796),
    .B(_01406_),
    .C(_01590_),
    .Y(_01672_));
 sky130_fd_sc_hd__a311oi_1 _22357_ (.A1(net3796),
    .A2(_01671_),
    .A3(_01489_),
    .B1(_01672_),
    .C1(net3780),
    .Y(_01673_));
 sky130_fd_sc_hd__nor4_1 _22358_ (.A(net3787),
    .B(_01409_),
    .C(_01506_),
    .D(_01494_),
    .Y(_01674_));
 sky130_fd_sc_hd__nor4_1 _22359_ (.A(net3781),
    .B(_01449_),
    .C(_01673_),
    .D(_01674_),
    .Y(_01675_));
 sky130_fd_sc_hd__a311oi_2 _22360_ (.A1(_01664_),
    .A2(_01616_),
    .A3(_01665_),
    .B1(_01670_),
    .C1(_01675_),
    .Y(_01676_));
 sky130_fd_sc_hd__nor2_2 _22361_ (.A(net3652),
    .B(_01379_),
    .Y(_01677_));
 sky130_fd_sc_hd__nand2_1 _22362_ (.A(_01349_),
    .B(_01677_),
    .Y(_01678_));
 sky130_fd_sc_hd__nor2_1 _22363_ (.A(net3802),
    .B(_01349_),
    .Y(_01679_));
 sky130_fd_sc_hd__nand2_2 _22364_ (.A(_01354_),
    .B(net3786),
    .Y(_01680_));
 sky130_fd_sc_hd__a32oi_1 _22365_ (.A1(net3802),
    .A2(_01379_),
    .A3(_01621_),
    .B1(_01679_),
    .B2(_01680_),
    .Y(_01681_));
 sky130_fd_sc_hd__a211oi_1 _22366_ (.A1(_01678_),
    .A2(_01681_),
    .B1(net3781),
    .C1(net3791),
    .Y(_01682_));
 sky130_fd_sc_hd__nand2b_4 _22367_ (.A_N(net3630),
    .B(net3788),
    .Y(_01683_));
 sky130_fd_sc_hd__nand3_1 _22368_ (.A(net3798),
    .B(_01399_),
    .C(_01683_),
    .Y(_01684_));
 sky130_fd_sc_hd__nand3_1 _22369_ (.A(_01354_),
    .B(_01400_),
    .C(_01438_),
    .Y(_01685_));
 sky130_fd_sc_hd__a21oi_1 _22370_ (.A1(_01684_),
    .A2(_01685_),
    .B1(_01599_),
    .Y(_01686_));
 sky130_fd_sc_hd__and3_1 _22371_ (.A(net3798),
    .B(_01530_),
    .C(_01651_),
    .X(_01687_));
 sky130_fd_sc_hd__a311oi_1 _22372_ (.A1(_01354_),
    .A2(_01429_),
    .A3(_01510_),
    .B1(_01552_),
    .C1(_01687_),
    .Y(_01688_));
 sky130_fd_sc_hd__nor3_1 _22373_ (.A(_01682_),
    .B(_01686_),
    .C(_01688_),
    .Y(_01689_));
 sky130_fd_sc_hd__nand2_1 _22374_ (.A(net3798),
    .B(net3786),
    .Y(_01690_));
 sky130_fd_sc_hd__a22oi_1 _22375_ (.A1(_12366_[0]),
    .A2(_01367_),
    .B1(_01444_),
    .B2(net3782),
    .Y(_01691_));
 sky130_fd_sc_hd__nor2_1 _22376_ (.A(_01427_),
    .B(_01463_),
    .Y(_01692_));
 sky130_fd_sc_hd__a21boi_2 _22377_ (.A1(_12374_[0]),
    .A2(_01692_),
    .B1_N(_01666_),
    .Y(_01693_));
 sky130_fd_sc_hd__o221ai_1 _22378_ (.A1(_01690_),
    .A2(_01691_),
    .B1(_01693_),
    .B2(_01599_),
    .C1(_01452_),
    .Y(_01694_));
 sky130_fd_sc_hd__a21oi_2 _22379_ (.A1(_01399_),
    .A2(_01411_),
    .B1(net3796),
    .Y(_01695_));
 sky130_fd_sc_hd__a311oi_1 _22380_ (.A1(net3796),
    .A2(_01683_),
    .A3(_01653_),
    .B1(_01695_),
    .C1(_01379_),
    .Y(_01696_));
 sky130_fd_sc_hd__o21ai_0 _22381_ (.A1(_12372_[0]),
    .A2(net3791),
    .B1(_01525_),
    .Y(_01697_));
 sky130_fd_sc_hd__a221oi_1 _22382_ (.A1(net3802),
    .A2(_01427_),
    .B1(_01697_),
    .B2(_01354_),
    .C1(net3780),
    .Y(_01698_));
 sky130_fd_sc_hd__nor3_1 _22383_ (.A(_01386_),
    .B(_01696_),
    .C(_01698_),
    .Y(_01699_));
 sky130_fd_sc_hd__nor2_2 _22384_ (.A(net3781),
    .B(_01452_),
    .Y(_01700_));
 sky130_fd_sc_hd__nand2_2 _22385_ (.A(net3652),
    .B(net3780),
    .Y(_01701_));
 sky130_fd_sc_hd__nor2_1 _22386_ (.A(net3796),
    .B(_01395_),
    .Y(_01702_));
 sky130_fd_sc_hd__nor2_1 _22387_ (.A(net3603),
    .B(_01702_),
    .Y(_01703_));
 sky130_fd_sc_hd__o22ai_1 _22388_ (.A1(_01343_),
    .A2(_01701_),
    .B1(_01703_),
    .B2(net3630),
    .Y(_01704_));
 sky130_fd_sc_hd__a31oi_1 _22389_ (.A1(net3791),
    .A2(_01700_),
    .A3(_01704_),
    .B1(_01448_),
    .Y(_01705_));
 sky130_fd_sc_hd__o221ai_1 _22390_ (.A1(_01452_),
    .A2(_01689_),
    .B1(_01694_),
    .B2(_01699_),
    .C1(_01705_),
    .Y(_01706_));
 sky130_fd_sc_hd__o311ai_0 _22391_ (.A1(_01657_),
    .A2(_01659_),
    .A3(_01663_),
    .B1(_01676_),
    .C1(_01706_),
    .Y(_00131_));
 sky130_fd_sc_hd__nor2_1 _22392_ (.A(net3786),
    .B(_01386_),
    .Y(_01707_));
 sky130_fd_sc_hd__o22ai_2 _22393_ (.A1(_12378_[0]),
    .A2(_01459_),
    .B1(_01549_),
    .B2(_01354_),
    .Y(_01708_));
 sky130_fd_sc_hd__nand2_1 _22394_ (.A(_01707_),
    .B(_01708_),
    .Y(_01709_));
 sky130_fd_sc_hd__a21oi_1 _22395_ (.A1(_01438_),
    .A2(_01538_),
    .B1(net3654),
    .Y(_01710_));
 sky130_fd_sc_hd__o22ai_1 _22396_ (.A1(net3784),
    .A2(_01523_),
    .B1(_01710_),
    .B2(_01512_),
    .Y(_01711_));
 sky130_fd_sc_hd__nand2_1 _22397_ (.A(_12369_[0]),
    .B(net3797),
    .Y(_01712_));
 sky130_fd_sc_hd__a21oi_1 _22398_ (.A1(_01498_),
    .A2(_01712_),
    .B1(net3792),
    .Y(_01713_));
 sky130_fd_sc_hd__nor3_2 _22399_ (.A(net3785),
    .B(_01388_),
    .C(_01713_),
    .Y(_01714_));
 sky130_fd_sc_hd__a21oi_1 _22400_ (.A1(net3786),
    .A2(_01711_),
    .B1(_01714_),
    .Y(_01715_));
 sky130_fd_sc_hd__a21oi_1 _22401_ (.A1(_01709_),
    .A2(_01715_),
    .B1(_01417_),
    .Y(_01716_));
 sky130_fd_sc_hd__nand2_1 _22402_ (.A(_12374_[0]),
    .B(_01463_),
    .Y(_01717_));
 sky130_fd_sc_hd__o21ai_0 _22403_ (.A1(_01401_),
    .A2(net3606),
    .B1(net3797),
    .Y(_01718_));
 sky130_fd_sc_hd__a31oi_1 _22404_ (.A1(_01717_),
    .A2(_01540_),
    .A3(_01718_),
    .B1(_01546_),
    .Y(_01719_));
 sky130_fd_sc_hd__a21oi_1 _22405_ (.A1(_01442_),
    .A2(_01547_),
    .B1(net3798),
    .Y(_01720_));
 sky130_fd_sc_hd__o311ai_0 _22406_ (.A1(_12366_[0]),
    .A2(_01354_),
    .A3(net3790),
    .B1(_01644_),
    .C1(_01707_),
    .Y(_01721_));
 sky130_fd_sc_hd__nor2_1 _22407_ (.A(_01720_),
    .B(_01721_),
    .Y(_01722_));
 sky130_fd_sc_hd__nor2_1 _22408_ (.A(net3656),
    .B(_01369_),
    .Y(_01723_));
 sky130_fd_sc_hd__a2111oi_1 _22409_ (.A1(net3655),
    .A2(_01660_),
    .B1(_01723_),
    .C1(_01552_),
    .D1(net3605),
    .Y(_01724_));
 sky130_fd_sc_hd__nor2_1 _22410_ (.A(_12376_[0]),
    .B(net3792),
    .Y(_01725_));
 sky130_fd_sc_hd__a21oi_1 _22411_ (.A1(net3792),
    .A2(_01558_),
    .B1(_01725_),
    .Y(_01726_));
 sky130_fd_sc_hd__o21ai_0 _22412_ (.A1(_01599_),
    .A2(_01726_),
    .B1(_01417_),
    .Y(_01727_));
 sky130_fd_sc_hd__o41ai_1 _22413_ (.A1(_01719_),
    .A2(_01722_),
    .A3(_01724_),
    .A4(_01727_),
    .B1(_01452_),
    .Y(_01728_));
 sky130_fd_sc_hd__a21oi_1 _22414_ (.A1(_01489_),
    .A2(_01660_),
    .B1(net3798),
    .Y(_01729_));
 sky130_fd_sc_hd__a311oi_1 _22415_ (.A1(net3798),
    .A2(_01644_),
    .A3(_01586_),
    .B1(_01729_),
    .C1(net3786),
    .Y(_01730_));
 sky130_fd_sc_hd__or3_1 _22416_ (.A(_12374_[0]),
    .B(net3654),
    .C(_01395_),
    .X(_01731_));
 sky130_fd_sc_hd__o21ai_0 _22417_ (.A1(_01568_),
    .A2(_01680_),
    .B1(_01731_),
    .Y(_01732_));
 sky130_fd_sc_hd__nor4_1 _22418_ (.A(net3784),
    .B(_01448_),
    .C(_01730_),
    .D(_01732_),
    .Y(_01733_));
 sky130_fd_sc_hd__nand3_1 _22419_ (.A(net3654),
    .B(_01547_),
    .C(_01507_),
    .Y(_01734_));
 sky130_fd_sc_hd__o211ai_1 _22420_ (.A1(net3654),
    .A2(_01461_),
    .B1(_01660_),
    .C1(net3786),
    .Y(_01735_));
 sky130_fd_sc_hd__nand3_1 _22421_ (.A(_01386_),
    .B(_01448_),
    .C(_01735_),
    .Y(_01736_));
 sky130_fd_sc_hd__a31oi_1 _22422_ (.A1(_01395_),
    .A2(_01621_),
    .A3(_01734_),
    .B1(_01736_),
    .Y(_01737_));
 sky130_fd_sc_hd__nand2b_2 _22423_ (.A_N(_12364_[0]),
    .B(net3798),
    .Y(_01738_));
 sky130_fd_sc_hd__a21oi_1 _22424_ (.A1(_01392_),
    .A2(_01738_),
    .B1(net3789),
    .Y(_01739_));
 sky130_fd_sc_hd__o211ai_1 _22425_ (.A1(_12369_[0]),
    .A2(net3793),
    .B1(_01644_),
    .C1(net3797),
    .Y(_01740_));
 sky130_fd_sc_hd__o311ai_0 _22426_ (.A1(net3797),
    .A2(_01375_),
    .A3(_01592_),
    .B1(_01740_),
    .C1(net3786),
    .Y(_01741_));
 sky130_fd_sc_hd__o2111a_4 _22427_ (.A1(_01468_),
    .A2(_01739_),
    .B1(_01741_),
    .C1(net3785),
    .D1(_01417_),
    .X(_01742_));
 sky130_fd_sc_hd__o21ai_0 _22428_ (.A1(net3796),
    .A2(_01379_),
    .B1(net3800),
    .Y(_01743_));
 sky130_fd_sc_hd__a21oi_1 _22429_ (.A1(_01343_),
    .A2(_01743_),
    .B1(net3604),
    .Y(_01744_));
 sky130_fd_sc_hd__a221oi_1 _22430_ (.A1(_01343_),
    .A2(net3603),
    .B1(_01702_),
    .B2(_12364_[0]),
    .C1(net3788),
    .Y(_01745_));
 sky130_fd_sc_hd__a21oi_1 _22431_ (.A1(net3788),
    .A2(_01744_),
    .B1(_01745_),
    .Y(_01746_));
 sky130_fd_sc_hd__a21oi_1 _22432_ (.A1(_01434_),
    .A2(_01690_),
    .B1(_01343_),
    .Y(_01747_));
 sky130_fd_sc_hd__nor4_1 _22433_ (.A(net3782),
    .B(_01417_),
    .C(_01746_),
    .D(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__nor4_1 _22434_ (.A(_01733_),
    .B(_01737_),
    .C(_01742_),
    .D(_01748_),
    .Y(_01749_));
 sky130_fd_sc_hd__o22ai_1 _22435_ (.A1(_01716_),
    .A2(_01728_),
    .B1(_01749_),
    .B2(_01452_),
    .Y(_00132_));
 sky130_fd_sc_hd__o21ai_0 _22436_ (.A1(_01349_),
    .A2(_01405_),
    .B1(_01666_),
    .Y(_01750_));
 sky130_fd_sc_hd__nand2_2 _22437_ (.A(_12369_[0]),
    .B(net3655),
    .Y(_01751_));
 sky130_fd_sc_hd__a21oi_1 _22438_ (.A1(_01621_),
    .A2(_01751_),
    .B1(net3793),
    .Y(_01752_));
 sky130_fd_sc_hd__nor3_1 _22439_ (.A(net3781),
    .B(_01388_),
    .C(_01752_),
    .Y(_01753_));
 sky130_fd_sc_hd__a21oi_1 _22440_ (.A1(_01385_),
    .A2(_01750_),
    .B1(_01753_),
    .Y(_01754_));
 sky130_fd_sc_hd__nor2_1 _22441_ (.A(net3796),
    .B(_01590_),
    .Y(_01755_));
 sky130_fd_sc_hd__a32oi_1 _22442_ (.A1(net3797),
    .A2(_01441_),
    .A3(_01525_),
    .B1(_01755_),
    .B2(_01644_),
    .Y(_01756_));
 sky130_fd_sc_hd__a21oi_1 _22443_ (.A1(_01488_),
    .A2(_01527_),
    .B1(net3797),
    .Y(_01757_));
 sky130_fd_sc_hd__a211oi_1 _22444_ (.A1(net3797),
    .A2(_01485_),
    .B1(_01757_),
    .C1(net3782),
    .Y(_01758_));
 sky130_fd_sc_hd__a21oi_1 _22445_ (.A1(net3782),
    .A2(_01756_),
    .B1(_01758_),
    .Y(_01759_));
 sky130_fd_sc_hd__nand2_1 _22446_ (.A(_01379_),
    .B(_01421_),
    .Y(_01760_));
 sky130_fd_sc_hd__o22ai_1 _22447_ (.A1(_01579_),
    .A2(_01754_),
    .B1(_01759_),
    .B2(_01760_),
    .Y(_01761_));
 sky130_fd_sc_hd__o21ai_0 _22448_ (.A1(net3656),
    .A2(net3651),
    .B1(_01540_),
    .Y(_01762_));
 sky130_fd_sc_hd__a21oi_1 _22449_ (.A1(_01385_),
    .A2(_01762_),
    .B1(_01448_),
    .Y(_01763_));
 sky130_fd_sc_hd__a21oi_1 _22450_ (.A1(_01343_),
    .A2(_01409_),
    .B1(_01401_),
    .Y(_01764_));
 sky130_fd_sc_hd__a22oi_1 _22451_ (.A1(net3800),
    .A2(net3607),
    .B1(_01463_),
    .B2(_12372_[0]),
    .Y(_01765_));
 sky130_fd_sc_hd__o21ai_1 _22452_ (.A1(net3800),
    .A2(_01764_),
    .B1(_01765_),
    .Y(_01766_));
 sky130_fd_sc_hd__a21oi_1 _22453_ (.A1(_01437_),
    .A2(_01429_),
    .B1(net3797),
    .Y(_01767_));
 sky130_fd_sc_hd__a211oi_1 _22454_ (.A1(net3802),
    .A2(net3607),
    .B1(_01546_),
    .C1(_01767_),
    .Y(_01768_));
 sky130_fd_sc_hd__o21ai_0 _22455_ (.A1(_12364_[0]),
    .A2(_01373_),
    .B1(_01527_),
    .Y(_01769_));
 sky130_fd_sc_hd__a211oi_1 _22456_ (.A1(net3655),
    .A2(_01769_),
    .B1(_01582_),
    .C1(_01481_),
    .Y(_01770_));
 sky130_fd_sc_hd__a211oi_1 _22457_ (.A1(_01616_),
    .A2(_01766_),
    .B1(_01768_),
    .C1(_01770_),
    .Y(_01771_));
 sky130_fd_sc_hd__nand2_1 _22458_ (.A(_01438_),
    .B(_01616_),
    .Y(_01772_));
 sky130_fd_sc_hd__a211oi_1 _22459_ (.A1(_12374_[0]),
    .A2(net3651),
    .B1(_01457_),
    .C1(_01772_),
    .Y(_01773_));
 sky130_fd_sc_hd__o311a_1 _22460_ (.A1(net3655),
    .A2(_01548_),
    .A3(_01461_),
    .B1(_01407_),
    .C1(_01385_),
    .X(_01774_));
 sky130_fd_sc_hd__nand2_2 _22461_ (.A(net3798),
    .B(_01561_),
    .Y(_01775_));
 sky130_fd_sc_hd__nor3_1 _22462_ (.A(net3800),
    .B(net3797),
    .C(_01373_),
    .Y(_01776_));
 sky130_fd_sc_hd__a311oi_1 _22463_ (.A1(net3797),
    .A2(_01489_),
    .A3(_01660_),
    .B1(_01776_),
    .C1(net3786),
    .Y(_01777_));
 sky130_fd_sc_hd__a311oi_1 _22464_ (.A1(net3786),
    .A2(_01644_),
    .A3(_01775_),
    .B1(_01777_),
    .C1(net3782),
    .Y(_01778_));
 sky130_fd_sc_hd__o41ai_1 _22465_ (.A1(_01417_),
    .A2(_01773_),
    .A3(_01774_),
    .A4(_01778_),
    .B1(_01420_),
    .Y(_01779_));
 sky130_fd_sc_hd__a21oi_1 _22466_ (.A1(_01763_),
    .A2(_01771_),
    .B1(_01779_),
    .Y(_01780_));
 sky130_fd_sc_hd__a31oi_1 _22467_ (.A1(net3797),
    .A2(_01489_),
    .A3(_01525_),
    .B1(_01757_),
    .Y(_01781_));
 sky130_fd_sc_hd__nand2_1 _22468_ (.A(_01373_),
    .B(_01751_),
    .Y(_01782_));
 sky130_fd_sc_hd__o211ai_1 _22469_ (.A1(net3592),
    .A2(_01479_),
    .B1(_01782_),
    .C1(net3782),
    .Y(_01783_));
 sky130_fd_sc_hd__o21ai_0 _22470_ (.A1(net3782),
    .A2(_01781_),
    .B1(_01783_),
    .Y(_01784_));
 sky130_fd_sc_hd__o32ai_1 _22471_ (.A1(_01400_),
    .A2(_01505_),
    .A3(_01506_),
    .B1(_01653_),
    .B2(net3652),
    .Y(_01785_));
 sky130_fd_sc_hd__a221oi_1 _22472_ (.A1(_12372_[0]),
    .A2(net3792),
    .B1(_01484_),
    .B2(_01427_),
    .C1(_01582_),
    .Y(_01786_));
 sky130_fd_sc_hd__nor2_1 _22473_ (.A(_01503_),
    .B(_01786_),
    .Y(_01787_));
 sky130_fd_sc_hd__o21ai_0 _22474_ (.A1(_01599_),
    .A2(_01785_),
    .B1(_01787_),
    .Y(_01788_));
 sky130_fd_sc_hd__a21oi_1 _22475_ (.A1(_01379_),
    .A2(_01784_),
    .B1(_01788_),
    .Y(_01789_));
 sky130_fd_sc_hd__nor3_1 _22476_ (.A(_01761_),
    .B(_01780_),
    .C(_01789_),
    .Y(_00133_));
 sky130_fd_sc_hd__a21oi_1 _22477_ (.A1(_01538_),
    .A2(_01660_),
    .B1(_01354_),
    .Y(_01790_));
 sky130_fd_sc_hd__a21oi_1 _22478_ (.A1(_12366_[0]),
    .A2(_01463_),
    .B1(_01790_),
    .Y(_01791_));
 sky130_fd_sc_hd__o211ai_1 _22479_ (.A1(net3788),
    .A2(_01613_),
    .B1(_01683_),
    .C1(net3652),
    .Y(_01792_));
 sky130_fd_sc_hd__nand3_1 _22480_ (.A(net3797),
    .B(_01510_),
    .C(_01660_),
    .Y(_01793_));
 sky130_fd_sc_hd__nand3_1 _22481_ (.A(net3784),
    .B(_01792_),
    .C(_01793_),
    .Y(_01794_));
 sky130_fd_sc_hd__o21ai_0 _22482_ (.A1(_01384_),
    .A2(_01791_),
    .B1(_01794_),
    .Y(_01795_));
 sky130_fd_sc_hd__o21ai_2 _22483_ (.A1(_01343_),
    .A2(_01354_),
    .B1(_01562_),
    .Y(_01796_));
 sky130_fd_sc_hd__o31ai_2 _22484_ (.A1(_12381_[0]),
    .A2(_12390_[0]),
    .A3(net3792),
    .B1(_01796_),
    .Y(_01797_));
 sky130_fd_sc_hd__nor3_1 _22485_ (.A(_01354_),
    .B(_01455_),
    .C(_01592_),
    .Y(_01798_));
 sky130_fd_sc_hd__nor3_1 _22486_ (.A(net3796),
    .B(_01521_),
    .C(_01590_),
    .Y(_01799_));
 sky130_fd_sc_hd__nor3_1 _22487_ (.A(net3781),
    .B(_01798_),
    .C(_01799_),
    .Y(_01800_));
 sky130_fd_sc_hd__a211oi_1 _22488_ (.A1(net3781),
    .A2(_01797_),
    .B1(_01800_),
    .C1(net3787),
    .Y(_01801_));
 sky130_fd_sc_hd__a211oi_1 _22489_ (.A1(net3787),
    .A2(_01795_),
    .B1(_01801_),
    .C1(_01417_),
    .Y(_01802_));
 sky130_fd_sc_hd__a21oi_1 _22490_ (.A1(net3788),
    .A2(_01613_),
    .B1(net3653),
    .Y(_01803_));
 sky130_fd_sc_hd__a32oi_1 _22491_ (.A1(net3653),
    .A2(_01442_),
    .A3(_01489_),
    .B1(_01803_),
    .B2(_01644_),
    .Y(_01804_));
 sky130_fd_sc_hd__nand2_1 _22492_ (.A(net3780),
    .B(_01804_),
    .Y(_01805_));
 sky130_fd_sc_hd__o21ai_0 _22493_ (.A1(net3802),
    .A2(net3604),
    .B1(net3795),
    .Y(_01806_));
 sky130_fd_sc_hd__nand2b_1 _22494_ (.A_N(_01460_),
    .B(_01806_),
    .Y(_01807_));
 sky130_fd_sc_hd__nor2_1 _22495_ (.A(net3630),
    .B(net3652),
    .Y(_01808_));
 sky130_fd_sc_hd__a21oi_1 _22496_ (.A1(net3652),
    .A2(_01679_),
    .B1(_01808_),
    .Y(_01809_));
 sky130_fd_sc_hd__nand2_1 _22497_ (.A(_12383_[0]),
    .B(net3791),
    .Y(_01810_));
 sky130_fd_sc_hd__o21ai_0 _22498_ (.A1(net3791),
    .A2(_01809_),
    .B1(_01810_),
    .Y(_01811_));
 sky130_fd_sc_hd__a311oi_1 _22499_ (.A1(_01683_),
    .A2(_01507_),
    .A3(_01677_),
    .B1(_01452_),
    .C1(net3784),
    .Y(_01812_));
 sky130_fd_sc_hd__o21ai_0 _22500_ (.A1(_01462_),
    .A2(_01701_),
    .B1(_01812_),
    .Y(_01813_));
 sky130_fd_sc_hd__a21oi_1 _22501_ (.A1(_01379_),
    .A2(_01811_),
    .B1(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__a311oi_1 _22502_ (.A1(_01700_),
    .A2(_01805_),
    .A3(_01807_),
    .B1(_01814_),
    .C1(_01664_),
    .Y(_01815_));
 sky130_fd_sc_hd__o211ai_1 _22503_ (.A1(net3656),
    .A2(net3780),
    .B1(_01434_),
    .C1(net3653),
    .Y(_01816_));
 sky130_fd_sc_hd__o21ai_0 _22504_ (.A1(_12374_[0]),
    .A2(net3787),
    .B1(net3791),
    .Y(_01817_));
 sky130_fd_sc_hd__o211ai_1 _22505_ (.A1(net3787),
    .A2(_01489_),
    .B1(_01817_),
    .C1(net3796),
    .Y(_01818_));
 sky130_fd_sc_hd__o2bb2ai_1 _22506_ (.A1_N(_01816_),
    .A2_N(_01818_),
    .B1(net3800),
    .B2(_01605_),
    .Y(_01819_));
 sky130_fd_sc_hd__a21boi_0 _22507_ (.A1(net3802),
    .A2(_01505_),
    .B1_N(_01411_),
    .Y(_01820_));
 sky130_fd_sc_hd__a21oi_1 _22508_ (.A1(net3802),
    .A2(net3606),
    .B1(_01506_),
    .Y(_01821_));
 sky130_fd_sc_hd__o21ai_0 _22509_ (.A1(_12378_[0]),
    .A2(_01820_),
    .B1(_01821_),
    .Y(_01822_));
 sky130_fd_sc_hd__a21oi_1 _22510_ (.A1(net3791),
    .A2(net3604),
    .B1(_01679_),
    .Y(_01823_));
 sky130_fd_sc_hd__o21ai_0 _22511_ (.A1(net3780),
    .A2(_01592_),
    .B1(_01622_),
    .Y(_01824_));
 sky130_fd_sc_hd__o2111ai_1 _22512_ (.A1(net3787),
    .A2(_01823_),
    .B1(_01824_),
    .C1(_01421_),
    .D1(net3781),
    .Y(_01825_));
 sky130_fd_sc_hd__a21oi_1 _22513_ (.A1(net3787),
    .A2(_01822_),
    .B1(_01825_),
    .Y(_01826_));
 sky130_fd_sc_hd__a31oi_1 _22514_ (.A1(_01384_),
    .A2(_01421_),
    .A3(_01819_),
    .B1(_01826_),
    .Y(_01827_));
 sky130_fd_sc_hd__nand2_1 _22515_ (.A(net3796),
    .B(_01671_),
    .Y(_01828_));
 sky130_fd_sc_hd__and3_4 _22516_ (.A(net3787),
    .B(_01652_),
    .C(_01828_),
    .X(_01829_));
 sky130_fd_sc_hd__a31oi_1 _22517_ (.A1(net3780),
    .A2(net393),
    .A3(_01467_),
    .B1(_01829_),
    .Y(_01830_));
 sky130_fd_sc_hd__a211oi_1 _22518_ (.A1(_12374_[0]),
    .A2(net3655),
    .B1(net3793),
    .C1(_01622_),
    .Y(_01831_));
 sky130_fd_sc_hd__a21oi_2 _22519_ (.A1(_12382_[0]),
    .A2(net3793),
    .B1(_01831_),
    .Y(_01832_));
 sky130_fd_sc_hd__nor3_1 _22520_ (.A(_01481_),
    .B(_01552_),
    .C(_01695_),
    .Y(_01833_));
 sky130_fd_sc_hd__nor2_1 _22521_ (.A(_01503_),
    .B(_01833_),
    .Y(_01834_));
 sky130_fd_sc_hd__o221ai_1 _22522_ (.A1(net3781),
    .A2(_01830_),
    .B1(_01832_),
    .B2(_01599_),
    .C1(_01834_),
    .Y(_01835_));
 sky130_fd_sc_hd__o211ai_1 _22523_ (.A1(_01802_),
    .A2(_01815_),
    .B1(_01827_),
    .C1(_01835_),
    .Y(_00134_));
 sky130_fd_sc_hd__o21ai_0 _22524_ (.A1(net3651),
    .A2(_01609_),
    .B1(_01349_),
    .Y(_01836_));
 sky130_fd_sc_hd__nand2_1 _22525_ (.A(_01505_),
    .B(_01606_),
    .Y(_01837_));
 sky130_fd_sc_hd__a21oi_1 _22526_ (.A1(_01836_),
    .A2(_01837_),
    .B1(net3802),
    .Y(_01838_));
 sky130_fd_sc_hd__o21ai_0 _22527_ (.A1(net3652),
    .A2(_01489_),
    .B1(_01701_),
    .Y(_01839_));
 sky130_fd_sc_hd__nor3_1 _22528_ (.A(net3781),
    .B(_01838_),
    .C(_01839_),
    .Y(_01840_));
 sky130_fd_sc_hd__a21oi_1 _22529_ (.A1(_01442_),
    .A2(_01459_),
    .B1(net3656),
    .Y(_01841_));
 sky130_fd_sc_hd__o21ai_0 _22530_ (.A1(net3605),
    .A2(_01841_),
    .B1(net3780),
    .Y(_01842_));
 sky130_fd_sc_hd__o21ai_0 _22531_ (.A1(net393),
    .A2(_01621_),
    .B1(_01479_),
    .Y(_01843_));
 sky130_fd_sc_hd__o21ai_0 _22532_ (.A1(_01349_),
    .A2(_01369_),
    .B1(_01411_),
    .Y(_01844_));
 sky130_fd_sc_hd__a22oi_1 _22533_ (.A1(net3656),
    .A2(_01843_),
    .B1(_01844_),
    .B2(net3787),
    .Y(_01845_));
 sky130_fd_sc_hd__a21oi_1 _22534_ (.A1(_01842_),
    .A2(_01845_),
    .B1(_01384_),
    .Y(_01846_));
 sky130_fd_sc_hd__nor3_2 _22535_ (.A(_01503_),
    .B(_01840_),
    .C(_01846_),
    .Y(_01847_));
 sky130_fd_sc_hd__nand2_1 _22536_ (.A(_12374_[0]),
    .B(net3797),
    .Y(_01848_));
 sky130_fd_sc_hd__a21oi_1 _22537_ (.A1(_01498_),
    .A2(_01848_),
    .B1(net3792),
    .Y(_01849_));
 sky130_fd_sc_hd__a211oi_1 _22538_ (.A1(_12390_[0]),
    .A2(net3794),
    .B1(_01849_),
    .C1(_01386_),
    .Y(_01850_));
 sky130_fd_sc_hd__nor2_1 _22539_ (.A(_12376_[0]),
    .B(net3789),
    .Y(_01851_));
 sky130_fd_sc_hd__a311oi_1 _22540_ (.A1(_12366_[0]),
    .A2(_01354_),
    .A3(net3789),
    .B1(_01851_),
    .C1(net3784),
    .Y(_01852_));
 sky130_fd_sc_hd__nor3_1 _22541_ (.A(net3786),
    .B(_01850_),
    .C(_01852_),
    .Y(_01853_));
 sky130_fd_sc_hd__a311oi_1 _22542_ (.A1(net3798),
    .A2(_01400_),
    .A3(_01525_),
    .B1(_01532_),
    .C1(_01546_),
    .Y(_01854_));
 sky130_fd_sc_hd__o21ai_0 _22543_ (.A1(_01400_),
    .A2(_01493_),
    .B1(_01616_),
    .Y(_01855_));
 sky130_fd_sc_hd__a31oi_1 _22544_ (.A1(net3794),
    .A2(_01392_),
    .A3(_01712_),
    .B1(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__nor4b_1 _22545_ (.A(_01853_),
    .B(_01854_),
    .C(_01856_),
    .D_N(_01453_),
    .Y(_01857_));
 sky130_fd_sc_hd__nor2_1 _22546_ (.A(_12365_[0]),
    .B(_01692_),
    .Y(_01858_));
 sky130_fd_sc_hd__and3_1 _22547_ (.A(net3797),
    .B(_01442_),
    .C(_01527_),
    .X(_01859_));
 sky130_fd_sc_hd__a211o_1 _22548_ (.A1(net3655),
    .A2(_01581_),
    .B1(_01859_),
    .C1(net3786),
    .X(_01860_));
 sky130_fd_sc_hd__o41ai_1 _22549_ (.A1(net3780),
    .A2(_01542_),
    .A3(_01638_),
    .A4(_01858_),
    .B1(_01860_),
    .Y(_01861_));
 sky130_fd_sc_hd__nor2_1 _22550_ (.A(_01549_),
    .B(_01776_),
    .Y(_01862_));
 sky130_fd_sc_hd__nor2_1 _22551_ (.A(net3802),
    .B(_01862_),
    .Y(_01863_));
 sky130_fd_sc_hd__a2111oi_0 _22552_ (.A1(_12364_[0]),
    .A2(_01409_),
    .B1(_01552_),
    .C1(_01542_),
    .D1(_01863_),
    .Y(_01864_));
 sky130_fd_sc_hd__o21ai_0 _22553_ (.A1(_12374_[0]),
    .A2(_01479_),
    .B1(_01385_),
    .Y(_01865_));
 sky130_fd_sc_hd__a31oi_1 _22554_ (.A1(net3797),
    .A2(_01507_),
    .A3(_01527_),
    .B1(_01865_),
    .Y(_01866_));
 sky130_fd_sc_hd__a2111oi_1 _22555_ (.A1(_01384_),
    .A2(_01861_),
    .B1(_01864_),
    .C1(_01866_),
    .D1(_01579_),
    .Y(_01867_));
 sky130_fd_sc_hd__nor3_1 _22556_ (.A(net3798),
    .B(_01443_),
    .C(_01485_),
    .Y(_01868_));
 sky130_fd_sc_hd__a311oi_1 _22557_ (.A1(net3798),
    .A2(_01525_),
    .A3(_01538_),
    .B1(_01868_),
    .C1(net3784),
    .Y(_01869_));
 sky130_fd_sc_hd__nand3b_1 _22558_ (.A_N(_01461_),
    .B(_01507_),
    .C(_01354_),
    .Y(_01870_));
 sky130_fd_sc_hd__a21oi_1 _22559_ (.A1(_01738_),
    .A2(_01870_),
    .B1(net3783),
    .Y(_01871_));
 sky130_fd_sc_hd__nand3_1 _22560_ (.A(_01354_),
    .B(_01510_),
    .C(_01660_),
    .Y(_01872_));
 sky130_fd_sc_hd__a21oi_1 _22561_ (.A1(_01614_),
    .A2(_01872_),
    .B1(_01401_),
    .Y(_01873_));
 sky130_fd_sc_hd__o211ai_1 _22562_ (.A1(_12369_[0]),
    .A2(net3794),
    .B1(_01796_),
    .C1(net3785),
    .Y(_01874_));
 sky130_fd_sc_hd__o2111ai_1 _22563_ (.A1(net3785),
    .A2(_01873_),
    .B1(_01874_),
    .C1(_01664_),
    .D1(net3786),
    .Y(_01875_));
 sky130_fd_sc_hd__o41ai_1 _22564_ (.A1(net3786),
    .A2(_01449_),
    .A3(_01869_),
    .A4(_01871_),
    .B1(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__nor4_1 _22565_ (.A(_01847_),
    .B(_01857_),
    .C(_01867_),
    .D(_01876_),
    .Y(_00135_));
 sky130_fd_sc_hd__xor3_1 _22566_ (.A(\sa01_sr[7] ),
    .B(net4228),
    .C(\sa21_sr[1] ),
    .X(_01877_));
 sky130_fd_sc_hd__xnor3_1 _22567_ (.A(_11059_),
    .B(_11060_),
    .C(_01877_),
    .X(_01878_));
 sky130_fd_sc_hd__nand2_1 _22568_ (.A(net4230),
    .B(\text_in_r[65] ),
    .Y(_01879_));
 sky130_fd_sc_hd__o21a_1 _22569_ (.A1(net398),
    .A2(_01878_),
    .B1(_01879_),
    .X(_01880_));
 sky130_fd_sc_hd__xor2_1 _22570_ (.A(net4153),
    .B(_01880_),
    .X(_01881_));
 sky130_fd_sc_hd__inv_16 _22571_ (.A(net3778),
    .Y(_01882_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_193 ();
 sky130_fd_sc_hd__xnor3_1 _22573_ (.A(\sa30_sub[7] ),
    .B(_06477_),
    .C(_06489_),
    .X(_01883_));
 sky130_fd_sc_hd__mux2i_2 _22574_ (.A0(\text_in_r[64] ),
    .A1(_01883_),
    .S(net4111),
    .Y(_01884_));
 sky130_fd_sc_hd__xor2_4 _22575_ (.A(net4157),
    .B(_01884_),
    .X(_01885_));
 sky130_fd_sc_hd__clkinv_8 _22576_ (.A(_01885_),
    .Y(_01886_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_191 ();
 sky130_fd_sc_hd__xor2_1 _22579_ (.A(\sa30_sub[1] ),
    .B(net4226),
    .X(_01888_));
 sky130_fd_sc_hd__xnor2_1 _22580_ (.A(_06495_),
    .B(_01888_),
    .Y(_01889_));
 sky130_fd_sc_hd__mux2i_2 _22581_ (.A0(\text_in_r[66] ),
    .A1(_01889_),
    .S(net4111),
    .Y(_01890_));
 sky130_fd_sc_hd__xnor2_4 _22582_ (.A(\u0.w[1][2] ),
    .B(_01890_),
    .Y(_01891_));
 sky130_fd_sc_hd__clkinv_16 _22583_ (.A(_01891_),
    .Y(_01892_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_184 ();
 sky130_fd_sc_hd__xnor2_2 _22591_ (.A(_06605_),
    .B(_11088_),
    .Y(_01897_));
 sky130_fd_sc_hd__nand2_2 _22592_ (.A(net4111),
    .B(_01897_),
    .Y(_01898_));
 sky130_fd_sc_hd__o21ai_4 _22593_ (.A1(net4112),
    .A2(\text_in_r[71] ),
    .B1(_01898_),
    .Y(_01899_));
 sky130_fd_sc_hd__xor2_2 _22594_ (.A(\u0.w[1][7] ),
    .B(_01899_),
    .X(_01900_));
 sky130_fd_sc_hd__xnor2_1 _22595_ (.A(\sa01_sr[5] ),
    .B(\sa21_sr[6] ),
    .Y(_01901_));
 sky130_fd_sc_hd__xnor2_1 _22596_ (.A(_11083_),
    .B(_01901_),
    .Y(_01902_));
 sky130_fd_sc_hd__nor2_2 _22597_ (.A(net398),
    .B(_01902_),
    .Y(_01903_));
 sky130_fd_sc_hd__a21oi_4 _22598_ (.A1(net398),
    .A2(\text_in_r[70] ),
    .B1(_01903_),
    .Y(_01904_));
 sky130_fd_sc_hd__xnor2_4 _22599_ (.A(net4142),
    .B(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__nor2_4 _22600_ (.A(_01900_),
    .B(_01905_),
    .Y(_01906_));
 sky130_fd_sc_hd__xor2_1 _22601_ (.A(net4187),
    .B(\sa01_sr[5] ),
    .X(_01907_));
 sky130_fd_sc_hd__xnor2_1 _22602_ (.A(_06560_),
    .B(_01907_),
    .Y(_01908_));
 sky130_fd_sc_hd__mux2i_4 _22603_ (.A0(\text_in_r[69] ),
    .A1(_01908_),
    .S(net4113),
    .Y(_01909_));
 sky130_fd_sc_hd__xnor2_4 _22604_ (.A(\u0.w[1][5] ),
    .B(_01909_),
    .Y(_01910_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_182 ();
 sky130_fd_sc_hd__nor2b_2 _22607_ (.A(net4230),
    .B_N(\u0.w[1][3] ),
    .Y(_01913_));
 sky130_fd_sc_hd__nor2_1 _22608_ (.A(\u0.w[1][3] ),
    .B(net4230),
    .Y(_01914_));
 sky130_fd_sc_hd__xnor3_1 _22609_ (.A(_06527_),
    .B(_11096_),
    .C(_11097_),
    .X(_01915_));
 sky130_fd_sc_hd__mux2i_4 _22610_ (.A0(_01913_),
    .A1(_01914_),
    .S(_01915_),
    .Y(_01916_));
 sky130_fd_sc_hd__nor2_2 _22611_ (.A(\u0.w[1][3] ),
    .B(net4112),
    .Y(_01917_));
 sky130_fd_sc_hd__nand2_1 _22612_ (.A(\u0.w[1][3] ),
    .B(net398),
    .Y(_01918_));
 sky130_fd_sc_hd__nor2_2 _22613_ (.A(\text_in_r[67] ),
    .B(_01918_),
    .Y(_01919_));
 sky130_fd_sc_hd__a21oi_4 _22614_ (.A1(\text_in_r[67] ),
    .A2(_01917_),
    .B1(_01919_),
    .Y(_01920_));
 sky130_fd_sc_hd__and2_4 _22615_ (.A(_01916_),
    .B(_01920_),
    .X(_01921_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_181 ();
 sky130_fd_sc_hd__nor2_4 _22617_ (.A(_01892_),
    .B(_01921_),
    .Y(_01923_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_177 ();
 sky130_fd_sc_hd__nand2_4 _22622_ (.A(net3771),
    .B(net3765),
    .Y(_01928_));
 sky130_fd_sc_hd__nand2_8 _22623_ (.A(_01916_),
    .B(_01920_),
    .Y(_01929_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_175 ();
 sky130_fd_sc_hd__nand2_2 _22626_ (.A(_01892_),
    .B(net3762),
    .Y(_01932_));
 sky130_fd_sc_hd__o21ai_0 _22627_ (.A1(net3778),
    .A2(_01928_),
    .B1(_01932_),
    .Y(_01933_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_174 ();
 sky130_fd_sc_hd__nor2_4 _22629_ (.A(_12398_[0]),
    .B(_12401_[0]),
    .Y(_01935_));
 sky130_fd_sc_hd__nor2_4 _22630_ (.A(net3775),
    .B(_01929_),
    .Y(_01936_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_173 ();
 sky130_fd_sc_hd__a222oi_1 _22632_ (.A1(_12396_[0]),
    .A2(_01923_),
    .B1(_01933_),
    .B2(net3777),
    .C1(_01935_),
    .C2(net3646),
    .Y(_01938_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_171 ();
 sky130_fd_sc_hd__nor2_4 _22635_ (.A(_12398_[0]),
    .B(net3762),
    .Y(_01941_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_170 ();
 sky130_fd_sc_hd__nor3_4 _22637_ (.A(net3779),
    .B(net3650),
    .C(net3765),
    .Y(_01943_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_169 ();
 sky130_fd_sc_hd__nor2_4 _22639_ (.A(net3771),
    .B(net3765),
    .Y(_01945_));
 sky130_fd_sc_hd__nand2_1 _22640_ (.A(_12406_[0]),
    .B(_01945_),
    .Y(_01946_));
 sky130_fd_sc_hd__o311ai_0 _22641_ (.A1(_01892_),
    .A2(_01941_),
    .A3(_01943_),
    .B1(_01946_),
    .C1(net3769),
    .Y(_01947_));
 sky130_fd_sc_hd__xor3_1 _22642_ (.A(_06512_),
    .B(_11117_),
    .C(_11118_),
    .X(_01948_));
 sky130_fd_sc_hd__mux2i_4 _22643_ (.A0(\text_in_r[68] ),
    .A1(_01948_),
    .S(net4113),
    .Y(_01949_));
 sky130_fd_sc_hd__xor2_4 _22644_ (.A(net4144),
    .B(_01949_),
    .X(_01950_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_167 ();
 sky130_fd_sc_hd__o211ai_1 _22647_ (.A1(net3769),
    .A2(_01938_),
    .B1(_01947_),
    .C1(net3758),
    .Y(_01953_));
 sky130_fd_sc_hd__xor2_4 _22648_ (.A(net4143),
    .B(_01909_),
    .X(_01954_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_164 ();
 sky130_fd_sc_hd__nand2_8 _22652_ (.A(net3649),
    .B(net3767),
    .Y(_01958_));
 sky130_fd_sc_hd__nor2_1 _22653_ (.A(_12404_[0]),
    .B(_01958_),
    .Y(_01959_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_163 ();
 sky130_fd_sc_hd__nand2_4 _22655_ (.A(_12398_[0]),
    .B(net3762),
    .Y(_01961_));
 sky130_fd_sc_hd__nor2_2 _22656_ (.A(net3778),
    .B(_01886_),
    .Y(_01962_));
 sky130_fd_sc_hd__o22ai_1 _22657_ (.A1(_01892_),
    .A2(_01961_),
    .B1(_01962_),
    .B2(_01928_),
    .Y(_01963_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_160 ();
 sky130_fd_sc_hd__a221o_1 _22661_ (.A1(_12417_[0]),
    .A2(net3762),
    .B1(net3646),
    .B2(_12397_[0]),
    .C1(net3769),
    .X(_01967_));
 sky130_fd_sc_hd__xnor2_4 _22662_ (.A(net4144),
    .B(_01949_),
    .Y(_01968_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_158 ();
 sky130_fd_sc_hd__o311ai_0 _22665_ (.A1(net3757),
    .A2(_01959_),
    .A3(_01963_),
    .B1(_01967_),
    .C1(net3752),
    .Y(_01971_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_156 ();
 sky130_fd_sc_hd__nor2_4 _22668_ (.A(_12397_[0]),
    .B(net3765),
    .Y(_01974_));
 sky130_fd_sc_hd__nor2_2 _22669_ (.A(_12406_[0]),
    .B(net3764),
    .Y(_01975_));
 sky130_fd_sc_hd__o21ai_0 _22670_ (.A1(_01974_),
    .A2(_01975_),
    .B1(net3771),
    .Y(_01976_));
 sky130_fd_sc_hd__o211ai_1 _22671_ (.A1(_12401_[0]),
    .A2(_01958_),
    .B1(net3757),
    .C1(_01976_),
    .Y(_01977_));
 sky130_fd_sc_hd__nor2_4 _22672_ (.A(_12401_[0]),
    .B(net3765),
    .Y(_01978_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_154 ();
 sky130_fd_sc_hd__o21ai_1 _22675_ (.A1(_01941_),
    .A2(_01978_),
    .B1(net3772),
    .Y(_01981_));
 sky130_fd_sc_hd__a21oi_1 _22676_ (.A1(_12396_[0]),
    .A2(net3646),
    .B1(net3757),
    .Y(_01982_));
 sky130_fd_sc_hd__a21oi_1 _22677_ (.A1(_01981_),
    .A2(_01982_),
    .B1(net3758),
    .Y(_01983_));
 sky130_fd_sc_hd__nand2_1 _22678_ (.A(_01977_),
    .B(_01983_),
    .Y(_01984_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_153 ();
 sky130_fd_sc_hd__nand2_2 _22680_ (.A(_12397_[0]),
    .B(_01892_),
    .Y(_01986_));
 sky130_fd_sc_hd__nand2_2 _22681_ (.A(_01882_),
    .B(net3771),
    .Y(_01987_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_151 ();
 sky130_fd_sc_hd__a31oi_2 _22684_ (.A1(net3765),
    .A2(_01986_),
    .A3(_01987_),
    .B1(net3752),
    .Y(_01990_));
 sky130_fd_sc_hd__nor2_4 _22685_ (.A(net3777),
    .B(_01892_),
    .Y(_01991_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_149 ();
 sky130_fd_sc_hd__nor2_1 _22688_ (.A(_12404_[0]),
    .B(net3771),
    .Y(_01994_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_148 ();
 sky130_fd_sc_hd__o21ai_0 _22690_ (.A1(net3601),
    .A2(_01994_),
    .B1(net3762),
    .Y(_01996_));
 sky130_fd_sc_hd__nand3_1 _22691_ (.A(net3769),
    .B(_01990_),
    .C(_01996_),
    .Y(_01997_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_146 ();
 sky130_fd_sc_hd__nand2_2 _22694_ (.A(net3777),
    .B(_01892_),
    .Y(_02000_));
 sky130_fd_sc_hd__nand2_1 _22695_ (.A(_01882_),
    .B(_01991_),
    .Y(_02001_));
 sky130_fd_sc_hd__a31oi_1 _22696_ (.A1(net3764),
    .A2(_02000_),
    .A3(_02001_),
    .B1(net3752),
    .Y(_02002_));
 sky130_fd_sc_hd__nand2_2 _22697_ (.A(_12401_[0]),
    .B(net3647),
    .Y(_02003_));
 sky130_fd_sc_hd__nand3_2 _22698_ (.A(_01954_),
    .B(_02002_),
    .C(_02003_),
    .Y(_02004_));
 sky130_fd_sc_hd__xnor2_4 _22699_ (.A(\u0.w[1][7] ),
    .B(_01899_),
    .Y(_02005_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_145 ();
 sky130_fd_sc_hd__nand2_8 _22701_ (.A(_02005_),
    .B(_01905_),
    .Y(_02007_));
 sky130_fd_sc_hd__a31oi_1 _22702_ (.A1(_01984_),
    .A2(_01997_),
    .A3(_02004_),
    .B1(_02007_),
    .Y(_02008_));
 sky130_fd_sc_hd__xnor2_4 _22703_ (.A(net3774),
    .B(net3763),
    .Y(_02009_));
 sky130_fd_sc_hd__nor2_1 _22704_ (.A(_12396_[0]),
    .B(_02009_),
    .Y(_02010_));
 sky130_fd_sc_hd__a211oi_1 _22705_ (.A1(_12397_[0]),
    .A2(_01923_),
    .B1(_01959_),
    .C1(_02010_),
    .Y(_02011_));
 sky130_fd_sc_hd__nor2_1 _22706_ (.A(net3779),
    .B(net3777),
    .Y(_02012_));
 sky130_fd_sc_hd__a22oi_1 _22707_ (.A1(_01882_),
    .A2(net3646),
    .B1(_01923_),
    .B2(_02012_),
    .Y(_02013_));
 sky130_fd_sc_hd__nand2_2 _22708_ (.A(net3777),
    .B(_01945_),
    .Y(_02014_));
 sky130_fd_sc_hd__o2111ai_1 _22709_ (.A1(_12398_[0]),
    .A2(_01928_),
    .B1(_02013_),
    .C1(_01905_),
    .D1(_02014_),
    .Y(_02015_));
 sky130_fd_sc_hd__o2111ai_1 _22710_ (.A1(_01905_),
    .A2(_02011_),
    .B1(net3758),
    .C1(net3757),
    .D1(_02015_),
    .Y(_02016_));
 sky130_fd_sc_hd__nand2_4 _22711_ (.A(net3779),
    .B(_01921_),
    .Y(_02017_));
 sky130_fd_sc_hd__nor2_4 _22712_ (.A(_12397_[0]),
    .B(net3771),
    .Y(_02018_));
 sky130_fd_sc_hd__nor2_2 _22713_ (.A(_01882_),
    .B(net3771),
    .Y(_02019_));
 sky130_fd_sc_hd__nand2_8 _22714_ (.A(_12397_[0]),
    .B(_01921_),
    .Y(_02020_));
 sky130_fd_sc_hd__nor2_1 _22715_ (.A(_02019_),
    .B(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hd__a21oi_1 _22716_ (.A1(_02017_),
    .A2(_02018_),
    .B1(_02021_),
    .Y(_02022_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_144 ();
 sky130_fd_sc_hd__nand2_2 _22718_ (.A(_12410_[0]),
    .B(net3763),
    .Y(_02024_));
 sky130_fd_sc_hd__nand2_4 _22719_ (.A(_01882_),
    .B(_01921_),
    .Y(_02025_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_143 ();
 sky130_fd_sc_hd__nor2_1 _22721_ (.A(net3650),
    .B(net3771),
    .Y(_02027_));
 sky130_fd_sc_hd__a32oi_1 _22722_ (.A1(net3771),
    .A2(_02024_),
    .A3(_02025_),
    .B1(_02017_),
    .B2(_02027_),
    .Y(_02028_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_142 ();
 sky130_fd_sc_hd__nand2_2 _22724_ (.A(net3756),
    .B(net3752),
    .Y(_02030_));
 sky130_fd_sc_hd__a21oi_1 _22725_ (.A1(_01905_),
    .A2(_02028_),
    .B1(_02030_),
    .Y(_02031_));
 sky130_fd_sc_hd__o21ai_2 _22726_ (.A1(_01905_),
    .A2(_02022_),
    .B1(_02031_),
    .Y(_02032_));
 sky130_fd_sc_hd__xor2_4 _22727_ (.A(\u0.w[1][6] ),
    .B(_01904_),
    .X(_02033_));
 sky130_fd_sc_hd__nand2_8 _22728_ (.A(net3774),
    .B(net3763),
    .Y(_02034_));
 sky130_fd_sc_hd__nor2_4 _22729_ (.A(_01882_),
    .B(net3765),
    .Y(_02035_));
 sky130_fd_sc_hd__o22ai_1 _22730_ (.A1(_12401_[0]),
    .A2(_02034_),
    .B1(_02035_),
    .B2(_02000_),
    .Y(_02036_));
 sky130_fd_sc_hd__nand2b_1 _22731_ (.A_N(_12410_[0]),
    .B(net3764),
    .Y(_02037_));
 sky130_fd_sc_hd__nand3_1 _22732_ (.A(_01892_),
    .B(_02025_),
    .C(_02037_),
    .Y(_02038_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_141 ();
 sky130_fd_sc_hd__nor2_4 _22734_ (.A(net3777),
    .B(net3763),
    .Y(_02040_));
 sky130_fd_sc_hd__a211oi_1 _22735_ (.A1(_12397_[0]),
    .A2(_01923_),
    .B1(_01950_),
    .C1(_02040_),
    .Y(_02041_));
 sky130_fd_sc_hd__a22oi_1 _22736_ (.A1(_01950_),
    .A2(_02036_),
    .B1(_02038_),
    .B2(_02041_),
    .Y(_02042_));
 sky130_fd_sc_hd__nand2_4 _22737_ (.A(net3649),
    .B(_01950_),
    .Y(_02043_));
 sky130_fd_sc_hd__nor2_1 _22738_ (.A(_01882_),
    .B(net3650),
    .Y(_02044_));
 sky130_fd_sc_hd__nand2_1 _22739_ (.A(net3753),
    .B(_02044_),
    .Y(_02045_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_140 ();
 sky130_fd_sc_hd__nor3_1 _22741_ (.A(_01905_),
    .B(net3767),
    .C(net3755),
    .Y(_02047_));
 sky130_fd_sc_hd__nand2_1 _22742_ (.A(_12404_[0]),
    .B(_01950_),
    .Y(_02048_));
 sky130_fd_sc_hd__o211ai_1 _22743_ (.A1(net3650),
    .A2(_01950_),
    .B1(_02048_),
    .C1(net3775),
    .Y(_02049_));
 sky130_fd_sc_hd__o2111ai_1 _22744_ (.A1(_12396_[0]),
    .A2(_02043_),
    .B1(_02045_),
    .C1(_02047_),
    .D1(_02049_),
    .Y(_02050_));
 sky130_fd_sc_hd__nand2_8 _22745_ (.A(_01882_),
    .B(net3650),
    .Y(_02051_));
 sky130_fd_sc_hd__nand2_2 _22746_ (.A(net3774),
    .B(_01968_),
    .Y(_02052_));
 sky130_fd_sc_hd__o22ai_1 _22747_ (.A1(_02051_),
    .A2(_02043_),
    .B1(_02052_),
    .B2(net3777),
    .Y(_02053_));
 sky130_fd_sc_hd__nand2_8 _22748_ (.A(net3779),
    .B(net3777),
    .Y(_02054_));
 sky130_fd_sc_hd__nand2_1 _22749_ (.A(net3774),
    .B(_01950_),
    .Y(_02055_));
 sky130_fd_sc_hd__o22ai_1 _22750_ (.A1(_01950_),
    .A2(_02054_),
    .B1(_02055_),
    .B2(_12397_[0]),
    .Y(_02056_));
 sky130_fd_sc_hd__nor2_2 _22751_ (.A(net3763),
    .B(net3755),
    .Y(_02057_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_139 ();
 sky130_fd_sc_hd__o211ai_1 _22753_ (.A1(_02053_),
    .A2(_02056_),
    .B1(_02057_),
    .C1(_02033_),
    .Y(_02059_));
 sky130_fd_sc_hd__o311a_4 _22754_ (.A1(_02033_),
    .A2(net3755),
    .A3(_02042_),
    .B1(_02050_),
    .C1(_02059_),
    .X(_02060_));
 sky130_fd_sc_hd__a31oi_1 _22755_ (.A1(_02016_),
    .A2(_02032_),
    .A3(_02060_),
    .B1(_02005_),
    .Y(_02061_));
 sky130_fd_sc_hd__a311oi_1 _22756_ (.A1(_01906_),
    .A2(_01953_),
    .A3(_01971_),
    .B1(_02008_),
    .C1(_02061_),
    .Y(_00136_));
 sky130_fd_sc_hd__nor3_2 _22757_ (.A(net3779),
    .B(net3777),
    .C(net3762),
    .Y(_02062_));
 sky130_fd_sc_hd__nor2_1 _22758_ (.A(_01882_),
    .B(_02034_),
    .Y(_02063_));
 sky130_fd_sc_hd__a211oi_1 _22759_ (.A1(net3649),
    .A2(_02024_),
    .B1(_02062_),
    .C1(_02063_),
    .Y(_02064_));
 sky130_fd_sc_hd__nor2_4 _22760_ (.A(net3650),
    .B(net3763),
    .Y(_02065_));
 sky130_fd_sc_hd__nand2_2 _22761_ (.A(_12397_[0]),
    .B(net3763),
    .Y(_02066_));
 sky130_fd_sc_hd__and3_4 _22762_ (.A(_12396_[0]),
    .B(_01916_),
    .C(_01920_),
    .X(_02067_));
 sky130_fd_sc_hd__nor2_1 _22763_ (.A(_01892_),
    .B(_02067_),
    .Y(_02068_));
 sky130_fd_sc_hd__nand2_1 _22764_ (.A(_02066_),
    .B(_02068_),
    .Y(_02069_));
 sky130_fd_sc_hd__o311ai_0 _22765_ (.A1(net3772),
    .A2(_01978_),
    .A3(_02065_),
    .B1(_02069_),
    .C1(net3757),
    .Y(_02070_));
 sky130_fd_sc_hd__o21ai_0 _22766_ (.A1(net3757),
    .A2(_02064_),
    .B1(_02070_),
    .Y(_02071_));
 sky130_fd_sc_hd__nor2_4 _22767_ (.A(net3777),
    .B(_01921_),
    .Y(_02072_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_138 ();
 sky130_fd_sc_hd__nor2_1 _22769_ (.A(net3650),
    .B(_02009_),
    .Y(_02073_));
 sky130_fd_sc_hd__a221oi_1 _22770_ (.A1(_12397_[0]),
    .A2(net3647),
    .B1(_02072_),
    .B2(net3779),
    .C1(_02073_),
    .Y(_02074_));
 sky130_fd_sc_hd__nand2b_4 _22771_ (.A_N(_12397_[0]),
    .B(net3763),
    .Y(_02075_));
 sky130_fd_sc_hd__nand2_2 _22772_ (.A(_12401_[0]),
    .B(net3765),
    .Y(_02076_));
 sky130_fd_sc_hd__a21oi_1 _22773_ (.A1(net3763),
    .A2(_02051_),
    .B1(net3774),
    .Y(_02077_));
 sky130_fd_sc_hd__a311oi_1 _22774_ (.A1(net3774),
    .A2(_02075_),
    .A3(_02076_),
    .B1(_02077_),
    .C1(net3755),
    .Y(_02078_));
 sky130_fd_sc_hd__a211oi_1 _22775_ (.A1(net3755),
    .A2(_02074_),
    .B1(_02078_),
    .C1(net3754),
    .Y(_02079_));
 sky130_fd_sc_hd__a21oi_1 _22776_ (.A1(_01968_),
    .A2(_02071_),
    .B1(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__nand2_1 _22777_ (.A(net3650),
    .B(_01892_),
    .Y(_02081_));
 sky130_fd_sc_hd__o21ai_0 _22778_ (.A1(_01945_),
    .A2(_02040_),
    .B1(net3779),
    .Y(_02082_));
 sky130_fd_sc_hd__a21oi_1 _22779_ (.A1(_02081_),
    .A2(_02082_),
    .B1(net3752),
    .Y(_02083_));
 sky130_fd_sc_hd__nand2_1 _22780_ (.A(net3779),
    .B(_01950_),
    .Y(_02084_));
 sky130_fd_sc_hd__a21oi_1 _22781_ (.A1(_02065_),
    .A2(_02084_),
    .B1(_02072_),
    .Y(_02085_));
 sky130_fd_sc_hd__nor2_1 _22782_ (.A(net3775),
    .B(_02085_),
    .Y(_02086_));
 sky130_fd_sc_hd__a21oi_1 _22783_ (.A1(_02066_),
    .A2(_02076_),
    .B1(_02052_),
    .Y(_02087_));
 sky130_fd_sc_hd__nor4_1 _22784_ (.A(_01954_),
    .B(_02083_),
    .C(_02086_),
    .D(_02087_),
    .Y(_02088_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_137 ();
 sky130_fd_sc_hd__nor2_4 _22786_ (.A(_12410_[0]),
    .B(net3765),
    .Y(_02090_));
 sky130_fd_sc_hd__nor3_4 _22787_ (.A(net3779),
    .B(net3650),
    .C(net3762),
    .Y(_02091_));
 sky130_fd_sc_hd__o21ai_0 _22788_ (.A1(_02090_),
    .A2(_02091_),
    .B1(net3772),
    .Y(_02092_));
 sky130_fd_sc_hd__nand3_1 _22789_ (.A(_01892_),
    .B(_02066_),
    .C(_02076_),
    .Y(_02093_));
 sky130_fd_sc_hd__o22ai_1 _22790_ (.A1(_12401_[0]),
    .A2(_01958_),
    .B1(_02009_),
    .B2(net3779),
    .Y(_02094_));
 sky130_fd_sc_hd__o21ai_0 _22791_ (.A1(net3758),
    .A2(_02094_),
    .B1(net3757),
    .Y(_02095_));
 sky130_fd_sc_hd__a31oi_1 _22792_ (.A1(net3760),
    .A2(_02092_),
    .A3(_02093_),
    .B1(_02095_),
    .Y(_02096_));
 sky130_fd_sc_hd__o21a_1 _22793_ (.A1(_02040_),
    .A2(_01978_),
    .B1(net3774),
    .X(_02097_));
 sky130_fd_sc_hd__nand2_4 _22794_ (.A(net3779),
    .B(net3762),
    .Y(_02098_));
 sky130_fd_sc_hd__a21oi_1 _22795_ (.A1(_02025_),
    .A2(_02098_),
    .B1(net3771),
    .Y(_02099_));
 sky130_fd_sc_hd__nor2_4 _22796_ (.A(net3769),
    .B(net3759),
    .Y(_02100_));
 sky130_fd_sc_hd__o21ai_0 _22797_ (.A1(_02097_),
    .A2(_02099_),
    .B1(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__nor2_4 _22798_ (.A(net3779),
    .B(net3767),
    .Y(_02102_));
 sky130_fd_sc_hd__nand2_1 _22799_ (.A(net3777),
    .B(net3775),
    .Y(_02103_));
 sky130_fd_sc_hd__and3_1 _22800_ (.A(_02102_),
    .B(_02081_),
    .C(_02103_),
    .X(_02104_));
 sky130_fd_sc_hd__nand2_1 _22801_ (.A(_12396_[0]),
    .B(net3649),
    .Y(_02105_));
 sky130_fd_sc_hd__a21oi_1 _22802_ (.A1(_02105_),
    .A2(_02103_),
    .B1(net3763),
    .Y(_02106_));
 sky130_fd_sc_hd__nor2_4 _22803_ (.A(_01954_),
    .B(net3760),
    .Y(_02107_));
 sky130_fd_sc_hd__o21ai_0 _22804_ (.A1(_02104_),
    .A2(_02106_),
    .B1(_02107_),
    .Y(_02108_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_136 ();
 sky130_fd_sc_hd__a21oi_1 _22806_ (.A1(_12404_[0]),
    .A2(_01892_),
    .B1(net3762),
    .Y(_02110_));
 sky130_fd_sc_hd__o21ai_0 _22807_ (.A1(_01892_),
    .A2(_02051_),
    .B1(_02110_),
    .Y(_02111_));
 sky130_fd_sc_hd__o311ai_1 _22808_ (.A1(_12420_[0]),
    .A2(net3766),
    .A3(net3769),
    .B1(net3759),
    .C1(_02111_),
    .Y(_02112_));
 sky130_fd_sc_hd__nand4_1 _22809_ (.A(_01900_),
    .B(_02101_),
    .C(_02108_),
    .D(_02112_),
    .Y(_02113_));
 sky130_fd_sc_hd__o311ai_0 _22810_ (.A1(_01900_),
    .A2(_02088_),
    .A3(_02096_),
    .B1(_02113_),
    .C1(_02033_),
    .Y(_02114_));
 sky130_fd_sc_hd__nor2_1 _22811_ (.A(_12396_[0]),
    .B(net3764),
    .Y(_02115_));
 sky130_fd_sc_hd__nor3_1 _22812_ (.A(net3772),
    .B(_02102_),
    .C(_02115_),
    .Y(_02116_));
 sky130_fd_sc_hd__a21oi_1 _22813_ (.A1(_12396_[0]),
    .A2(net3764),
    .B1(_01941_),
    .Y(_02117_));
 sky130_fd_sc_hd__o21ai_2 _22814_ (.A1(_01974_),
    .A2(_02065_),
    .B1(_01892_),
    .Y(_02118_));
 sky130_fd_sc_hd__o211ai_1 _22815_ (.A1(_01892_),
    .A2(_02117_),
    .B1(_02118_),
    .C1(net3752),
    .Y(_02119_));
 sky130_fd_sc_hd__o31ai_1 _22816_ (.A1(net3752),
    .A2(_02097_),
    .A3(_02116_),
    .B1(_02119_),
    .Y(_02120_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_135 ();
 sky130_fd_sc_hd__nand2_1 _22818_ (.A(net3777),
    .B(net3647),
    .Y(_02122_));
 sky130_fd_sc_hd__o21ai_0 _22819_ (.A1(_01974_),
    .A2(_02062_),
    .B1(net3774),
    .Y(_02123_));
 sky130_fd_sc_hd__a21oi_1 _22820_ (.A1(_02122_),
    .A2(_02123_),
    .B1(net3754),
    .Y(_02124_));
 sky130_fd_sc_hd__a21oi_1 _22821_ (.A1(net3762),
    .A2(_02012_),
    .B1(_01941_),
    .Y(_02125_));
 sky130_fd_sc_hd__nor3_2 _22822_ (.A(net3771),
    .B(net3758),
    .C(_02125_),
    .Y(_02126_));
 sky130_fd_sc_hd__nor2_1 _22823_ (.A(net3649),
    .B(_01950_),
    .Y(_02127_));
 sky130_fd_sc_hd__nand2_4 _22824_ (.A(_12410_[0]),
    .B(net3768),
    .Y(_02128_));
 sky130_fd_sc_hd__and3_4 _22825_ (.A(_02127_),
    .B(_02075_),
    .C(_02128_),
    .X(_02129_));
 sky130_fd_sc_hd__nor2_4 _22826_ (.A(_02005_),
    .B(_02033_),
    .Y(_02130_));
 sky130_fd_sc_hd__o41ai_1 _22827_ (.A1(_01910_),
    .A2(_02124_),
    .A3(_02126_),
    .A4(_02129_),
    .B1(_02130_),
    .Y(_02131_));
 sky130_fd_sc_hd__a21o_1 _22828_ (.A1(_01910_),
    .A2(_02120_),
    .B1(_02131_),
    .X(_02132_));
 sky130_fd_sc_hd__o211a_4 _22829_ (.A1(_02007_),
    .A2(_02080_),
    .B1(_02114_),
    .C1(_02132_),
    .X(_00137_));
 sky130_fd_sc_hd__nand2_2 _22830_ (.A(_12406_[0]),
    .B(_01921_),
    .Y(_02133_));
 sky130_fd_sc_hd__nand2_1 _22831_ (.A(net3771),
    .B(_02133_),
    .Y(_02134_));
 sky130_fd_sc_hd__o221ai_1 _22832_ (.A1(_12401_[0]),
    .A2(net3771),
    .B1(_02102_),
    .B2(_02134_),
    .C1(net3756),
    .Y(_02135_));
 sky130_fd_sc_hd__nor2_1 _22833_ (.A(net3650),
    .B(_01921_),
    .Y(_02136_));
 sky130_fd_sc_hd__nor3_1 _22834_ (.A(_01892_),
    .B(_02136_),
    .C(_01975_),
    .Y(_02137_));
 sky130_fd_sc_hd__nor2_1 _22835_ (.A(_12410_[0]),
    .B(net3764),
    .Y(_02138_));
 sky130_fd_sc_hd__nor3_1 _22836_ (.A(net3776),
    .B(_01978_),
    .C(net3577),
    .Y(_02139_));
 sky130_fd_sc_hd__nor3_2 _22837_ (.A(net3760),
    .B(_02137_),
    .C(_02139_),
    .Y(_02140_));
 sky130_fd_sc_hd__a21oi_1 _22838_ (.A1(net3759),
    .A2(_02135_),
    .B1(_02140_),
    .Y(_02141_));
 sky130_fd_sc_hd__nand2_1 _22839_ (.A(net3648),
    .B(_02133_),
    .Y(_02142_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_134 ();
 sky130_fd_sc_hd__o21ai_0 _22841_ (.A1(_01974_),
    .A2(_02065_),
    .B1(net3776),
    .Y(_02144_));
 sky130_fd_sc_hd__o21ai_1 _22842_ (.A1(_01974_),
    .A2(_02142_),
    .B1(_02144_),
    .Y(_02145_));
 sky130_fd_sc_hd__nand2_4 _22843_ (.A(_01910_),
    .B(_01968_),
    .Y(_02146_));
 sky130_fd_sc_hd__nand2_2 _22844_ (.A(net3650),
    .B(_01921_),
    .Y(_02147_));
 sky130_fd_sc_hd__nand2_4 _22845_ (.A(_12406_[0]),
    .B(net3762),
    .Y(_02148_));
 sky130_fd_sc_hd__a21oi_1 _22846_ (.A1(_12410_[0]),
    .A2(net3766),
    .B1(net3771),
    .Y(_02149_));
 sky130_fd_sc_hd__a32oi_1 _22847_ (.A1(net3771),
    .A2(_02147_),
    .A3(_02148_),
    .B1(_02149_),
    .B2(_02098_),
    .Y(_02150_));
 sky130_fd_sc_hd__o21ai_0 _22848_ (.A1(_02146_),
    .A2(_02150_),
    .B1(_02130_),
    .Y(_02151_));
 sky130_fd_sc_hd__a31oi_1 _22849_ (.A1(net3759),
    .A2(_02135_),
    .A3(_02145_),
    .B1(_02151_),
    .Y(_02152_));
 sky130_fd_sc_hd__o21ai_0 _22850_ (.A1(_01910_),
    .A2(_02141_),
    .B1(_02152_),
    .Y(_02153_));
 sky130_fd_sc_hd__nor3_4 _22851_ (.A(net3778),
    .B(_01886_),
    .C(_01892_),
    .Y(_02154_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_133 ();
 sky130_fd_sc_hd__nand2_1 _22853_ (.A(_12417_[0]),
    .B(net3765),
    .Y(_02156_));
 sky130_fd_sc_hd__nor2_4 _22854_ (.A(net3757),
    .B(net3752),
    .Y(_02157_));
 sky130_fd_sc_hd__o311ai_0 _22855_ (.A1(net3765),
    .A2(_02018_),
    .A3(_02154_),
    .B1(_02156_),
    .C1(_02157_),
    .Y(_02158_));
 sky130_fd_sc_hd__nor2_1 _22856_ (.A(_12420_[0]),
    .B(net3762),
    .Y(_02159_));
 sky130_fd_sc_hd__nand2_4 _22857_ (.A(_01954_),
    .B(_01950_),
    .Y(_02160_));
 sky130_fd_sc_hd__a311o_1 _22858_ (.A1(net3762),
    .A2(_02054_),
    .A3(_01987_),
    .B1(_02159_),
    .C1(_02160_),
    .X(_02161_));
 sky130_fd_sc_hd__nor2_4 _22859_ (.A(net3779),
    .B(net3762),
    .Y(_02162_));
 sky130_fd_sc_hd__o21a_1 _22860_ (.A1(_02162_),
    .A2(_02019_),
    .B1(_12397_[0]),
    .X(_02163_));
 sky130_fd_sc_hd__o22ai_1 _22861_ (.A1(net3601),
    .A2(_02098_),
    .B1(_01987_),
    .B2(_02072_),
    .Y(_02164_));
 sky130_fd_sc_hd__nor2_2 _22862_ (.A(_01974_),
    .B(_02067_),
    .Y(_02165_));
 sky130_fd_sc_hd__nand2b_2 _22863_ (.A_N(_12404_[0]),
    .B(net3764),
    .Y(_02166_));
 sky130_fd_sc_hd__nand3_2 _22864_ (.A(net3771),
    .B(_02025_),
    .C(_02166_),
    .Y(_02167_));
 sky130_fd_sc_hd__o211ai_1 _22865_ (.A1(net3773),
    .A2(_02165_),
    .B1(_02167_),
    .C1(net3756),
    .Y(_02168_));
 sky130_fd_sc_hd__o311ai_0 _22866_ (.A1(net3757),
    .A2(_02163_),
    .A3(_02164_),
    .B1(_02168_),
    .C1(net3752),
    .Y(_02169_));
 sky130_fd_sc_hd__nand4_1 _22867_ (.A(_02005_),
    .B(_02158_),
    .C(_02161_),
    .D(_02169_),
    .Y(_02170_));
 sky130_fd_sc_hd__nor2_1 _22868_ (.A(_12401_[0]),
    .B(net3771),
    .Y(_02171_));
 sky130_fd_sc_hd__o21ai_2 _22869_ (.A1(_02171_),
    .A2(_02154_),
    .B1(net3762),
    .Y(_02172_));
 sky130_fd_sc_hd__nand2_2 _22870_ (.A(_01990_),
    .B(_02172_),
    .Y(_02173_));
 sky130_fd_sc_hd__nand2_2 _22871_ (.A(net3768),
    .B(_01968_),
    .Y(_02174_));
 sky130_fd_sc_hd__and2_4 _22872_ (.A(_12410_[0]),
    .B(_01892_),
    .X(_02175_));
 sky130_fd_sc_hd__and2_0 _22873_ (.A(_12401_[0]),
    .B(net3771),
    .X(_02176_));
 sky130_fd_sc_hd__nor2_1 _22874_ (.A(_02175_),
    .B(_02176_),
    .Y(_02177_));
 sky130_fd_sc_hd__nand2_2 _22875_ (.A(net3762),
    .B(_01968_),
    .Y(_02178_));
 sky130_fd_sc_hd__nor2_2 _22876_ (.A(net3777),
    .B(net3776),
    .Y(_02179_));
 sky130_fd_sc_hd__nor2_2 _22877_ (.A(net3779),
    .B(_02179_),
    .Y(_02180_));
 sky130_fd_sc_hd__o221a_1 _22878_ (.A1(_02174_),
    .A2(_02177_),
    .B1(_02178_),
    .B2(_02180_),
    .C1(net3756),
    .X(_02181_));
 sky130_fd_sc_hd__nand2_4 _22879_ (.A(_01910_),
    .B(_01950_),
    .Y(_02182_));
 sky130_fd_sc_hd__nand2_2 _22880_ (.A(_01882_),
    .B(net3649),
    .Y(_02183_));
 sky130_fd_sc_hd__o32a_1 _22881_ (.A1(_02040_),
    .A2(_02136_),
    .A3(_02183_),
    .B1(_02034_),
    .B2(_12410_[0]),
    .X(_02184_));
 sky130_fd_sc_hd__nand3_1 _22882_ (.A(_12397_[0]),
    .B(net3775),
    .C(net3767),
    .Y(_02185_));
 sky130_fd_sc_hd__o211ai_1 _22883_ (.A1(net3777),
    .A2(_02034_),
    .B1(_02107_),
    .C1(_02185_),
    .Y(_02186_));
 sky130_fd_sc_hd__o21ai_0 _22884_ (.A1(_12398_[0]),
    .A2(net3765),
    .B1(_01892_),
    .Y(_02187_));
 sky130_fd_sc_hd__nor2_1 _22885_ (.A(_02162_),
    .B(_02187_),
    .Y(_02188_));
 sky130_fd_sc_hd__o22ai_1 _22886_ (.A1(_02182_),
    .A2(_02184_),
    .B1(_02186_),
    .B2(_02188_),
    .Y(_02189_));
 sky130_fd_sc_hd__a21oi_1 _22887_ (.A1(_02173_),
    .A2(_02181_),
    .B1(_02189_),
    .Y(_02190_));
 sky130_fd_sc_hd__o21ai_0 _22888_ (.A1(_02005_),
    .A2(_02190_),
    .B1(net3645),
    .Y(_02191_));
 sky130_fd_sc_hd__nor2_1 _22889_ (.A(_12404_[0]),
    .B(net3764),
    .Y(_02192_));
 sky130_fd_sc_hd__o21ai_2 _22890_ (.A1(net3779),
    .A2(net3777),
    .B1(net3764),
    .Y(_02193_));
 sky130_fd_sc_hd__nand3b_1 _22891_ (.A_N(_02192_),
    .B(net3648),
    .C(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__nor2_1 _22892_ (.A(net3766),
    .B(_01935_),
    .Y(_02195_));
 sky130_fd_sc_hd__a21oi_1 _22893_ (.A1(net3766),
    .A2(_02051_),
    .B1(_02195_),
    .Y(_02196_));
 sky130_fd_sc_hd__nand2_1 _22894_ (.A(net3773),
    .B(_02196_),
    .Y(_02197_));
 sky130_fd_sc_hd__nand2_1 _22895_ (.A(_01892_),
    .B(_01962_),
    .Y(_02198_));
 sky130_fd_sc_hd__nand2_1 _22896_ (.A(_12415_[0]),
    .B(net3762),
    .Y(_02199_));
 sky130_fd_sc_hd__o21ai_0 _22897_ (.A1(net3762),
    .A2(_02198_),
    .B1(_02199_),
    .Y(_02200_));
 sky130_fd_sc_hd__a221oi_1 _22898_ (.A1(_12401_[0]),
    .A2(_01945_),
    .B1(_02165_),
    .B2(net3773),
    .C1(net3756),
    .Y(_02201_));
 sky130_fd_sc_hd__a211oi_1 _22899_ (.A1(net3756),
    .A2(_02200_),
    .B1(_02201_),
    .C1(net3752),
    .Y(_02202_));
 sky130_fd_sc_hd__a31oi_1 _22900_ (.A1(_02107_),
    .A2(_02194_),
    .A3(_02197_),
    .B1(_02202_),
    .Y(_02203_));
 sky130_fd_sc_hd__nand2_1 _22901_ (.A(_12424_[0]),
    .B(net3768),
    .Y(_02204_));
 sky130_fd_sc_hd__o21ai_0 _22902_ (.A1(net3768),
    .A2(_02180_),
    .B1(_02204_),
    .Y(_02205_));
 sky130_fd_sc_hd__nand2_4 _22903_ (.A(_02005_),
    .B(net3645),
    .Y(_02206_));
 sky130_fd_sc_hd__a21oi_1 _22904_ (.A1(_02100_),
    .A2(_02205_),
    .B1(_02206_),
    .Y(_02207_));
 sky130_fd_sc_hd__a32oi_1 _22905_ (.A1(_02153_),
    .A2(_02170_),
    .A3(_02191_),
    .B1(_02203_),
    .B2(_02207_),
    .Y(_00138_));
 sky130_fd_sc_hd__nor3b_1 _22906_ (.A(_01978_),
    .B(net3776),
    .C_N(_02017_),
    .Y(_02208_));
 sky130_fd_sc_hd__a31oi_1 _22907_ (.A1(net3776),
    .A2(_02020_),
    .A3(_02037_),
    .B1(_02208_),
    .Y(_02209_));
 sky130_fd_sc_hd__nor2_1 _22908_ (.A(_12396_[0]),
    .B(_01921_),
    .Y(_02210_));
 sky130_fd_sc_hd__nand3_1 _22909_ (.A(net3648),
    .B(_02147_),
    .C(_02075_),
    .Y(_02211_));
 sky130_fd_sc_hd__o311ai_0 _22910_ (.A1(net3648),
    .A2(_02192_),
    .A3(_02210_),
    .B1(_02211_),
    .C1(net3753),
    .Y(_02212_));
 sky130_fd_sc_hd__o21ai_0 _22911_ (.A1(net3753),
    .A2(_02209_),
    .B1(_02212_),
    .Y(_02213_));
 sky130_fd_sc_hd__o21ai_0 _22912_ (.A1(net3779),
    .A2(_02043_),
    .B1(_02052_),
    .Y(_02214_));
 sky130_fd_sc_hd__a21oi_1 _22913_ (.A1(_12397_[0]),
    .A2(_02043_),
    .B1(_02214_),
    .Y(_02215_));
 sky130_fd_sc_hd__nor2_1 _22914_ (.A(net3650),
    .B(net3753),
    .Y(_02216_));
 sky130_fd_sc_hd__o22ai_1 _22915_ (.A1(_01991_),
    .A2(_02084_),
    .B1(_02183_),
    .B2(_02216_),
    .Y(_02217_));
 sky130_fd_sc_hd__a22oi_1 _22916_ (.A1(net3650),
    .A2(_02127_),
    .B1(_02217_),
    .B2(net3767),
    .Y(_02218_));
 sky130_fd_sc_hd__o211ai_1 _22917_ (.A1(net3767),
    .A2(_02215_),
    .B1(_02218_),
    .C1(net3755),
    .Y(_02219_));
 sky130_fd_sc_hd__o21ai_2 _22918_ (.A1(net3756),
    .A2(_02213_),
    .B1(_02219_),
    .Y(_02220_));
 sky130_fd_sc_hd__nor3_1 _22919_ (.A(net3775),
    .B(_02090_),
    .C(_01975_),
    .Y(_02221_));
 sky130_fd_sc_hd__a31oi_1 _22920_ (.A1(net3775),
    .A2(_02020_),
    .A3(_02098_),
    .B1(_02221_),
    .Y(_02222_));
 sky130_fd_sc_hd__o41ai_1 _22921_ (.A1(_01923_),
    .A2(net3753),
    .A3(_02044_),
    .A4(_02179_),
    .B1(net3756),
    .Y(_02223_));
 sky130_fd_sc_hd__a21oi_1 _22922_ (.A1(net3753),
    .A2(_02222_),
    .B1(_02223_),
    .Y(_02224_));
 sky130_fd_sc_hd__nand2_1 _22923_ (.A(net3765),
    .B(_01991_),
    .Y(_02225_));
 sky130_fd_sc_hd__a21oi_2 _22924_ (.A1(_02014_),
    .A2(_02225_),
    .B1(net3779),
    .Y(_02226_));
 sky130_fd_sc_hd__o21ai_2 _22925_ (.A1(_12397_[0]),
    .A2(_01958_),
    .B1(_02157_),
    .Y(_02227_));
 sky130_fd_sc_hd__a211oi_4 _22926_ (.A1(_12404_[0]),
    .A2(_01923_),
    .B1(_02226_),
    .C1(_02227_),
    .Y(_02228_));
 sky130_fd_sc_hd__nor2_1 _22927_ (.A(_01921_),
    .B(_02054_),
    .Y(_02229_));
 sky130_fd_sc_hd__a311oi_1 _22928_ (.A1(_12404_[0]),
    .A2(net3648),
    .A3(_01921_),
    .B1(_02186_),
    .C1(_02229_),
    .Y(_02230_));
 sky130_fd_sc_hd__nor3_2 _22929_ (.A(_02224_),
    .B(_02228_),
    .C(_02230_),
    .Y(_02231_));
 sky130_fd_sc_hd__nor3_1 _22930_ (.A(net3774),
    .B(net3767),
    .C(_01910_),
    .Y(_02232_));
 sky130_fd_sc_hd__a21oi_1 _22931_ (.A1(net3774),
    .A2(_02057_),
    .B1(_02232_),
    .Y(_02233_));
 sky130_fd_sc_hd__o21ai_2 _22932_ (.A1(_01910_),
    .A2(_02017_),
    .B1(_01961_),
    .Y(_02234_));
 sky130_fd_sc_hd__o31ai_1 _22933_ (.A1(_12404_[0]),
    .A2(_01958_),
    .A3(_01910_),
    .B1(net3754),
    .Y(_02235_));
 sky130_fd_sc_hd__a21oi_1 _22934_ (.A1(net3774),
    .A2(_02234_),
    .B1(_02235_),
    .Y(_02236_));
 sky130_fd_sc_hd__o21ai_2 _22935_ (.A1(_12397_[0]),
    .A2(_02233_),
    .B1(_02236_),
    .Y(_02237_));
 sky130_fd_sc_hd__a221oi_1 _22936_ (.A1(_01921_),
    .A2(net3602),
    .B1(_02009_),
    .B2(_12406_[0]),
    .C1(_02182_),
    .Y(_02238_));
 sky130_fd_sc_hd__nor3_2 _22937_ (.A(net3775),
    .B(_02090_),
    .C(_02065_),
    .Y(_02239_));
 sky130_fd_sc_hd__nor2_2 _22938_ (.A(_12397_[0]),
    .B(net3762),
    .Y(_02240_));
 sky130_fd_sc_hd__a211oi_1 _22939_ (.A1(net3762),
    .A2(_01935_),
    .B1(_02240_),
    .C1(_01892_),
    .Y(_02241_));
 sky130_fd_sc_hd__nor3_1 _22940_ (.A(_02160_),
    .B(_02239_),
    .C(_02241_),
    .Y(_02242_));
 sky130_fd_sc_hd__nor4_1 _22941_ (.A(_02005_),
    .B(_01905_),
    .C(_02238_),
    .D(_02242_),
    .Y(_02243_));
 sky130_fd_sc_hd__nand3_2 _22942_ (.A(net3771),
    .B(_02020_),
    .C(_02148_),
    .Y(_02244_));
 sky130_fd_sc_hd__o21ai_0 _22943_ (.A1(_02072_),
    .A2(net3577),
    .B1(_01892_),
    .Y(_02245_));
 sky130_fd_sc_hd__a21oi_1 _22944_ (.A1(_02244_),
    .A2(_02245_),
    .B1(_02146_),
    .Y(_02246_));
 sky130_fd_sc_hd__a21oi_1 _22945_ (.A1(net3776),
    .A2(_02017_),
    .B1(net3777),
    .Y(_02247_));
 sky130_fd_sc_hd__o22ai_1 _22946_ (.A1(net3779),
    .A2(_01958_),
    .B1(_02034_),
    .B2(_12396_[0]),
    .Y(_02248_));
 sky130_fd_sc_hd__nor3_1 _22947_ (.A(_02182_),
    .B(_02247_),
    .C(_02248_),
    .Y(_02249_));
 sky130_fd_sc_hd__o41ai_1 _22948_ (.A1(net3602),
    .A2(_01910_),
    .A3(_02175_),
    .A4(_02174_),
    .B1(_02130_),
    .Y(_02250_));
 sky130_fd_sc_hd__o21ai_0 _22949_ (.A1(_12406_[0]),
    .A2(net3771),
    .B1(net3762),
    .Y(_02251_));
 sky130_fd_sc_hd__a21oi_1 _22950_ (.A1(net3771),
    .A2(_01935_),
    .B1(_02251_),
    .Y(_02252_));
 sky130_fd_sc_hd__nor3b_1 _22951_ (.A(_02252_),
    .B(_02160_),
    .C_N(_02111_),
    .Y(_02253_));
 sky130_fd_sc_hd__nor4_1 _22952_ (.A(_02246_),
    .B(_02249_),
    .C(_02250_),
    .D(_02253_),
    .Y(_02254_));
 sky130_fd_sc_hd__a21oi_1 _22953_ (.A1(_02237_),
    .A2(_02243_),
    .B1(_02254_),
    .Y(_02255_));
 sky130_fd_sc_hd__o221ai_4 _22954_ (.A1(_02206_),
    .A2(_02220_),
    .B1(_02231_),
    .B2(_02007_),
    .C1(_02255_),
    .Y(_00139_));
 sky130_fd_sc_hd__nor3_1 _22955_ (.A(net3771),
    .B(_02102_),
    .C(_02067_),
    .Y(_02256_));
 sky130_fd_sc_hd__a21oi_1 _22956_ (.A1(_01892_),
    .A2(_02148_),
    .B1(_01941_),
    .Y(_02257_));
 sky130_fd_sc_hd__o32ai_1 _22957_ (.A1(net3602),
    .A2(_02182_),
    .A3(_02256_),
    .B1(_02257_),
    .B2(_02146_),
    .Y(_02258_));
 sky130_fd_sc_hd__o22ai_1 _22958_ (.A1(net3779),
    .A2(_02055_),
    .B1(_02105_),
    .B2(net3761),
    .Y(_02259_));
 sky130_fd_sc_hd__nand2_1 _22959_ (.A(net3763),
    .B(_02259_),
    .Y(_02260_));
 sky130_fd_sc_hd__a21oi_1 _22960_ (.A1(net3777),
    .A2(_02043_),
    .B1(net3779),
    .Y(_02261_));
 sky130_fd_sc_hd__o21ai_0 _22961_ (.A1(_01991_),
    .A2(_02261_),
    .B1(net3767),
    .Y(_02262_));
 sky130_fd_sc_hd__nor3_2 _22962_ (.A(net3650),
    .B(net3767),
    .C(_01968_),
    .Y(_02263_));
 sky130_fd_sc_hd__o21ai_0 _22963_ (.A1(_02127_),
    .A2(_02263_),
    .B1(net3779),
    .Y(_02264_));
 sky130_fd_sc_hd__a31oi_2 _22964_ (.A1(_02260_),
    .A2(_02262_),
    .A3(_02264_),
    .B1(_01910_),
    .Y(_02265_));
 sky130_fd_sc_hd__or3_1 _22965_ (.A(_02007_),
    .B(_02258_),
    .C(_02265_),
    .X(_02266_));
 sky130_fd_sc_hd__o21ai_1 _22966_ (.A1(_02018_),
    .A2(_02176_),
    .B1(net3766),
    .Y(_02267_));
 sky130_fd_sc_hd__a211oi_1 _22967_ (.A1(_02002_),
    .A2(_02267_),
    .B1(_02126_),
    .C1(_01954_),
    .Y(_02268_));
 sky130_fd_sc_hd__o221ai_1 _22968_ (.A1(_12410_[0]),
    .A2(_01958_),
    .B1(_02065_),
    .B2(_01892_),
    .C1(net3761),
    .Y(_02269_));
 sky130_fd_sc_hd__o21ai_0 _22969_ (.A1(_02162_),
    .A2(_02035_),
    .B1(_01892_),
    .Y(_02270_));
 sky130_fd_sc_hd__o21ai_0 _22970_ (.A1(_01978_),
    .A2(_02067_),
    .B1(net3774),
    .Y(_02271_));
 sky130_fd_sc_hd__nand3_1 _22971_ (.A(_01968_),
    .B(_02270_),
    .C(_02271_),
    .Y(_02272_));
 sky130_fd_sc_hd__a21oi_1 _22972_ (.A1(_02269_),
    .A2(_02272_),
    .B1(_01910_),
    .Y(_02273_));
 sky130_fd_sc_hd__o21ai_1 _22973_ (.A1(_02268_),
    .A2(_02273_),
    .B1(_02130_),
    .Y(_02274_));
 sky130_fd_sc_hd__nor2_4 _22974_ (.A(_02005_),
    .B(_01905_),
    .Y(_02275_));
 sky130_fd_sc_hd__nand2_1 _22975_ (.A(net3762),
    .B(_01962_),
    .Y(_02276_));
 sky130_fd_sc_hd__o21ai_0 _22976_ (.A1(_02072_),
    .A2(_02067_),
    .B1(_01892_),
    .Y(_02277_));
 sky130_fd_sc_hd__o2111ai_1 _22977_ (.A1(_12398_[0]),
    .A2(_01928_),
    .B1(net3757),
    .C1(_02276_),
    .D1(_02277_),
    .Y(_02278_));
 sky130_fd_sc_hd__nand2_1 _22978_ (.A(_12408_[0]),
    .B(net3765),
    .Y(_02279_));
 sky130_fd_sc_hd__o211ai_1 _22979_ (.A1(net3765),
    .A2(_01986_),
    .B1(_02279_),
    .C1(net3769),
    .Y(_02280_));
 sky130_fd_sc_hd__nand3_4 _22980_ (.A(net3758),
    .B(_02278_),
    .C(_02280_),
    .Y(_02281_));
 sky130_fd_sc_hd__nand2b_1 _22981_ (.A_N(_12406_[0]),
    .B(net3763),
    .Y(_02282_));
 sky130_fd_sc_hd__nor2b_1 _22982_ (.A(_02057_),
    .B_N(_02282_),
    .Y(_02283_));
 sky130_fd_sc_hd__a21oi_1 _22983_ (.A1(_01923_),
    .A2(_01910_),
    .B1(net3647),
    .Y(_02284_));
 sky130_fd_sc_hd__a31oi_1 _22984_ (.A1(net3762),
    .A2(_01991_),
    .A3(net3755),
    .B1(_02091_),
    .Y(_02285_));
 sky130_fd_sc_hd__o221ai_1 _22985_ (.A1(net3774),
    .A2(_02283_),
    .B1(_02284_),
    .B2(_01882_),
    .C1(_02285_),
    .Y(_02286_));
 sky130_fd_sc_hd__nand2_1 _22986_ (.A(net3754),
    .B(_02286_),
    .Y(_02287_));
 sky130_fd_sc_hd__nand3_2 _22987_ (.A(_02275_),
    .B(_02281_),
    .C(_02287_),
    .Y(_02288_));
 sky130_fd_sc_hd__o21ai_1 _22988_ (.A1(_12406_[0]),
    .A2(_01892_),
    .B1(_02093_),
    .Y(_02289_));
 sky130_fd_sc_hd__a21boi_0 _22989_ (.A1(_12410_[0]),
    .A2(net3771),
    .B1_N(_01986_),
    .Y(_02290_));
 sky130_fd_sc_hd__o22ai_1 _22990_ (.A1(_02154_),
    .A2(_02251_),
    .B1(_02290_),
    .B2(net3762),
    .Y(_02291_));
 sky130_fd_sc_hd__o21ai_0 _22991_ (.A1(_02182_),
    .A2(_02291_),
    .B1(_01906_),
    .Y(_02292_));
 sky130_fd_sc_hd__nor2_1 _22992_ (.A(_12401_[0]),
    .B(net3762),
    .Y(_02293_));
 sky130_fd_sc_hd__nand2_1 _22993_ (.A(_12396_[0]),
    .B(net3762),
    .Y(_02294_));
 sky130_fd_sc_hd__nand2_1 _22994_ (.A(net3771),
    .B(_02294_),
    .Y(_02295_));
 sky130_fd_sc_hd__o32ai_1 _22995_ (.A1(net3771),
    .A2(_02035_),
    .A3(_02293_),
    .B1(_02295_),
    .B2(_02091_),
    .Y(_02296_));
 sky130_fd_sc_hd__nor3_1 _22996_ (.A(_02019_),
    .B(_02154_),
    .C(_02178_),
    .Y(_02297_));
 sky130_fd_sc_hd__o21ai_0 _22997_ (.A1(_02174_),
    .A2(_02177_),
    .B1(_01954_),
    .Y(_02298_));
 sky130_fd_sc_hd__a211oi_1 _22998_ (.A1(net3759),
    .A2(_02296_),
    .B1(_02297_),
    .C1(_02298_),
    .Y(_02299_));
 sky130_fd_sc_hd__a211o_1 _22999_ (.A1(_02107_),
    .A2(_02289_),
    .B1(_02292_),
    .C1(_02299_),
    .X(_02300_));
 sky130_fd_sc_hd__nand4_1 _23000_ (.A(_02266_),
    .B(_02274_),
    .C(_02288_),
    .D(_02300_),
    .Y(_00140_));
 sky130_fd_sc_hd__a221oi_1 _23001_ (.A1(_12401_[0]),
    .A2(net3762),
    .B1(net3646),
    .B2(_12406_[0]),
    .C1(_01963_),
    .Y(_02301_));
 sky130_fd_sc_hd__nor2_4 _23002_ (.A(_02033_),
    .B(_01968_),
    .Y(_02302_));
 sky130_fd_sc_hd__o21ai_0 _23003_ (.A1(_02162_),
    .A2(_02090_),
    .B1(_01892_),
    .Y(_02303_));
 sky130_fd_sc_hd__a31oi_1 _23004_ (.A1(_01981_),
    .A2(_02302_),
    .A3(_02303_),
    .B1(net3757),
    .Y(_02304_));
 sky130_fd_sc_hd__nor2_1 _23005_ (.A(_01892_),
    .B(net3764),
    .Y(_02305_));
 sky130_fd_sc_hd__a22oi_1 _23006_ (.A1(_12404_[0]),
    .A2(_01945_),
    .B1(_02305_),
    .B2(net3777),
    .Y(_02306_));
 sky130_fd_sc_hd__nor2_2 _23007_ (.A(_01921_),
    .B(net3753),
    .Y(_02307_));
 sky130_fd_sc_hd__o21ai_0 _23008_ (.A1(_02305_),
    .A2(_02307_),
    .B1(net3779),
    .Y(_02308_));
 sky130_fd_sc_hd__a211oi_1 _23009_ (.A1(_02034_),
    .A2(_01968_),
    .B1(_02307_),
    .C1(net3779),
    .Y(_02309_));
 sky130_fd_sc_hd__nor2_1 _23010_ (.A(_01882_),
    .B(_02174_),
    .Y(_02310_));
 sky130_fd_sc_hd__o21ai_0 _23011_ (.A1(_02309_),
    .A2(_02310_),
    .B1(net3650),
    .Y(_02311_));
 sky130_fd_sc_hd__o2111ai_1 _23012_ (.A1(net3760),
    .A2(_02306_),
    .B1(_02308_),
    .C1(_02311_),
    .D1(_02033_),
    .Y(_02312_));
 sky130_fd_sc_hd__o311a_1 _23013_ (.A1(net3645),
    .A2(net3758),
    .A3(_02301_),
    .B1(_02304_),
    .C1(_02312_),
    .X(_02313_));
 sky130_fd_sc_hd__nand2_2 _23014_ (.A(_02033_),
    .B(net3758),
    .Y(_02314_));
 sky130_fd_sc_hd__o21ai_0 _23015_ (.A1(_12396_[0]),
    .A2(net3767),
    .B1(_02128_),
    .Y(_02315_));
 sky130_fd_sc_hd__nor2_1 _23016_ (.A(_12397_[0]),
    .B(_02034_),
    .Y(_02316_));
 sky130_fd_sc_hd__a21oi_2 _23017_ (.A1(net3649),
    .A2(_02315_),
    .B1(_02316_),
    .Y(_02317_));
 sky130_fd_sc_hd__a21oi_1 _23018_ (.A1(net3772),
    .A2(_02076_),
    .B1(_01943_),
    .Y(_02318_));
 sky130_fd_sc_hd__nand2_1 _23019_ (.A(_12398_[0]),
    .B(net3765),
    .Y(_02319_));
 sky130_fd_sc_hd__a21oi_1 _23020_ (.A1(_02319_),
    .A2(_02066_),
    .B1(net3772),
    .Y(_02320_));
 sky130_fd_sc_hd__o21ai_0 _23021_ (.A1(_01882_),
    .A2(_01928_),
    .B1(_02033_),
    .Y(_02321_));
 sky130_fd_sc_hd__o221ai_1 _23022_ (.A1(_02033_),
    .A2(_02318_),
    .B1(_02320_),
    .B2(_02321_),
    .C1(net3752),
    .Y(_02322_));
 sky130_fd_sc_hd__o211ai_1 _23023_ (.A1(net3777),
    .A2(_01932_),
    .B1(_02244_),
    .C1(_02302_),
    .Y(_02323_));
 sky130_fd_sc_hd__o2111ai_1 _23024_ (.A1(_02314_),
    .A2(_02317_),
    .B1(net3757),
    .C1(_02322_),
    .D1(_02323_),
    .Y(_02324_));
 sky130_fd_sc_hd__nand2_1 _23025_ (.A(_02005_),
    .B(_02324_),
    .Y(_02325_));
 sky130_fd_sc_hd__a21oi_1 _23026_ (.A1(net3650),
    .A2(_01928_),
    .B1(_02091_),
    .Y(_02326_));
 sky130_fd_sc_hd__o221ai_1 _23027_ (.A1(_12401_[0]),
    .A2(_01958_),
    .B1(_02034_),
    .B2(_02051_),
    .C1(net3755),
    .Y(_02327_));
 sky130_fd_sc_hd__o221ai_1 _23028_ (.A1(net3755),
    .A2(_02326_),
    .B1(_02327_),
    .B2(_02073_),
    .C1(net3761),
    .Y(_02328_));
 sky130_fd_sc_hd__a21oi_1 _23029_ (.A1(_02128_),
    .A2(_02166_),
    .B1(net3775),
    .Y(_02329_));
 sky130_fd_sc_hd__a21oi_1 _23030_ (.A1(_02305_),
    .A2(_02051_),
    .B1(_02329_),
    .Y(_02330_));
 sky130_fd_sc_hd__nor3_1 _23031_ (.A(net3771),
    .B(_01943_),
    .C(_01975_),
    .Y(_02331_));
 sky130_fd_sc_hd__a311oi_1 _23032_ (.A1(net3771),
    .A2(_02017_),
    .A3(_02075_),
    .B1(_02331_),
    .C1(_02146_),
    .Y(_02332_));
 sky130_fd_sc_hd__a21oi_1 _23033_ (.A1(_02100_),
    .A2(_02330_),
    .B1(_02332_),
    .Y(_02333_));
 sky130_fd_sc_hd__a311oi_1 _23034_ (.A1(net3774),
    .A2(_02020_),
    .A3(_02075_),
    .B1(_02329_),
    .C1(_01910_),
    .Y(_02334_));
 sky130_fd_sc_hd__o21ai_0 _23035_ (.A1(_12410_[0]),
    .A2(net3774),
    .B1(net3763),
    .Y(_02335_));
 sky130_fd_sc_hd__a31o_1 _23036_ (.A1(_01910_),
    .A2(_02003_),
    .A3(_02335_),
    .B1(net3761),
    .X(_02336_));
 sky130_fd_sc_hd__a32oi_1 _23037_ (.A1(_02162_),
    .A2(_02081_),
    .A3(_02103_),
    .B1(_01935_),
    .B2(_01923_),
    .Y(_02337_));
 sky130_fd_sc_hd__nor2_1 _23038_ (.A(net3779),
    .B(net3649),
    .Y(_02338_));
 sky130_fd_sc_hd__a221oi_1 _23039_ (.A1(_12404_[0]),
    .A2(net3763),
    .B1(_02040_),
    .B2(_02338_),
    .C1(_01910_),
    .Y(_02339_));
 sky130_fd_sc_hd__a21oi_1 _23040_ (.A1(_01910_),
    .A2(_02337_),
    .B1(_02339_),
    .Y(_02340_));
 sky130_fd_sc_hd__o22ai_1 _23041_ (.A1(_02334_),
    .A2(_02336_),
    .B1(_02340_),
    .B2(_01968_),
    .Y(_02341_));
 sky130_fd_sc_hd__a32oi_1 _23042_ (.A1(_02130_),
    .A2(_02328_),
    .A3(_02333_),
    .B1(_02341_),
    .B2(_02275_),
    .Y(_02342_));
 sky130_fd_sc_hd__o21ai_0 _23043_ (.A1(_02313_),
    .A2(_02325_),
    .B1(_02342_),
    .Y(_00141_));
 sky130_fd_sc_hd__o21a_1 _23044_ (.A1(_12397_[0]),
    .A2(_01892_),
    .B1(_02198_),
    .X(_02343_));
 sky130_fd_sc_hd__o211ai_1 _23045_ (.A1(net3762),
    .A2(_02343_),
    .B1(_02199_),
    .C1(net3752),
    .Y(_02344_));
 sky130_fd_sc_hd__o21ai_1 _23046_ (.A1(_01941_),
    .A2(_01943_),
    .B1(_01892_),
    .Y(_02345_));
 sky130_fd_sc_hd__o311ai_0 _23047_ (.A1(_01892_),
    .A2(_02102_),
    .A3(_02240_),
    .B1(_02345_),
    .C1(net3759),
    .Y(_02346_));
 sky130_fd_sc_hd__nand3_1 _23048_ (.A(net3769),
    .B(_02344_),
    .C(_02346_),
    .Y(_02347_));
 sky130_fd_sc_hd__nand2_1 _23049_ (.A(_12404_[0]),
    .B(_01968_),
    .Y(_02348_));
 sky130_fd_sc_hd__nand2_1 _23050_ (.A(_12397_[0]),
    .B(net3761),
    .Y(_02349_));
 sky130_fd_sc_hd__nor3_1 _23051_ (.A(net3649),
    .B(_01968_),
    .C(_01935_),
    .Y(_02350_));
 sky130_fd_sc_hd__a31oi_1 _23052_ (.A1(net3649),
    .A2(_02348_),
    .A3(_02349_),
    .B1(_02350_),
    .Y(_02351_));
 sky130_fd_sc_hd__o21ai_0 _23053_ (.A1(net3777),
    .A2(net3754),
    .B1(net3779),
    .Y(_02352_));
 sky130_fd_sc_hd__o21ai_0 _23054_ (.A1(net3650),
    .A2(_02043_),
    .B1(_02352_),
    .Y(_02353_));
 sky130_fd_sc_hd__o21ai_0 _23055_ (.A1(_01991_),
    .A2(_02353_),
    .B1(net3763),
    .Y(_02354_));
 sky130_fd_sc_hd__o211ai_1 _23056_ (.A1(net3763),
    .A2(_02351_),
    .B1(_02354_),
    .C1(net3755),
    .Y(_02355_));
 sky130_fd_sc_hd__nand3_1 _23057_ (.A(net3650),
    .B(net3768),
    .C(_01968_),
    .Y(_02356_));
 sky130_fd_sc_hd__a21oi_1 _23058_ (.A1(_02020_),
    .A2(_02148_),
    .B1(_01968_),
    .Y(_02357_));
 sky130_fd_sc_hd__nand2_1 _23059_ (.A(net3771),
    .B(_02178_),
    .Y(_02358_));
 sky130_fd_sc_hd__o21ai_0 _23060_ (.A1(_01882_),
    .A2(net3759),
    .B1(net3648),
    .Y(_02359_));
 sky130_fd_sc_hd__o22ai_1 _23061_ (.A1(_02357_),
    .A2(_02358_),
    .B1(_02359_),
    .B2(_02263_),
    .Y(_02360_));
 sky130_fd_sc_hd__a41o_1 _23062_ (.A1(_01905_),
    .A2(net3756),
    .A3(_02356_),
    .A4(_02360_),
    .B1(_02005_),
    .X(_02361_));
 sky130_fd_sc_hd__or2_0 _23063_ (.A(_02316_),
    .B(_02239_),
    .X(_02362_));
 sky130_fd_sc_hd__nand2_1 _23064_ (.A(_12404_[0]),
    .B(net3765),
    .Y(_02363_));
 sky130_fd_sc_hd__a21oi_1 _23065_ (.A1(_02282_),
    .A2(_02363_),
    .B1(net3774),
    .Y(_02364_));
 sky130_fd_sc_hd__o311ai_2 _23066_ (.A1(_01910_),
    .A2(_02063_),
    .A3(_02364_),
    .B1(net3754),
    .C1(_02033_),
    .Y(_02365_));
 sky130_fd_sc_hd__a21oi_2 _23067_ (.A1(_01910_),
    .A2(_02362_),
    .B1(_02365_),
    .Y(_02366_));
 sky130_fd_sc_hd__a21oi_1 _23068_ (.A1(_12406_[0]),
    .A2(_01892_),
    .B1(net3762),
    .Y(_02367_));
 sky130_fd_sc_hd__a221oi_1 _23069_ (.A1(_12414_[0]),
    .A2(net3762),
    .B1(_01987_),
    .B2(_02367_),
    .C1(net3757),
    .Y(_02368_));
 sky130_fd_sc_hd__a211oi_2 _23070_ (.A1(net3757),
    .A2(_02172_),
    .B1(_02314_),
    .C1(_02368_),
    .Y(_02369_));
 sky130_fd_sc_hd__nand2_1 _23071_ (.A(_01991_),
    .B(_02307_),
    .Y(_02370_));
 sky130_fd_sc_hd__o21a_1 _23072_ (.A1(_01950_),
    .A2(_02138_),
    .B1(net3775),
    .X(_02371_));
 sky130_fd_sc_hd__o21ai_0 _23073_ (.A1(_02216_),
    .A2(_02371_),
    .B1(_01882_),
    .Y(_02372_));
 sky130_fd_sc_hd__nand3_1 _23074_ (.A(net3779),
    .B(net3777),
    .C(net3775),
    .Y(_02373_));
 sky130_fd_sc_hd__a21oi_1 _23075_ (.A1(_02147_),
    .A2(_02373_),
    .B1(_12410_[0]),
    .Y(_02374_));
 sky130_fd_sc_hd__o31ai_1 _23076_ (.A1(_02179_),
    .A2(_02229_),
    .A3(_02374_),
    .B1(net3753),
    .Y(_02375_));
 sky130_fd_sc_hd__a311oi_2 _23077_ (.A1(_02370_),
    .A2(_02372_),
    .A3(_02375_),
    .B1(net3756),
    .C1(_02033_),
    .Y(_02376_));
 sky130_fd_sc_hd__nor4_1 _23078_ (.A(_02361_),
    .B(_02366_),
    .C(_02369_),
    .D(_02376_),
    .Y(_02377_));
 sky130_fd_sc_hd__a31o_1 _23079_ (.A1(_01892_),
    .A2(_02193_),
    .A3(_02133_),
    .B1(_01910_),
    .X(_02378_));
 sky130_fd_sc_hd__a31oi_1 _23080_ (.A1(net3771),
    .A2(_01961_),
    .A3(_02128_),
    .B1(_02378_),
    .Y(_02379_));
 sky130_fd_sc_hd__a21oi_1 _23081_ (.A1(net3779),
    .A2(net3771),
    .B1(_02193_),
    .Y(_02380_));
 sky130_fd_sc_hd__nor3_1 _23082_ (.A(_12413_[0]),
    .B(_12422_[0]),
    .C(net3762),
    .Y(_02381_));
 sky130_fd_sc_hd__nor3_1 _23083_ (.A(net3757),
    .B(_02380_),
    .C(_02381_),
    .Y(_02382_));
 sky130_fd_sc_hd__nor3_1 _23084_ (.A(net3752),
    .B(_02379_),
    .C(_02382_),
    .Y(_02383_));
 sky130_fd_sc_hd__nand2_1 _23085_ (.A(net3777),
    .B(net3766),
    .Y(_02384_));
 sky130_fd_sc_hd__nor3_1 _23086_ (.A(net3773),
    .B(_02195_),
    .C(_02240_),
    .Y(_02385_));
 sky130_fd_sc_hd__a31oi_1 _23087_ (.A1(net3773),
    .A2(_02384_),
    .A3(_02148_),
    .B1(_02385_),
    .Y(_02386_));
 sky130_fd_sc_hd__nor2_1 _23088_ (.A(_02030_),
    .B(_02386_),
    .Y(_02387_));
 sky130_fd_sc_hd__o21ai_0 _23089_ (.A1(_12396_[0]),
    .A2(net3762),
    .B1(_02148_),
    .Y(_02388_));
 sky130_fd_sc_hd__a221oi_1 _23090_ (.A1(_12398_[0]),
    .A2(_01945_),
    .B1(_02388_),
    .B2(net3773),
    .C1(_02146_),
    .Y(_02389_));
 sky130_fd_sc_hd__nor4_1 _23091_ (.A(_02007_),
    .B(_02383_),
    .C(_02387_),
    .D(_02389_),
    .Y(_02390_));
 sky130_fd_sc_hd__a311o_1 _23092_ (.A1(_01906_),
    .A2(_02347_),
    .A3(_02355_),
    .B1(_02377_),
    .C1(_02390_),
    .X(_00142_));
 sky130_fd_sc_hd__nor2_1 _23093_ (.A(_12408_[0]),
    .B(net3765),
    .Y(_02391_));
 sky130_fd_sc_hd__a31oi_1 _23094_ (.A1(_12398_[0]),
    .A2(_01892_),
    .A3(net3765),
    .B1(_02391_),
    .Y(_02392_));
 sky130_fd_sc_hd__a21oi_1 _23095_ (.A1(_02157_),
    .A2(_02392_),
    .B1(_02206_),
    .Y(_02393_));
 sky130_fd_sc_hd__nor2_1 _23096_ (.A(_12401_[0]),
    .B(_01892_),
    .Y(_02394_));
 sky130_fd_sc_hd__o21ai_0 _23097_ (.A1(_02019_),
    .A2(_02394_),
    .B1(net3762),
    .Y(_02395_));
 sky130_fd_sc_hd__o21ai_0 _23098_ (.A1(net3602),
    .A2(_02025_),
    .B1(_02395_),
    .Y(_02396_));
 sky130_fd_sc_hd__o31ai_1 _23099_ (.A1(_01892_),
    .A2(_02162_),
    .A3(_01974_),
    .B1(_02118_),
    .Y(_02397_));
 sky130_fd_sc_hd__a21oi_1 _23100_ (.A1(_12406_[0]),
    .A2(net3771),
    .B1(_02018_),
    .Y(_02398_));
 sky130_fd_sc_hd__nor2_1 _23101_ (.A(net3762),
    .B(_02398_),
    .Y(_02399_));
 sky130_fd_sc_hd__a211oi_2 _23102_ (.A1(_12422_[0]),
    .A2(net3762),
    .B1(_02160_),
    .C1(_02399_),
    .Y(_02400_));
 sky130_fd_sc_hd__a221oi_1 _23103_ (.A1(_02107_),
    .A2(_02396_),
    .B1(_02397_),
    .B2(_02100_),
    .C1(_02400_),
    .Y(_02401_));
 sky130_fd_sc_hd__o21ai_0 _23104_ (.A1(net3647),
    .A2(_02307_),
    .B1(net3650),
    .Y(_02402_));
 sky130_fd_sc_hd__nand3_1 _23105_ (.A(net3777),
    .B(_01923_),
    .C(_01968_),
    .Y(_02403_));
 sky130_fd_sc_hd__a21oi_1 _23106_ (.A1(_02402_),
    .A2(_02403_),
    .B1(net3779),
    .Y(_02404_));
 sky130_fd_sc_hd__nand3_1 _23107_ (.A(_02043_),
    .B(_02185_),
    .C(_02275_),
    .Y(_02405_));
 sky130_fd_sc_hd__a211oi_1 _23108_ (.A1(net3777),
    .A2(_01936_),
    .B1(net3760),
    .C1(_02033_),
    .Y(_02406_));
 sky130_fd_sc_hd__o221ai_1 _23109_ (.A1(_12410_[0]),
    .A2(_02034_),
    .B1(_02009_),
    .B2(_12397_[0]),
    .C1(_02406_),
    .Y(_02407_));
 sky130_fd_sc_hd__nand2_1 _23110_ (.A(net3776),
    .B(_02128_),
    .Y(_02408_));
 sky130_fd_sc_hd__o221ai_1 _23111_ (.A1(_02102_),
    .A2(_02142_),
    .B1(_02408_),
    .B2(_02072_),
    .C1(_02302_),
    .Y(_02409_));
 sky130_fd_sc_hd__and3_1 _23112_ (.A(net3756),
    .B(_02407_),
    .C(_02409_),
    .X(_02410_));
 sky130_fd_sc_hd__o22ai_2 _23113_ (.A1(_02404_),
    .A2(_02405_),
    .B1(_02410_),
    .B2(_02005_),
    .Y(_02411_));
 sky130_fd_sc_hd__a21oi_1 _23114_ (.A1(_01892_),
    .A2(_02072_),
    .B1(_02065_),
    .Y(_02412_));
 sky130_fd_sc_hd__nand2_1 _23115_ (.A(_12396_[0]),
    .B(_01923_),
    .Y(_02413_));
 sky130_fd_sc_hd__o211ai_1 _23116_ (.A1(net3779),
    .A2(_02412_),
    .B1(_02406_),
    .C1(_02413_),
    .Y(_02414_));
 sky130_fd_sc_hd__o21ai_0 _23117_ (.A1(_02035_),
    .A2(net3577),
    .B1(net3771),
    .Y(_02415_));
 sky130_fd_sc_hd__o211ai_1 _23118_ (.A1(_12406_[0]),
    .A2(_01932_),
    .B1(_02302_),
    .C1(_02415_),
    .Y(_02416_));
 sky130_fd_sc_hd__a21oi_1 _23119_ (.A1(_01932_),
    .A2(_02225_),
    .B1(net3779),
    .Y(_02417_));
 sky130_fd_sc_hd__nand2_1 _23120_ (.A(_01882_),
    .B(_02065_),
    .Y(_02418_));
 sky130_fd_sc_hd__o21ai_0 _23121_ (.A1(_01936_),
    .A2(_02072_),
    .B1(net3779),
    .Y(_02419_));
 sky130_fd_sc_hd__a211oi_1 _23122_ (.A1(net3777),
    .A2(_01923_),
    .B1(net3760),
    .C1(_02040_),
    .Y(_02420_));
 sky130_fd_sc_hd__a31oi_1 _23123_ (.A1(_01950_),
    .A2(_02418_),
    .A3(_02419_),
    .B1(_02420_),
    .Y(_02421_));
 sky130_fd_sc_hd__o21ai_0 _23124_ (.A1(_02417_),
    .A2(_02421_),
    .B1(net3645),
    .Y(_02422_));
 sky130_fd_sc_hd__nand4_1 _23125_ (.A(net3769),
    .B(_02414_),
    .C(_02416_),
    .D(_02422_),
    .Y(_02423_));
 sky130_fd_sc_hd__a21oi_1 _23126_ (.A1(_01882_),
    .A2(_02000_),
    .B1(net3764),
    .Y(_02424_));
 sky130_fd_sc_hd__nor3_1 _23127_ (.A(_02146_),
    .B(_02252_),
    .C(_02424_),
    .Y(_02425_));
 sky130_fd_sc_hd__a211o_1 _23128_ (.A1(_12404_[0]),
    .A2(net3762),
    .B1(_02062_),
    .C1(net3771),
    .X(_02426_));
 sky130_fd_sc_hd__and3_4 _23129_ (.A(_02157_),
    .B(_02069_),
    .C(_02426_),
    .X(_02427_));
 sky130_fd_sc_hd__nor2_1 _23130_ (.A(_12396_[0]),
    .B(_01892_),
    .Y(_02428_));
 sky130_fd_sc_hd__nor3_1 _23131_ (.A(net3771),
    .B(_01941_),
    .C(_02102_),
    .Y(_02429_));
 sky130_fd_sc_hd__o21ai_0 _23132_ (.A1(_02428_),
    .A2(_02429_),
    .B1(net3759),
    .Y(_02430_));
 sky130_fd_sc_hd__o311ai_0 _23133_ (.A1(net3759),
    .A2(_02293_),
    .A3(_02380_),
    .B1(_02430_),
    .C1(net3757),
    .Y(_02431_));
 sky130_fd_sc_hd__nor4b_1 _23134_ (.A(_02007_),
    .B(_02425_),
    .C(_02427_),
    .D_N(_02431_),
    .Y(_02432_));
 sky130_fd_sc_hd__a221o_1 _23135_ (.A1(_02393_),
    .A2(_02401_),
    .B1(_02411_),
    .B2(_02423_),
    .C1(_02432_),
    .X(_00143_));
 sky130_fd_sc_hd__xor3_1 _23136_ (.A(\sa02_sr[7] ),
    .B(\sa02_sr[0] ),
    .C(\sa20_sub[1] ),
    .X(_02433_));
 sky130_fd_sc_hd__xnor3_1 _23137_ (.A(_11612_),
    .B(_11613_),
    .C(_02433_),
    .X(_02434_));
 sky130_fd_sc_hd__nand2_1 _23138_ (.A(net4230),
    .B(\text_in_r[33] ),
    .Y(_02435_));
 sky130_fd_sc_hd__o21a_4 _23139_ (.A1(net4230),
    .A2(_02434_),
    .B1(_02435_),
    .X(_02436_));
 sky130_fd_sc_hd__xor2_4 _23140_ (.A(\u0.w[2][1] ),
    .B(_02436_),
    .X(_02437_));
 sky130_fd_sc_hd__clkinvlp_4 _23141_ (.A(_02437_),
    .Y(_02438_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_131 ();
 sky130_fd_sc_hd__xnor3_1 _23144_ (.A(\sa12_sr[0] ),
    .B(net4201),
    .C(net4182),
    .X(_02440_));
 sky130_fd_sc_hd__xor2_1 _23145_ (.A(_07074_),
    .B(_02440_),
    .X(_02441_));
 sky130_fd_sc_hd__mux2i_2 _23146_ (.A0(\text_in_r[32] ),
    .A1(_02441_),
    .S(net4111),
    .Y(_02442_));
 sky130_fd_sc_hd__xor2_4 _23147_ (.A(\u0.w[2][0] ),
    .B(_02442_),
    .X(_02443_));
 sky130_fd_sc_hd__clkinv_16 _23148_ (.A(net3748),
    .Y(_02444_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_130 ();
 sky130_fd_sc_hd__xor2_1 _23150_ (.A(net4185),
    .B(net4224),
    .X(_02445_));
 sky130_fd_sc_hd__xnor2_1 _23151_ (.A(_07094_),
    .B(_02445_),
    .Y(_02446_));
 sky130_fd_sc_hd__mux2i_4 _23152_ (.A0(\text_in_r[34] ),
    .A1(_02446_),
    .S(net4114),
    .Y(_02447_));
 sky130_fd_sc_hd__xnor2_4 _23153_ (.A(\u0.w[2][2] ),
    .B(_02447_),
    .Y(_02448_));
 sky130_fd_sc_hd__clkinv_16 _23154_ (.A(_02448_),
    .Y(_02449_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_124 ();
 sky130_fd_sc_hd__xnor3_1 _23161_ (.A(net4196),
    .B(_07084_),
    .C(_09455_),
    .X(_02453_));
 sky130_fd_sc_hd__nor2_2 _23162_ (.A(net4231),
    .B(_02453_),
    .Y(_02454_));
 sky130_fd_sc_hd__a21oi_4 _23163_ (.A1(net4231),
    .A2(\text_in_r[39] ),
    .B1(_02454_),
    .Y(_02455_));
 sky130_fd_sc_hd__xnor2_4 _23164_ (.A(\u0.w[2][7] ),
    .B(_02455_),
    .Y(_02456_));
 sky130_fd_sc_hd__xnor2_1 _23165_ (.A(\sa31_sub[5] ),
    .B(\sa02_sr[6] ),
    .Y(_02457_));
 sky130_fd_sc_hd__xnor2_1 _23166_ (.A(_07116_),
    .B(_02457_),
    .Y(_02458_));
 sky130_fd_sc_hd__nand2_1 _23167_ (.A(net4231),
    .B(\text_in_r[38] ),
    .Y(_02459_));
 sky130_fd_sc_hd__o21ai_2 _23168_ (.A1(net4231),
    .A2(_02458_),
    .B1(_02459_),
    .Y(_02460_));
 sky130_fd_sc_hd__xor2_4 _23169_ (.A(\u0.w[2][6] ),
    .B(_02460_),
    .X(_02461_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_123 ();
 sky130_fd_sc_hd__xnor2_1 _23171_ (.A(\sa02_sr[4] ),
    .B(net4197),
    .Y(_02463_));
 sky130_fd_sc_hd__xnor2_1 _23172_ (.A(_11635_),
    .B(_02463_),
    .Y(_02464_));
 sky130_fd_sc_hd__nor2_2 _23173_ (.A(net4230),
    .B(_02464_),
    .Y(_02465_));
 sky130_fd_sc_hd__a21oi_4 _23174_ (.A1(net398),
    .A2(\text_in_r[37] ),
    .B1(_02465_),
    .Y(_02466_));
 sky130_fd_sc_hd__xnor2_4 _23175_ (.A(\u0.w[2][5] ),
    .B(_02466_),
    .Y(_02467_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_121 ();
 sky130_fd_sc_hd__xor3_1 _23178_ (.A(_07135_),
    .B(_11665_),
    .C(_11666_),
    .X(_02470_));
 sky130_fd_sc_hd__mux2i_4 _23179_ (.A0(\text_in_r[36] ),
    .A1(_02470_),
    .S(net4114),
    .Y(_02471_));
 sky130_fd_sc_hd__xor2_4 _23180_ (.A(\u0.w[2][4] ),
    .B(_02471_),
    .X(_02472_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_119 ();
 sky130_fd_sc_hd__xnor3_1 _23183_ (.A(_07148_),
    .B(_11646_),
    .C(_11647_),
    .X(_02475_));
 sky130_fd_sc_hd__nand2b_1 _23184_ (.A_N(\text_in_r[35] ),
    .B(net4230),
    .Y(_02476_));
 sky130_fd_sc_hd__o211a_4 _23185_ (.A1(net398),
    .A2(_02475_),
    .B1(_02476_),
    .C1(\u0.w[2][3] ),
    .X(_02477_));
 sky130_fd_sc_hd__and2_4 _23186_ (.A(net4230),
    .B(\text_in_r[35] ),
    .X(_02478_));
 sky130_fd_sc_hd__a211oi_4 _23187_ (.A1(net4115),
    .A2(_02475_),
    .B1(_02478_),
    .C1(\u0.w[2][3] ),
    .Y(_02479_));
 sky130_fd_sc_hd__or2_4 _23188_ (.A(_02477_),
    .B(_02479_),
    .X(_02480_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_116 ();
 sky130_fd_sc_hd__nand2_2 _23192_ (.A(net3751),
    .B(net3749),
    .Y(_02484_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_115 ();
 sky130_fd_sc_hd__nand2_8 _23194_ (.A(_02444_),
    .B(net3746),
    .Y(_02486_));
 sky130_fd_sc_hd__nand2_2 _23195_ (.A(_02484_),
    .B(_02486_),
    .Y(_02487_));
 sky130_fd_sc_hd__xnor2_1 _23196_ (.A(_02480_),
    .B(_02487_),
    .Y(_02488_));
 sky130_fd_sc_hd__nor2_4 _23197_ (.A(_02477_),
    .B(_02479_),
    .Y(_02489_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_113 ();
 sky130_fd_sc_hd__a21oi_4 _23200_ (.A1(net3643),
    .A2(_02444_),
    .B1(net3734),
    .Y(_02492_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_111 ();
 sky130_fd_sc_hd__nor2_1 _23203_ (.A(_12428_[0]),
    .B(_02480_),
    .Y(_02495_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_108 ();
 sky130_fd_sc_hd__nand2_8 _23207_ (.A(_12429_[0]),
    .B(_02480_),
    .Y(_02499_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_107 ();
 sky130_fd_sc_hd__o211ai_1 _23209_ (.A1(_12436_[0]),
    .A2(_02480_),
    .B1(_02499_),
    .C1(net3745),
    .Y(_02501_));
 sky130_fd_sc_hd__o311ai_0 _23210_ (.A1(net3745),
    .A2(_02492_),
    .A3(_02495_),
    .B1(net3740),
    .C1(_02501_),
    .Y(_02502_));
 sky130_fd_sc_hd__o21ai_0 _23211_ (.A1(net3740),
    .A2(_02488_),
    .B1(_02502_),
    .Y(_02503_));
 sky130_fd_sc_hd__xnor2_4 _23212_ (.A(\u0.w[2][4] ),
    .B(_02471_),
    .Y(_02504_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_105 ();
 sky130_fd_sc_hd__nand2_8 _23215_ (.A(net3751),
    .B(net3737),
    .Y(_02507_));
 sky130_fd_sc_hd__nor2_2 _23216_ (.A(_12429_[0]),
    .B(net3746),
    .Y(_02508_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 ();
 sky130_fd_sc_hd__nor2_1 _23219_ (.A(net3643),
    .B(net3746),
    .Y(_02511_));
 sky130_fd_sc_hd__nor2_1 _23220_ (.A(_02511_),
    .B(_02499_),
    .Y(_02512_));
 sky130_fd_sc_hd__a21oi_2 _23221_ (.A1(_02507_),
    .A2(_02508_),
    .B1(_02512_),
    .Y(_02513_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 ();
 sky130_fd_sc_hd__nand2_8 _23223_ (.A(_02449_),
    .B(net3736),
    .Y(_02515_));
 sky130_fd_sc_hd__xnor2_2 _23224_ (.A(net3745),
    .B(net3734),
    .Y(_02516_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 ();
 sky130_fd_sc_hd__nand3_2 _23227_ (.A(_12429_[0]),
    .B(net3745),
    .C(net3734),
    .Y(_02519_));
 sky130_fd_sc_hd__o221ai_1 _23228_ (.A1(_12436_[0]),
    .A2(_02515_),
    .B1(_02516_),
    .B2(_12428_[0]),
    .C1(_02519_),
    .Y(_02520_));
 sky130_fd_sc_hd__nor2_1 _23229_ (.A(net3729),
    .B(_02520_),
    .Y(_02521_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_99 ();
 sky130_fd_sc_hd__a211oi_1 _23231_ (.A1(net3729),
    .A2(_02513_),
    .B1(_02521_),
    .C1(_02467_),
    .Y(_02523_));
 sky130_fd_sc_hd__a21oi_1 _23232_ (.A1(_02467_),
    .A2(_02503_),
    .B1(_02523_),
    .Y(_02524_));
 sky130_fd_sc_hd__xor2_4 _23233_ (.A(\u0.w[2][5] ),
    .B(_02466_),
    .X(_02525_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_93 ();
 sky130_fd_sc_hd__nand2_8 _23240_ (.A(net3746),
    .B(_02489_),
    .Y(_02532_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_90 ();
 sky130_fd_sc_hd__nand2_2 _23244_ (.A(net3749),
    .B(_02449_),
    .Y(_02536_));
 sky130_fd_sc_hd__nor2_4 _23245_ (.A(net3643),
    .B(net3737),
    .Y(_02537_));
 sky130_fd_sc_hd__o22ai_1 _23246_ (.A1(_12433_[0]),
    .A2(_02532_),
    .B1(_02536_),
    .B2(_02537_),
    .Y(_02538_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_88 ();
 sky130_fd_sc_hd__nor2_1 _23249_ (.A(net3751),
    .B(net3732),
    .Y(_02541_));
 sky130_fd_sc_hd__nor2_1 _23250_ (.A(_12442_[0]),
    .B(_02480_),
    .Y(_02542_));
 sky130_fd_sc_hd__nand2_8 _23251_ (.A(_02444_),
    .B(net3737),
    .Y(_02543_));
 sky130_fd_sc_hd__o311ai_0 _23252_ (.A1(net3746),
    .A2(_02541_),
    .A3(net3576),
    .B1(_02519_),
    .C1(_02543_),
    .Y(_02544_));
 sky130_fd_sc_hd__nor2_1 _23253_ (.A(net3742),
    .B(_02544_),
    .Y(_02545_));
 sky130_fd_sc_hd__a21oi_1 _23254_ (.A1(net3742),
    .A2(_02538_),
    .B1(_02545_),
    .Y(_02546_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_85 ();
 sky130_fd_sc_hd__nand2_2 _23258_ (.A(net3746),
    .B(_02480_),
    .Y(_02550_));
 sky130_fd_sc_hd__nor2_4 _23259_ (.A(net3746),
    .B(net3732),
    .Y(_02551_));
 sky130_fd_sc_hd__nor3_1 _23260_ (.A(net3749),
    .B(_02449_),
    .C(_02480_),
    .Y(_02552_));
 sky130_fd_sc_hd__o21ai_0 _23261_ (.A1(_02551_),
    .A2(_02552_),
    .B1(net3644),
    .Y(_02553_));
 sky130_fd_sc_hd__nand3_4 _23262_ (.A(net3749),
    .B(_02449_),
    .C(net3732),
    .Y(_02554_));
 sky130_fd_sc_hd__o2111ai_1 _23263_ (.A1(_12430_[0]),
    .A2(_02550_),
    .B1(_02553_),
    .C1(_02554_),
    .D1(net3742),
    .Y(_02555_));
 sky130_fd_sc_hd__nor2_4 _23264_ (.A(net3643),
    .B(net3732),
    .Y(_02556_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_83 ();
 sky130_fd_sc_hd__nand2_4 _23267_ (.A(_12442_[0]),
    .B(net3732),
    .Y(_02559_));
 sky130_fd_sc_hd__nand2_4 _23268_ (.A(net3643),
    .B(_02480_),
    .Y(_02560_));
 sky130_fd_sc_hd__nand3_1 _23269_ (.A(net3746),
    .B(_02559_),
    .C(_02560_),
    .Y(_02561_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_81 ();
 sky130_fd_sc_hd__o211ai_1 _23272_ (.A1(_02556_),
    .A2(_02536_),
    .B1(_02561_),
    .C1(_02504_),
    .Y(_02564_));
 sky130_fd_sc_hd__xor2_4 _23273_ (.A(\u0.w[2][7] ),
    .B(_02455_),
    .X(_02565_));
 sky130_fd_sc_hd__nand2_8 _23274_ (.A(_02565_),
    .B(net3744),
    .Y(_02566_));
 sky130_fd_sc_hd__a31oi_1 _23275_ (.A1(net3640),
    .A2(_02555_),
    .A3(_02564_),
    .B1(_02566_),
    .Y(_02567_));
 sky130_fd_sc_hd__o21ai_2 _23276_ (.A1(net3640),
    .A2(_02546_),
    .B1(_02567_),
    .Y(_02568_));
 sky130_fd_sc_hd__inv_2 _23277_ (.A(_02461_),
    .Y(_02569_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_80 ();
 sky130_fd_sc_hd__o21ai_0 _23279_ (.A1(net3751),
    .A2(_02449_),
    .B1(net3736),
    .Y(_02571_));
 sky130_fd_sc_hd__nor2_4 _23280_ (.A(_12430_[0]),
    .B(_12433_[0]),
    .Y(_02572_));
 sky130_fd_sc_hd__nor2_4 _23281_ (.A(_02449_),
    .B(net3736),
    .Y(_02573_));
 sky130_fd_sc_hd__a221oi_1 _23282_ (.A1(net3749),
    .A2(_02571_),
    .B1(_02572_),
    .B2(_02551_),
    .C1(_02573_),
    .Y(_02574_));
 sky130_fd_sc_hd__o21ai_0 _23283_ (.A1(_12428_[0]),
    .A2(_02532_),
    .B1(_02472_),
    .Y(_02575_));
 sky130_fd_sc_hd__a221o_1 _23284_ (.A1(_12449_[0]),
    .A2(net3732),
    .B1(_02551_),
    .B2(_12429_[0]),
    .C1(net3742),
    .X(_02576_));
 sky130_fd_sc_hd__o211ai_1 _23285_ (.A1(_02574_),
    .A2(_02575_),
    .B1(net3640),
    .C1(_02576_),
    .Y(_02577_));
 sky130_fd_sc_hd__a21oi_1 _23286_ (.A1(_02569_),
    .A2(_02577_),
    .B1(_02565_),
    .Y(_02578_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_79 ();
 sky130_fd_sc_hd__nor2_2 _23288_ (.A(_12430_[0]),
    .B(net3732),
    .Y(_02580_));
 sky130_fd_sc_hd__nor3_4 _23289_ (.A(net3750),
    .B(_02444_),
    .C(net3738),
    .Y(_02581_));
 sky130_fd_sc_hd__nor3_2 _23290_ (.A(_02449_),
    .B(_02580_),
    .C(_02581_),
    .Y(_02582_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_78 ();
 sky130_fd_sc_hd__nor2_4 _23292_ (.A(net3746),
    .B(net3737),
    .Y(_02584_));
 sky130_fd_sc_hd__nand2_2 _23293_ (.A(_12438_[0]),
    .B(_02584_),
    .Y(_02585_));
 sky130_fd_sc_hd__nand2_1 _23294_ (.A(net3741),
    .B(_02585_),
    .Y(_02586_));
 sky130_fd_sc_hd__nand3_2 _23295_ (.A(net3643),
    .B(net3749),
    .C(net3738),
    .Y(_02587_));
 sky130_fd_sc_hd__o211ai_1 _23296_ (.A1(_12430_[0]),
    .A2(net3739),
    .B1(_02587_),
    .C1(net3745),
    .Y(_02588_));
 sky130_fd_sc_hd__o211ai_1 _23297_ (.A1(_12436_[0]),
    .A2(_02515_),
    .B1(_02588_),
    .C1(net3729),
    .Y(_02589_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_77 ();
 sky130_fd_sc_hd__nor2_1 _23299_ (.A(_02565_),
    .B(_02525_),
    .Y(_02591_));
 sky130_fd_sc_hd__o211a_4 _23300_ (.A1(_02582_),
    .A2(_02586_),
    .B1(_02589_),
    .C1(_02591_),
    .X(_02592_));
 sky130_fd_sc_hd__nor2_4 _23301_ (.A(net3749),
    .B(net3736),
    .Y(_02593_));
 sky130_fd_sc_hd__nand2b_4 _23302_ (.A_N(_12429_[0]),
    .B(_02480_),
    .Y(_02594_));
 sky130_fd_sc_hd__o211ai_1 _23303_ (.A1(_12436_[0]),
    .A2(_02480_),
    .B1(_02594_),
    .C1(_02449_),
    .Y(_02595_));
 sky130_fd_sc_hd__o311a_1 _23304_ (.A1(_02449_),
    .A2(_02556_),
    .A3(_02593_),
    .B1(_02595_),
    .C1(net3740),
    .X(_02596_));
 sky130_fd_sc_hd__nand2_4 _23305_ (.A(_12430_[0]),
    .B(net3738),
    .Y(_02597_));
 sky130_fd_sc_hd__nand2_4 _23306_ (.A(_12433_[0]),
    .B(net3734),
    .Y(_02598_));
 sky130_fd_sc_hd__and3_4 _23307_ (.A(net3745),
    .B(_02597_),
    .C(_02598_),
    .X(_02599_));
 sky130_fd_sc_hd__a211oi_2 _23308_ (.A1(_12428_[0]),
    .A2(_02551_),
    .B1(_02599_),
    .C1(net3741),
    .Y(_02600_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_76 ();
 sky130_fd_sc_hd__a21oi_1 _23310_ (.A1(net3643),
    .A2(_02444_),
    .B1(net3738),
    .Y(_02602_));
 sky130_fd_sc_hd__o221ai_1 _23311_ (.A1(net3591),
    .A2(net3734),
    .B1(_02602_),
    .B2(_02449_),
    .C1(_02554_),
    .Y(_02603_));
 sky130_fd_sc_hd__o21ai_0 _23312_ (.A1(net3591),
    .A2(_02515_),
    .B1(net3729),
    .Y(_02604_));
 sky130_fd_sc_hd__nor3_2 _23313_ (.A(_12429_[0]),
    .B(_02477_),
    .C(net4070),
    .Y(_02605_));
 sky130_fd_sc_hd__nor2_4 _23314_ (.A(_12438_[0]),
    .B(net3734),
    .Y(_02606_));
 sky130_fd_sc_hd__o21a_1 _23315_ (.A1(_02605_),
    .A2(_02606_),
    .B1(net3745),
    .X(_02607_));
 sky130_fd_sc_hd__o221ai_1 _23316_ (.A1(net3729),
    .A2(_02603_),
    .B1(_02604_),
    .B2(_02607_),
    .C1(net3640),
    .Y(_02608_));
 sky130_fd_sc_hd__o31a_1 _23317_ (.A1(net3640),
    .A2(_02596_),
    .A3(_02600_),
    .B1(_02608_),
    .X(_02609_));
 sky130_fd_sc_hd__o22ai_1 _23318_ (.A1(_02578_),
    .A2(_02592_),
    .B1(_02609_),
    .B2(_02569_),
    .Y(_02610_));
 sky130_fd_sc_hd__o311ai_1 _23319_ (.A1(_02456_),
    .A2(_02461_),
    .A3(_02524_),
    .B1(_02568_),
    .C1(_02610_),
    .Y(_00144_));
 sky130_fd_sc_hd__nor2_4 _23320_ (.A(_02456_),
    .B(_02461_),
    .Y(_02611_));
 sky130_fd_sc_hd__nand2_8 _23321_ (.A(net3643),
    .B(net3732),
    .Y(_02612_));
 sky130_fd_sc_hd__nor2_1 _23322_ (.A(_02444_),
    .B(_02449_),
    .Y(_02613_));
 sky130_fd_sc_hd__nor2_4 _23323_ (.A(net3749),
    .B(net3746),
    .Y(_02614_));
 sky130_fd_sc_hd__mux2i_1 _23324_ (.A0(_12428_[0]),
    .A1(net3749),
    .S(net3746),
    .Y(_02615_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_75 ();
 sky130_fd_sc_hd__o32ai_1 _23326_ (.A1(_02612_),
    .A2(_02613_),
    .A3(_02614_),
    .B1(_02615_),
    .B2(net3732),
    .Y(_02617_));
 sky130_fd_sc_hd__nand2_1 _23327_ (.A(net3751),
    .B(net3732),
    .Y(_02618_));
 sky130_fd_sc_hd__nor3_4 _23328_ (.A(_12433_[0]),
    .B(_02477_),
    .C(net4070),
    .Y(_02619_));
 sky130_fd_sc_hd__a211oi_1 _23329_ (.A1(_02444_),
    .A2(_02480_),
    .B1(_02619_),
    .C1(_02449_),
    .Y(_02620_));
 sky130_fd_sc_hd__a311oi_1 _23330_ (.A1(_02449_),
    .A2(_02560_),
    .A3(_02618_),
    .B1(_02620_),
    .C1(net3642),
    .Y(_02621_));
 sky130_fd_sc_hd__a21oi_1 _23331_ (.A1(net3642),
    .A2(_02617_),
    .B1(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__nand3_2 _23332_ (.A(net3643),
    .B(_02444_),
    .C(net3746),
    .Y(_02623_));
 sky130_fd_sc_hd__nand2_1 _23333_ (.A(_12436_[0]),
    .B(_02449_),
    .Y(_02624_));
 sky130_fd_sc_hd__nor3_1 _23334_ (.A(_12452_[0]),
    .B(net3642),
    .C(net3737),
    .Y(_02625_));
 sky130_fd_sc_hd__a311o_1 _23335_ (.A1(net3737),
    .A2(_02623_),
    .A3(_02624_),
    .B1(_02625_),
    .C1(_02504_),
    .X(_02626_));
 sky130_fd_sc_hd__o21ai_2 _23336_ (.A1(net3743),
    .A2(_02622_),
    .B1(_02626_),
    .Y(_02627_));
 sky130_fd_sc_hd__nand2_1 _23337_ (.A(_12442_[0]),
    .B(_02584_),
    .Y(_02628_));
 sky130_fd_sc_hd__nor2_1 _23338_ (.A(net3751),
    .B(net3736),
    .Y(_02629_));
 sky130_fd_sc_hd__o21ai_0 _23339_ (.A1(_02492_),
    .A2(_02629_),
    .B1(net3745),
    .Y(_02630_));
 sky130_fd_sc_hd__nand2_1 _23340_ (.A(_02467_),
    .B(net3729),
    .Y(_02631_));
 sky130_fd_sc_hd__a21oi_1 _23341_ (.A1(_02628_),
    .A2(_02630_),
    .B1(_02631_),
    .Y(_02632_));
 sky130_fd_sc_hd__nand2_8 _23342_ (.A(_02456_),
    .B(_02461_),
    .Y(_02633_));
 sky130_fd_sc_hd__nand2_1 _23343_ (.A(_02525_),
    .B(net3729),
    .Y(_02634_));
 sky130_fd_sc_hd__nand2_4 _23344_ (.A(_12429_[0]),
    .B(net3734),
    .Y(_02635_));
 sky130_fd_sc_hd__nand2_4 _23345_ (.A(_12428_[0]),
    .B(_02480_),
    .Y(_02636_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_74 ();
 sky130_fd_sc_hd__a21oi_2 _23347_ (.A1(_02635_),
    .A2(_02636_),
    .B1(_02449_),
    .Y(_02638_));
 sky130_fd_sc_hd__and3_1 _23348_ (.A(_02449_),
    .B(_02598_),
    .C(_02543_),
    .X(_02639_));
 sky130_fd_sc_hd__a211o_1 _23349_ (.A1(net3591),
    .A2(net3738),
    .B1(_02605_),
    .C1(_02449_),
    .X(_02640_));
 sky130_fd_sc_hd__o21ai_0 _23350_ (.A1(net3745),
    .A2(_02602_),
    .B1(_02640_),
    .Y(_02641_));
 sky130_fd_sc_hd__nand2_2 _23351_ (.A(net3642),
    .B(_02472_),
    .Y(_02642_));
 sky130_fd_sc_hd__o32ai_1 _23352_ (.A1(_02634_),
    .A2(_02638_),
    .A3(_02639_),
    .B1(_02641_),
    .B2(_02642_),
    .Y(_02643_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_73 ();
 sky130_fd_sc_hd__nand2_2 _23354_ (.A(_12429_[0]),
    .B(_02449_),
    .Y(_02644_));
 sky130_fd_sc_hd__o22ai_1 _23355_ (.A1(_02489_),
    .A2(_02644_),
    .B1(_02516_),
    .B2(_02444_),
    .Y(_02645_));
 sky130_fd_sc_hd__nand2_8 _23356_ (.A(_02525_),
    .B(net3740),
    .Y(_02646_));
 sky130_fd_sc_hd__a211oi_1 _23357_ (.A1(net3751),
    .A2(_02593_),
    .B1(_02645_),
    .C1(_02646_),
    .Y(_02647_));
 sky130_fd_sc_hd__nor4_1 _23358_ (.A(_02632_),
    .B(_02633_),
    .C(_02643_),
    .D(_02647_),
    .Y(_02648_));
 sky130_fd_sc_hd__a21oi_2 _23359_ (.A1(_02611_),
    .A2(_02627_),
    .B1(_02648_),
    .Y(_02649_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_72 ();
 sky130_fd_sc_hd__or3_4 _23361_ (.A(_12429_[0]),
    .B(_02477_),
    .C(net4070),
    .X(_02651_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_71 ();
 sky130_fd_sc_hd__o21ai_4 _23363_ (.A1(_12433_[0]),
    .A2(net3732),
    .B1(_02651_),
    .Y(_02653_));
 sky130_fd_sc_hd__nor2_1 _23364_ (.A(net3746),
    .B(_02653_),
    .Y(_02654_));
 sky130_fd_sc_hd__nand2_8 _23365_ (.A(net3749),
    .B(net3736),
    .Y(_02655_));
 sky130_fd_sc_hd__nor2_1 _23366_ (.A(net3751),
    .B(_02655_),
    .Y(_02656_));
 sky130_fd_sc_hd__nor3_1 _23367_ (.A(_02449_),
    .B(_02656_),
    .C(net3576),
    .Y(_02657_));
 sky130_fd_sc_hd__o22ai_1 _23368_ (.A1(_12433_[0]),
    .A2(_02515_),
    .B1(_02516_),
    .B2(net3751),
    .Y(_02658_));
 sky130_fd_sc_hd__nand2_1 _23369_ (.A(_02504_),
    .B(_02658_),
    .Y(_02659_));
 sky130_fd_sc_hd__o311ai_2 _23370_ (.A1(_02504_),
    .A2(_02654_),
    .A3(_02657_),
    .B1(_02659_),
    .C1(net3640),
    .Y(_02660_));
 sky130_fd_sc_hd__nor2_2 _23371_ (.A(_02565_),
    .B(_02461_),
    .Y(_02661_));
 sky130_fd_sc_hd__nor2_4 _23372_ (.A(_02525_),
    .B(net3740),
    .Y(_02662_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_70 ();
 sky130_fd_sc_hd__nand2_2 _23374_ (.A(net3749),
    .B(net3732),
    .Y(_02664_));
 sky130_fd_sc_hd__nand3_1 _23375_ (.A(_02449_),
    .B(_02664_),
    .C(_02543_),
    .Y(_02665_));
 sky130_fd_sc_hd__o21ai_0 _23376_ (.A1(_02449_),
    .A2(_02653_),
    .B1(_02665_),
    .Y(_02666_));
 sky130_fd_sc_hd__nand2_1 _23377_ (.A(_02662_),
    .B(_02666_),
    .Y(_02667_));
 sky130_fd_sc_hd__nor2_4 _23378_ (.A(_02525_),
    .B(net3729),
    .Y(_02668_));
 sky130_fd_sc_hd__nor2_4 _23379_ (.A(_02444_),
    .B(_02480_),
    .Y(_02669_));
 sky130_fd_sc_hd__o21ai_0 _23380_ (.A1(net3745),
    .A2(_02669_),
    .B1(net3644),
    .Y(_02670_));
 sky130_fd_sc_hd__o2111ai_1 _23381_ (.A1(net3644),
    .A2(_02655_),
    .B1(_02668_),
    .C1(_02670_),
    .D1(_02532_),
    .Y(_02671_));
 sky130_fd_sc_hd__nand4_1 _23382_ (.A(_02660_),
    .B(_02661_),
    .C(_02667_),
    .D(_02671_),
    .Y(_02672_));
 sky130_fd_sc_hd__nand3_4 _23383_ (.A(net3644),
    .B(_02444_),
    .C(net3738),
    .Y(_02673_));
 sky130_fd_sc_hd__a21oi_1 _23384_ (.A1(_02651_),
    .A2(_02673_),
    .B1(_02449_),
    .Y(_02674_));
 sky130_fd_sc_hd__nor2_1 _23385_ (.A(_02444_),
    .B(_02515_),
    .Y(_02675_));
 sky130_fd_sc_hd__o211ai_1 _23386_ (.A1(_12428_[0]),
    .A2(net3735),
    .B1(_02612_),
    .C1(_02449_),
    .Y(_02676_));
 sky130_fd_sc_hd__nand3_1 _23387_ (.A(net3745),
    .B(_02655_),
    .C(_02598_),
    .Y(_02677_));
 sky130_fd_sc_hd__a31oi_1 _23388_ (.A1(_02668_),
    .A2(_02676_),
    .A3(_02677_),
    .B1(_02566_),
    .Y(_02678_));
 sky130_fd_sc_hd__a21oi_2 _23389_ (.A1(_02655_),
    .A2(_02651_),
    .B1(net3746),
    .Y(_02679_));
 sky130_fd_sc_hd__nand2b_2 _23390_ (.A_N(_12430_[0]),
    .B(_02480_),
    .Y(_02680_));
 sky130_fd_sc_hd__nand2_1 _23391_ (.A(_12428_[0]),
    .B(net3732),
    .Y(_02681_));
 sky130_fd_sc_hd__a21oi_1 _23392_ (.A1(_02680_),
    .A2(_02681_),
    .B1(_02449_),
    .Y(_02682_));
 sky130_fd_sc_hd__nor3_1 _23393_ (.A(net3641),
    .B(_02679_),
    .C(_02682_),
    .Y(_02683_));
 sky130_fd_sc_hd__nand2_4 _23394_ (.A(_12442_[0]),
    .B(net3738),
    .Y(_02684_));
 sky130_fd_sc_hd__nand3_1 _23395_ (.A(net3643),
    .B(_02444_),
    .C(net3732),
    .Y(_02685_));
 sky130_fd_sc_hd__a21oi_1 _23396_ (.A1(_02680_),
    .A2(_02685_),
    .B1(net3746),
    .Y(_02686_));
 sky130_fd_sc_hd__a311oi_1 _23397_ (.A1(net3746),
    .A2(_02651_),
    .A3(_02684_),
    .B1(_02686_),
    .C1(net3642),
    .Y(_02687_));
 sky130_fd_sc_hd__o21ai_1 _23398_ (.A1(_02683_),
    .A2(_02687_),
    .B1(net3731),
    .Y(_02688_));
 sky130_fd_sc_hd__o311ai_0 _23399_ (.A1(_02646_),
    .A2(_02674_),
    .A3(_02675_),
    .B1(_02678_),
    .C1(_02688_),
    .Y(_02689_));
 sky130_fd_sc_hd__and3_4 _23400_ (.A(_02649_),
    .B(_02672_),
    .C(_02689_),
    .X(_00145_));
 sky130_fd_sc_hd__nand2_4 _23401_ (.A(_12430_[0]),
    .B(net3735),
    .Y(_02690_));
 sky130_fd_sc_hd__nand2_1 _23402_ (.A(_02690_),
    .B(_02507_),
    .Y(_02691_));
 sky130_fd_sc_hd__nand2_4 _23403_ (.A(_02444_),
    .B(net3732),
    .Y(_02692_));
 sky130_fd_sc_hd__a21oi_2 _23404_ (.A1(_02692_),
    .A2(_02499_),
    .B1(_02449_),
    .Y(_02693_));
 sky130_fd_sc_hd__a21oi_1 _23405_ (.A1(_02449_),
    .A2(_02691_),
    .B1(_02693_),
    .Y(_02694_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_69 ();
 sky130_fd_sc_hd__nand4_1 _23407_ (.A(net3644),
    .B(_02449_),
    .C(_02664_),
    .D(_02543_),
    .Y(_02696_));
 sky130_fd_sc_hd__o211ai_1 _23408_ (.A1(_12442_[0]),
    .A2(_02532_),
    .B1(_02696_),
    .C1(_02472_),
    .Y(_02697_));
 sky130_fd_sc_hd__o21ai_0 _23409_ (.A1(_02472_),
    .A2(_02694_),
    .B1(_02697_),
    .Y(_02698_));
 sky130_fd_sc_hd__nand2_2 _23410_ (.A(net3643),
    .B(net3746),
    .Y(_02699_));
 sky130_fd_sc_hd__nand2_4 _23411_ (.A(net3643),
    .B(net3749),
    .Y(_02700_));
 sky130_fd_sc_hd__nand2b_1 _23412_ (.A_N(_12433_[0]),
    .B(_02449_),
    .Y(_02701_));
 sky130_fd_sc_hd__o221ai_2 _23413_ (.A1(_02532_),
    .A2(_02700_),
    .B1(_02701_),
    .B2(_02480_),
    .C1(_02472_),
    .Y(_02702_));
 sky130_fd_sc_hd__a31oi_2 _23414_ (.A1(_02480_),
    .A2(_02644_),
    .A3(_02699_),
    .B1(_02702_),
    .Y(_02703_));
 sky130_fd_sc_hd__nor2_4 _23415_ (.A(_02449_),
    .B(net3734),
    .Y(_02704_));
 sky130_fd_sc_hd__a21oi_1 _23416_ (.A1(_02692_),
    .A2(_02684_),
    .B1(net3747),
    .Y(_02705_));
 sky130_fd_sc_hd__a211oi_1 _23417_ (.A1(_12433_[0]),
    .A2(_02704_),
    .B1(_02705_),
    .C1(_02537_),
    .Y(_02706_));
 sky130_fd_sc_hd__o21ai_0 _23418_ (.A1(_02472_),
    .A2(_02706_),
    .B1(net3641),
    .Y(_02707_));
 sky130_fd_sc_hd__o22ai_1 _23419_ (.A1(net3641),
    .A2(_02698_),
    .B1(_02703_),
    .B2(_02707_),
    .Y(_02708_));
 sky130_fd_sc_hd__nand2_2 _23420_ (.A(_12438_[0]),
    .B(net3738),
    .Y(_02709_));
 sky130_fd_sc_hd__a21oi_1 _23421_ (.A1(_02651_),
    .A2(_02709_),
    .B1(net3747),
    .Y(_02710_));
 sky130_fd_sc_hd__a31oi_1 _23422_ (.A1(net3747),
    .A2(_02655_),
    .A3(_02651_),
    .B1(_02710_),
    .Y(_02711_));
 sky130_fd_sc_hd__nor3_1 _23423_ (.A(_02449_),
    .B(_02669_),
    .C(_02606_),
    .Y(_02712_));
 sky130_fd_sc_hd__nor2_4 _23424_ (.A(_12442_[0]),
    .B(net3732),
    .Y(_02713_));
 sky130_fd_sc_hd__nor3_1 _23425_ (.A(net3746),
    .B(_02619_),
    .C(_02713_),
    .Y(_02714_));
 sky130_fd_sc_hd__o21ai_0 _23426_ (.A1(_02712_),
    .A2(_02714_),
    .B1(_02504_),
    .Y(_02715_));
 sky130_fd_sc_hd__nand3_1 _23427_ (.A(net3747),
    .B(_02612_),
    .C(_02709_),
    .Y(_02716_));
 sky130_fd_sc_hd__a31oi_1 _23428_ (.A1(_02472_),
    .A2(_02716_),
    .A3(_02701_),
    .B1(net3642),
    .Y(_02717_));
 sky130_fd_sc_hd__nand2b_4 _23429_ (.A_N(_12442_[0]),
    .B(_02480_),
    .Y(_02718_));
 sky130_fd_sc_hd__nor2_4 _23430_ (.A(_02444_),
    .B(_02489_),
    .Y(_02719_));
 sky130_fd_sc_hd__nor2_1 _23431_ (.A(_12438_[0]),
    .B(_02480_),
    .Y(_02720_));
 sky130_fd_sc_hd__nor3_1 _23432_ (.A(_02449_),
    .B(_02719_),
    .C(_02720_),
    .Y(_02721_));
 sky130_fd_sc_hd__a31oi_1 _23433_ (.A1(_02449_),
    .A2(_02612_),
    .A3(_02718_),
    .B1(_02721_),
    .Y(_02722_));
 sky130_fd_sc_hd__a222oi_1 _23434_ (.A1(_02668_),
    .A2(_02711_),
    .B1(_02715_),
    .B2(_02717_),
    .C1(_02722_),
    .C2(_02662_),
    .Y(_02723_));
 sky130_fd_sc_hd__nand2_4 _23435_ (.A(net3732),
    .B(_02572_),
    .Y(_02724_));
 sky130_fd_sc_hd__a21oi_1 _23436_ (.A1(_02673_),
    .A2(_02724_),
    .B1(_02449_),
    .Y(_02725_));
 sky130_fd_sc_hd__nand2_1 _23437_ (.A(_12436_[0]),
    .B(_02480_),
    .Y(_02726_));
 sky130_fd_sc_hd__a21oi_1 _23438_ (.A1(_02685_),
    .A2(_02726_),
    .B1(net3746),
    .Y(_02727_));
 sky130_fd_sc_hd__o21ai_0 _23439_ (.A1(_02725_),
    .A2(_02727_),
    .B1(_02504_),
    .Y(_02728_));
 sky130_fd_sc_hd__a32oi_1 _23440_ (.A1(net3746),
    .A2(_02651_),
    .A3(_02636_),
    .B1(_02584_),
    .B2(_12433_[0]),
    .Y(_02729_));
 sky130_fd_sc_hd__nand2_1 _23441_ (.A(net3743),
    .B(_02729_),
    .Y(_02730_));
 sky130_fd_sc_hd__a21oi_1 _23442_ (.A1(_12447_[0]),
    .A2(net3732),
    .B1(net3730),
    .Y(_02731_));
 sky130_fd_sc_hd__o21ai_0 _23443_ (.A1(_02515_),
    .A2(_02700_),
    .B1(_02731_),
    .Y(_02732_));
 sky130_fd_sc_hd__o221ai_1 _23444_ (.A1(_12456_[0]),
    .A2(net3732),
    .B1(_02612_),
    .B2(_02614_),
    .C1(net3730),
    .Y(_02733_));
 sky130_fd_sc_hd__a21oi_1 _23445_ (.A1(_02732_),
    .A2(_02733_),
    .B1(net3642),
    .Y(_02734_));
 sky130_fd_sc_hd__nand2_4 _23446_ (.A(_02456_),
    .B(_02569_),
    .Y(_02735_));
 sky130_fd_sc_hd__a311o_1 _23447_ (.A1(net3642),
    .A2(_02728_),
    .A3(_02730_),
    .B1(_02734_),
    .C1(_02735_),
    .X(_02736_));
 sky130_fd_sc_hd__o21ai_0 _23448_ (.A1(_02566_),
    .A2(_02723_),
    .B1(_02736_),
    .Y(_02737_));
 sky130_fd_sc_hd__a311oi_1 _23449_ (.A1(net3643),
    .A2(net3749),
    .A3(net3746),
    .B1(net3737),
    .C1(_02508_),
    .Y(_02738_));
 sky130_fd_sc_hd__a21oi_1 _23450_ (.A1(_12449_[0]),
    .A2(net3737),
    .B1(_02738_),
    .Y(_02739_));
 sky130_fd_sc_hd__a2bb2oi_1 _23451_ (.A1_N(_02699_),
    .A2_N(_02593_),
    .B1(_02537_),
    .B2(_02486_),
    .Y(_02740_));
 sky130_fd_sc_hd__o21ai_0 _23452_ (.A1(_02541_),
    .A2(_02511_),
    .B1(_12429_[0]),
    .Y(_02741_));
 sky130_fd_sc_hd__a21oi_1 _23453_ (.A1(_02740_),
    .A2(_02741_),
    .B1(net3742),
    .Y(_02742_));
 sky130_fd_sc_hd__a211oi_1 _23454_ (.A1(net3742),
    .A2(_02739_),
    .B1(_02742_),
    .C1(net3640),
    .Y(_02743_));
 sky130_fd_sc_hd__nand2_1 _23455_ (.A(_12436_[0]),
    .B(net3732),
    .Y(_02744_));
 sky130_fd_sc_hd__nand3_1 _23456_ (.A(net3746),
    .B(_02507_),
    .C(_02744_),
    .Y(_02745_));
 sky130_fd_sc_hd__nand3_1 _23457_ (.A(_02449_),
    .B(_02651_),
    .C(_02636_),
    .Y(_02746_));
 sky130_fd_sc_hd__o21ai_1 _23458_ (.A1(_12452_[0]),
    .A2(net3733),
    .B1(net3743),
    .Y(_02747_));
 sky130_fd_sc_hd__a31oi_1 _23459_ (.A1(net3732),
    .A2(_02699_),
    .A3(_02484_),
    .B1(_02747_),
    .Y(_02748_));
 sky130_fd_sc_hd__a311oi_1 _23460_ (.A1(_02504_),
    .A2(_02745_),
    .A3(_02746_),
    .B1(_02748_),
    .C1(net3642),
    .Y(_02749_));
 sky130_fd_sc_hd__nor3_1 _23461_ (.A(_02633_),
    .B(_02743_),
    .C(_02749_),
    .Y(_02750_));
 sky130_fd_sc_hd__a211oi_1 _23462_ (.A1(_02611_),
    .A2(_02708_),
    .B1(_02737_),
    .C1(_02750_),
    .Y(_00146_));
 sky130_fd_sc_hd__nor2_1 _23463_ (.A(_12436_[0]),
    .B(net3734),
    .Y(_02751_));
 sky130_fd_sc_hd__nor3_1 _23464_ (.A(net3745),
    .B(_02605_),
    .C(_02751_),
    .Y(_02752_));
 sky130_fd_sc_hd__a311oi_1 _23465_ (.A1(net3745),
    .A2(_02690_),
    .A3(_02507_),
    .B1(_02752_),
    .C1(_02467_),
    .Y(_02753_));
 sky130_fd_sc_hd__a211oi_1 _23466_ (.A1(_02690_),
    .A2(_02594_),
    .B1(_02449_),
    .C1(_02525_),
    .Y(_02754_));
 sky130_fd_sc_hd__nand2_1 _23467_ (.A(_12438_[0]),
    .B(_02516_),
    .Y(_02755_));
 sky130_fd_sc_hd__nand2_2 _23468_ (.A(_02444_),
    .B(_02704_),
    .Y(_02756_));
 sky130_fd_sc_hd__nor3_1 _23469_ (.A(net3745),
    .B(_02719_),
    .C(net3576),
    .Y(_02757_));
 sky130_fd_sc_hd__a311oi_1 _23470_ (.A1(net3745),
    .A2(_02594_),
    .A3(_02724_),
    .B1(_02757_),
    .C1(_02646_),
    .Y(_02758_));
 sky130_fd_sc_hd__a311oi_1 _23471_ (.A1(_02668_),
    .A2(_02755_),
    .A3(_02756_),
    .B1(_02758_),
    .C1(_02461_),
    .Y(_02759_));
 sky130_fd_sc_hd__o31ai_1 _23472_ (.A1(net3740),
    .A2(_02753_),
    .A3(_02754_),
    .B1(_02759_),
    .Y(_02760_));
 sky130_fd_sc_hd__o21ai_2 _23473_ (.A1(_12438_[0]),
    .A2(_02480_),
    .B1(_02726_),
    .Y(_02761_));
 sky130_fd_sc_hd__a21oi_1 _23474_ (.A1(_02449_),
    .A2(_02761_),
    .B1(_02725_),
    .Y(_02762_));
 sky130_fd_sc_hd__o211ai_1 _23475_ (.A1(_02525_),
    .A2(_02692_),
    .B1(_02718_),
    .C1(_02449_),
    .Y(_02763_));
 sky130_fd_sc_hd__nand2_8 _23476_ (.A(_12438_[0]),
    .B(_02489_),
    .Y(_02764_));
 sky130_fd_sc_hd__nand3_1 _23477_ (.A(_02467_),
    .B(_02499_),
    .C(_02764_),
    .Y(_02765_));
 sky130_fd_sc_hd__o211ai_1 _23478_ (.A1(net3642),
    .A2(_02655_),
    .B1(_02765_),
    .C1(net3746),
    .Y(_02766_));
 sky130_fd_sc_hd__a21oi_1 _23479_ (.A1(net3746),
    .A2(_02507_),
    .B1(net3749),
    .Y(_02767_));
 sky130_fd_sc_hd__a2111oi_0 _23480_ (.A1(net3644),
    .A2(_02551_),
    .B1(_02575_),
    .C1(_02767_),
    .D1(net3640),
    .Y(_02768_));
 sky130_fd_sc_hd__a31oi_1 _23481_ (.A1(_02504_),
    .A2(_02763_),
    .A3(_02766_),
    .B1(_02768_),
    .Y(_02769_));
 sky130_fd_sc_hd__o211ai_1 _23482_ (.A1(_02646_),
    .A2(_02762_),
    .B1(_02769_),
    .C1(_02461_),
    .Y(_02770_));
 sky130_fd_sc_hd__nand2_1 _23483_ (.A(_12436_[0]),
    .B(_02573_),
    .Y(_02771_));
 sky130_fd_sc_hd__o21ai_0 _23484_ (.A1(_12429_[0]),
    .A2(_02515_),
    .B1(_02771_),
    .Y(_02772_));
 sky130_fd_sc_hd__a21oi_1 _23485_ (.A1(_02554_),
    .A2(_02756_),
    .B1(net3750),
    .Y(_02773_));
 sky130_fd_sc_hd__a221o_1 _23486_ (.A1(_12436_[0]),
    .A2(_02551_),
    .B1(_02669_),
    .B2(net3750),
    .C1(net3741),
    .X(_02774_));
 sky130_fd_sc_hd__o32ai_1 _23487_ (.A1(net3729),
    .A2(_02772_),
    .A3(_02773_),
    .B1(_02774_),
    .B2(_02693_),
    .Y(_02775_));
 sky130_fd_sc_hd__o21ai_0 _23488_ (.A1(_02606_),
    .A2(net3576),
    .B1(_02449_),
    .Y(_02776_));
 sky130_fd_sc_hd__nand3_4 _23489_ (.A(net3745),
    .B(_02594_),
    .C(_02612_),
    .Y(_02777_));
 sky130_fd_sc_hd__nand3_1 _23490_ (.A(net3729),
    .B(_02776_),
    .C(_02777_),
    .Y(_02778_));
 sky130_fd_sc_hd__nor2_1 _23491_ (.A(net3643),
    .B(_02444_),
    .Y(_02779_));
 sky130_fd_sc_hd__o31ai_1 _23492_ (.A1(_02573_),
    .A2(_02779_),
    .A3(_02614_),
    .B1(net3741),
    .Y(_02780_));
 sky130_fd_sc_hd__a21oi_1 _23493_ (.A1(_02778_),
    .A2(_02780_),
    .B1(_02467_),
    .Y(_02781_));
 sky130_fd_sc_hd__a211oi_1 _23494_ (.A1(_02467_),
    .A2(_02775_),
    .B1(_02781_),
    .C1(_02633_),
    .Y(_02782_));
 sky130_fd_sc_hd__nand3_1 _23495_ (.A(_02449_),
    .B(_02651_),
    .C(_02543_),
    .Y(_02783_));
 sky130_fd_sc_hd__o311ai_0 _23496_ (.A1(_02449_),
    .A2(_02495_),
    .A3(_02751_),
    .B1(_02783_),
    .C1(_02662_),
    .Y(_02784_));
 sky130_fd_sc_hd__nor2_4 _23497_ (.A(_02467_),
    .B(net3741),
    .Y(_02785_));
 sky130_fd_sc_hd__o21ai_0 _23498_ (.A1(_02556_),
    .A2(_02605_),
    .B1(_02449_),
    .Y(_02786_));
 sky130_fd_sc_hd__nand2_1 _23499_ (.A(net3749),
    .B(_02704_),
    .Y(_02787_));
 sky130_fd_sc_hd__a31oi_1 _23500_ (.A1(_02785_),
    .A2(_02786_),
    .A3(_02787_),
    .B1(_02735_),
    .Y(_02788_));
 sky130_fd_sc_hd__nand2_1 _23501_ (.A(_02784_),
    .B(_02788_),
    .Y(_02789_));
 sky130_fd_sc_hd__a32oi_1 _23502_ (.A1(net3644),
    .A2(_02449_),
    .A3(_02655_),
    .B1(_02556_),
    .B2(_02486_),
    .Y(_02790_));
 sky130_fd_sc_hd__a21oi_1 _23503_ (.A1(_02519_),
    .A2(_02790_),
    .B1(_02646_),
    .Y(_02791_));
 sky130_fd_sc_hd__o211ai_1 _23504_ (.A1(_12442_[0]),
    .A2(net3736),
    .B1(_02499_),
    .C1(net3745),
    .Y(_02792_));
 sky130_fd_sc_hd__or3_1 _23505_ (.A(net3745),
    .B(_02556_),
    .C(_02619_),
    .X(_02793_));
 sky130_fd_sc_hd__a21oi_1 _23506_ (.A1(_02792_),
    .A2(_02793_),
    .B1(_02642_),
    .Y(_02794_));
 sky130_fd_sc_hd__nor3_2 _23507_ (.A(_02789_),
    .B(_02791_),
    .C(_02794_),
    .Y(_02795_));
 sky130_fd_sc_hd__a311oi_1 _23508_ (.A1(_02565_),
    .A2(_02760_),
    .A3(_02770_),
    .B1(_02782_),
    .C1(_02795_),
    .Y(_00147_));
 sky130_fd_sc_hd__nand3_1 _23509_ (.A(_12429_[0]),
    .B(_02449_),
    .C(net3733),
    .Y(_02796_));
 sky130_fd_sc_hd__nand2_1 _23510_ (.A(_12440_[0]),
    .B(net3737),
    .Y(_02797_));
 sky130_fd_sc_hd__nor2_1 _23511_ (.A(net3643),
    .B(_02532_),
    .Y(_02798_));
 sky130_fd_sc_hd__a2111oi_1 _23512_ (.A1(_02449_),
    .A2(_02764_),
    .B1(_02798_),
    .C1(net3743),
    .D1(_02656_),
    .Y(_02799_));
 sky130_fd_sc_hd__a31oi_2 _23513_ (.A1(net3743),
    .A2(_02796_),
    .A3(_02797_),
    .B1(_02799_),
    .Y(_02800_));
 sky130_fd_sc_hd__a21oi_1 _23514_ (.A1(_02597_),
    .A2(_02692_),
    .B1(_02449_),
    .Y(_02801_));
 sky130_fd_sc_hd__o22ai_1 _23515_ (.A1(_12428_[0]),
    .A2(_02515_),
    .B1(_02664_),
    .B2(net3643),
    .Y(_02802_));
 sky130_fd_sc_hd__o21ai_1 _23516_ (.A1(_02669_),
    .A2(_02556_),
    .B1(net3746),
    .Y(_02803_));
 sky130_fd_sc_hd__nand4_1 _23517_ (.A(_02504_),
    .B(_02585_),
    .C(_02673_),
    .D(_02803_),
    .Y(_02804_));
 sky130_fd_sc_hd__o311ai_0 _23518_ (.A1(net3731),
    .A2(_02801_),
    .A3(_02802_),
    .B1(_02804_),
    .C1(net3641),
    .Y(_02805_));
 sky130_fd_sc_hd__o21ai_0 _23519_ (.A1(net3641),
    .A2(_02800_),
    .B1(_02805_),
    .Y(_02806_));
 sky130_fd_sc_hd__a21oi_1 _23520_ (.A1(_02449_),
    .A2(_02764_),
    .B1(_02580_),
    .Y(_02807_));
 sky130_fd_sc_hd__nand3_1 _23521_ (.A(_02449_),
    .B(_02612_),
    .C(_02636_),
    .Y(_02808_));
 sky130_fd_sc_hd__nand3_1 _23522_ (.A(net3743),
    .B(_02486_),
    .C(_02808_),
    .Y(_02809_));
 sky130_fd_sc_hd__o21ai_0 _23523_ (.A1(net3743),
    .A2(_02807_),
    .B1(_02809_),
    .Y(_02810_));
 sky130_fd_sc_hd__nor2_2 _23524_ (.A(net3747),
    .B(net3731),
    .Y(_02811_));
 sky130_fd_sc_hd__nor2_2 _23525_ (.A(net3747),
    .B(net3743),
    .Y(_02812_));
 sky130_fd_sc_hd__a32oi_1 _23526_ (.A1(_02499_),
    .A2(_02764_),
    .A3(_02811_),
    .B1(_02812_),
    .B2(_02653_),
    .Y(_02813_));
 sky130_fd_sc_hd__a21oi_1 _23527_ (.A1(_12438_[0]),
    .A2(net3731),
    .B1(_02449_),
    .Y(_02814_));
 sky130_fd_sc_hd__o31ai_1 _23528_ (.A1(net3731),
    .A2(_02581_),
    .A3(_02713_),
    .B1(_02814_),
    .Y(_02815_));
 sky130_fd_sc_hd__a21oi_1 _23529_ (.A1(_02813_),
    .A2(_02815_),
    .B1(_02461_),
    .Y(_02816_));
 sky130_fd_sc_hd__a2111oi_0 _23530_ (.A1(_02461_),
    .A2(_02810_),
    .B1(net3641),
    .C1(_02565_),
    .D1(_02816_),
    .Y(_02817_));
 sky130_fd_sc_hd__a21oi_2 _23531_ (.A1(_12433_[0]),
    .A2(net3746),
    .B1(_02508_),
    .Y(_02818_));
 sky130_fd_sc_hd__nand3_1 _23532_ (.A(net3732),
    .B(_02536_),
    .C(_02623_),
    .Y(_02819_));
 sky130_fd_sc_hd__o211ai_1 _23533_ (.A1(net3732),
    .A2(_02818_),
    .B1(_02819_),
    .C1(net3743),
    .Y(_02820_));
 sky130_fd_sc_hd__o21ai_4 _23534_ (.A1(net3751),
    .A2(net3749),
    .B1(net3732),
    .Y(_02821_));
 sky130_fd_sc_hd__nand3_1 _23535_ (.A(_02597_),
    .B(_02821_),
    .C(_02812_),
    .Y(_02822_));
 sky130_fd_sc_hd__a211oi_1 _23536_ (.A1(_12428_[0]),
    .A2(_02480_),
    .B1(_02619_),
    .C1(_02449_),
    .Y(_02823_));
 sky130_fd_sc_hd__a311oi_1 _23537_ (.A1(_02449_),
    .A2(_02560_),
    .A3(_02618_),
    .B1(_02823_),
    .C1(net3743),
    .Y(_02824_));
 sky130_fd_sc_hd__a221oi_1 _23538_ (.A1(net3749),
    .A2(_02704_),
    .B1(_02718_),
    .B2(_02449_),
    .C1(net3731),
    .Y(_02825_));
 sky130_fd_sc_hd__nor3_1 _23539_ (.A(net3642),
    .B(_02824_),
    .C(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__a31oi_1 _23540_ (.A1(net3642),
    .A2(_02820_),
    .A3(_02822_),
    .B1(_02826_),
    .Y(_02827_));
 sky130_fd_sc_hd__o21ai_0 _23541_ (.A1(_02444_),
    .A2(_02811_),
    .B1(net3643),
    .Y(_02828_));
 sky130_fd_sc_hd__and3_1 _23542_ (.A(_02480_),
    .B(_02486_),
    .C(_02828_),
    .X(_02829_));
 sky130_fd_sc_hd__nor2_1 _23543_ (.A(_02449_),
    .B(net3731),
    .Y(_02830_));
 sky130_fd_sc_hd__a221oi_1 _23544_ (.A1(net3643),
    .A2(_02830_),
    .B1(_02812_),
    .B2(_12428_[0]),
    .C1(_02480_),
    .Y(_02831_));
 sky130_fd_sc_hd__nor2_1 _23545_ (.A(_02504_),
    .B(_02664_),
    .Y(_02832_));
 sky130_fd_sc_hd__a21oi_1 _23546_ (.A1(net3747),
    .A2(net3731),
    .B1(_02832_),
    .Y(_02833_));
 sky130_fd_sc_hd__nor2_1 _23547_ (.A(net3642),
    .B(_02633_),
    .Y(_02834_));
 sky130_fd_sc_hd__o221ai_1 _23548_ (.A1(_02829_),
    .A2(_02831_),
    .B1(_02833_),
    .B2(net3643),
    .C1(_02834_),
    .Y(_02835_));
 sky130_fd_sc_hd__nor3_1 _23549_ (.A(_12433_[0]),
    .B(_02830_),
    .C(_02812_),
    .Y(_02836_));
 sky130_fd_sc_hd__nor3_1 _23550_ (.A(_02449_),
    .B(net3730),
    .C(_02700_),
    .Y(_02837_));
 sky130_fd_sc_hd__nor3_1 _23551_ (.A(_12442_[0]),
    .B(net3746),
    .C(net3743),
    .Y(_02838_));
 sky130_fd_sc_hd__a21oi_1 _23552_ (.A1(net3643),
    .A2(net3749),
    .B1(_02472_),
    .Y(_02839_));
 sky130_fd_sc_hd__nor2_1 _23553_ (.A(_12428_[0]),
    .B(_02504_),
    .Y(_02840_));
 sky130_fd_sc_hd__nand2_1 _23554_ (.A(net3751),
    .B(_02449_),
    .Y(_02841_));
 sky130_fd_sc_hd__o311ai_0 _23555_ (.A1(_02449_),
    .A2(_02839_),
    .A3(_02840_),
    .B1(net3732),
    .C1(_02841_),
    .Y(_02842_));
 sky130_fd_sc_hd__o41ai_1 _23556_ (.A1(net3732),
    .A2(_02836_),
    .A3(_02837_),
    .A4(_02838_),
    .B1(_02842_),
    .Y(_02843_));
 sky130_fd_sc_hd__nand3_1 _23557_ (.A(net3641),
    .B(_02661_),
    .C(_02843_),
    .Y(_02844_));
 sky130_fd_sc_hd__o211ai_1 _23558_ (.A1(_02566_),
    .A2(_02827_),
    .B1(_02835_),
    .C1(_02844_),
    .Y(_02845_));
 sky130_fd_sc_hd__a211o_1 _23559_ (.A1(_02611_),
    .A2(_02806_),
    .B1(_02817_),
    .C1(_02845_),
    .X(_00148_));
 sky130_fd_sc_hd__nand2_1 _23560_ (.A(_12438_[0]),
    .B(_02551_),
    .Y(_02846_));
 sky130_fd_sc_hd__nand4_1 _23561_ (.A(_02588_),
    .B(_02598_),
    .C(_02662_),
    .D(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__a32oi_1 _23562_ (.A1(net3745),
    .A2(_02499_),
    .A3(_02764_),
    .B1(_02584_),
    .B2(_02444_),
    .Y(_02848_));
 sky130_fd_sc_hd__a311oi_1 _23563_ (.A1(_02449_),
    .A2(_02507_),
    .A3(_02559_),
    .B1(_02599_),
    .C1(_02525_),
    .Y(_02849_));
 sky130_fd_sc_hd__a211o_1 _23564_ (.A1(_02525_),
    .A2(_02848_),
    .B1(_02849_),
    .C1(net3729),
    .X(_02850_));
 sky130_fd_sc_hd__a21oi_1 _23565_ (.A1(net3591),
    .A2(net3739),
    .B1(_02467_),
    .Y(_02851_));
 sky130_fd_sc_hd__o211ai_1 _23566_ (.A1(net3745),
    .A2(_02581_),
    .B1(_02851_),
    .C1(net3729),
    .Y(_02852_));
 sky130_fd_sc_hd__a31oi_1 _23567_ (.A1(_02847_),
    .A2(_02850_),
    .A3(_02852_),
    .B1(_02633_),
    .Y(_02853_));
 sky130_fd_sc_hd__o21ai_1 _23568_ (.A1(_12436_[0]),
    .A2(net3739),
    .B1(_02684_),
    .Y(_02854_));
 sky130_fd_sc_hd__mux2i_1 _23569_ (.A0(_02492_),
    .A1(_02854_),
    .S(_02449_),
    .Y(_02855_));
 sky130_fd_sc_hd__nor3_1 _23570_ (.A(net3745),
    .B(_02581_),
    .C(_02606_),
    .Y(_02856_));
 sky130_fd_sc_hd__a311oi_1 _23571_ (.A1(net3745),
    .A2(_02507_),
    .A3(_02651_),
    .B1(_02856_),
    .C1(_02525_),
    .Y(_02857_));
 sky130_fd_sc_hd__a21oi_1 _23572_ (.A1(_02525_),
    .A2(_02855_),
    .B1(_02857_),
    .Y(_02858_));
 sky130_fd_sc_hd__nor2_1 _23573_ (.A(net3749),
    .B(_02516_),
    .Y(_02859_));
 sky130_fd_sc_hd__a221oi_1 _23574_ (.A1(net3591),
    .A2(_02551_),
    .B1(_02602_),
    .B2(net3745),
    .C1(_02859_),
    .Y(_02860_));
 sky130_fd_sc_hd__o21ai_0 _23575_ (.A1(net3749),
    .A2(_02704_),
    .B1(_02587_),
    .Y(_02861_));
 sky130_fd_sc_hd__a21oi_1 _23576_ (.A1(_02668_),
    .A2(_02861_),
    .B1(_02566_),
    .Y(_02862_));
 sky130_fd_sc_hd__o21ai_0 _23577_ (.A1(_02646_),
    .A2(_02860_),
    .B1(_02862_),
    .Y(_02863_));
 sky130_fd_sc_hd__a21oi_1 _23578_ (.A1(net3729),
    .A2(_02858_),
    .B1(_02863_),
    .Y(_02864_));
 sky130_fd_sc_hd__nand2_2 _23579_ (.A(_02449_),
    .B(net3735),
    .Y(_02865_));
 sky130_fd_sc_hd__nor2_1 _23580_ (.A(_12442_[0]),
    .B(_02865_),
    .Y(_02866_));
 sky130_fd_sc_hd__a21oi_1 _23581_ (.A1(net3591),
    .A2(_02449_),
    .B1(net3735),
    .Y(_02867_));
 sky130_fd_sc_hd__o21ai_0 _23582_ (.A1(_02866_),
    .A2(_02867_),
    .B1(_02467_),
    .Y(_02868_));
 sky130_fd_sc_hd__a21oi_1 _23583_ (.A1(_02594_),
    .A2(_02635_),
    .B1(_02449_),
    .Y(_02869_));
 sky130_fd_sc_hd__a21oi_1 _23584_ (.A1(_02449_),
    .A2(_02854_),
    .B1(_02869_),
    .Y(_02870_));
 sky130_fd_sc_hd__nand2_1 _23585_ (.A(_02525_),
    .B(_02870_),
    .Y(_02871_));
 sky130_fd_sc_hd__o32ai_1 _23586_ (.A1(_02560_),
    .A2(_02613_),
    .A3(_02614_),
    .B1(_02724_),
    .B2(_02449_),
    .Y(_02872_));
 sky130_fd_sc_hd__nor2_4 _23587_ (.A(net3642),
    .B(net3731),
    .Y(_02873_));
 sky130_fd_sc_hd__o211ai_1 _23588_ (.A1(net3732),
    .A2(_02623_),
    .B1(_02744_),
    .C1(_02873_),
    .Y(_02874_));
 sky130_fd_sc_hd__o211ai_1 _23589_ (.A1(_02642_),
    .A2(_02872_),
    .B1(_02874_),
    .C1(_02611_),
    .Y(_02875_));
 sky130_fd_sc_hd__a31oi_1 _23590_ (.A1(net3729),
    .A2(_02868_),
    .A3(_02871_),
    .B1(_02875_),
    .Y(_02876_));
 sky130_fd_sc_hd__nand2_4 _23591_ (.A(net3741),
    .B(net3734),
    .Y(_02877_));
 sky130_fd_sc_hd__a21oi_1 _23592_ (.A1(_02550_),
    .A2(_02877_),
    .B1(net3644),
    .Y(_02878_));
 sky130_fd_sc_hd__nand2_1 _23593_ (.A(_12436_[0]),
    .B(_02584_),
    .Y(_02879_));
 sky130_fd_sc_hd__a21oi_1 _23594_ (.A1(_02787_),
    .A2(_02879_),
    .B1(net3741),
    .Y(_02880_));
 sky130_fd_sc_hd__o2111ai_1 _23595_ (.A1(net3741),
    .A2(_02573_),
    .B1(_02877_),
    .C1(_02444_),
    .D1(net3644),
    .Y(_02881_));
 sky130_fd_sc_hd__o31ai_1 _23596_ (.A1(net3749),
    .A2(net3741),
    .A3(_02507_),
    .B1(_02881_),
    .Y(_02882_));
 sky130_fd_sc_hd__nor4_1 _23597_ (.A(net3641),
    .B(_02878_),
    .C(_02880_),
    .D(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__a21oi_1 _23598_ (.A1(_02597_),
    .A2(_02635_),
    .B1(net3745),
    .Y(_02884_));
 sky130_fd_sc_hd__a211oi_1 _23599_ (.A1(net3750),
    .A2(_02704_),
    .B1(_02884_),
    .C1(net3741),
    .Y(_02885_));
 sky130_fd_sc_hd__o21ai_0 _23600_ (.A1(_12428_[0]),
    .A2(net3739),
    .B1(_02684_),
    .Y(_02886_));
 sky130_fd_sc_hd__nor2_1 _23601_ (.A(_12429_[0]),
    .B(_02532_),
    .Y(_02887_));
 sky130_fd_sc_hd__a211oi_1 _23602_ (.A1(_02449_),
    .A2(_02886_),
    .B1(_02887_),
    .C1(net3729),
    .Y(_02888_));
 sky130_fd_sc_hd__nor3_1 _23603_ (.A(_02467_),
    .B(_02885_),
    .C(_02888_),
    .Y(_02889_));
 sky130_fd_sc_hd__nor3_1 _23604_ (.A(_02735_),
    .B(_02883_),
    .C(_02889_),
    .Y(_02890_));
 sky130_fd_sc_hd__nor4_1 _23605_ (.A(_02853_),
    .B(_02864_),
    .C(_02876_),
    .D(_02890_),
    .Y(_00149_));
 sky130_fd_sc_hd__o21ai_0 _23606_ (.A1(_02580_),
    .A2(_02581_),
    .B1(_02449_),
    .Y(_02891_));
 sky130_fd_sc_hd__nor2_1 _23607_ (.A(net3746),
    .B(_02700_),
    .Y(_02892_));
 sky130_fd_sc_hd__o21ai_0 _23608_ (.A1(_12429_[0]),
    .A2(_02449_),
    .B1(_02480_),
    .Y(_02893_));
 sky130_fd_sc_hd__o22ai_2 _23609_ (.A1(_12447_[0]),
    .A2(_02480_),
    .B1(_02892_),
    .B2(_02893_),
    .Y(_02894_));
 sky130_fd_sc_hd__a32oi_1 _23610_ (.A1(_02668_),
    .A2(_02777_),
    .A3(_02891_),
    .B1(_02894_),
    .B2(_02662_),
    .Y(_02895_));
 sky130_fd_sc_hd__o211ai_1 _23611_ (.A1(net3732),
    .A2(_02818_),
    .B1(_02554_),
    .C1(_02472_),
    .Y(_02896_));
 sky130_fd_sc_hd__nor2_1 _23612_ (.A(net3749),
    .B(_02449_),
    .Y(_02897_));
 sky130_fd_sc_hd__o21ai_2 _23613_ (.A1(net3751),
    .A2(_02897_),
    .B1(net3733),
    .Y(_02898_));
 sky130_fd_sc_hd__o211ai_1 _23614_ (.A1(_12436_[0]),
    .A2(_02515_),
    .B1(_02898_),
    .C1(net3730),
    .Y(_02899_));
 sky130_fd_sc_hd__o211ai_1 _23615_ (.A1(_02582_),
    .A2(_02896_),
    .B1(_02899_),
    .C1(net3641),
    .Y(_02900_));
 sky130_fd_sc_hd__nor2_1 _23616_ (.A(net3643),
    .B(_02472_),
    .Y(_02901_));
 sky130_fd_sc_hd__o21ai_1 _23617_ (.A1(_02832_),
    .A2(_02901_),
    .B1(_02449_),
    .Y(_02902_));
 sky130_fd_sc_hd__a21oi_1 _23618_ (.A1(_12429_[0]),
    .A2(net3742),
    .B1(net3732),
    .Y(_02903_));
 sky130_fd_sc_hd__nor2_1 _23619_ (.A(_02449_),
    .B(_02903_),
    .Y(_02904_));
 sky130_fd_sc_hd__o21ai_0 _23620_ (.A1(_12438_[0]),
    .A2(_02877_),
    .B1(_02904_),
    .Y(_02905_));
 sky130_fd_sc_hd__o2111ai_1 _23621_ (.A1(net3742),
    .A2(_02543_),
    .B1(_02902_),
    .C1(_02905_),
    .D1(net3640),
    .Y(_02906_));
 sky130_fd_sc_hd__o21a_1 _23622_ (.A1(_02449_),
    .A2(_02484_),
    .B1(_02543_),
    .X(_02907_));
 sky130_fd_sc_hd__a21oi_1 _23623_ (.A1(net3751),
    .A2(_02669_),
    .B1(_02614_),
    .Y(_02908_));
 sky130_fd_sc_hd__o21ai_0 _23624_ (.A1(_12442_[0]),
    .A2(_02907_),
    .B1(_02908_),
    .Y(_02909_));
 sky130_fd_sc_hd__a2bb2oi_1 _23625_ (.A1_N(_02504_),
    .A2_N(_02614_),
    .B1(_02713_),
    .B2(net3746),
    .Y(_02910_));
 sky130_fd_sc_hd__o22ai_1 _23626_ (.A1(_02486_),
    .A2(_02877_),
    .B1(_02910_),
    .B2(net3751),
    .Y(_02911_));
 sky130_fd_sc_hd__a22oi_1 _23627_ (.A1(_02662_),
    .A2(_02909_),
    .B1(_02911_),
    .B2(net3642),
    .Y(_02912_));
 sky130_fd_sc_hd__a211o_1 _23628_ (.A1(_02449_),
    .A2(_02761_),
    .B1(_02798_),
    .C1(net3743),
    .X(_02913_));
 sky130_fd_sc_hd__o32ai_1 _23629_ (.A1(net3746),
    .A2(_02719_),
    .A3(_02542_),
    .B1(_02532_),
    .B2(_12429_[0]),
    .Y(_02914_));
 sky130_fd_sc_hd__a21oi_1 _23630_ (.A1(_12438_[0]),
    .A2(_02449_),
    .B1(_02489_),
    .Y(_02915_));
 sky130_fd_sc_hd__a221oi_1 _23631_ (.A1(_12446_[0]),
    .A2(_02489_),
    .B1(_02699_),
    .B2(_02915_),
    .C1(_02504_),
    .Y(_02916_));
 sky130_fd_sc_hd__a211oi_1 _23632_ (.A1(_02504_),
    .A2(_02914_),
    .B1(_02916_),
    .C1(net3640),
    .Y(_02917_));
 sky130_fd_sc_hd__a311oi_1 _23633_ (.A1(net3640),
    .A2(_02702_),
    .A3(_02913_),
    .B1(_02917_),
    .C1(_02461_),
    .Y(_02918_));
 sky130_fd_sc_hd__a311oi_2 _23634_ (.A1(_02461_),
    .A2(_02906_),
    .A3(_02912_),
    .B1(_02918_),
    .C1(_02456_),
    .Y(_02919_));
 sky130_fd_sc_hd__o21ai_0 _23635_ (.A1(_12428_[0]),
    .A2(net3732),
    .B1(_02764_),
    .Y(_02920_));
 sky130_fd_sc_hd__a22oi_1 _23636_ (.A1(_12430_[0]),
    .A2(_02584_),
    .B1(_02920_),
    .B2(net3746),
    .Y(_02921_));
 sky130_fd_sc_hd__a21oi_2 _23637_ (.A1(net3751),
    .A2(net3746),
    .B1(_02821_),
    .Y(_02922_));
 sky130_fd_sc_hd__o31ai_4 _23638_ (.A1(_12445_[0]),
    .A2(_12454_[0]),
    .A3(net3733),
    .B1(net3743),
    .Y(_02923_));
 sky130_fd_sc_hd__o22ai_2 _23639_ (.A1(net3743),
    .A2(_02921_),
    .B1(_02922_),
    .B2(_02923_),
    .Y(_02924_));
 sky130_fd_sc_hd__nand3_1 _23640_ (.A(_02449_),
    .B(_02821_),
    .C(_02709_),
    .Y(_02925_));
 sky130_fd_sc_hd__nand3_1 _23641_ (.A(net3745),
    .B(_02690_),
    .C(_02684_),
    .Y(_02926_));
 sky130_fd_sc_hd__o21ai_0 _23642_ (.A1(net3591),
    .A2(net3739),
    .B1(_02499_),
    .Y(_02927_));
 sky130_fd_sc_hd__and3_1 _23643_ (.A(net3745),
    .B(_02655_),
    .C(_02764_),
    .X(_02928_));
 sky130_fd_sc_hd__a31oi_1 _23644_ (.A1(_02449_),
    .A2(_02690_),
    .A3(_02927_),
    .B1(_02928_),
    .Y(_02929_));
 sky130_fd_sc_hd__a32o_1 _23645_ (.A1(_02873_),
    .A2(_02925_),
    .A3(_02926_),
    .B1(_02929_),
    .B2(_02785_),
    .X(_02930_));
 sky130_fd_sc_hd__a211oi_1 _23646_ (.A1(net3642),
    .A2(_02924_),
    .B1(_02930_),
    .C1(_02633_),
    .Y(_02931_));
 sky130_fd_sc_hd__a311oi_1 _23647_ (.A1(_02661_),
    .A2(_02895_),
    .A3(_02900_),
    .B1(_02919_),
    .C1(_02931_),
    .Y(_00150_));
 sky130_fd_sc_hd__a21oi_1 _23648_ (.A1(_02449_),
    .A2(_02593_),
    .B1(_02719_),
    .Y(_02932_));
 sky130_fd_sc_hd__a21oi_1 _23649_ (.A1(_12428_[0]),
    .A2(_02573_),
    .B1(_02631_),
    .Y(_02933_));
 sky130_fd_sc_hd__o21ai_1 _23650_ (.A1(net3751),
    .A2(_02932_),
    .B1(_02933_),
    .Y(_02934_));
 sky130_fd_sc_hd__o221ai_1 _23651_ (.A1(_12442_[0]),
    .A2(_02532_),
    .B1(_02516_),
    .B2(_12429_[0]),
    .C1(_02785_),
    .Y(_02935_));
 sky130_fd_sc_hd__a21oi_1 _23652_ (.A1(_02934_),
    .A2(_02935_),
    .B1(_02675_),
    .Y(_02936_));
 sky130_fd_sc_hd__nand3_1 _23653_ (.A(net3747),
    .B(_02692_),
    .C(_02684_),
    .Y(_02937_));
 sky130_fd_sc_hd__nand3_1 _23654_ (.A(_02449_),
    .B(_02612_),
    .C(_02709_),
    .Y(_02938_));
 sky130_fd_sc_hd__nand3_1 _23655_ (.A(_02873_),
    .B(_02937_),
    .C(_02938_),
    .Y(_02939_));
 sky130_fd_sc_hd__o21ai_0 _23656_ (.A1(_02537_),
    .A2(_02713_),
    .B1(net3747),
    .Y(_02940_));
 sky130_fd_sc_hd__o211ai_1 _23657_ (.A1(_12438_[0]),
    .A2(_02865_),
    .B1(_02668_),
    .C1(_02940_),
    .Y(_02941_));
 sky130_fd_sc_hd__nand2_1 _23658_ (.A(_02939_),
    .B(_02941_),
    .Y(_02942_));
 sky130_fd_sc_hd__nand2b_1 _23659_ (.A_N(_12433_[0]),
    .B(net3746),
    .Y(_02943_));
 sky130_fd_sc_hd__a21oi_1 _23660_ (.A1(_02841_),
    .A2(_02943_),
    .B1(net3737),
    .Y(_02944_));
 sky130_fd_sc_hd__o21ai_0 _23661_ (.A1(_02560_),
    .A2(_02897_),
    .B1(_02504_),
    .Y(_02945_));
 sky130_fd_sc_hd__nor2_1 _23662_ (.A(_12440_[0]),
    .B(net3737),
    .Y(_02946_));
 sky130_fd_sc_hd__a31oi_1 _23663_ (.A1(_12430_[0]),
    .A2(_02449_),
    .A3(net3737),
    .B1(_02946_),
    .Y(_02947_));
 sky130_fd_sc_hd__o22ai_1 _23664_ (.A1(_02944_),
    .A2(_02945_),
    .B1(_02947_),
    .B2(_02504_),
    .Y(_02948_));
 sky130_fd_sc_hd__nor2_1 _23665_ (.A(_12454_[0]),
    .B(net3737),
    .Y(_02949_));
 sky130_fd_sc_hd__a211oi_1 _23666_ (.A1(_12438_[0]),
    .A2(net3746),
    .B1(_02489_),
    .C1(_02508_),
    .Y(_02950_));
 sky130_fd_sc_hd__o31ai_1 _23667_ (.A1(_02504_),
    .A2(_02949_),
    .A3(_02950_),
    .B1(net3640),
    .Y(_02951_));
 sky130_fd_sc_hd__a311oi_1 _23668_ (.A1(net3746),
    .A2(_02651_),
    .A3(_02560_),
    .B1(_02679_),
    .C1(net3743),
    .Y(_02952_));
 sky130_fd_sc_hd__o22ai_1 _23669_ (.A1(net3640),
    .A2(_02948_),
    .B1(_02951_),
    .B2(_02952_),
    .Y(_02953_));
 sky130_fd_sc_hd__a21oi_1 _23670_ (.A1(_02673_),
    .A2(_02744_),
    .B1(net3746),
    .Y(_02954_));
 sky130_fd_sc_hd__o21ai_0 _23671_ (.A1(_02638_),
    .A2(_02954_),
    .B1(_02472_),
    .Y(_02955_));
 sky130_fd_sc_hd__nand2_1 _23672_ (.A(_02449_),
    .B(_02543_),
    .Y(_02956_));
 sky130_fd_sc_hd__nor2_1 _23673_ (.A(net3743),
    .B(_02556_),
    .Y(_02957_));
 sky130_fd_sc_hd__o221ai_1 _23674_ (.A1(_02532_),
    .A2(_02572_),
    .B1(_02956_),
    .B2(_02720_),
    .C1(_02957_),
    .Y(_02958_));
 sky130_fd_sc_hd__nand4_1 _23675_ (.A(_02461_),
    .B(net3642),
    .C(_02955_),
    .D(_02958_),
    .Y(_02959_));
 sky130_fd_sc_hd__nor2_1 _23676_ (.A(_12428_[0]),
    .B(_02449_),
    .Y(_02960_));
 sky130_fd_sc_hd__a31oi_1 _23677_ (.A1(_02449_),
    .A2(_02680_),
    .A3(_02612_),
    .B1(_02960_),
    .Y(_02961_));
 sky130_fd_sc_hd__o21ai_0 _23678_ (.A1(_12433_[0]),
    .A2(net3732),
    .B1(net3730),
    .Y(_02962_));
 sky130_fd_sc_hd__o22ai_1 _23679_ (.A1(net3730),
    .A2(_02961_),
    .B1(_02962_),
    .B2(_02922_),
    .Y(_02963_));
 sky130_fd_sc_hd__a31oi_1 _23680_ (.A1(_02461_),
    .A2(net3640),
    .A3(_02963_),
    .B1(_02565_),
    .Y(_02964_));
 sky130_fd_sc_hd__o211ai_1 _23681_ (.A1(_02461_),
    .A2(_02953_),
    .B1(_02959_),
    .C1(_02964_),
    .Y(_02965_));
 sky130_fd_sc_hd__o21ai_0 _23682_ (.A1(_02444_),
    .A2(_02532_),
    .B1(_02543_),
    .Y(_02966_));
 sky130_fd_sc_hd__o21ai_1 _23683_ (.A1(_02551_),
    .A2(_02593_),
    .B1(net3750),
    .Y(_02967_));
 sky130_fd_sc_hd__a21oi_1 _23684_ (.A1(_02587_),
    .A2(_02967_),
    .B1(net3729),
    .Y(_02968_));
 sky130_fd_sc_hd__a21oi_1 _23685_ (.A1(_02865_),
    .A2(_02756_),
    .B1(net3750),
    .Y(_02969_));
 sky130_fd_sc_hd__a211oi_1 _23686_ (.A1(net3729),
    .A2(_02966_),
    .B1(_02968_),
    .C1(_02969_),
    .Y(_02970_));
 sky130_fd_sc_hd__a21oi_1 _23687_ (.A1(_02515_),
    .A2(_02877_),
    .B1(net3749),
    .Y(_02971_));
 sky130_fd_sc_hd__a31oi_1 _23688_ (.A1(net3749),
    .A2(_02504_),
    .A3(_02573_),
    .B1(_02971_),
    .Y(_02972_));
 sky130_fd_sc_hd__nor2_1 _23689_ (.A(_02467_),
    .B(_02811_),
    .Y(_02973_));
 sky130_fd_sc_hd__o221ai_1 _23690_ (.A1(_02449_),
    .A2(_02499_),
    .B1(_02972_),
    .B2(net3750),
    .C1(_02973_),
    .Y(_02974_));
 sky130_fd_sc_hd__o211ai_1 _23691_ (.A1(net3641),
    .A2(_02970_),
    .B1(_02974_),
    .C1(_02611_),
    .Y(_02975_));
 sky130_fd_sc_hd__o311a_4 _23692_ (.A1(_02566_),
    .A2(_02936_),
    .A3(_02942_),
    .B1(_02965_),
    .C1(_02975_),
    .X(_00151_));
 sky130_fd_sc_hd__xor3_1 _23693_ (.A(\sa03_sr[7] ),
    .B(\sa03_sr[0] ),
    .C(\sa21_sub[1] ),
    .X(_02976_));
 sky130_fd_sc_hd__xnor3_1 _23694_ (.A(_00771_),
    .B(_00772_),
    .C(_02976_),
    .X(_02977_));
 sky130_fd_sc_hd__nand2_1 _23695_ (.A(net4230),
    .B(\text_in_r[1] ),
    .Y(_02978_));
 sky130_fd_sc_hd__o21a_4 _23696_ (.A1(net4230),
    .A2(_02977_),
    .B1(_02978_),
    .X(_02979_));
 sky130_fd_sc_hd__xor2_4 _23697_ (.A(net4134),
    .B(_02979_),
    .X(_02980_));
 sky130_fd_sc_hd__inv_16 _23698_ (.A(_02980_),
    .Y(_02981_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_67 ();
 sky130_fd_sc_hd__xnor3_1 _23701_ (.A(net4211),
    .B(net4195),
    .C(net4179),
    .X(_02983_));
 sky130_fd_sc_hd__xor2_1 _23702_ (.A(_07657_),
    .B(_02983_),
    .X(_02984_));
 sky130_fd_sc_hd__mux2i_2 _23703_ (.A0(\text_in_r[0] ),
    .A1(_02984_),
    .S(_05879_),
    .Y(_02985_));
 sky130_fd_sc_hd__xor2_4 _23704_ (.A(\u0.tmp_w[0] ),
    .B(_02985_),
    .X(_02986_));
 sky130_fd_sc_hd__clkinv_16 _23705_ (.A(_02986_),
    .Y(_02987_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_65 ();
 sky130_fd_sc_hd__xor2_1 _23708_ (.A(net4181),
    .B(net4222),
    .X(_02989_));
 sky130_fd_sc_hd__xnor2_1 _23709_ (.A(_07678_),
    .B(_02989_),
    .Y(_02990_));
 sky130_fd_sc_hd__mux2i_2 _23710_ (.A0(\text_in_r[2] ),
    .A1(_02990_),
    .S(_05879_),
    .Y(_02991_));
 sky130_fd_sc_hd__xnor2_4 _23711_ (.A(\u0.tmp_w[2] ),
    .B(_02991_),
    .Y(_02992_));
 sky130_fd_sc_hd__clkinv_16 _23712_ (.A(_02992_),
    .Y(_02993_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_56 ();
 sky130_fd_sc_hd__xnor3_1 _23722_ (.A(_07701_),
    .B(_07712_),
    .C(_00818_),
    .X(_03000_));
 sky130_fd_sc_hd__nand2_1 _23723_ (.A(net398),
    .B(\text_in_r[4] ),
    .Y(_03001_));
 sky130_fd_sc_hd__o21a_4 _23724_ (.A1(net398),
    .A2(_03000_),
    .B1(_03001_),
    .X(_03002_));
 sky130_fd_sc_hd__xnor2_1 _23725_ (.A(\u0.tmp_w[4] ),
    .B(_03002_),
    .Y(_03003_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_53 ();
 sky130_fd_sc_hd__xnor3_1 _23729_ (.A(_07723_),
    .B(_00825_),
    .C(_00826_),
    .X(_03007_));
 sky130_fd_sc_hd__nand2b_1 _23730_ (.A_N(\text_in_r[3] ),
    .B(net4230),
    .Y(_03008_));
 sky130_fd_sc_hd__o211a_4 _23731_ (.A1(net4230),
    .A2(_03007_),
    .B1(_03008_),
    .C1(\u0.tmp_w[3] ),
    .X(_03009_));
 sky130_fd_sc_hd__and2_0 _23732_ (.A(net4230),
    .B(\text_in_r[3] ),
    .X(_03010_));
 sky130_fd_sc_hd__a211oi_2 _23733_ (.A1(net4115),
    .A2(_03007_),
    .B1(_03010_),
    .C1(\u0.tmp_w[3] ),
    .Y(_03011_));
 sky130_fd_sc_hd__nor2_4 _23734_ (.A(_03009_),
    .B(_03011_),
    .Y(_03012_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_50 ();
 sky130_fd_sc_hd__nor2_1 _23738_ (.A(_02981_),
    .B(net3721),
    .Y(_03016_));
 sky130_fd_sc_hd__or2_4 _23739_ (.A(_03009_),
    .B(_03011_),
    .X(_03017_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_47 ();
 sky130_fd_sc_hd__nor2_2 _23743_ (.A(net3590),
    .B(_03017_),
    .Y(_03021_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_45 ();
 sky130_fd_sc_hd__o21ai_0 _23746_ (.A1(_03016_),
    .A2(_03021_),
    .B1(net3724),
    .Y(_03024_));
 sky130_fd_sc_hd__nor2_4 _23747_ (.A(net3724),
    .B(net3719),
    .Y(_03025_));
 sky130_fd_sc_hd__nand2_1 _23748_ (.A(net3725),
    .B(_03025_),
    .Y(_03026_));
 sky130_fd_sc_hd__nor2_4 _23749_ (.A(_02987_),
    .B(net3717),
    .Y(_03027_));
 sky130_fd_sc_hd__nor2_4 _23750_ (.A(net3728),
    .B(_03012_),
    .Y(_03028_));
 sky130_fd_sc_hd__o21ai_0 _23751_ (.A1(_03027_),
    .A2(_03028_),
    .B1(_02993_),
    .Y(_03029_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_42 ();
 sky130_fd_sc_hd__nand2_8 _23755_ (.A(net3724),
    .B(net3717),
    .Y(_03033_));
 sky130_fd_sc_hd__nor2_2 _23756_ (.A(_12462_[0]),
    .B(_03033_),
    .Y(_03034_));
 sky130_fd_sc_hd__nor2_1 _23757_ (.A(net3723),
    .B(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__a32oi_1 _23758_ (.A1(net3723),
    .A2(_03024_),
    .A3(_03026_),
    .B1(_03029_),
    .B2(_03035_),
    .Y(_03036_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_37 ();
 sky130_fd_sc_hd__nand2_8 _23764_ (.A(net3639),
    .B(net3724),
    .Y(_03041_));
 sky130_fd_sc_hd__a211oi_1 _23765_ (.A1(_12462_[0]),
    .A2(net3719),
    .B1(_03041_),
    .C1(net3723),
    .Y(_03042_));
 sky130_fd_sc_hd__a31oi_1 _23766_ (.A1(net3725),
    .A2(_02993_),
    .A3(net3723),
    .B1(_03042_),
    .Y(_03043_));
 sky130_fd_sc_hd__xnor3_1 _23767_ (.A(\sa32_sub[4] ),
    .B(\sa03_sr[4] ),
    .C(\sa03_sr[5] ),
    .X(_03044_));
 sky130_fd_sc_hd__xor2_1 _23768_ (.A(_07700_),
    .B(_03044_),
    .X(_03045_));
 sky130_fd_sc_hd__mux2i_4 _23769_ (.A0(\text_in_r[5] ),
    .A1(_03045_),
    .S(net4116),
    .Y(_03046_));
 sky130_fd_sc_hd__xnor2_4 _23770_ (.A(net4127),
    .B(_03046_),
    .Y(_03047_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_35 ();
 sky130_fd_sc_hd__xnor2_1 _23773_ (.A(\sa32_sub[5] ),
    .B(\sa03_sr[6] ),
    .Y(_03050_));
 sky130_fd_sc_hd__xnor2_1 _23774_ (.A(_07705_),
    .B(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hd__nand2_1 _23775_ (.A(net398),
    .B(\text_in_r[6] ),
    .Y(_03052_));
 sky130_fd_sc_hd__o21ai_2 _23776_ (.A1(net398),
    .A2(_03051_),
    .B1(_03052_),
    .Y(_03053_));
 sky130_fd_sc_hd__xnor2_4 _23777_ (.A(\u0.tmp_w[6] ),
    .B(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_34 ();
 sky130_fd_sc_hd__xnor2_1 _23779_ (.A(_07670_),
    .B(_09941_),
    .Y(_03056_));
 sky130_fd_sc_hd__xnor2_1 _23780_ (.A(net4191),
    .B(_03056_),
    .Y(_03057_));
 sky130_fd_sc_hd__mux2i_4 _23781_ (.A0(\text_in_r[7] ),
    .A1(_03057_),
    .S(net4116),
    .Y(_03058_));
 sky130_fd_sc_hd__xor2_4 _23782_ (.A(\u0.tmp_w[7] ),
    .B(_03058_),
    .X(_03059_));
 sky130_fd_sc_hd__nand2b_4 _23783_ (.A_N(_03054_),
    .B(_03059_),
    .Y(_03060_));
 sky130_fd_sc_hd__nor2_1 _23784_ (.A(net3715),
    .B(_03060_),
    .Y(_03061_));
 sky130_fd_sc_hd__o21ai_0 _23785_ (.A1(net3728),
    .A2(_03043_),
    .B1(_03061_),
    .Y(_03062_));
 sky130_fd_sc_hd__nand2_4 _23786_ (.A(net3727),
    .B(_03017_),
    .Y(_03063_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_32 ();
 sky130_fd_sc_hd__nand2_2 _23789_ (.A(net3590),
    .B(net3721),
    .Y(_03066_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_30 ();
 sky130_fd_sc_hd__a21oi_1 _23792_ (.A1(_03063_),
    .A2(_03066_),
    .B1(net3724),
    .Y(_03069_));
 sky130_fd_sc_hd__nand2_4 _23793_ (.A(_02987_),
    .B(net3719),
    .Y(_03070_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_28 ();
 sky130_fd_sc_hd__nand3_2 _23796_ (.A(_12461_[0]),
    .B(net3724),
    .C(net3721),
    .Y(_03073_));
 sky130_fd_sc_hd__nand3_1 _23797_ (.A(net3723),
    .B(_03070_),
    .C(_03073_),
    .Y(_03074_));
 sky130_fd_sc_hd__xor2_4 _23798_ (.A(\u0.tmp_w[4] ),
    .B(_03002_),
    .X(_03075_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__nor2_1 _23802_ (.A(_02981_),
    .B(net3719),
    .Y(_03079_));
 sky130_fd_sc_hd__nand2_8 _23803_ (.A(net3724),
    .B(_03012_),
    .Y(_03080_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_22 ();
 sky130_fd_sc_hd__o32ai_1 _23807_ (.A1(_02987_),
    .A2(net3724),
    .A3(_03079_),
    .B1(_03080_),
    .B2(_12465_[0]),
    .Y(_03084_));
 sky130_fd_sc_hd__nand2_1 _23808_ (.A(net3714),
    .B(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hd__xor2_4 _23809_ (.A(net4127),
    .B(_03046_),
    .X(_03086_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_20 ();
 sky130_fd_sc_hd__nor2_2 _23812_ (.A(net3712),
    .B(_03060_),
    .Y(_03089_));
 sky130_fd_sc_hd__o211ai_1 _23813_ (.A1(_03069_),
    .A2(_03074_),
    .B1(_03085_),
    .C1(_03089_),
    .Y(_03090_));
 sky130_fd_sc_hd__o21ai_0 _23814_ (.A1(_03036_),
    .A2(_03062_),
    .B1(_03090_),
    .Y(_03091_));
 sky130_fd_sc_hd__nor3_4 _23815_ (.A(net3727),
    .B(_02987_),
    .C(_02993_),
    .Y(_03092_));
 sky130_fd_sc_hd__nor2_4 _23816_ (.A(_12465_[0]),
    .B(net3724),
    .Y(_03093_));
 sky130_fd_sc_hd__o31ai_2 _23817_ (.A1(net3721),
    .A2(_03092_),
    .A3(_03093_),
    .B1(net3714),
    .Y(_03094_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_19 ();
 sky130_fd_sc_hd__nor2_4 _23819_ (.A(net3725),
    .B(_03017_),
    .Y(_03096_));
 sky130_fd_sc_hd__a21oi_1 _23820_ (.A1(_12462_[0]),
    .A2(_03017_),
    .B1(_03096_),
    .Y(_03097_));
 sky130_fd_sc_hd__o22ai_1 _23821_ (.A1(_12460_[0]),
    .A2(_03080_),
    .B1(_03097_),
    .B2(net3724),
    .Y(_03098_));
 sky130_fd_sc_hd__or2_4 _23822_ (.A(_03094_),
    .B(_03098_),
    .X(_03099_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_18 ();
 sky130_fd_sc_hd__xnor2_4 _23824_ (.A(\u0.tmp_w[7] ),
    .B(_03058_),
    .Y(_03101_));
 sky130_fd_sc_hd__nand2_8 _23825_ (.A(_03054_),
    .B(_03101_),
    .Y(_03102_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_17 ();
 sky130_fd_sc_hd__nor2_2 _23827_ (.A(net3724),
    .B(net3722),
    .Y(_03104_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_14 ();
 sky130_fd_sc_hd__a221oi_1 _23831_ (.A1(_12481_[0]),
    .A2(net3721),
    .B1(_03104_),
    .B2(_12461_[0]),
    .C1(net3714),
    .Y(_03108_));
 sky130_fd_sc_hd__nor3_1 _23832_ (.A(net3716),
    .B(_03102_),
    .C(_03108_),
    .Y(_03109_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__nor2_4 _23837_ (.A(_12462_[0]),
    .B(net3721),
    .Y(_03114_));
 sky130_fd_sc_hd__nor3_4 _23838_ (.A(net3727),
    .B(net3639),
    .C(net3720),
    .Y(_03115_));
 sky130_fd_sc_hd__nor3_1 _23839_ (.A(_02993_),
    .B(_03114_),
    .C(_03115_),
    .Y(_03116_));
 sky130_fd_sc_hd__a211oi_1 _23840_ (.A1(_12470_[0]),
    .A2(_03025_),
    .B1(_03116_),
    .C1(net3723),
    .Y(_03117_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__nand2_2 _23842_ (.A(_02993_),
    .B(_03017_),
    .Y(_03119_));
 sky130_fd_sc_hd__nor2_1 _23843_ (.A(_12468_[0]),
    .B(net3600),
    .Y(_03120_));
 sky130_fd_sc_hd__nand2_1 _23844_ (.A(_12462_[0]),
    .B(net3721),
    .Y(_03121_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__o21ai_0 _23846_ (.A1(net3727),
    .A2(net3639),
    .B1(net3720),
    .Y(_03123_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__a21oi_1 _23848_ (.A1(_03121_),
    .A2(_03123_),
    .B1(net3638),
    .Y(_03125_));
 sky130_fd_sc_hd__nor3_2 _23849_ (.A(_03075_),
    .B(_03120_),
    .C(_03125_),
    .Y(_03126_));
 sky130_fd_sc_hd__nor4_2 _23850_ (.A(net3712),
    .B(_03102_),
    .C(_03117_),
    .D(_03126_),
    .Y(_03127_));
 sky130_fd_sc_hd__a21oi_2 _23851_ (.A1(_03099_),
    .A2(_03109_),
    .B1(_03127_),
    .Y(_03128_));
 sky130_fd_sc_hd__nand2_2 _23852_ (.A(_12461_[0]),
    .B(_02993_),
    .Y(_03129_));
 sky130_fd_sc_hd__nand2_8 _23853_ (.A(_02981_),
    .B(net3724),
    .Y(_03130_));
 sky130_fd_sc_hd__a31oi_1 _23854_ (.A1(_03017_),
    .A2(_03129_),
    .A3(_03130_),
    .B1(net3723),
    .Y(_03131_));
 sky130_fd_sc_hd__nor2_1 _23855_ (.A(net3725),
    .B(_02993_),
    .Y(_03132_));
 sky130_fd_sc_hd__nor2_1 _23856_ (.A(_12468_[0]),
    .B(net3724),
    .Y(_03133_));
 sky130_fd_sc_hd__o21ai_0 _23857_ (.A1(net3599),
    .A2(_03133_),
    .B1(net3721),
    .Y(_03134_));
 sky130_fd_sc_hd__nand2_1 _23858_ (.A(_12460_[0]),
    .B(_03104_),
    .Y(_03135_));
 sky130_fd_sc_hd__nor2_4 _23859_ (.A(_12465_[0]),
    .B(net3719),
    .Y(_03136_));
 sky130_fd_sc_hd__o21ai_0 _23860_ (.A1(_03136_),
    .A2(_03114_),
    .B1(net3724),
    .Y(_03137_));
 sky130_fd_sc_hd__a21oi_1 _23861_ (.A1(_03135_),
    .A2(_03137_),
    .B1(net3714),
    .Y(_03138_));
 sky130_fd_sc_hd__a21oi_1 _23862_ (.A1(_03131_),
    .A2(_03134_),
    .B1(_03138_),
    .Y(_03139_));
 sky130_fd_sc_hd__a21oi_2 _23863_ (.A1(_02981_),
    .A2(_02987_),
    .B1(net3718),
    .Y(_03140_));
 sky130_fd_sc_hd__nor2_4 _23864_ (.A(_12465_[0]),
    .B(net3722),
    .Y(_03141_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__a211oi_1 _23866_ (.A1(net3725),
    .A2(_03025_),
    .B1(_03141_),
    .C1(net3723),
    .Y(_03143_));
 sky130_fd_sc_hd__o21ai_0 _23867_ (.A1(_02993_),
    .A2(_03140_),
    .B1(_03143_),
    .Y(_03144_));
 sky130_fd_sc_hd__nor2_2 _23868_ (.A(_12461_[0]),
    .B(_03017_),
    .Y(_03145_));
 sky130_fd_sc_hd__nor2_2 _23869_ (.A(_12470_[0]),
    .B(net3721),
    .Y(_03146_));
 sky130_fd_sc_hd__o21ai_0 _23870_ (.A1(_03145_),
    .A2(_03146_),
    .B1(net3724),
    .Y(_03147_));
 sky130_fd_sc_hd__o211ai_1 _23871_ (.A1(_12465_[0]),
    .A2(net3600),
    .B1(_03147_),
    .C1(net3723),
    .Y(_03148_));
 sky130_fd_sc_hd__nand2b_4 _23872_ (.A_N(_03054_),
    .B(_03101_),
    .Y(_03149_));
 sky130_fd_sc_hd__a31oi_1 _23873_ (.A1(net3712),
    .A2(_03144_),
    .A3(_03148_),
    .B1(_03149_),
    .Y(_03150_));
 sky130_fd_sc_hd__o21ai_2 _23874_ (.A1(net3712),
    .A2(_03139_),
    .B1(_03150_),
    .Y(_03151_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__a21oi_1 _23876_ (.A1(net3726),
    .A2(_03047_),
    .B1(net3638),
    .Y(_03153_));
 sky130_fd_sc_hd__nor2_4 _23877_ (.A(net3638),
    .B(_03047_),
    .Y(_03154_));
 sky130_fd_sc_hd__nor2_4 _23878_ (.A(net3726),
    .B(net3724),
    .Y(_03155_));
 sky130_fd_sc_hd__a22oi_1 _23879_ (.A1(net3629),
    .A2(_03154_),
    .B1(_03155_),
    .B2(_03047_),
    .Y(_03156_));
 sky130_fd_sc_hd__o21ai_1 _23880_ (.A1(net3727),
    .A2(_03153_),
    .B1(_03156_),
    .Y(_03157_));
 sky130_fd_sc_hd__o31ai_1 _23881_ (.A1(net3629),
    .A2(net3724),
    .A3(_03047_),
    .B1(net3721),
    .Y(_03158_));
 sky130_fd_sc_hd__nand2_1 _23882_ (.A(net3727),
    .B(net3726),
    .Y(_03159_));
 sky130_fd_sc_hd__a21oi_2 _23883_ (.A1(_03041_),
    .A2(_03159_),
    .B1(_03086_),
    .Y(_03160_));
 sky130_fd_sc_hd__o22ai_4 _23884_ (.A1(net3721),
    .A2(_03157_),
    .B1(_03158_),
    .B2(_03160_),
    .Y(_03161_));
 sky130_fd_sc_hd__nand2_8 _23885_ (.A(_02993_),
    .B(net3722),
    .Y(_03162_));
 sky130_fd_sc_hd__and2_0 _23886_ (.A(_03033_),
    .B(_03162_),
    .X(_03163_));
 sky130_fd_sc_hd__o221ai_1 _23887_ (.A1(_12468_[0]),
    .A2(net3600),
    .B1(_03163_),
    .B2(_12460_[0]),
    .C1(_03073_),
    .Y(_03164_));
 sky130_fd_sc_hd__a21oi_1 _23888_ (.A1(net3713),
    .A2(_03164_),
    .B1(net3723),
    .Y(_03165_));
 sky130_fd_sc_hd__nand2_4 _23889_ (.A(_12468_[0]),
    .B(net3721),
    .Y(_03166_));
 sky130_fd_sc_hd__o21ai_0 _23890_ (.A1(_12461_[0]),
    .A2(net3721),
    .B1(_03166_),
    .Y(_03167_));
 sky130_fd_sc_hd__nand3_4 _23891_ (.A(_02981_),
    .B(net3639),
    .C(_03017_),
    .Y(_03168_));
 sky130_fd_sc_hd__nand2_2 _23892_ (.A(_12460_[0]),
    .B(net3721),
    .Y(_03169_));
 sky130_fd_sc_hd__nand3_1 _23893_ (.A(_02993_),
    .B(_03168_),
    .C(_03169_),
    .Y(_03170_));
 sky130_fd_sc_hd__o21ai_0 _23894_ (.A1(_02993_),
    .A2(_03167_),
    .B1(_03170_),
    .Y(_03171_));
 sky130_fd_sc_hd__nand2_1 _23895_ (.A(net3715),
    .B(_03171_),
    .Y(_03172_));
 sky130_fd_sc_hd__nand2_8 _23896_ (.A(_03054_),
    .B(_03059_),
    .Y(_03173_));
 sky130_fd_sc_hd__a221o_1 _23897_ (.A1(net3723),
    .A2(_03161_),
    .B1(_03165_),
    .B2(_03172_),
    .C1(_03173_),
    .X(_03174_));
 sky130_fd_sc_hd__nand4b_1 _23898_ (.A_N(_03091_),
    .B(_03128_),
    .C(_03151_),
    .D(_03174_),
    .Y(_00152_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__o211ai_1 _23900_ (.A1(_12462_[0]),
    .A2(net3721),
    .B1(_03169_),
    .C1(net3724),
    .Y(_03176_));
 sky130_fd_sc_hd__inv_4 _23901_ (.A(_12461_[0]),
    .Y(_03177_));
 sky130_fd_sc_hd__nand2_8 _23902_ (.A(_03177_),
    .B(_03012_),
    .Y(_03178_));
 sky130_fd_sc_hd__nand2_4 _23903_ (.A(net3725),
    .B(_03017_),
    .Y(_03179_));
 sky130_fd_sc_hd__nand3_1 _23904_ (.A(_02993_),
    .B(_03178_),
    .C(_03179_),
    .Y(_03180_));
 sky130_fd_sc_hd__nand2_1 _23905_ (.A(_12465_[0]),
    .B(net3721),
    .Y(_03181_));
 sky130_fd_sc_hd__a21oi_1 _23906_ (.A1(net3637),
    .A2(_03181_),
    .B1(_02993_),
    .Y(_03182_));
 sky130_fd_sc_hd__nand2_4 _23907_ (.A(_02981_),
    .B(net3721),
    .Y(_03183_));
 sky130_fd_sc_hd__nand2b_1 _23908_ (.A_N(_12460_[0]),
    .B(_03017_),
    .Y(_03184_));
 sky130_fd_sc_hd__a21oi_1 _23909_ (.A1(_03183_),
    .A2(_03184_),
    .B1(net3724),
    .Y(_03185_));
 sky130_fd_sc_hd__nor3_1 _23910_ (.A(net3723),
    .B(_03182_),
    .C(_03185_),
    .Y(_03186_));
 sky130_fd_sc_hd__a31oi_1 _23911_ (.A1(net3723),
    .A2(_03176_),
    .A3(_03180_),
    .B1(_03186_),
    .Y(_03187_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__a21oi_1 _23913_ (.A1(net3590),
    .A2(net3719),
    .B1(_02993_),
    .Y(_03189_));
 sky130_fd_sc_hd__a21oi_1 _23914_ (.A1(_03178_),
    .A2(_03189_),
    .B1(net3714),
    .Y(_03190_));
 sky130_fd_sc_hd__nand2_8 _23915_ (.A(net3639),
    .B(net3721),
    .Y(_03191_));
 sky130_fd_sc_hd__nor2_2 _23916_ (.A(net3728),
    .B(_03191_),
    .Y(_03192_));
 sky130_fd_sc_hd__o21ai_0 _23917_ (.A1(_03114_),
    .A2(_03192_),
    .B1(_02993_),
    .Y(_03193_));
 sky130_fd_sc_hd__nand3_2 _23918_ (.A(net3725),
    .B(_02993_),
    .C(net3717),
    .Y(_03194_));
 sky130_fd_sc_hd__nand2_1 _23919_ (.A(net3714),
    .B(_03194_),
    .Y(_03195_));
 sky130_fd_sc_hd__a21oi_1 _23920_ (.A1(_03168_),
    .A2(_03178_),
    .B1(_02993_),
    .Y(_03196_));
 sky130_fd_sc_hd__o2bb2ai_1 _23921_ (.A1_N(_03190_),
    .A2_N(_03193_),
    .B1(_03195_),
    .B2(_03196_),
    .Y(_03197_));
 sky130_fd_sc_hd__a22oi_1 _23922_ (.A1(_03089_),
    .A2(_03187_),
    .B1(_03197_),
    .B2(_03061_),
    .Y(_03198_));
 sky130_fd_sc_hd__nor2_1 _23923_ (.A(net3639),
    .B(_02993_),
    .Y(_03199_));
 sky130_fd_sc_hd__a21oi_1 _23924_ (.A1(_12460_[0]),
    .A2(_02993_),
    .B1(_03199_),
    .Y(_03200_));
 sky130_fd_sc_hd__o32ai_1 _23925_ (.A1(_03155_),
    .A2(_03183_),
    .A3(_03199_),
    .B1(_03200_),
    .B2(net3721),
    .Y(_03201_));
 sky130_fd_sc_hd__a21oi_1 _23926_ (.A1(_03063_),
    .A2(_03183_),
    .B1(net3724),
    .Y(_03202_));
 sky130_fd_sc_hd__nor3_1 _23927_ (.A(net3715),
    .B(_03182_),
    .C(_03202_),
    .Y(_03203_));
 sky130_fd_sc_hd__a21oi_1 _23928_ (.A1(net3715),
    .A2(_03201_),
    .B1(_03203_),
    .Y(_03204_));
 sky130_fd_sc_hd__nand2_2 _23929_ (.A(_12468_[0]),
    .B(net3638),
    .Y(_03205_));
 sky130_fd_sc_hd__nor2_4 _23930_ (.A(net3727),
    .B(net3726),
    .Y(_03206_));
 sky130_fd_sc_hd__nand2_1 _23931_ (.A(net3724),
    .B(_03206_),
    .Y(_03207_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__nor3_1 _23933_ (.A(_12484_[0]),
    .B(_03047_),
    .C(net3720),
    .Y(_03209_));
 sky130_fd_sc_hd__a31oi_2 _23934_ (.A1(net3720),
    .A2(_03205_),
    .A3(_03207_),
    .B1(_03209_),
    .Y(_03210_));
 sky130_fd_sc_hd__a21oi_1 _23935_ (.A1(_03075_),
    .A2(_03210_),
    .B1(_03173_),
    .Y(_03211_));
 sky130_fd_sc_hd__o21ai_2 _23936_ (.A1(_03075_),
    .A2(_03204_),
    .B1(_03211_),
    .Y(_03212_));
 sky130_fd_sc_hd__nand2_1 _23937_ (.A(_12465_[0]),
    .B(net3718),
    .Y(_03213_));
 sky130_fd_sc_hd__nand3_1 _23938_ (.A(net3724),
    .B(_03178_),
    .C(_03213_),
    .Y(_03214_));
 sky130_fd_sc_hd__o211ai_1 _23939_ (.A1(net3724),
    .A2(_03140_),
    .B1(_03214_),
    .C1(net3714),
    .Y(_03215_));
 sky130_fd_sc_hd__nand2_1 _23940_ (.A(_12474_[0]),
    .B(_02993_),
    .Y(_03216_));
 sky130_fd_sc_hd__a21oi_1 _23941_ (.A1(_03130_),
    .A2(_03216_),
    .B1(net3718),
    .Y(_03217_));
 sky130_fd_sc_hd__nor2_1 _23942_ (.A(_12465_[0]),
    .B(net3723),
    .Y(_03218_));
 sky130_fd_sc_hd__nor3_1 _23943_ (.A(_03206_),
    .B(_03033_),
    .C(_03218_),
    .Y(_03219_));
 sky130_fd_sc_hd__a21oi_1 _23944_ (.A1(net3723),
    .A2(_03217_),
    .B1(_03219_),
    .Y(_03220_));
 sky130_fd_sc_hd__nand3_1 _23945_ (.A(net3716),
    .B(_03215_),
    .C(_03220_),
    .Y(_03221_));
 sky130_fd_sc_hd__xnor2_1 _23946_ (.A(_02993_),
    .B(_03012_),
    .Y(_03222_));
 sky130_fd_sc_hd__a222oi_1 _23947_ (.A1(_12461_[0]),
    .A2(_03104_),
    .B1(_03222_),
    .B2(net3725),
    .C1(_03096_),
    .C2(net3728),
    .Y(_03223_));
 sky130_fd_sc_hd__nand2_1 _23948_ (.A(net3714),
    .B(_03223_),
    .Y(_03224_));
 sky130_fd_sc_hd__nor3_1 _23949_ (.A(_03177_),
    .B(_03009_),
    .C(_03011_),
    .Y(_03225_));
 sky130_fd_sc_hd__and2_4 _23950_ (.A(_12460_[0]),
    .B(_03017_),
    .X(_03226_));
 sky130_fd_sc_hd__o21ai_1 _23951_ (.A1(net3575),
    .A2(_03226_),
    .B1(net3724),
    .Y(_03227_));
 sky130_fd_sc_hd__nor2_4 _23952_ (.A(_02987_),
    .B(net3721),
    .Y(_03228_));
 sky130_fd_sc_hd__o21ai_0 _23953_ (.A1(_03136_),
    .A2(_03228_),
    .B1(_02993_),
    .Y(_03229_));
 sky130_fd_sc_hd__nand3_1 _23954_ (.A(net3723),
    .B(_03227_),
    .C(_03229_),
    .Y(_03230_));
 sky130_fd_sc_hd__a31oi_1 _23955_ (.A1(net3712),
    .A2(_03224_),
    .A3(_03230_),
    .B1(_03149_),
    .Y(_03231_));
 sky130_fd_sc_hd__nand2_1 _23956_ (.A(_12474_[0]),
    .B(net3724),
    .Y(_03232_));
 sky130_fd_sc_hd__a21oi_1 _23957_ (.A1(_03129_),
    .A2(_03232_),
    .B1(net3718),
    .Y(_03233_));
 sky130_fd_sc_hd__a2bb2oi_1 _23958_ (.A1_N(_12465_[0]),
    .A2_N(net3600),
    .B1(_03222_),
    .B2(_02981_),
    .Y(_03234_));
 sky130_fd_sc_hd__o22ai_1 _23959_ (.A1(_03094_),
    .A2(_03233_),
    .B1(_03234_),
    .B2(net3714),
    .Y(_03235_));
 sky130_fd_sc_hd__a21oi_1 _23960_ (.A1(_03070_),
    .A2(_03162_),
    .B1(_02981_),
    .Y(_03236_));
 sky130_fd_sc_hd__o21ai_1 _23961_ (.A1(_03155_),
    .A2(_03236_),
    .B1(net3714),
    .Y(_03237_));
 sky130_fd_sc_hd__nor2_1 _23962_ (.A(_02981_),
    .B(net3723),
    .Y(_03238_));
 sky130_fd_sc_hd__o21ai_0 _23963_ (.A1(_03179_),
    .A2(_03238_),
    .B1(_03191_),
    .Y(_03239_));
 sky130_fd_sc_hd__a21oi_1 _23964_ (.A1(_12465_[0]),
    .A2(net3717),
    .B1(net3575),
    .Y(_03240_));
 sky130_fd_sc_hd__o31ai_1 _23965_ (.A1(_02993_),
    .A2(net3714),
    .A3(_03240_),
    .B1(net3716),
    .Y(_03241_));
 sky130_fd_sc_hd__a21oi_1 _23966_ (.A1(_02993_),
    .A2(_03239_),
    .B1(_03241_),
    .Y(_03242_));
 sky130_fd_sc_hd__a221oi_1 _23967_ (.A1(net3712),
    .A2(_03235_),
    .B1(_03237_),
    .B2(_03242_),
    .C1(_03102_),
    .Y(_03243_));
 sky130_fd_sc_hd__a21oi_2 _23968_ (.A1(_03221_),
    .A2(_03231_),
    .B1(_03243_),
    .Y(_03244_));
 sky130_fd_sc_hd__nand3_1 _23969_ (.A(_03198_),
    .B(_03212_),
    .C(_03244_),
    .Y(_00153_));
 sky130_fd_sc_hd__nor2_2 _23970_ (.A(_12462_[0]),
    .B(_12465_[0]),
    .Y(_03245_));
 sky130_fd_sc_hd__nand2_2 _23971_ (.A(net3721),
    .B(_03245_),
    .Y(_03246_));
 sky130_fd_sc_hd__a211oi_1 _23972_ (.A1(_12468_[0]),
    .A2(_03017_),
    .B1(_03192_),
    .C1(net3724),
    .Y(_03247_));
 sky130_fd_sc_hd__a311o_1 _23973_ (.A1(net3724),
    .A2(_03168_),
    .A3(_03246_),
    .B1(_03247_),
    .C1(_03075_),
    .X(_03248_));
 sky130_fd_sc_hd__nand2_1 _23974_ (.A(_12465_[0]),
    .B(_03025_),
    .Y(_03249_));
 sky130_fd_sc_hd__o311ai_0 _23975_ (.A1(_02993_),
    .A2(_03145_),
    .A3(_03226_),
    .B1(_03249_),
    .C1(_03075_),
    .Y(_03250_));
 sky130_fd_sc_hd__o32a_1 _23976_ (.A1(_02981_),
    .A2(_03017_),
    .A3(net3599),
    .B1(_03130_),
    .B2(_03096_),
    .X(_03251_));
 sky130_fd_sc_hd__nor2_1 _23977_ (.A(_02981_),
    .B(net3724),
    .Y(_03252_));
 sky130_fd_sc_hd__o21ai_0 _23978_ (.A1(_03028_),
    .A2(_03252_),
    .B1(_12461_[0]),
    .Y(_03253_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__a21oi_1 _23980_ (.A1(_03251_),
    .A2(_03253_),
    .B1(net3714),
    .Y(_03255_));
 sky130_fd_sc_hd__nor2_4 _23981_ (.A(_12461_[0]),
    .B(net3724),
    .Y(_03256_));
 sky130_fd_sc_hd__nor3_1 _23982_ (.A(_03017_),
    .B(_03092_),
    .C(_03256_),
    .Y(_03257_));
 sky130_fd_sc_hd__a211oi_1 _23983_ (.A1(_12481_[0]),
    .A2(_03017_),
    .B1(_03257_),
    .C1(net3723),
    .Y(_03258_));
 sky130_fd_sc_hd__nor2_1 _23984_ (.A(_03059_),
    .B(net3712),
    .Y(_03259_));
 sky130_fd_sc_hd__o31ai_1 _23985_ (.A1(_03054_),
    .A2(_03255_),
    .A3(_03258_),
    .B1(_03259_),
    .Y(_03260_));
 sky130_fd_sc_hd__a31oi_1 _23986_ (.A1(_03054_),
    .A2(_03248_),
    .A3(_03250_),
    .B1(_03260_),
    .Y(_03261_));
 sky130_fd_sc_hd__mux2i_1 _23987_ (.A0(_12474_[0]),
    .A1(_12465_[0]),
    .S(net3724),
    .Y(_03262_));
 sky130_fd_sc_hd__nand2_2 _23988_ (.A(_03017_),
    .B(_03262_),
    .Y(_03263_));
 sky130_fd_sc_hd__nand2_1 _23989_ (.A(net3639),
    .B(net3638),
    .Y(_03264_));
 sky130_fd_sc_hd__nor2_4 _23990_ (.A(net3727),
    .B(_03017_),
    .Y(_03265_));
 sky130_fd_sc_hd__nand2_2 _23991_ (.A(_03264_),
    .B(_03265_),
    .Y(_03266_));
 sky130_fd_sc_hd__o21ai_2 _23992_ (.A1(_03092_),
    .A2(_03093_),
    .B1(net3721),
    .Y(_03267_));
 sky130_fd_sc_hd__a32oi_1 _23993_ (.A1(net3723),
    .A2(_03263_),
    .A3(_03266_),
    .B1(_03131_),
    .B2(_03267_),
    .Y(_03268_));
 sky130_fd_sc_hd__nor2_1 _23994_ (.A(net3716),
    .B(_03268_),
    .Y(_03269_));
 sky130_fd_sc_hd__nand2_8 _23995_ (.A(net3629),
    .B(net3720),
    .Y(_03270_));
 sky130_fd_sc_hd__a21oi_1 _23996_ (.A1(_03270_),
    .A2(_03191_),
    .B1(_02993_),
    .Y(_03271_));
 sky130_fd_sc_hd__nor2_1 _23997_ (.A(_12462_[0]),
    .B(_03017_),
    .Y(_03272_));
 sky130_fd_sc_hd__nor3_1 _23998_ (.A(net3724),
    .B(_03028_),
    .C(_03272_),
    .Y(_03273_));
 sky130_fd_sc_hd__nor2_1 _23999_ (.A(net3590),
    .B(_03080_),
    .Y(_03274_));
 sky130_fd_sc_hd__nand2_4 _24000_ (.A(_02981_),
    .B(_02993_),
    .Y(_03275_));
 sky130_fd_sc_hd__a21oi_1 _24001_ (.A1(_03191_),
    .A2(net3637),
    .B1(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__o21ai_0 _24002_ (.A1(_03274_),
    .A2(_03276_),
    .B1(net3714),
    .Y(_03277_));
 sky130_fd_sc_hd__o311a_1 _24003_ (.A1(net3714),
    .A2(_03271_),
    .A3(_03273_),
    .B1(_03277_),
    .C1(net3716),
    .X(_03278_));
 sky130_fd_sc_hd__nor3_1 _24004_ (.A(_03173_),
    .B(_03269_),
    .C(_03278_),
    .Y(_03279_));
 sky130_fd_sc_hd__a21oi_1 _24005_ (.A1(_12470_[0]),
    .A2(_03017_),
    .B1(_03145_),
    .Y(_03280_));
 sky130_fd_sc_hd__nand3_1 _24006_ (.A(net3724),
    .B(_03178_),
    .C(net3637),
    .Y(_03281_));
 sky130_fd_sc_hd__o21ai_0 _24007_ (.A1(net3724),
    .A2(_03280_),
    .B1(_03281_),
    .Y(_03282_));
 sky130_fd_sc_hd__nand2_8 _24008_ (.A(_12470_[0]),
    .B(net3721),
    .Y(_03283_));
 sky130_fd_sc_hd__nand2b_4 _24009_ (.A_N(_12474_[0]),
    .B(_03017_),
    .Y(_03284_));
 sky130_fd_sc_hd__a21oi_1 _24010_ (.A1(_03183_),
    .A2(_03284_),
    .B1(net3724),
    .Y(_03285_));
 sky130_fd_sc_hd__a311oi_1 _24011_ (.A1(net3724),
    .A2(_03070_),
    .A3(_03283_),
    .B1(_03285_),
    .C1(_03075_),
    .Y(_03286_));
 sky130_fd_sc_hd__a21oi_1 _24012_ (.A1(_03075_),
    .A2(_03282_),
    .B1(_03286_),
    .Y(_03287_));
 sky130_fd_sc_hd__a21oi_1 _24013_ (.A1(_12470_[0]),
    .A2(_03017_),
    .B1(_02993_),
    .Y(_03288_));
 sky130_fd_sc_hd__a2111oi_0 _24014_ (.A1(_03183_),
    .A2(_03288_),
    .B1(net3723),
    .C1(net3716),
    .D1(_03093_),
    .Y(_03289_));
 sky130_fd_sc_hd__nor2_1 _24015_ (.A(_03060_),
    .B(_03289_),
    .Y(_03290_));
 sky130_fd_sc_hd__nor3_1 _24016_ (.A(_02993_),
    .B(_03027_),
    .C(_03146_),
    .Y(_03291_));
 sky130_fd_sc_hd__nor2_2 _24017_ (.A(net3590),
    .B(net3721),
    .Y(_03292_));
 sky130_fd_sc_hd__nor3_1 _24018_ (.A(net3724),
    .B(_03136_),
    .C(_03292_),
    .Y(_03293_));
 sky130_fd_sc_hd__o211ai_1 _24019_ (.A1(_03291_),
    .A2(_03293_),
    .B1(net3723),
    .C1(net3712),
    .Y(_03294_));
 sky130_fd_sc_hd__o211a_1 _24020_ (.A1(net3712),
    .A2(_03287_),
    .B1(_03290_),
    .C1(_03294_),
    .X(_03295_));
 sky130_fd_sc_hd__o21ai_0 _24021_ (.A1(_12488_[0]),
    .A2(net3721),
    .B1(_03266_),
    .Y(_03296_));
 sky130_fd_sc_hd__a21oi_1 _24022_ (.A1(_12479_[0]),
    .A2(net3721),
    .B1(net3723),
    .Y(_03297_));
 sky130_fd_sc_hd__o41ai_1 _24023_ (.A1(net3727),
    .A2(net3639),
    .A3(net3724),
    .A4(net3721),
    .B1(_03297_),
    .Y(_03298_));
 sky130_fd_sc_hd__o21ai_0 _24024_ (.A1(_03075_),
    .A2(_03296_),
    .B1(_03298_),
    .Y(_03299_));
 sky130_fd_sc_hd__nor3_1 _24025_ (.A(net3724),
    .B(_03145_),
    .C(_03226_),
    .Y(_03300_));
 sky130_fd_sc_hd__a311oi_1 _24026_ (.A1(net3724),
    .A2(_03166_),
    .A3(_03063_),
    .B1(_03300_),
    .C1(_03075_),
    .Y(_03301_));
 sky130_fd_sc_hd__o21ai_0 _24027_ (.A1(_12484_[0]),
    .A2(net3721),
    .B1(_03075_),
    .Y(_03302_));
 sky130_fd_sc_hd__a31oi_1 _24028_ (.A1(net3721),
    .A2(_03159_),
    .A3(_03130_),
    .B1(_03302_),
    .Y(_03303_));
 sky130_fd_sc_hd__nor3_1 _24029_ (.A(_03054_),
    .B(_03301_),
    .C(_03303_),
    .Y(_03304_));
 sky130_fd_sc_hd__a2111oi_0 _24030_ (.A1(_03054_),
    .A2(_03299_),
    .B1(_03304_),
    .C1(net3716),
    .D1(_03059_),
    .Y(_03305_));
 sky130_fd_sc_hd__nor4_1 _24031_ (.A(_03261_),
    .B(_03279_),
    .C(_03295_),
    .D(_03305_),
    .Y(_00154_));
 sky130_fd_sc_hd__nor2_2 _24032_ (.A(_12470_[0]),
    .B(_03017_),
    .Y(_03306_));
 sky130_fd_sc_hd__a211oi_2 _24033_ (.A1(_12468_[0]),
    .A2(_03017_),
    .B1(_03306_),
    .C1(net3724),
    .Y(_03307_));
 sky130_fd_sc_hd__a31oi_1 _24034_ (.A1(net3724),
    .A2(_03168_),
    .A3(_03246_),
    .B1(_03307_),
    .Y(_03308_));
 sky130_fd_sc_hd__o22ai_1 _24035_ (.A1(_12460_[0]),
    .A2(_03080_),
    .B1(net3600),
    .B2(net3727),
    .Y(_03309_));
 sky130_fd_sc_hd__a21oi_1 _24036_ (.A1(net3724),
    .A2(_03063_),
    .B1(net3726),
    .Y(_03310_));
 sky130_fd_sc_hd__o21ai_0 _24037_ (.A1(_03309_),
    .A2(_03310_),
    .B1(net3715),
    .Y(_03311_));
 sky130_fd_sc_hd__o21ai_0 _24038_ (.A1(net3715),
    .A2(_03308_),
    .B1(_03311_),
    .Y(_03312_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__nor2_2 _24040_ (.A(_03047_),
    .B(net3721),
    .Y(_03314_));
 sky130_fd_sc_hd__a32oi_1 _24041_ (.A1(net3716),
    .A2(_03270_),
    .A3(_03283_),
    .B1(_03314_),
    .B2(net3726),
    .Y(_03315_));
 sky130_fd_sc_hd__a311oi_1 _24042_ (.A1(net3639),
    .A2(net3716),
    .A3(net3721),
    .B1(_03292_),
    .C1(net3724),
    .Y(_03316_));
 sky130_fd_sc_hd__a21oi_2 _24043_ (.A1(net3724),
    .A2(_03315_),
    .B1(_03316_),
    .Y(_03317_));
 sky130_fd_sc_hd__a21oi_1 _24044_ (.A1(net3723),
    .A2(_03317_),
    .B1(_03060_),
    .Y(_03318_));
 sky130_fd_sc_hd__o21ai_0 _24045_ (.A1(net3723),
    .A2(_03312_),
    .B1(_03318_),
    .Y(_03319_));
 sky130_fd_sc_hd__a21oi_1 _24046_ (.A1(_12461_[0]),
    .A2(_03017_),
    .B1(_03021_),
    .Y(_03320_));
 sky130_fd_sc_hd__nor3_1 _24047_ (.A(net3724),
    .B(_03016_),
    .C(_03136_),
    .Y(_03321_));
 sky130_fd_sc_hd__a21oi_1 _24048_ (.A1(net3724),
    .A2(_03320_),
    .B1(_03321_),
    .Y(_03322_));
 sky130_fd_sc_hd__o221ai_1 _24049_ (.A1(net3599),
    .A2(_03063_),
    .B1(_03228_),
    .B2(_03275_),
    .C1(_03073_),
    .Y(_03323_));
 sky130_fd_sc_hd__nor2_1 _24050_ (.A(net3715),
    .B(_03323_),
    .Y(_03324_));
 sky130_fd_sc_hd__a21oi_1 _24051_ (.A1(net3715),
    .A2(_03322_),
    .B1(_03324_),
    .Y(_03325_));
 sky130_fd_sc_hd__nor2_2 _24052_ (.A(net3724),
    .B(net3713),
    .Y(_03326_));
 sky130_fd_sc_hd__o21ai_0 _24053_ (.A1(_03154_),
    .A2(_03326_),
    .B1(net3726),
    .Y(_03327_));
 sky130_fd_sc_hd__nand3_1 _24054_ (.A(_12468_[0]),
    .B(net3724),
    .C(_03047_),
    .Y(_03328_));
 sky130_fd_sc_hd__nor2_1 _24055_ (.A(net3724),
    .B(_03047_),
    .Y(_03329_));
 sky130_fd_sc_hd__nand2_1 _24056_ (.A(net3727),
    .B(_03329_),
    .Y(_03330_));
 sky130_fd_sc_hd__nand4_1 _24057_ (.A(net3720),
    .B(_03327_),
    .C(_03328_),
    .D(_03330_),
    .Y(_03331_));
 sky130_fd_sc_hd__xnor2_1 _24058_ (.A(net3629),
    .B(net3712),
    .Y(_03332_));
 sky130_fd_sc_hd__nand3_1 _24059_ (.A(_12460_[0]),
    .B(net3724),
    .C(net3716),
    .Y(_03333_));
 sky130_fd_sc_hd__o211ai_1 _24060_ (.A1(net3724),
    .A2(_03332_),
    .B1(_03333_),
    .C1(net3721),
    .Y(_03334_));
 sky130_fd_sc_hd__a31oi_1 _24061_ (.A1(net3723),
    .A2(_03331_),
    .A3(_03334_),
    .B1(_03102_),
    .Y(_03335_));
 sky130_fd_sc_hd__o21ai_0 _24062_ (.A1(net3723),
    .A2(_03325_),
    .B1(_03335_),
    .Y(_03336_));
 sky130_fd_sc_hd__nor2_4 _24063_ (.A(_03054_),
    .B(_03059_),
    .Y(_03337_));
 sky130_fd_sc_hd__a211oi_1 _24064_ (.A1(_12470_[0]),
    .A2(_03017_),
    .B1(_03047_),
    .C1(net3724),
    .Y(_03338_));
 sky130_fd_sc_hd__nand2_1 _24065_ (.A(net3727),
    .B(net3721),
    .Y(_03339_));
 sky130_fd_sc_hd__a21boi_0 _24066_ (.A1(_03270_),
    .A2(_03339_),
    .B1_N(_03154_),
    .Y(_03340_));
 sky130_fd_sc_hd__nand2b_1 _24067_ (.A_N(_12468_[0]),
    .B(net3720),
    .Y(_03341_));
 sky130_fd_sc_hd__a21oi_1 _24068_ (.A1(_03191_),
    .A2(_03341_),
    .B1(net3724),
    .Y(_03342_));
 sky130_fd_sc_hd__nor2_1 _24069_ (.A(net3629),
    .B(_03033_),
    .Y(_03343_));
 sky130_fd_sc_hd__nor4_1 _24070_ (.A(net3713),
    .B(_03115_),
    .C(_03342_),
    .D(_03343_),
    .Y(_03344_));
 sky130_fd_sc_hd__a2111oi_0 _24071_ (.A1(_03066_),
    .A2(_03338_),
    .B1(_03340_),
    .C1(_03344_),
    .D1(_03075_),
    .Y(_03345_));
 sky130_fd_sc_hd__nor2_2 _24072_ (.A(_03086_),
    .B(net3721),
    .Y(_03346_));
 sky130_fd_sc_hd__nand3_1 _24073_ (.A(_02981_),
    .B(_03080_),
    .C(_03264_),
    .Y(_03347_));
 sky130_fd_sc_hd__a21oi_1 _24074_ (.A1(net3716),
    .A2(_03228_),
    .B1(_03347_),
    .Y(_03348_));
 sky130_fd_sc_hd__nand3_1 _24075_ (.A(_12468_[0]),
    .B(_03047_),
    .C(net3721),
    .Y(_03349_));
 sky130_fd_sc_hd__nand2_1 _24076_ (.A(net3639),
    .B(_03314_),
    .Y(_03350_));
 sky130_fd_sc_hd__a21oi_2 _24077_ (.A1(_03349_),
    .A2(_03350_),
    .B1(net3638),
    .Y(_03351_));
 sky130_fd_sc_hd__nand2_1 _24078_ (.A(_03075_),
    .B(_03337_),
    .Y(_03352_));
 sky130_fd_sc_hd__a2111oi_2 _24079_ (.A1(_03256_),
    .A2(_03346_),
    .B1(_03348_),
    .C1(_03351_),
    .D1(_03352_),
    .Y(_03353_));
 sky130_fd_sc_hd__a21oi_1 _24080_ (.A1(_03337_),
    .A2(_03345_),
    .B1(_03353_),
    .Y(_03354_));
 sky130_fd_sc_hd__o211ai_1 _24081_ (.A1(net3629),
    .A2(net3721),
    .B1(_03246_),
    .C1(net3724),
    .Y(_03355_));
 sky130_fd_sc_hd__o311ai_0 _24082_ (.A1(net3724),
    .A2(_03021_),
    .A3(_03228_),
    .B1(_03355_),
    .C1(net3713),
    .Y(_03356_));
 sky130_fd_sc_hd__a221oi_1 _24083_ (.A1(_12470_[0]),
    .A2(_03163_),
    .B1(net3599),
    .B2(_03017_),
    .C1(net3713),
    .Y(_03357_));
 sky130_fd_sc_hd__nor3_1 _24084_ (.A(_03173_),
    .B(net3723),
    .C(_03357_),
    .Y(_03358_));
 sky130_fd_sc_hd__nor2_4 _24085_ (.A(_02981_),
    .B(_03033_),
    .Y(_03359_));
 sky130_fd_sc_hd__nand2_1 _24086_ (.A(_03178_),
    .B(_03341_),
    .Y(_03360_));
 sky130_fd_sc_hd__o31ai_1 _24087_ (.A1(net3629),
    .A2(_03086_),
    .A3(net3721),
    .B1(_03121_),
    .Y(_03361_));
 sky130_fd_sc_hd__a222oi_1 _24088_ (.A1(_03086_),
    .A2(_03359_),
    .B1(_03360_),
    .B2(_03329_),
    .C1(_03361_),
    .C2(net3724),
    .Y(_03362_));
 sky130_fd_sc_hd__nor3_1 _24089_ (.A(_03173_),
    .B(_03075_),
    .C(_03362_),
    .Y(_03363_));
 sky130_fd_sc_hd__a21oi_1 _24090_ (.A1(_03356_),
    .A2(_03358_),
    .B1(_03363_),
    .Y(_03364_));
 sky130_fd_sc_hd__nand4_1 _24091_ (.A(_03319_),
    .B(_03336_),
    .C(_03354_),
    .D(_03364_),
    .Y(_00155_));
 sky130_fd_sc_hd__nor2_2 _24092_ (.A(_03003_),
    .B(_03086_),
    .Y(_03365_));
 sky130_fd_sc_hd__o21ai_0 _24093_ (.A1(_03115_),
    .A2(_03292_),
    .B1(net3724),
    .Y(_03366_));
 sky130_fd_sc_hd__nand3_1 _24094_ (.A(_02993_),
    .B(_03270_),
    .C(_03283_),
    .Y(_03367_));
 sky130_fd_sc_hd__a31oi_1 _24095_ (.A1(_03365_),
    .A2(_03366_),
    .A3(_03367_),
    .B1(_03102_),
    .Y(_03368_));
 sky130_fd_sc_hd__nand2_1 _24096_ (.A(_12470_[0]),
    .B(net3724),
    .Y(_03369_));
 sky130_fd_sc_hd__o21ai_0 _24097_ (.A1(net3724),
    .A2(_03240_),
    .B1(_03369_),
    .Y(_03370_));
 sky130_fd_sc_hd__nor2_4 _24098_ (.A(_03075_),
    .B(_03086_),
    .Y(_03371_));
 sky130_fd_sc_hd__nor2_2 _24099_ (.A(net3728),
    .B(_03179_),
    .Y(_03372_));
 sky130_fd_sc_hd__nand2_1 _24100_ (.A(net3724),
    .B(_03169_),
    .Y(_03373_));
 sky130_fd_sc_hd__o32a_1 _24101_ (.A1(net3724),
    .A2(_03079_),
    .A3(_03141_),
    .B1(_03372_),
    .B2(_03373_),
    .X(_03374_));
 sky130_fd_sc_hd__o21ai_0 _24102_ (.A1(_03092_),
    .A2(_03252_),
    .B1(net3721),
    .Y(_03375_));
 sky130_fd_sc_hd__a21oi_1 _24103_ (.A1(_03263_),
    .A2(_03375_),
    .B1(net3714),
    .Y(_03376_));
 sky130_fd_sc_hd__a211oi_1 _24104_ (.A1(net3714),
    .A2(_03374_),
    .B1(_03376_),
    .C1(net3716),
    .Y(_03377_));
 sky130_fd_sc_hd__a21oi_1 _24105_ (.A1(_03370_),
    .A2(_03371_),
    .B1(_03377_),
    .Y(_03378_));
 sky130_fd_sc_hd__o211ai_1 _24106_ (.A1(_02993_),
    .A2(_03114_),
    .B1(_03283_),
    .C1(net3723),
    .Y(_03379_));
 sky130_fd_sc_hd__o311ai_0 _24107_ (.A1(net3724),
    .A2(_03265_),
    .A3(_03226_),
    .B1(net3714),
    .C1(_03041_),
    .Y(_03380_));
 sky130_fd_sc_hd__nand3_1 _24108_ (.A(net3716),
    .B(_03379_),
    .C(_03380_),
    .Y(_03381_));
 sky130_fd_sc_hd__nand2_1 _24109_ (.A(_02993_),
    .B(net3714),
    .Y(_03382_));
 sky130_fd_sc_hd__a21oi_1 _24110_ (.A1(net3725),
    .A2(_03382_),
    .B1(net3728),
    .Y(_03383_));
 sky130_fd_sc_hd__nor3_1 _24111_ (.A(net3722),
    .B(_03132_),
    .C(_03383_),
    .Y(_03384_));
 sky130_fd_sc_hd__nor2_1 _24112_ (.A(net3723),
    .B(_03130_),
    .Y(_03385_));
 sky130_fd_sc_hd__a311oi_1 _24113_ (.A1(_12460_[0]),
    .A2(_02993_),
    .A3(net3723),
    .B1(_03017_),
    .C1(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__nor2_1 _24114_ (.A(_02993_),
    .B(net3714),
    .Y(_03387_));
 sky130_fd_sc_hd__a21oi_1 _24115_ (.A1(net3714),
    .A2(_03027_),
    .B1(_03387_),
    .Y(_03388_));
 sky130_fd_sc_hd__o221ai_1 _24116_ (.A1(_03384_),
    .A2(_03386_),
    .B1(_03388_),
    .B2(_02981_),
    .C1(net3712),
    .Y(_03389_));
 sky130_fd_sc_hd__o21a_4 _24117_ (.A1(_03096_),
    .A2(_03226_),
    .B1(_02993_),
    .X(_03390_));
 sky130_fd_sc_hd__nand2_1 _24118_ (.A(_12472_[0]),
    .B(_03017_),
    .Y(_03391_));
 sky130_fd_sc_hd__o211ai_1 _24119_ (.A1(_03017_),
    .A2(_03129_),
    .B1(_03391_),
    .C1(net3716),
    .Y(_03392_));
 sky130_fd_sc_hd__o41ai_1 _24120_ (.A1(net3716),
    .A2(_03034_),
    .A3(_03115_),
    .A4(_03390_),
    .B1(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__o21ai_1 _24121_ (.A1(_03306_),
    .A2(_03346_),
    .B1(net3638),
    .Y(_03394_));
 sky130_fd_sc_hd__nand3_1 _24122_ (.A(net3724),
    .B(_03047_),
    .C(net3722),
    .Y(_03395_));
 sky130_fd_sc_hd__a21oi_1 _24123_ (.A1(_03119_),
    .A2(_03395_),
    .B1(_02981_),
    .Y(_03396_));
 sky130_fd_sc_hd__a2111oi_0 _24124_ (.A1(_03154_),
    .A2(_03096_),
    .B1(_03396_),
    .C1(_03372_),
    .D1(net3714),
    .Y(_03397_));
 sky130_fd_sc_hd__a221oi_1 _24125_ (.A1(net3714),
    .A2(_03393_),
    .B1(_03394_),
    .B2(_03397_),
    .C1(_03173_),
    .Y(_03398_));
 sky130_fd_sc_hd__a31o_1 _24126_ (.A1(_03337_),
    .A2(_03381_),
    .A3(_03389_),
    .B1(_03398_),
    .X(_03399_));
 sky130_fd_sc_hd__nand3b_1 _24127_ (.A_N(_03027_),
    .B(_02993_),
    .C(_03270_),
    .Y(_03400_));
 sky130_fd_sc_hd__o311ai_0 _24128_ (.A1(_02993_),
    .A2(_03141_),
    .A3(_03192_),
    .B1(_03400_),
    .C1(net3715),
    .Y(_03401_));
 sky130_fd_sc_hd__o22ai_1 _24129_ (.A1(net3590),
    .A2(net3600),
    .B1(_03228_),
    .B2(_02993_),
    .Y(_03402_));
 sky130_fd_sc_hd__a21oi_1 _24130_ (.A1(net3712),
    .A2(_03402_),
    .B1(net3723),
    .Y(_03403_));
 sky130_fd_sc_hd__nor3_1 _24131_ (.A(_02993_),
    .B(_03136_),
    .C(_03226_),
    .Y(_03404_));
 sky130_fd_sc_hd__o21ai_0 _24132_ (.A1(_03114_),
    .A2(_03192_),
    .B1(_03326_),
    .Y(_03405_));
 sky130_fd_sc_hd__o311a_4 _24133_ (.A1(net3715),
    .A2(_03202_),
    .A3(_03404_),
    .B1(_03405_),
    .C1(net3723),
    .X(_03406_));
 sky130_fd_sc_hd__a211oi_2 _24134_ (.A1(_03401_),
    .A2(_03403_),
    .B1(_03406_),
    .C1(_03060_),
    .Y(_03407_));
 sky130_fd_sc_hd__a211oi_2 _24135_ (.A1(_03368_),
    .A2(_03378_),
    .B1(_03399_),
    .C1(_03407_),
    .Y(_00156_));
 sky130_fd_sc_hd__inv_1 _24136_ (.A(_12470_[0]),
    .Y(_03408_));
 sky130_fd_sc_hd__o211ai_1 _24137_ (.A1(_03408_),
    .A2(net3600),
    .B1(_03181_),
    .C1(net3715),
    .Y(_03409_));
 sky130_fd_sc_hd__a21oi_1 _24138_ (.A1(_12465_[0]),
    .A2(net3720),
    .B1(net3638),
    .Y(_03410_));
 sky130_fd_sc_hd__o21ai_0 _24139_ (.A1(_03115_),
    .A2(_03410_),
    .B1(_03086_),
    .Y(_03411_));
 sky130_fd_sc_hd__o21ai_0 _24140_ (.A1(_03125_),
    .A2(_03409_),
    .B1(_03411_),
    .Y(_03412_));
 sky130_fd_sc_hd__a31oi_1 _24141_ (.A1(_03101_),
    .A2(net3723),
    .A3(_03412_),
    .B1(_03054_),
    .Y(_03413_));
 sky130_fd_sc_hd__o21ai_0 _24142_ (.A1(_03028_),
    .A2(net3575),
    .B1(net3724),
    .Y(_03414_));
 sky130_fd_sc_hd__o311ai_0 _24143_ (.A1(net3724),
    .A2(_03146_),
    .A3(_03115_),
    .B1(_03414_),
    .C1(net3716),
    .Y(_03415_));
 sky130_fd_sc_hd__a31oi_2 _24144_ (.A1(_02993_),
    .A2(_03166_),
    .A3(_03284_),
    .B1(net3715),
    .Y(_03416_));
 sky130_fd_sc_hd__o21ai_0 _24145_ (.A1(_03206_),
    .A2(_03033_),
    .B1(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__nand2_1 _24146_ (.A(_03415_),
    .B(_03417_),
    .Y(_03418_));
 sky130_fd_sc_hd__nand3_1 _24147_ (.A(_03059_),
    .B(net3723),
    .C(_03418_),
    .Y(_03419_));
 sky130_fd_sc_hd__nand2_1 _24148_ (.A(_03270_),
    .B(_03283_),
    .Y(_03420_));
 sky130_fd_sc_hd__o22ai_1 _24149_ (.A1(net3726),
    .A2(_03162_),
    .B1(_03420_),
    .B2(net3638),
    .Y(_03421_));
 sky130_fd_sc_hd__o211ai_1 _24150_ (.A1(_12462_[0]),
    .A2(_02993_),
    .B1(_03017_),
    .C1(_03275_),
    .Y(_03422_));
 sky130_fd_sc_hd__o21ai_0 _24151_ (.A1(_03017_),
    .A2(_03262_),
    .B1(_03422_),
    .Y(_03423_));
 sky130_fd_sc_hd__a21oi_1 _24152_ (.A1(_03259_),
    .A2(_03423_),
    .B1(net3723),
    .Y(_03424_));
 sky130_fd_sc_hd__a211oi_1 _24153_ (.A1(net3712),
    .A2(_03265_),
    .B1(_03346_),
    .C1(net3726),
    .Y(_03425_));
 sky130_fd_sc_hd__o21ai_0 _24154_ (.A1(net3639),
    .A2(_03314_),
    .B1(net3724),
    .Y(_03426_));
 sky130_fd_sc_hd__o21ai_0 _24155_ (.A1(net3712),
    .A2(_03028_),
    .B1(_03162_),
    .Y(_03427_));
 sky130_fd_sc_hd__a221oi_1 _24156_ (.A1(_03093_),
    .A2(_03314_),
    .B1(_03427_),
    .B2(net3726),
    .C1(_03101_),
    .Y(_03428_));
 sky130_fd_sc_hd__o21ai_0 _24157_ (.A1(_03425_),
    .A2(_03426_),
    .B1(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__o311ai_0 _24158_ (.A1(_03059_),
    .A2(net3716),
    .A3(_03421_),
    .B1(_03424_),
    .C1(_03429_),
    .Y(_03430_));
 sky130_fd_sc_hd__o21ai_0 _24159_ (.A1(net3727),
    .A2(net3714),
    .B1(_03017_),
    .Y(_03431_));
 sky130_fd_sc_hd__a21oi_1 _24160_ (.A1(net3727),
    .A2(_03365_),
    .B1(_03431_),
    .Y(_03432_));
 sky130_fd_sc_hd__a21oi_1 _24161_ (.A1(_03265_),
    .A2(_03387_),
    .B1(_03432_),
    .Y(_03433_));
 sky130_fd_sc_hd__nand4_1 _24162_ (.A(net3723),
    .B(_03047_),
    .C(net3721),
    .D(_03205_),
    .Y(_03434_));
 sky130_fd_sc_hd__o22ai_1 _24163_ (.A1(net3639),
    .A2(_03033_),
    .B1(_03205_),
    .B2(net3720),
    .Y(_03435_));
 sky130_fd_sc_hd__a32oi_1 _24164_ (.A1(net3727),
    .A2(net3600),
    .A3(_03434_),
    .B1(_03435_),
    .B2(net3723),
    .Y(_03436_));
 sky130_fd_sc_hd__o211ai_1 _24165_ (.A1(net3726),
    .A2(_03433_),
    .B1(_03436_),
    .C1(net3716),
    .Y(_03437_));
 sky130_fd_sc_hd__a21oi_1 _24166_ (.A1(_12462_[0]),
    .A2(_03017_),
    .B1(net3575),
    .Y(_03438_));
 sky130_fd_sc_hd__nor2_1 _24167_ (.A(net3724),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__nor2_1 _24168_ (.A(_12460_[0]),
    .B(_03017_),
    .Y(_03440_));
 sky130_fd_sc_hd__a21oi_1 _24169_ (.A1(_12474_[0]),
    .A2(_03017_),
    .B1(_03440_),
    .Y(_03441_));
 sky130_fd_sc_hd__o221ai_1 _24170_ (.A1(net3629),
    .A2(_03080_),
    .B1(_03441_),
    .B2(net3724),
    .C1(net3714),
    .Y(_03442_));
 sky130_fd_sc_hd__o311ai_0 _24171_ (.A1(net3714),
    .A2(_03359_),
    .A3(_03439_),
    .B1(_03442_),
    .C1(_03086_),
    .Y(_03443_));
 sky130_fd_sc_hd__nand3_1 _24172_ (.A(net3724),
    .B(_03270_),
    .C(_03178_),
    .Y(_03444_));
 sky130_fd_sc_hd__nand4_1 _24173_ (.A(_03059_),
    .B(net3723),
    .C(_03416_),
    .D(_03444_),
    .Y(_03445_));
 sky130_fd_sc_hd__nand2_1 _24174_ (.A(_03054_),
    .B(_03445_),
    .Y(_03446_));
 sky130_fd_sc_hd__nor2_1 _24175_ (.A(_12474_[0]),
    .B(_03162_),
    .Y(_03447_));
 sky130_fd_sc_hd__a21oi_1 _24176_ (.A1(_12465_[0]),
    .A2(net3638),
    .B1(net3721),
    .Y(_03448_));
 sky130_fd_sc_hd__o21ai_0 _24177_ (.A1(_03447_),
    .A2(_03448_),
    .B1(_03371_),
    .Y(_03449_));
 sky130_fd_sc_hd__nor4_1 _24178_ (.A(net3727),
    .B(net3721),
    .C(_03155_),
    .D(_03199_),
    .Y(_03450_));
 sky130_fd_sc_hd__o21ai_0 _24179_ (.A1(_02993_),
    .A2(_03246_),
    .B1(net3715),
    .Y(_03451_));
 sky130_fd_sc_hd__o211ai_1 _24180_ (.A1(_02993_),
    .A2(_03168_),
    .B1(_03166_),
    .C1(net3713),
    .Y(_03452_));
 sky130_fd_sc_hd__o211ai_1 _24181_ (.A1(_03450_),
    .A2(_03451_),
    .B1(_03075_),
    .C1(_03452_),
    .Y(_03453_));
 sky130_fd_sc_hd__a21oi_1 _24182_ (.A1(_03449_),
    .A2(_03453_),
    .B1(_03101_),
    .Y(_03454_));
 sky130_fd_sc_hd__a311oi_1 _24183_ (.A1(_03101_),
    .A2(_03437_),
    .A3(_03443_),
    .B1(_03446_),
    .C1(_03454_),
    .Y(_03455_));
 sky130_fd_sc_hd__a31o_4 _24184_ (.A1(_03413_),
    .A2(_03419_),
    .A3(_03430_),
    .B1(_03455_),
    .X(_00157_));
 sky130_fd_sc_hd__a211oi_1 _24185_ (.A1(net3720),
    .A2(_03245_),
    .B1(_03115_),
    .C1(_02993_),
    .Y(_03456_));
 sky130_fd_sc_hd__a311oi_1 _24186_ (.A1(_02993_),
    .A2(_03270_),
    .A3(_03191_),
    .B1(_03456_),
    .C1(net3723),
    .Y(_03457_));
 sky130_fd_sc_hd__a21oi_1 _24187_ (.A1(_02981_),
    .A2(_03041_),
    .B1(net3720),
    .Y(_03458_));
 sky130_fd_sc_hd__nor3_1 _24188_ (.A(_03075_),
    .B(_03120_),
    .C(_03458_),
    .Y(_03459_));
 sky130_fd_sc_hd__nor3_1 _24189_ (.A(net3727),
    .B(net3639),
    .C(net3724),
    .Y(_03460_));
 sky130_fd_sc_hd__o21ai_0 _24190_ (.A1(net3629),
    .A2(_02993_),
    .B1(net3720),
    .Y(_03461_));
 sky130_fd_sc_hd__o22ai_1 _24191_ (.A1(_12479_[0]),
    .A2(net3720),
    .B1(_03460_),
    .B2(_03461_),
    .Y(_03462_));
 sky130_fd_sc_hd__o21ai_0 _24192_ (.A1(_03075_),
    .A2(_03462_),
    .B1(_03047_),
    .Y(_03463_));
 sky130_fd_sc_hd__nor3_1 _24193_ (.A(net3724),
    .B(_03114_),
    .C(_03115_),
    .Y(_03464_));
 sky130_fd_sc_hd__a311oi_1 _24194_ (.A1(net3724),
    .A2(_03270_),
    .A3(_03339_),
    .B1(_03464_),
    .C1(net3723),
    .Y(_03465_));
 sky130_fd_sc_hd__o32ai_2 _24195_ (.A1(_03047_),
    .A2(_03457_),
    .A3(_03459_),
    .B1(_03463_),
    .B2(_03465_),
    .Y(_03466_));
 sky130_fd_sc_hd__o32ai_1 _24196_ (.A1(net3724),
    .A2(_03021_),
    .A3(_03228_),
    .B1(_03080_),
    .B2(_12461_[0]),
    .Y(_03467_));
 sky130_fd_sc_hd__a21oi_1 _24197_ (.A1(_12470_[0]),
    .A2(_02993_),
    .B1(net3722),
    .Y(_03468_));
 sky130_fd_sc_hd__a221oi_2 _24198_ (.A1(_12478_[0]),
    .A2(net3722),
    .B1(_03130_),
    .B2(_03468_),
    .C1(net3723),
    .Y(_03469_));
 sky130_fd_sc_hd__a21oi_1 _24199_ (.A1(net3723),
    .A2(_03467_),
    .B1(_03469_),
    .Y(_03470_));
 sky130_fd_sc_hd__o21ai_0 _24200_ (.A1(_02993_),
    .A2(_03079_),
    .B1(net3723),
    .Y(_03471_));
 sky130_fd_sc_hd__o221ai_1 _24201_ (.A1(net3723),
    .A2(_03267_),
    .B1(_03307_),
    .B2(_03471_),
    .C1(net3712),
    .Y(_03472_));
 sky130_fd_sc_hd__o21ai_0 _24202_ (.A1(net3712),
    .A2(_03470_),
    .B1(_03472_),
    .Y(_03473_));
 sky130_fd_sc_hd__o22ai_1 _24203_ (.A1(_03102_),
    .A2(_03466_),
    .B1(_03473_),
    .B2(_03173_),
    .Y(_03474_));
 sky130_fd_sc_hd__mux2i_1 _24204_ (.A0(_03408_),
    .A1(_12460_[0]),
    .S(net3719),
    .Y(_03475_));
 sky130_fd_sc_hd__a32o_1 _24205_ (.A1(net3724),
    .A2(net3715),
    .A3(_03475_),
    .B1(_03025_),
    .B2(_12462_[0]),
    .X(_03476_));
 sky130_fd_sc_hd__nand2_1 _24206_ (.A(net3723),
    .B(_03476_),
    .Y(_03477_));
 sky130_fd_sc_hd__o21ai_0 _24207_ (.A1(_02981_),
    .A2(_02993_),
    .B1(_03140_),
    .Y(_03478_));
 sky130_fd_sc_hd__o311ai_0 _24208_ (.A1(_12477_[0]),
    .A2(_12486_[0]),
    .A3(net3722),
    .B1(_03478_),
    .C1(net3714),
    .Y(_03479_));
 sky130_fd_sc_hd__nand2_1 _24209_ (.A(_03477_),
    .B(_03479_),
    .Y(_03480_));
 sky130_fd_sc_hd__nand2_1 _24210_ (.A(net3715),
    .B(_03337_),
    .Y(_03481_));
 sky130_fd_sc_hd__nor2_2 _24211_ (.A(net3723),
    .B(net3717),
    .Y(_03482_));
 sky130_fd_sc_hd__nor2_1 _24212_ (.A(_02981_),
    .B(net3714),
    .Y(_03483_));
 sky130_fd_sc_hd__a211oi_1 _24213_ (.A1(_02987_),
    .A2(_02993_),
    .B1(net3723),
    .C1(net3728),
    .Y(_03484_));
 sky130_fd_sc_hd__nor4_1 _24214_ (.A(net3590),
    .B(_02993_),
    .C(net3714),
    .D(net3721),
    .Y(_03485_));
 sky130_fd_sc_hd__a211o_1 _24215_ (.A1(_03027_),
    .A2(_03483_),
    .B1(_03484_),
    .C1(_03485_),
    .X(_03486_));
 sky130_fd_sc_hd__a221o_1 _24216_ (.A1(net3723),
    .A2(_03155_),
    .B1(_03482_),
    .B2(net3599),
    .C1(_03486_),
    .X(_03487_));
 sky130_fd_sc_hd__nand2_1 _24217_ (.A(_03089_),
    .B(_03487_),
    .Y(_03488_));
 sky130_fd_sc_hd__a211oi_1 _24218_ (.A1(net3714),
    .A2(_03027_),
    .B1(_03483_),
    .C1(net3724),
    .Y(_03489_));
 sky130_fd_sc_hd__o21ai_0 _24219_ (.A1(_12470_[0]),
    .A2(net3723),
    .B1(net3721),
    .Y(_03490_));
 sky130_fd_sc_hd__o21ai_0 _24220_ (.A1(net3723),
    .A2(_03270_),
    .B1(_03490_),
    .Y(_03491_));
 sky130_fd_sc_hd__nor2_1 _24221_ (.A(_02993_),
    .B(_03491_),
    .Y(_03492_));
 sky130_fd_sc_hd__o221ai_1 _24222_ (.A1(net3714),
    .A2(_03070_),
    .B1(_03489_),
    .B2(_03492_),
    .C1(_03061_),
    .Y(_03493_));
 sky130_fd_sc_hd__a21oi_1 _24223_ (.A1(_12461_[0]),
    .A2(net3719),
    .B1(_03136_),
    .Y(_03494_));
 sky130_fd_sc_hd__a21oi_1 _24224_ (.A1(net3637),
    .A2(_03283_),
    .B1(_02993_),
    .Y(_03495_));
 sky130_fd_sc_hd__a2111oi_0 _24225_ (.A1(_02993_),
    .A2(_03494_),
    .B1(_03495_),
    .C1(_03476_),
    .D1(net3714),
    .Y(_03496_));
 sky130_fd_sc_hd__mux2i_1 _24226_ (.A0(_12474_[0]),
    .A1(_12470_[0]),
    .S(_02993_),
    .Y(_03497_));
 sky130_fd_sc_hd__o21ai_1 _24227_ (.A1(net3721),
    .A2(_03497_),
    .B1(_03086_),
    .Y(_03498_));
 sky130_fd_sc_hd__o21ai_0 _24228_ (.A1(_12462_[0]),
    .A2(net3638),
    .B1(net3721),
    .Y(_03499_));
 sky130_fd_sc_hd__a21oi_1 _24229_ (.A1(net3638),
    .A2(_03206_),
    .B1(_03499_),
    .Y(_03500_));
 sky130_fd_sc_hd__nor3_2 _24230_ (.A(net3723),
    .B(_03498_),
    .C(_03500_),
    .Y(_03501_));
 sky130_fd_sc_hd__o21ai_1 _24231_ (.A1(_03496_),
    .A2(_03501_),
    .B1(_03337_),
    .Y(_03502_));
 sky130_fd_sc_hd__o2111ai_1 _24232_ (.A1(_03480_),
    .A2(_03481_),
    .B1(_03488_),
    .C1(_03493_),
    .D1(_03502_),
    .Y(_03503_));
 sky130_fd_sc_hd__nor2_1 _24233_ (.A(_03474_),
    .B(_03503_),
    .Y(_00158_));
 sky130_fd_sc_hd__o21ai_0 _24234_ (.A1(_03028_),
    .A2(_03145_),
    .B1(net3724),
    .Y(_03504_));
 sky130_fd_sc_hd__a211oi_1 _24235_ (.A1(_03180_),
    .A2(_03504_),
    .B1(net3714),
    .C1(net3715),
    .Y(_03505_));
 sky130_fd_sc_hd__nor2_1 _24236_ (.A(_12465_[0]),
    .B(_02993_),
    .Y(_03506_));
 sky130_fd_sc_hd__o21ai_0 _24237_ (.A1(_03252_),
    .A2(_03506_),
    .B1(_03012_),
    .Y(_03507_));
 sky130_fd_sc_hd__nand2_1 _24238_ (.A(_03041_),
    .B(_03028_),
    .Y(_03508_));
 sky130_fd_sc_hd__nand3_1 _24239_ (.A(_12462_[0]),
    .B(_02993_),
    .C(_03017_),
    .Y(_03509_));
 sky130_fd_sc_hd__o21ai_0 _24240_ (.A1(_12472_[0]),
    .A2(_03017_),
    .B1(_03509_),
    .Y(_03510_));
 sky130_fd_sc_hd__a32o_1 _24241_ (.A1(_03371_),
    .A2(_03507_),
    .A3(_03508_),
    .B1(_03510_),
    .B2(_03365_),
    .X(_03511_));
 sky130_fd_sc_hd__a21oi_1 _24242_ (.A1(_12470_[0]),
    .A2(net3724),
    .B1(_03256_),
    .Y(_03512_));
 sky130_fd_sc_hd__nor2_1 _24243_ (.A(_12486_[0]),
    .B(net3717),
    .Y(_03513_));
 sky130_fd_sc_hd__a2111oi_0 _24244_ (.A1(net3719),
    .A2(_03512_),
    .B1(_03513_),
    .C1(net3715),
    .D1(net3723),
    .Y(_03514_));
 sky130_fd_sc_hd__nor3_1 _24245_ (.A(_03505_),
    .B(_03511_),
    .C(_03514_),
    .Y(_03515_));
 sky130_fd_sc_hd__a21oi_1 _24246_ (.A1(_03166_),
    .A2(_03168_),
    .B1(net3724),
    .Y(_03516_));
 sky130_fd_sc_hd__nand2_1 _24247_ (.A(net3714),
    .B(_03227_),
    .Y(_03517_));
 sky130_fd_sc_hd__a21oi_1 _24248_ (.A1(net3637),
    .A2(_03283_),
    .B1(net3724),
    .Y(_03518_));
 sky130_fd_sc_hd__o21ai_0 _24249_ (.A1(_03080_),
    .A2(_03245_),
    .B1(_03063_),
    .Y(_03519_));
 sky130_fd_sc_hd__o21ai_0 _24250_ (.A1(_03518_),
    .A2(_03519_),
    .B1(net3723),
    .Y(_03520_));
 sky130_fd_sc_hd__o21a_1 _24251_ (.A1(_03516_),
    .A2(_03517_),
    .B1(_03520_),
    .X(_03521_));
 sky130_fd_sc_hd__o21ai_0 _24252_ (.A1(net3714),
    .A2(_03080_),
    .B1(net3725),
    .Y(_03522_));
 sky130_fd_sc_hd__o311ai_0 _24253_ (.A1(net3725),
    .A2(_03104_),
    .A3(_03482_),
    .B1(_03522_),
    .C1(_02981_),
    .Y(_03523_));
 sky130_fd_sc_hd__nor2_1 _24254_ (.A(_03173_),
    .B(net3716),
    .Y(_03524_));
 sky130_fd_sc_hd__o2111ai_1 _24255_ (.A1(_02993_),
    .A2(_03270_),
    .B1(_03382_),
    .C1(_03523_),
    .D1(_03524_),
    .Y(_03525_));
 sky130_fd_sc_hd__o221ai_1 _24256_ (.A1(_03102_),
    .A2(_03515_),
    .B1(_03521_),
    .B2(_03481_),
    .C1(_03525_),
    .Y(_03526_));
 sky130_fd_sc_hd__a21oi_1 _24257_ (.A1(_03041_),
    .A2(_03275_),
    .B1(net3720),
    .Y(_03527_));
 sky130_fd_sc_hd__nor2_1 _24258_ (.A(_12470_[0]),
    .B(_03162_),
    .Y(_03528_));
 sky130_fd_sc_hd__a21oi_1 _24259_ (.A1(_03339_),
    .A2(_03284_),
    .B1(_02993_),
    .Y(_03529_));
 sky130_fd_sc_hd__o21ai_0 _24260_ (.A1(_03528_),
    .A2(_03529_),
    .B1(_03047_),
    .Y(_03530_));
 sky130_fd_sc_hd__o211ai_1 _24261_ (.A1(_03498_),
    .A2(_03527_),
    .B1(_03530_),
    .C1(_03075_),
    .Y(_03531_));
 sky130_fd_sc_hd__o21ai_0 _24262_ (.A1(net3724),
    .A2(_03191_),
    .B1(_03179_),
    .Y(_03532_));
 sky130_fd_sc_hd__nand3_1 _24263_ (.A(_12460_[0]),
    .B(net3724),
    .C(net3722),
    .Y(_03533_));
 sky130_fd_sc_hd__nand3_1 _24264_ (.A(net3716),
    .B(_03194_),
    .C(_03533_),
    .Y(_03534_));
 sky130_fd_sc_hd__a21oi_1 _24265_ (.A1(_02981_),
    .A2(_03532_),
    .B1(_03534_),
    .Y(_03535_));
 sky130_fd_sc_hd__o21ai_0 _24266_ (.A1(_12474_[0]),
    .A2(_03080_),
    .B1(_03194_),
    .Y(_03536_));
 sky130_fd_sc_hd__a211oi_1 _24267_ (.A1(_03177_),
    .A2(_03222_),
    .B1(_03536_),
    .C1(net3716),
    .Y(_03537_));
 sky130_fd_sc_hd__o21ai_1 _24268_ (.A1(_03535_),
    .A2(_03537_),
    .B1(net3723),
    .Y(_03538_));
 sky130_fd_sc_hd__a21oi_1 _24269_ (.A1(_03531_),
    .A2(_03538_),
    .B1(_03060_),
    .Y(_03539_));
 sky130_fd_sc_hd__nand2_1 _24270_ (.A(_12460_[0]),
    .B(net3724),
    .Y(_03540_));
 sky130_fd_sc_hd__o21ai_2 _24271_ (.A1(_03114_),
    .A2(_03265_),
    .B1(_02993_),
    .Y(_03541_));
 sky130_fd_sc_hd__nor2_1 _24272_ (.A(net3714),
    .B(_03141_),
    .Y(_03542_));
 sky130_fd_sc_hd__a32oi_1 _24273_ (.A1(net3714),
    .A2(_03540_),
    .A3(_03541_),
    .B1(_03542_),
    .B2(_03478_),
    .Y(_03543_));
 sky130_fd_sc_hd__nor3_1 _24274_ (.A(net3716),
    .B(_03149_),
    .C(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__a21oi_1 _24275_ (.A1(net3600),
    .A2(_03191_),
    .B1(_02981_),
    .Y(_03545_));
 sky130_fd_sc_hd__o21ai_0 _24276_ (.A1(_03372_),
    .A2(_03545_),
    .B1(net3714),
    .Y(_03546_));
 sky130_fd_sc_hd__o21ai_0 _24277_ (.A1(net3725),
    .A2(_03033_),
    .B1(_03162_),
    .Y(_03547_));
 sky130_fd_sc_hd__o21ai_0 _24278_ (.A1(_02987_),
    .A2(_03080_),
    .B1(_03070_),
    .Y(_03548_));
 sky130_fd_sc_hd__a22oi_1 _24279_ (.A1(_02981_),
    .A2(_03547_),
    .B1(_03548_),
    .B2(net3723),
    .Y(_03549_));
 sky130_fd_sc_hd__a211oi_1 _24280_ (.A1(_03546_),
    .A2(_03549_),
    .B1(_03173_),
    .C1(net3712),
    .Y(_03550_));
 sky130_fd_sc_hd__or4_4 _24281_ (.A(_03526_),
    .B(_03539_),
    .C(_03544_),
    .D(_03550_),
    .X(_00159_));
 sky130_fd_sc_hd__nor3_1 _24282_ (.A(\dcnt[1] ),
    .B(\dcnt[3] ),
    .C(\dcnt[2] ),
    .Y(_03551_));
 sky130_fd_sc_hd__and3b_1 _24283_ (.A_N(net4232),
    .B(\dcnt[0] ),
    .C(_03551_),
    .X(_00160_));
 sky130_fd_sc_hd__xor2_1 _24284_ (.A(net4170),
    .B(\sa00_sr[0] ),
    .X(_00185_));
 sky130_fd_sc_hd__xor2_1 _24285_ (.A(net4169),
    .B(\sa00_sr[1] ),
    .X(_00186_));
 sky130_fd_sc_hd__xor2_1 _24286_ (.A(net4168),
    .B(\sa00_sr[2] ),
    .X(_00187_));
 sky130_fd_sc_hd__xor2_1 _24287_ (.A(net4167),
    .B(\sa00_sr[3] ),
    .X(_00188_));
 sky130_fd_sc_hd__xor2_1 _24288_ (.A(net4166),
    .B(\sa00_sr[4] ),
    .X(_00189_));
 sky130_fd_sc_hd__xor2_1 _24289_ (.A(net4165),
    .B(\sa00_sr[5] ),
    .X(_00190_));
 sky130_fd_sc_hd__xor2_1 _24290_ (.A(\u0.w[0][30] ),
    .B(\sa00_sr[6] ),
    .X(_00191_));
 sky130_fd_sc_hd__xor2_1 _24291_ (.A(\u0.w[0][31] ),
    .B(net4229),
    .X(_00192_));
 sky130_fd_sc_hd__xor2_1 _24292_ (.A(net4151),
    .B(\sa01_sr[0] ),
    .X(_00281_));
 sky130_fd_sc_hd__xor2_1 _24293_ (.A(\u0.w[1][25] ),
    .B(net4227),
    .X(_00282_));
 sky130_fd_sc_hd__xor2_1 _24294_ (.A(net4149),
    .B(net4226),
    .X(_00283_));
 sky130_fd_sc_hd__xor2_1 _24295_ (.A(net4148),
    .B(net4225),
    .X(_00284_));
 sky130_fd_sc_hd__xor2_1 _24296_ (.A(\u0.w[1][28] ),
    .B(\sa01_sr[4] ),
    .X(_00285_));
 sky130_fd_sc_hd__xor2_1 _24297_ (.A(net4146),
    .B(\sa01_sr[5] ),
    .X(_00286_));
 sky130_fd_sc_hd__xor2_1 _24298_ (.A(net4145),
    .B(\sa01_sr[6] ),
    .X(_00287_));
 sky130_fd_sc_hd__xor2_1 _24299_ (.A(\u0.w[1][31] ),
    .B(\sa01_sr[7] ),
    .X(_00288_));
 sky130_fd_sc_hd__xor2_1 _24300_ (.A(\u0.w[2][24] ),
    .B(\sa02_sr[0] ),
    .X(_00241_));
 sky130_fd_sc_hd__xor2_1 _24301_ (.A(net4137),
    .B(\sa02_sr[1] ),
    .X(_00242_));
 sky130_fd_sc_hd__xor2_1 _24302_ (.A(\u0.w[2][26] ),
    .B(net4224),
    .X(_00243_));
 sky130_fd_sc_hd__xor2_1 _24303_ (.A(\u0.w[2][27] ),
    .B(\sa02_sr[3] ),
    .X(_00244_));
 sky130_fd_sc_hd__xor2_1 _24304_ (.A(\u0.w[2][28] ),
    .B(\sa02_sr[4] ),
    .X(_00245_));
 sky130_fd_sc_hd__xor2_1 _24305_ (.A(\u0.w[2][29] ),
    .B(\sa02_sr[5] ),
    .X(_00246_));
 sky130_fd_sc_hd__xor2_1 _24306_ (.A(\u0.w[2][30] ),
    .B(\sa02_sr[6] ),
    .X(_00247_));
 sky130_fd_sc_hd__xor2_1 _24307_ (.A(\u0.w[2][31] ),
    .B(\sa02_sr[7] ),
    .X(_00248_));
 sky130_fd_sc_hd__xor2_1 _24308_ (.A(net4131),
    .B(\sa03_sr[0] ),
    .X(_00209_));
 sky130_fd_sc_hd__xor2_1 _24309_ (.A(net4130),
    .B(\sa03_sr[1] ),
    .X(_00210_));
 sky130_fd_sc_hd__xor2_1 _24310_ (.A(\u0.tmp_w[26] ),
    .B(net4222),
    .X(_00211_));
 sky130_fd_sc_hd__xor2_1 _24311_ (.A(\u0.tmp_w[27] ),
    .B(\sa03_sr[3] ),
    .X(_00212_));
 sky130_fd_sc_hd__xor2_1 _24312_ (.A(net4129),
    .B(\sa03_sr[4] ),
    .X(_00213_));
 sky130_fd_sc_hd__xor2_1 _24313_ (.A(net4128),
    .B(\sa03_sr[5] ),
    .X(_00214_));
 sky130_fd_sc_hd__xor2_1 _24314_ (.A(\u0.tmp_w[30] ),
    .B(\sa03_sr[6] ),
    .X(_00215_));
 sky130_fd_sc_hd__xor2_1 _24315_ (.A(\u0.tmp_w[31] ),
    .B(net4221),
    .X(_00216_));
 sky130_fd_sc_hd__xor2_1 _24316_ (.A(\u0.w[0][16] ),
    .B(net4220),
    .X(_00177_));
 sky130_fd_sc_hd__xor2_1 _24317_ (.A(\u0.w[0][17] ),
    .B(\sa10_sr[1] ),
    .X(_00178_));
 sky130_fd_sc_hd__xor2_1 _24318_ (.A(\u0.w[0][18] ),
    .B(net4219),
    .X(_00179_));
 sky130_fd_sc_hd__xor2_1 _24319_ (.A(\u0.w[0][19] ),
    .B(\sa10_sr[3] ),
    .X(_00180_));
 sky130_fd_sc_hd__xor2_1 _24320_ (.A(\u0.w[0][20] ),
    .B(net4217),
    .X(_00181_));
 sky130_fd_sc_hd__xor2_1 _24321_ (.A(net4172),
    .B(\sa10_sr[5] ),
    .X(_00182_));
 sky130_fd_sc_hd__xor2_1 _24322_ (.A(net4171),
    .B(\sa10_sr[6] ),
    .X(_00183_));
 sky130_fd_sc_hd__xor2_1 _24323_ (.A(\u0.w[0][23] ),
    .B(net4216),
    .X(_00184_));
 sky130_fd_sc_hd__xor2_1 _24324_ (.A(net4155),
    .B(\sa11_sr[0] ),
    .X(_00273_));
 sky130_fd_sc_hd__xor2_1 _24325_ (.A(net4154),
    .B(\sa11_sr[1] ),
    .X(_00274_));
 sky130_fd_sc_hd__xor2_1 _24326_ (.A(\u0.w[1][18] ),
    .B(\sa11_sr[2] ),
    .X(_00275_));
 sky130_fd_sc_hd__xor2_1 _24327_ (.A(\u0.w[1][19] ),
    .B(\sa11_sr[3] ),
    .X(_00276_));
 sky130_fd_sc_hd__xor2_1 _24328_ (.A(\u0.w[1][20] ),
    .B(\sa11_sr[4] ),
    .X(_00277_));
 sky130_fd_sc_hd__xor2_1 _24329_ (.A(\u0.w[1][21] ),
    .B(\sa11_sr[5] ),
    .X(_00278_));
 sky130_fd_sc_hd__xor2_1 _24330_ (.A(net4152),
    .B(\sa11_sr[6] ),
    .X(_00279_));
 sky130_fd_sc_hd__xor2_1 _24331_ (.A(\u0.w[1][23] ),
    .B(net4214),
    .X(_00280_));
 sky130_fd_sc_hd__xor2_1 _24332_ (.A(\u0.w[2][16] ),
    .B(\sa12_sr[0] ),
    .X(_00233_));
 sky130_fd_sc_hd__xor2_1 _24333_ (.A(net4139),
    .B(\sa12_sr[1] ),
    .X(_00234_));
 sky130_fd_sc_hd__xor2_1 _24334_ (.A(\u0.w[2][18] ),
    .B(net4213),
    .X(_00235_));
 sky130_fd_sc_hd__xor2_1 _24335_ (.A(\u0.w[2][19] ),
    .B(\sa12_sr[3] ),
    .X(_00236_));
 sky130_fd_sc_hd__xor2_1 _24336_ (.A(net4138),
    .B(\sa12_sr[4] ),
    .X(_00237_));
 sky130_fd_sc_hd__xor2_1 _24337_ (.A(\u0.w[2][21] ),
    .B(\sa12_sr[5] ),
    .X(_00238_));
 sky130_fd_sc_hd__xor2_1 _24338_ (.A(\u0.w[2][22] ),
    .B(\sa12_sr[6] ),
    .X(_00239_));
 sky130_fd_sc_hd__xor2_1 _24339_ (.A(\u0.w[2][23] ),
    .B(\sa12_sr[7] ),
    .X(_00240_));
 sky130_fd_sc_hd__xor2_1 _24340_ (.A(\u0.tmp_w[16] ),
    .B(net4211),
    .X(_00201_));
 sky130_fd_sc_hd__xor2_1 _24341_ (.A(\u0.tmp_w[17] ),
    .B(net4210),
    .X(_00202_));
 sky130_fd_sc_hd__xor2_1 _24342_ (.A(\u0.tmp_w[18] ),
    .B(net4209),
    .X(_00203_));
 sky130_fd_sc_hd__xor2_1 _24343_ (.A(\u0.tmp_w[19] ),
    .B(\sa10_sub[3] ),
    .X(_00204_));
 sky130_fd_sc_hd__xor2_1 _24344_ (.A(\u0.tmp_w[20] ),
    .B(\sa10_sub[4] ),
    .X(_00205_));
 sky130_fd_sc_hd__xor2_1 _24345_ (.A(net4133),
    .B(\sa10_sub[5] ),
    .X(_00206_));
 sky130_fd_sc_hd__xor2_1 _24346_ (.A(net4132),
    .B(\sa10_sub[6] ),
    .X(_00207_));
 sky130_fd_sc_hd__xor2_1 _24347_ (.A(\u0.tmp_w[23] ),
    .B(\sa10_sub[7] ),
    .X(_00208_));
 sky130_fd_sc_hd__xor2_1 _24348_ (.A(\u0.w[0][8] ),
    .B(\sa20_sr[0] ),
    .X(_00169_));
 sky130_fd_sc_hd__xor2_1 _24349_ (.A(net4158),
    .B(\sa20_sr[1] ),
    .X(_00170_));
 sky130_fd_sc_hd__xor2_1 _24350_ (.A(\u0.w[0][10] ),
    .B(\sa20_sr[2] ),
    .X(_00171_));
 sky130_fd_sc_hd__xor2_1 _24351_ (.A(net4177),
    .B(\sa20_sr[3] ),
    .X(_00172_));
 sky130_fd_sc_hd__xor2_1 _24352_ (.A(net4176),
    .B(\sa20_sr[4] ),
    .X(_00173_));
 sky130_fd_sc_hd__xor2_1 _24353_ (.A(net4175),
    .B(net4208),
    .X(_00174_));
 sky130_fd_sc_hd__xor2_1 _24354_ (.A(net4174),
    .B(\sa20_sr[6] ),
    .X(_00175_));
 sky130_fd_sc_hd__xor2_1 _24355_ (.A(\u0.w[0][15] ),
    .B(net4207),
    .X(_00176_));
 sky130_fd_sc_hd__xor2_1 _24356_ (.A(\u0.w[1][8] ),
    .B(net4206),
    .X(_00257_));
 sky130_fd_sc_hd__xor2_1 _24357_ (.A(\u0.w[1][9] ),
    .B(\sa21_sr[1] ),
    .X(_00258_));
 sky130_fd_sc_hd__xor2_1 _24358_ (.A(\u0.w[1][10] ),
    .B(net4205),
    .X(_00259_));
 sky130_fd_sc_hd__xor2_1 _24359_ (.A(\u0.w[1][11] ),
    .B(\sa21_sr[3] ),
    .X(_00260_));
 sky130_fd_sc_hd__xor2_1 _24360_ (.A(\u0.w[1][12] ),
    .B(\sa21_sr[4] ),
    .X(_00261_));
 sky130_fd_sc_hd__xor2_1 _24361_ (.A(net4156),
    .B(net4203),
    .X(_00262_));
 sky130_fd_sc_hd__xor2_1 _24362_ (.A(\u0.w[1][14] ),
    .B(\sa21_sr[6] ),
    .X(_00263_));
 sky130_fd_sc_hd__xor2_1 _24363_ (.A(\u0.w[1][15] ),
    .B(\sa21_sr[7] ),
    .X(_00264_));
 sky130_fd_sc_hd__xor2_1 _24364_ (.A(\u0.w[2][8] ),
    .B(net4201),
    .X(_00225_));
 sky130_fd_sc_hd__xor2_1 _24365_ (.A(\u0.w[2][9] ),
    .B(\sa20_sub[1] ),
    .X(_00226_));
 sky130_fd_sc_hd__xor2_1 _24366_ (.A(\u0.w[2][10] ),
    .B(net4200),
    .X(_00227_));
 sky130_fd_sc_hd__xor2_1 _24367_ (.A(net4141),
    .B(\sa20_sub[3] ),
    .X(_00228_));
 sky130_fd_sc_hd__xor2_1 _24368_ (.A(net4140),
    .B(net4198),
    .X(_00229_));
 sky130_fd_sc_hd__xor2_1 _24369_ (.A(\u0.w[2][13] ),
    .B(net4197),
    .X(_00230_));
 sky130_fd_sc_hd__xor2_1 _24370_ (.A(\u0.w[2][14] ),
    .B(\sa20_sub[6] ),
    .X(_00231_));
 sky130_fd_sc_hd__xor2_1 _24371_ (.A(\u0.w[2][15] ),
    .B(net4196),
    .X(_00232_));
 sky130_fd_sc_hd__xor2_1 _24372_ (.A(net4126),
    .B(net4195),
    .X(_00193_));
 sky130_fd_sc_hd__xor2_1 _24373_ (.A(\u0.tmp_w[9] ),
    .B(net4194),
    .X(_00194_));
 sky130_fd_sc_hd__xor2_1 _24374_ (.A(\u0.tmp_w[10] ),
    .B(net4193),
    .X(_00195_));
 sky130_fd_sc_hd__xor2_1 _24375_ (.A(\u0.tmp_w[11] ),
    .B(net4192),
    .X(_00196_));
 sky130_fd_sc_hd__xor2_1 _24376_ (.A(\u0.tmp_w[12] ),
    .B(\sa21_sub[4] ),
    .X(_00197_));
 sky130_fd_sc_hd__xor2_1 _24377_ (.A(\u0.tmp_w[13] ),
    .B(\sa21_sub[5] ),
    .X(_00198_));
 sky130_fd_sc_hd__xor2_1 _24378_ (.A(\u0.tmp_w[14] ),
    .B(\sa21_sub[6] ),
    .X(_00199_));
 sky130_fd_sc_hd__xor2_1 _24379_ (.A(\u0.tmp_w[15] ),
    .B(net4191),
    .X(_00200_));
 sky130_fd_sc_hd__xor2_1 _24380_ (.A(net4178),
    .B(\sa30_sr[0] ),
    .X(_00161_));
 sky130_fd_sc_hd__xor2_1 _24381_ (.A(net4173),
    .B(\sa30_sr[1] ),
    .X(_00162_));
 sky130_fd_sc_hd__xor2_1 _24382_ (.A(\u0.w[0][2] ),
    .B(\sa30_sr[2] ),
    .X(_00163_));
 sky130_fd_sc_hd__xor2_1 _24383_ (.A(net4163),
    .B(\sa30_sr[3] ),
    .X(_00164_));
 sky130_fd_sc_hd__xor2_1 _24384_ (.A(\u0.w[0][4] ),
    .B(net4190),
    .X(_00165_));
 sky130_fd_sc_hd__xor2_1 _24385_ (.A(net4161),
    .B(\sa30_sr[5] ),
    .X(_00166_));
 sky130_fd_sc_hd__xor2_1 _24386_ (.A(net4160),
    .B(\sa30_sr[6] ),
    .X(_00167_));
 sky130_fd_sc_hd__xor2_1 _24387_ (.A(net4159),
    .B(net4189),
    .X(_00168_));
 sky130_fd_sc_hd__xor2_1 _24388_ (.A(net4157),
    .B(\sa30_sub[0] ),
    .X(_00249_));
 sky130_fd_sc_hd__xor2_1 _24389_ (.A(net4153),
    .B(\sa30_sub[1] ),
    .X(_00250_));
 sky130_fd_sc_hd__xor2_1 _24390_ (.A(\u0.w[1][2] ),
    .B(\sa30_sub[2] ),
    .X(_00251_));
 sky130_fd_sc_hd__xor2_1 _24391_ (.A(\u0.w[1][3] ),
    .B(net4188),
    .X(_00252_));
 sky130_fd_sc_hd__xor2_1 _24392_ (.A(net4144),
    .B(net4187),
    .X(_00253_));
 sky130_fd_sc_hd__xor2_1 _24393_ (.A(net4143),
    .B(\sa30_sub[5] ),
    .X(_00254_));
 sky130_fd_sc_hd__xor2_1 _24394_ (.A(net4142),
    .B(\sa30_sub[6] ),
    .X(_00255_));
 sky130_fd_sc_hd__xor2_1 _24395_ (.A(\u0.w[1][7] ),
    .B(\sa30_sub[7] ),
    .X(_00256_));
 sky130_fd_sc_hd__xor2_1 _24396_ (.A(\u0.w[2][0] ),
    .B(\sa31_sub[0] ),
    .X(_00217_));
 sky130_fd_sc_hd__xor2_1 _24397_ (.A(\u0.w[2][1] ),
    .B(net4185),
    .X(_00218_));
 sky130_fd_sc_hd__xor2_1 _24398_ (.A(\u0.w[2][2] ),
    .B(net4184),
    .X(_00219_));
 sky130_fd_sc_hd__xor2_1 _24399_ (.A(\u0.w[2][3] ),
    .B(net4183),
    .X(_00220_));
 sky130_fd_sc_hd__xor2_1 _24400_ (.A(\u0.w[2][4] ),
    .B(\sa31_sub[4] ),
    .X(_00221_));
 sky130_fd_sc_hd__xor2_1 _24401_ (.A(\u0.w[2][5] ),
    .B(\sa31_sub[5] ),
    .X(_00222_));
 sky130_fd_sc_hd__xor2_1 _24402_ (.A(\u0.w[2][6] ),
    .B(\sa31_sub[6] ),
    .X(_00223_));
 sky130_fd_sc_hd__xor2_1 _24403_ (.A(\u0.w[2][7] ),
    .B(net4182),
    .X(_00224_));
 sky130_fd_sc_hd__xor2_1 _24404_ (.A(\u0.tmp_w[0] ),
    .B(\sa32_sub[0] ),
    .X(_00265_));
 sky130_fd_sc_hd__xor2_1 _24405_ (.A(net4134),
    .B(net4181),
    .X(_00266_));
 sky130_fd_sc_hd__xor2_1 _24406_ (.A(\u0.tmp_w[2] ),
    .B(\sa32_sub[2] ),
    .X(_00267_));
 sky130_fd_sc_hd__xor2_1 _24407_ (.A(\u0.tmp_w[3] ),
    .B(net4180),
    .X(_00268_));
 sky130_fd_sc_hd__xor2_1 _24408_ (.A(\u0.tmp_w[4] ),
    .B(\sa32_sub[4] ),
    .X(_00269_));
 sky130_fd_sc_hd__xor2_1 _24409_ (.A(net4127),
    .B(\sa32_sub[5] ),
    .X(_00270_));
 sky130_fd_sc_hd__xor2_1 _24410_ (.A(\u0.tmp_w[6] ),
    .B(\sa32_sub[6] ),
    .X(_00271_));
 sky130_fd_sc_hd__xor2_1 _24411_ (.A(\u0.tmp_w[7] ),
    .B(net4179),
    .X(_00272_));
 sky130_fd_sc_hd__inv_1 _24412_ (.A(\u0.r0.rcnt[0] ),
    .Y(\u0.r0.rcnt_next[0] ));
 sky130_fd_sc_hd__inv_1 _24413_ (.A(\u0.r0.rcnt[1] ),
    .Y(_12490_[0]));
 sky130_fd_sc_hd__nor2b_1 _24414_ (.A(\dcnt[2] ),
    .B_N(\dcnt[3] ),
    .Y(_03552_));
 sky130_fd_sc_hd__nor2_1 _24415_ (.A(\dcnt[1] ),
    .B(\dcnt[0] ),
    .Y(_03553_));
 sky130_fd_sc_hd__mux2i_1 _24416_ (.A0(\dcnt[2] ),
    .A1(_03552_),
    .S(_03553_),
    .Y(_03554_));
 sky130_fd_sc_hd__nor3b_1 _24417_ (.A(net4232),
    .B(_03554_),
    .C_N(net130),
    .Y(_00407_));
 sky130_fd_sc_hd__xnor2_1 _24418_ (.A(\u0.r0.rcnt[2] ),
    .B(_12498_[0]),
    .Y(_03555_));
 sky130_fd_sc_hd__a21o_1 _24419_ (.A1(_12496_[0]),
    .A2(_03555_),
    .B1(net4235),
    .X(_00409_));
 sky130_fd_sc_hd__xor2_1 _24420_ (.A(\u0.r0.rcnt[2] ),
    .B(_12498_[0]),
    .X(_03556_));
 sky130_fd_sc_hd__nand3_1 _24421_ (.A(\u0.r0.rcnt[2] ),
    .B(\u0.r0.rcnt[1] ),
    .C(\u0.r0.rcnt[0] ),
    .Y(_03557_));
 sky130_fd_sc_hd__xor2_2 _24422_ (.A(\u0.r0.rcnt[3] ),
    .B(_03557_),
    .X(_03558_));
 sky130_fd_sc_hd__nor2_1 _24423_ (.A(\u0.r0.rcnt_next[1] ),
    .B(_03558_),
    .Y(_03559_));
 sky130_fd_sc_hd__a21oi_1 _24424_ (.A1(_12491_[0]),
    .A2(_03558_),
    .B1(_03559_),
    .Y(_03560_));
 sky130_fd_sc_hd__nor3_1 _24425_ (.A(net4235),
    .B(_03556_),
    .C(_03560_),
    .Y(_00410_));
 sky130_fd_sc_hd__mux2i_1 _24426_ (.A0(_12491_[0]),
    .A1(_12494_[0]),
    .S(_03558_),
    .Y(_03561_));
 sky130_fd_sc_hd__nor3_1 _24427_ (.A(net4235),
    .B(_03556_),
    .C(_03561_),
    .Y(_00411_));
 sky130_fd_sc_hd__mux2i_1 _24428_ (.A0(_12496_[0]),
    .A1(_12492_[0]),
    .S(_03558_),
    .Y(_03562_));
 sky130_fd_sc_hd__nor3_1 _24429_ (.A(net4235),
    .B(_03556_),
    .C(_03562_),
    .Y(_00412_));
 sky130_fd_sc_hd__nor3_1 _24430_ (.A(\u0.r0.rcnt_next[1] ),
    .B(_03556_),
    .C(_03558_),
    .Y(_03563_));
 sky130_fd_sc_hd__a31oi_1 _24431_ (.A1(_12496_[0]),
    .A2(_03556_),
    .A3(_03558_),
    .B1(_03563_),
    .Y(_03564_));
 sky130_fd_sc_hd__nor2_1 _24432_ (.A(net4235),
    .B(_03564_),
    .Y(_00413_));
 sky130_fd_sc_hd__xnor2_1 _24433_ (.A(_03555_),
    .B(_03558_),
    .Y(_03565_));
 sky130_fd_sc_hd__nor3b_1 _24434_ (.A(net4235),
    .B(_03565_),
    .C_N(_12491_[0]),
    .Y(_00414_));
 sky130_fd_sc_hd__nor2_1 _24435_ (.A(net4235),
    .B(_03555_),
    .Y(_00419_));
 sky130_fd_sc_hd__and3_1 _24436_ (.A(_12494_[0]),
    .B(_03558_),
    .C(_00419_),
    .X(_00415_));
 sky130_fd_sc_hd__and3_1 _24437_ (.A(_12492_[0]),
    .B(_03558_),
    .C(_00419_),
    .X(_00416_));
 sky130_fd_sc_hd__nor2_1 _24438_ (.A(net4235),
    .B(\u0.r0.rcnt[0] ),
    .Y(_00417_));
 sky130_fd_sc_hd__nor2b_1 _24439_ (.A(net4235),
    .B_N(\u0.r0.rcnt_next[1] ),
    .Y(_00418_));
 sky130_fd_sc_hd__nor2_1 _24440_ (.A(net4235),
    .B(_03558_),
    .Y(_00420_));
 sky130_fd_sc_hd__nor2_1 _24441_ (.A(\dcnt[0] ),
    .B(_03551_),
    .Y(_03566_));
 sky130_fd_sc_hd__o21a_1 _24442_ (.A1(net4232),
    .A2(_03566_),
    .B1(net130),
    .X(_00405_));
 sky130_fd_sc_hd__a21oi_1 _24443_ (.A1(\dcnt[1] ),
    .A2(\dcnt[0] ),
    .B1(net4232),
    .Y(_03567_));
 sky130_fd_sc_hd__o21ai_0 _24444_ (.A1(\dcnt[3] ),
    .A2(\dcnt[2] ),
    .B1(_03553_),
    .Y(_03568_));
 sky130_fd_sc_hd__a21boi_0 _24445_ (.A1(_03567_),
    .A2(_03568_),
    .B1_N(net130),
    .Y(_00406_));
 sky130_fd_sc_hd__o31a_1 _24446_ (.A1(\dcnt[1] ),
    .A2(\dcnt[0] ),
    .A3(\dcnt[2] ),
    .B1(\dcnt[3] ),
    .X(_03569_));
 sky130_fd_sc_hd__o21a_1 _24447_ (.A1(net4232),
    .A2(_03569_),
    .B1(net130),
    .X(_00408_));
 sky130_fd_sc_hd__ha_4 _24448_ (.A(_03592_),
    .B(_03585_),
    .COUT(_11828_[0]),
    .SUM(_11829_[0]));
 sky130_fd_sc_hd__ha_4 _24449_ (.A(net4105),
    .B(net4106),
    .COUT(_11830_[0]),
    .SUM(_11831_[0]));
 sky130_fd_sc_hd__ha_4 _24450_ (.A(net4105),
    .B(_03586_),
    .COUT(_11833_[0]),
    .SUM(_11834_[0]));
 sky130_fd_sc_hd__ha_4 _24451_ (.A(net4105),
    .B(_03586_),
    .COUT(_11835_[0]),
    .SUM(_11836_[0]));
 sky130_fd_sc_hd__ha_4 _24452_ (.A(_03593_),
    .B(net4106),
    .COUT(_11838_[0]),
    .SUM(_11839_[0]));
 sky130_fd_sc_hd__ha_4 _24453_ (.A(_03593_),
    .B(net4106),
    .COUT(_11840_[0]),
    .SUM(_11841_[0]));
 sky130_fd_sc_hd__ha_4 _24454_ (.A(_03593_),
    .B(_03586_),
    .COUT(_11842_[0]),
    .SUM(_11843_[0]));
 sky130_fd_sc_hd__ha_4 _24455_ (.A(_03593_),
    .B(_03586_),
    .COUT(_11844_[0]),
    .SUM(_11845_[0]));
 sky130_fd_sc_hd__ha_1 _24456_ (.A(net4105),
    .B(net4100),
    .COUT(_11847_[0]),
    .SUM(_11848_[0]));
 sky130_fd_sc_hd__ha_4 _24457_ (.A(net4105),
    .B(_03617_),
    .COUT(_11849_[0]),
    .SUM(_11850_[0]));
 sky130_fd_sc_hd__ha_1 _24458_ (.A(net4105),
    .B(_03618_),
    .COUT(_11852_[0]),
    .SUM(_11853_[0]));
 sky130_fd_sc_hd__ha_4 _24459_ (.A(net4105),
    .B(_03618_),
    .COUT(_11854_[0]),
    .SUM(_11855_[0]));
 sky130_fd_sc_hd__ha_1 _24460_ (.A(_03593_),
    .B(_03617_),
    .COUT(_11856_[0]),
    .SUM(_11857_[0]));
 sky130_fd_sc_hd__ha_1 _24461_ (.A(_03593_),
    .B(_03617_),
    .COUT(_11858_[0]),
    .SUM(_11859_[0]));
 sky130_fd_sc_hd__ha_4 _24462_ (.A(_11860_[0]),
    .B(_03690_),
    .COUT(_11862_[0]),
    .SUM(_11863_[0]));
 sky130_fd_sc_hd__ha_4 _24463_ (.A(_11860_[0]),
    .B(net4090),
    .COUT(_11864_[0]),
    .SUM(_11865_[0]));
 sky130_fd_sc_hd__ha_4 _24464_ (.A(_11860_[0]),
    .B(_03691_),
    .COUT(_11867_[0]),
    .SUM(_11868_[0]));
 sky130_fd_sc_hd__ha_4 _24465_ (.A(_11860_[0]),
    .B(_03691_),
    .COUT(_11869_[0]),
    .SUM(_11870_[0]));
 sky130_fd_sc_hd__ha_4 _24466_ (.A(_03696_),
    .B(net4090),
    .COUT(_11872_[0]),
    .SUM(_11873_[0]));
 sky130_fd_sc_hd__ha_4 _24467_ (.A(_03696_),
    .B(net4090),
    .COUT(_11874_[0]),
    .SUM(_11875_[0]));
 sky130_fd_sc_hd__ha_4 _24468_ (.A(_03696_),
    .B(_03691_),
    .COUT(_11876_[0]),
    .SUM(_11877_[0]));
 sky130_fd_sc_hd__ha_4 _24469_ (.A(_03696_),
    .B(net4063),
    .COUT(_11878_[0]),
    .SUM(_11879_[0]));
 sky130_fd_sc_hd__ha_1 _24470_ (.A(net4089),
    .B(net4088),
    .COUT(_11881_[0]),
    .SUM(_11882_[0]));
 sky130_fd_sc_hd__ha_4 _24471_ (.A(net4089),
    .B(net4088),
    .COUT(_11883_[0]),
    .SUM(_11884_[0]));
 sky130_fd_sc_hd__ha_1 _24472_ (.A(net4089),
    .B(_03704_),
    .COUT(_11886_[0]),
    .SUM(_11887_[0]));
 sky130_fd_sc_hd__ha_1 _24473_ (.A(net4089),
    .B(_03704_),
    .COUT(_11888_[0]),
    .SUM(_11889_[0]));
 sky130_fd_sc_hd__ha_1 _24474_ (.A(_03696_),
    .B(_03702_),
    .COUT(_11890_[0]),
    .SUM(_11891_[0]));
 sky130_fd_sc_hd__ha_1 _24475_ (.A(_03696_),
    .B(_03702_),
    .COUT(_11892_[0]),
    .SUM(_11893_[0]));
 sky130_fd_sc_hd__ha_4 _24476_ (.A(_03630_),
    .B(_03624_),
    .COUT(_11896_[0]),
    .SUM(_11897_[0]));
 sky130_fd_sc_hd__ha_4 _24477_ (.A(net4094),
    .B(net4097),
    .COUT(_11898_[0]),
    .SUM(_11899_[0]));
 sky130_fd_sc_hd__ha_4 _24478_ (.A(net4095),
    .B(_03625_),
    .COUT(_11901_[0]),
    .SUM(_11902_[0]));
 sky130_fd_sc_hd__ha_4 _24479_ (.A(_03630_),
    .B(_03625_),
    .COUT(_11903_[0]),
    .SUM(_11904_[0]));
 sky130_fd_sc_hd__ha_4 _24480_ (.A(_03631_),
    .B(net4099),
    .COUT(_11906_[0]),
    .SUM(_11907_[0]));
 sky130_fd_sc_hd__ha_4 _24481_ (.A(_03631_),
    .B(net4097),
    .COUT(_11908_[0]),
    .SUM(_11909_[0]));
 sky130_fd_sc_hd__ha_4 _24482_ (.A(_03631_),
    .B(_03625_),
    .COUT(_11910_[0]),
    .SUM(_11911_[0]));
 sky130_fd_sc_hd__ha_4 _24483_ (.A(_03631_),
    .B(_03625_),
    .COUT(_11912_[0]),
    .SUM(_11913_[0]));
 sky130_fd_sc_hd__ha_1 _24484_ (.A(net4094),
    .B(_03637_),
    .COUT(_11915_[0]),
    .SUM(_11916_[0]));
 sky130_fd_sc_hd__ha_4 _24485_ (.A(net4096),
    .B(net4093),
    .COUT(_11917_[0]),
    .SUM(_11918_[0]));
 sky130_fd_sc_hd__ha_1 _24486_ (.A(net4096),
    .B(_03639_),
    .COUT(_11920_[0]),
    .SUM(_11921_[0]));
 sky130_fd_sc_hd__ha_1 _24487_ (.A(net4096),
    .B(_03639_),
    .COUT(_11922_[0]),
    .SUM(_11923_[0]));
 sky130_fd_sc_hd__ha_1 _24488_ (.A(_03631_),
    .B(net4093),
    .COUT(_11924_[0]),
    .SUM(_11925_[0]));
 sky130_fd_sc_hd__ha_1 _24489_ (.A(_03631_),
    .B(net4093),
    .COUT(_11926_[0]),
    .SUM(_11927_[0]));
 sky130_fd_sc_hd__ha_4 _24490_ (.A(_03772_),
    .B(_03777_),
    .COUT(_11930_[0]),
    .SUM(_11931_[0]));
 sky130_fd_sc_hd__ha_4 _24491_ (.A(_03777_),
    .B(_03772_),
    .COUT(_11932_[0]),
    .SUM(_11933_[0]));
 sky130_fd_sc_hd__ha_4 _24492_ (.A(_03777_),
    .B(_03773_),
    .COUT(_11935_[0]),
    .SUM(_11936_[0]));
 sky130_fd_sc_hd__ha_4 _24493_ (.A(_03777_),
    .B(_03773_),
    .COUT(_11937_[0]),
    .SUM(_11938_[0]));
 sky130_fd_sc_hd__ha_4 _24494_ (.A(_03778_),
    .B(_03772_),
    .COUT(_11940_[0]),
    .SUM(_11941_[0]));
 sky130_fd_sc_hd__ha_4 _24495_ (.A(_03778_),
    .B(_03772_),
    .COUT(_11942_[0]),
    .SUM(_11943_[0]));
 sky130_fd_sc_hd__ha_4 _24496_ (.A(_03778_),
    .B(_03773_),
    .COUT(_11944_[0]),
    .SUM(_11945_[0]));
 sky130_fd_sc_hd__ha_4 _24497_ (.A(_03778_),
    .B(_03773_),
    .COUT(_11946_[0]),
    .SUM(_11947_[0]));
 sky130_fd_sc_hd__ha_1 _24498_ (.A(net4078),
    .B(net4082),
    .COUT(_11949_[0]),
    .SUM(_11950_[0]));
 sky130_fd_sc_hd__ha_4 _24499_ (.A(net4080),
    .B(net4082),
    .COUT(_11951_[0]),
    .SUM(_11952_[0]));
 sky130_fd_sc_hd__ha_1 _24500_ (.A(_03784_),
    .B(net4082),
    .COUT(_11954_[0]),
    .SUM(_11955_[0]));
 sky130_fd_sc_hd__ha_1 _24501_ (.A(_03784_),
    .B(net4082),
    .COUT(_11956_[0]),
    .SUM(_11957_[0]));
 sky130_fd_sc_hd__ha_1 _24502_ (.A(_03784_),
    .B(_03778_),
    .COUT(_11958_[0]),
    .SUM(_11959_[0]));
 sky130_fd_sc_hd__ha_1 _24503_ (.A(_03784_),
    .B(_03778_),
    .COUT(_11960_[0]),
    .SUM(_11961_[0]));
 sky130_fd_sc_hd__ha_4 _24504_ (.A(_05890_),
    .B(_05883_),
    .COUT(_11964_[0]),
    .SUM(_11965_[0]));
 sky130_fd_sc_hd__ha_4 _24505_ (.A(_05890_),
    .B(net4059),
    .COUT(_11966_[0]),
    .SUM(_11967_[0]));
 sky130_fd_sc_hd__ha_4 _24506_ (.A(_05890_),
    .B(_05884_),
    .COUT(_11969_[0]),
    .SUM(_11970_[0]));
 sky130_fd_sc_hd__ha_4 _24507_ (.A(_05891_),
    .B(_05883_),
    .COUT(_11972_[0]),
    .SUM(_11973_[0]));
 sky130_fd_sc_hd__ha_4 _24508_ (.A(_05891_),
    .B(_05883_),
    .COUT(_11974_[0]),
    .SUM(_11975_[0]));
 sky130_fd_sc_hd__ha_1 _24509_ (.A(_05891_),
    .B(net3710),
    .COUT(_11976_[0]),
    .SUM(_11977_[0]));
 sky130_fd_sc_hd__ha_4 _24510_ (.A(_05891_),
    .B(_05884_),
    .COUT(_11978_[0]),
    .SUM(_11979_[0]));
 sky130_fd_sc_hd__ha_1 _24511_ (.A(net4054),
    .B(net4057),
    .COUT(_11981_[0]),
    .SUM(_11982_[0]));
 sky130_fd_sc_hd__ha_1 _24512_ (.A(net4054),
    .B(net3710),
    .COUT(_11983_[0]),
    .SUM(_11984_[0]));
 sky130_fd_sc_hd__ha_1 _24513_ (.A(net4054),
    .B(_05884_),
    .COUT(_11985_[0]),
    .SUM(_11986_[0]));
 sky130_fd_sc_hd__ha_1 _24514_ (.A(_05900_),
    .B(net4057),
    .COUT(_11988_[0]),
    .SUM(_11989_[0]));
 sky130_fd_sc_hd__ha_1 _24515_ (.A(net3709),
    .B(net4057),
    .COUT(_11990_[0]),
    .SUM(_11991_[0]));
 sky130_fd_sc_hd__ha_1 _24516_ (.A(_05900_),
    .B(net3710),
    .COUT(_11992_[0]),
    .SUM(_11993_[0]));
 sky130_fd_sc_hd__ha_4 _24517_ (.A(_06493_),
    .B(_06486_),
    .COUT(_11996_[0]),
    .SUM(_11997_[0]));
 sky130_fd_sc_hd__ha_4 _24518_ (.A(_06493_),
    .B(net4037),
    .COUT(_11998_[0]),
    .SUM(_11999_[0]));
 sky130_fd_sc_hd__ha_4 _24519_ (.A(_06493_),
    .B(_06487_),
    .COUT(_12001_[0]),
    .SUM(_12002_[0]));
 sky130_fd_sc_hd__ha_4 _24520_ (.A(_06494_),
    .B(net4037),
    .COUT(_12004_[0]),
    .SUM(_12005_[0]));
 sky130_fd_sc_hd__ha_4 _24521_ (.A(_06494_),
    .B(net4037),
    .COUT(_12006_[0]),
    .SUM(_12007_[0]));
 sky130_fd_sc_hd__ha_1 _24522_ (.A(_06494_),
    .B(net3703),
    .COUT(_12008_[0]),
    .SUM(_12009_[0]));
 sky130_fd_sc_hd__ha_4 _24523_ (.A(_06494_),
    .B(net3703),
    .COUT(_12010_[0]),
    .SUM(_12011_[0]));
 sky130_fd_sc_hd__ha_1 _24524_ (.A(net4033),
    .B(net4037),
    .COUT(_12013_[0]),
    .SUM(_12014_[0]));
 sky130_fd_sc_hd__ha_1 _24525_ (.A(net4033),
    .B(net3703),
    .COUT(_12015_[0]),
    .SUM(_12016_[0]));
 sky130_fd_sc_hd__ha_1 _24526_ (.A(net4033),
    .B(net3704),
    .COUT(_12017_[0]),
    .SUM(_12018_[0]));
 sky130_fd_sc_hd__ha_1 _24527_ (.A(net3702),
    .B(net4037),
    .COUT(_12020_[0]),
    .SUM(_12021_[0]));
 sky130_fd_sc_hd__ha_1 _24528_ (.A(_06505_),
    .B(net4037),
    .COUT(_12022_[0]),
    .SUM(_12023_[0]));
 sky130_fd_sc_hd__ha_1 _24529_ (.A(_06505_),
    .B(net3703),
    .COUT(_12024_[0]),
    .SUM(_12025_[0]));
 sky130_fd_sc_hd__ha_4 _24530_ (.A(net4012),
    .B(_07081_),
    .COUT(_12028_[0]),
    .SUM(_12029_[0]));
 sky130_fd_sc_hd__ha_4 _24531_ (.A(net4013),
    .B(_07081_),
    .COUT(_12030_[0]),
    .SUM(_12031_[0]));
 sky130_fd_sc_hd__ha_4 _24532_ (.A(net4013),
    .B(_07082_),
    .COUT(_12033_[0]),
    .SUM(_12034_[0]));
 sky130_fd_sc_hd__ha_4 _24533_ (.A(_07090_),
    .B(net406),
    .COUT(_12036_[0]),
    .SUM(_12037_[0]));
 sky130_fd_sc_hd__ha_4 _24534_ (.A(_07090_),
    .B(net405),
    .COUT(_12038_[0]),
    .SUM(_12039_[0]));
 sky130_fd_sc_hd__ha_1 _24535_ (.A(_07090_),
    .B(_07082_),
    .COUT(_12040_[0]),
    .SUM(_12041_[0]));
 sky130_fd_sc_hd__ha_4 _24536_ (.A(_07090_),
    .B(_07082_),
    .COUT(_12042_[0]),
    .SUM(_12043_[0]));
 sky130_fd_sc_hd__ha_1 _24537_ (.A(net4010),
    .B(net4014),
    .COUT(_12045_[0]),
    .SUM(_12046_[0]));
 sky130_fd_sc_hd__ha_1 _24538_ (.A(net4010),
    .B(_07082_),
    .COUT(_12047_[0]),
    .SUM(_12048_[0]));
 sky130_fd_sc_hd__ha_1 _24539_ (.A(net4011),
    .B(_07082_),
    .COUT(_12049_[0]),
    .SUM(_12050_[0]));
 sky130_fd_sc_hd__ha_1 _24540_ (.A(_07100_),
    .B(net4015),
    .COUT(_12052_[0]),
    .SUM(_12053_[0]));
 sky130_fd_sc_hd__ha_1 _24541_ (.A(_07100_),
    .B(net4014),
    .COUT(_12054_[0]),
    .SUM(_12055_[0]));
 sky130_fd_sc_hd__ha_1 _24542_ (.A(_07100_),
    .B(_07082_),
    .COUT(_12056_[0]),
    .SUM(_12057_[0]));
 sky130_fd_sc_hd__ha_4 _24543_ (.A(_07675_),
    .B(_07667_),
    .COUT(_12060_[0]),
    .SUM(_12061_[0]));
 sky130_fd_sc_hd__ha_4 _24544_ (.A(_07675_),
    .B(_07667_),
    .COUT(_12062_[0]),
    .SUM(_12063_[0]));
 sky130_fd_sc_hd__ha_4 _24545_ (.A(_07675_),
    .B(_07668_),
    .COUT(_12065_[0]),
    .SUM(_12066_[0]));
 sky130_fd_sc_hd__ha_4 _24546_ (.A(_07676_),
    .B(_07667_),
    .COUT(_12068_[0]),
    .SUM(_12069_[0]));
 sky130_fd_sc_hd__ha_4 _24547_ (.A(_07676_),
    .B(_07667_),
    .COUT(_12070_[0]),
    .SUM(_12071_[0]));
 sky130_fd_sc_hd__ha_1 _24548_ (.A(_07676_),
    .B(net3696),
    .COUT(_12072_[0]),
    .SUM(_12073_[0]));
 sky130_fd_sc_hd__ha_4 _24549_ (.A(_07676_),
    .B(_07668_),
    .COUT(_12074_[0]),
    .SUM(_12075_[0]));
 sky130_fd_sc_hd__ha_1 _24550_ (.A(net3995),
    .B(net3999),
    .COUT(_12077_[0]),
    .SUM(_12078_[0]));
 sky130_fd_sc_hd__ha_1 _24551_ (.A(net3995),
    .B(net3696),
    .COUT(_12079_[0]),
    .SUM(_12080_[0]));
 sky130_fd_sc_hd__ha_4 _24552_ (.A(net3995),
    .B(net3696),
    .COUT(_12081_[0]),
    .SUM(_12082_[0]));
 sky130_fd_sc_hd__ha_1 _24553_ (.A(_07684_),
    .B(net3999),
    .COUT(_12084_[0]),
    .SUM(_12085_[0]));
 sky130_fd_sc_hd__ha_1 _24554_ (.A(_07684_),
    .B(net3999),
    .COUT(_12086_[0]),
    .SUM(_12087_[0]));
 sky130_fd_sc_hd__ha_1 _24555_ (.A(net3693),
    .B(net3696),
    .COUT(_12088_[0]),
    .SUM(_12089_[0]));
 sky130_fd_sc_hd__ha_4 _24556_ (.A(_08243_),
    .B(_08237_),
    .COUT(_12092_[0]),
    .SUM(_12093_[0]));
 sky130_fd_sc_hd__ha_4 _24557_ (.A(net3980),
    .B(net3981),
    .COUT(_12094_[0]),
    .SUM(_12095_[0]));
 sky130_fd_sc_hd__ha_4 _24558_ (.A(net3980),
    .B(_08238_),
    .COUT(_12097_[0]),
    .SUM(_12098_[0]));
 sky130_fd_sc_hd__ha_4 _24559_ (.A(_08244_),
    .B(net3981),
    .COUT(_12100_[0]),
    .SUM(_12101_[0]));
 sky130_fd_sc_hd__ha_4 _24560_ (.A(_08244_),
    .B(net3981),
    .COUT(_12102_[0]),
    .SUM(_12103_[0]));
 sky130_fd_sc_hd__ha_1 _24561_ (.A(net3688),
    .B(net3690),
    .COUT(_12104_[0]),
    .SUM(_12105_[0]));
 sky130_fd_sc_hd__ha_4 _24562_ (.A(_08244_),
    .B(_08238_),
    .COUT(_12106_[0]),
    .SUM(_12107_[0]));
 sky130_fd_sc_hd__ha_1 _24563_ (.A(net3978),
    .B(net3981),
    .COUT(_12109_[0]),
    .SUM(_12110_[0]));
 sky130_fd_sc_hd__ha_1 _24564_ (.A(net3978),
    .B(net3690),
    .COUT(_12111_[0]),
    .SUM(_12112_[0]));
 sky130_fd_sc_hd__ha_1 _24565_ (.A(net3978),
    .B(_08238_),
    .COUT(_12113_[0]),
    .SUM(_12114_[0]));
 sky130_fd_sc_hd__ha_1 _24566_ (.A(_08250_),
    .B(net3982),
    .COUT(_12116_[0]),
    .SUM(_12117_[0]));
 sky130_fd_sc_hd__ha_1 _24567_ (.A(_08250_),
    .B(net3981),
    .COUT(_12118_[0]),
    .SUM(_12119_[0]));
 sky130_fd_sc_hd__ha_1 _24568_ (.A(_08250_),
    .B(net3690),
    .COUT(_12120_[0]),
    .SUM(_12121_[0]));
 sky130_fd_sc_hd__ha_4 _24569_ (.A(_08811_),
    .B(_08805_),
    .COUT(_12124_[0]),
    .SUM(_12125_[0]));
 sky130_fd_sc_hd__ha_4 _24570_ (.A(_08811_),
    .B(_08805_),
    .COUT(_12126_[0]),
    .SUM(_12127_[0]));
 sky130_fd_sc_hd__ha_4 _24571_ (.A(_08811_),
    .B(_08806_),
    .COUT(_12129_[0]),
    .SUM(_12130_[0]));
 sky130_fd_sc_hd__ha_4 _24572_ (.A(_08812_),
    .B(net3958),
    .COUT(_12132_[0]),
    .SUM(_12133_[0]));
 sky130_fd_sc_hd__ha_4 _24573_ (.A(_08812_),
    .B(net3958),
    .COUT(_12134_[0]),
    .SUM(_12135_[0]));
 sky130_fd_sc_hd__ha_1 _24574_ (.A(net3683),
    .B(_08806_),
    .COUT(_12136_[0]),
    .SUM(_12137_[0]));
 sky130_fd_sc_hd__ha_4 _24575_ (.A(_08812_),
    .B(_08806_),
    .COUT(_12138_[0]),
    .SUM(_12139_[0]));
 sky130_fd_sc_hd__ha_1 _24576_ (.A(net3956),
    .B(net3958),
    .COUT(_12141_[0]),
    .SUM(_12142_[0]));
 sky130_fd_sc_hd__ha_1 _24577_ (.A(net3956),
    .B(_08806_),
    .COUT(_12143_[0]),
    .SUM(_12144_[0]));
 sky130_fd_sc_hd__ha_1 _24578_ (.A(net3956),
    .B(net3686),
    .COUT(_12145_[0]),
    .SUM(_12146_[0]));
 sky130_fd_sc_hd__ha_1 _24579_ (.A(_08818_),
    .B(net3959),
    .COUT(_12148_[0]),
    .SUM(_12149_[0]));
 sky130_fd_sc_hd__ha_1 _24580_ (.A(_08818_),
    .B(net3958),
    .COUT(_12150_[0]),
    .SUM(_12151_[0]));
 sky130_fd_sc_hd__ha_1 _24581_ (.A(_08818_),
    .B(net3686),
    .COUT(_12152_[0]),
    .SUM(_12153_[0]));
 sky130_fd_sc_hd__ha_4 _24582_ (.A(net3932),
    .B(_09363_),
    .COUT(_12156_[0]),
    .SUM(_12157_[0]));
 sky130_fd_sc_hd__ha_4 _24583_ (.A(net3932),
    .B(_09363_),
    .COUT(_12158_[0]),
    .SUM(_12159_[0]));
 sky130_fd_sc_hd__ha_4 _24584_ (.A(net3932),
    .B(_09364_),
    .COUT(_12161_[0]),
    .SUM(_12162_[0]));
 sky130_fd_sc_hd__ha_4 _24585_ (.A(_09370_),
    .B(_09363_),
    .COUT(_12164_[0]),
    .SUM(_12165_[0]));
 sky130_fd_sc_hd__ha_4 _24586_ (.A(_09370_),
    .B(_09363_),
    .COUT(_12166_[0]),
    .SUM(_12167_[0]));
 sky130_fd_sc_hd__ha_2 _24587_ (.A(_09370_),
    .B(net3678),
    .COUT(_12168_[0]),
    .SUM(_12169_[0]));
 sky130_fd_sc_hd__ha_4 _24588_ (.A(_09370_),
    .B(_09364_),
    .COUT(_12170_[0]),
    .SUM(_12171_[0]));
 sky130_fd_sc_hd__ha_1 _24589_ (.A(net3931),
    .B(net3936),
    .COUT(_12173_[0]),
    .SUM(_12174_[0]));
 sky130_fd_sc_hd__ha_1 _24590_ (.A(net3931),
    .B(net3678),
    .COUT(_12175_[0]),
    .SUM(_12176_[0]));
 sky130_fd_sc_hd__ha_1 _24591_ (.A(net3931),
    .B(net3678),
    .COUT(_12177_[0]),
    .SUM(_12178_[0]));
 sky130_fd_sc_hd__ha_1 _24592_ (.A(_09375_),
    .B(net3935),
    .COUT(_12180_[0]),
    .SUM(_12181_[0]));
 sky130_fd_sc_hd__ha_1 _24593_ (.A(_09375_),
    .B(net3936),
    .COUT(_12182_[0]),
    .SUM(_12183_[0]));
 sky130_fd_sc_hd__ha_1 _24594_ (.A(_09375_),
    .B(_09364_),
    .COUT(_12184_[0]),
    .SUM(_12185_[0]));
 sky130_fd_sc_hd__ha_4 _24595_ (.A(net409),
    .B(net3907),
    .COUT(_12188_[0]),
    .SUM(_12189_[0]));
 sky130_fd_sc_hd__ha_4 _24596_ (.A(net3906),
    .B(net3908),
    .COUT(_12190_[0]),
    .SUM(_12191_[0]));
 sky130_fd_sc_hd__ha_4 _24597_ (.A(net409),
    .B(_09923_),
    .COUT(_12193_[0]),
    .SUM(_12194_[0]));
 sky130_fd_sc_hd__ha_4 _24598_ (.A(_09929_),
    .B(net3908),
    .COUT(_12196_[0]),
    .SUM(_12197_[0]));
 sky130_fd_sc_hd__ha_4 _24599_ (.A(_09929_),
    .B(_09922_),
    .COUT(_12198_[0]),
    .SUM(_12199_[0]));
 sky130_fd_sc_hd__ha_1 _24600_ (.A(_09929_),
    .B(_09923_),
    .COUT(_12200_[0]),
    .SUM(_12201_[0]));
 sky130_fd_sc_hd__ha_4 _24601_ (.A(_09929_),
    .B(_09923_),
    .COUT(_12202_[0]),
    .SUM(_12203_[0]));
 sky130_fd_sc_hd__ha_1 _24602_ (.A(net3904),
    .B(net3908),
    .COUT(_12205_[0]),
    .SUM(_12206_[0]));
 sky130_fd_sc_hd__ha_1 _24603_ (.A(net3904),
    .B(_09923_),
    .COUT(_12207_[0]),
    .SUM(_12208_[0]));
 sky130_fd_sc_hd__ha_1 _24604_ (.A(net3904),
    .B(_09923_),
    .COUT(_12209_[0]),
    .SUM(_12210_[0]));
 sky130_fd_sc_hd__ha_1 _24605_ (.A(_09936_),
    .B(net3908),
    .COUT(_12212_[0]),
    .SUM(_12213_[0]));
 sky130_fd_sc_hd__ha_1 _24606_ (.A(_09936_),
    .B(net3908),
    .COUT(_12214_[0]),
    .SUM(_12215_[0]));
 sky130_fd_sc_hd__ha_1 _24607_ (.A(_09936_),
    .B(_09923_),
    .COUT(_12216_[0]),
    .SUM(_12217_[0]));
 sky130_fd_sc_hd__ha_4 _24608_ (.A(net388),
    .B(net3885),
    .COUT(_12220_[0]),
    .SUM(_12221_[0]));
 sky130_fd_sc_hd__ha_4 _24609_ (.A(net3885),
    .B(net3888),
    .COUT(_12222_[0]),
    .SUM(_12223_[0]));
 sky130_fd_sc_hd__ha_4 _24610_ (.A(net3885),
    .B(_10495_),
    .COUT(_12225_[0]),
    .SUM(_12226_[0]));
 sky130_fd_sc_hd__ha_4 _24611_ (.A(_10495_),
    .B(net3885),
    .COUT(_12227_[0]),
    .SUM(_12228_[0]));
 sky130_fd_sc_hd__ha_4 _24612_ (.A(_10500_),
    .B(net3888),
    .COUT(_12230_[0]),
    .SUM(_12231_[0]));
 sky130_fd_sc_hd__ha_4 _24613_ (.A(_10500_),
    .B(net3888),
    .COUT(_12232_[0]),
    .SUM(_12233_[0]));
 sky130_fd_sc_hd__ha_4 _24614_ (.A(_10500_),
    .B(_10495_),
    .COUT(_12234_[0]),
    .SUM(_12235_[0]));
 sky130_fd_sc_hd__ha_4 _24615_ (.A(_10500_),
    .B(_10495_),
    .COUT(_12236_[0]),
    .SUM(_12237_[0]));
 sky130_fd_sc_hd__ha_1 _24616_ (.A(net3883),
    .B(net3888),
    .COUT(_12239_[0]),
    .SUM(_12240_[0]));
 sky130_fd_sc_hd__ha_1 _24617_ (.A(net3883),
    .B(_10495_),
    .COUT(_12241_[0]),
    .SUM(_12242_[0]));
 sky130_fd_sc_hd__ha_1 _24618_ (.A(net3883),
    .B(_10495_),
    .COUT(_12243_[0]),
    .SUM(_12244_[0]));
 sky130_fd_sc_hd__ha_1 _24619_ (.A(_10509_),
    .B(net3888),
    .COUT(_12246_[0]),
    .SUM(_12247_[0]));
 sky130_fd_sc_hd__ha_1 _24620_ (.A(_10509_),
    .B(net3888),
    .COUT(_12248_[0]),
    .SUM(_12249_[0]));
 sky130_fd_sc_hd__ha_1 _24621_ (.A(_10509_),
    .B(_10495_),
    .COUT(_12250_[0]),
    .SUM(_12251_[0]));
 sky130_fd_sc_hd__ha_1 _24622_ (.A(net3675),
    .B(_10495_),
    .COUT(_12252_[0]),
    .SUM(_12253_[0]));
 sky130_fd_sc_hd__ha_4 _24623_ (.A(net3865),
    .B(net3867),
    .COUT(_12256_[0]),
    .SUM(_12257_[0]));
 sky130_fd_sc_hd__ha_4 _24624_ (.A(net3866),
    .B(net3867),
    .COUT(_12258_[0]),
    .SUM(_12259_[0]));
 sky130_fd_sc_hd__ha_4 _24625_ (.A(net3865),
    .B(_11065_),
    .COUT(_12261_[0]),
    .SUM(_12262_[0]));
 sky130_fd_sc_hd__ha_4 _24626_ (.A(net3865),
    .B(_11065_),
    .COUT(_12263_[0]),
    .SUM(_12264_[0]));
 sky130_fd_sc_hd__ha_4 _24627_ (.A(_11071_),
    .B(net3868),
    .COUT(_12266_[0]),
    .SUM(_12267_[0]));
 sky130_fd_sc_hd__ha_4 _24628_ (.A(_11071_),
    .B(net3867),
    .COUT(_12268_[0]),
    .SUM(_12269_[0]));
 sky130_fd_sc_hd__ha_4 _24629_ (.A(_11071_),
    .B(_11065_),
    .COUT(_12270_[0]),
    .SUM(_12271_[0]));
 sky130_fd_sc_hd__ha_4 _24630_ (.A(_11071_),
    .B(_11065_),
    .COUT(_12272_[0]),
    .SUM(_12273_[0]));
 sky130_fd_sc_hd__ha_1 _24631_ (.A(net3863),
    .B(net3868),
    .COUT(_12275_[0]),
    .SUM(_12276_[0]));
 sky130_fd_sc_hd__ha_1 _24632_ (.A(net3863),
    .B(_11065_),
    .COUT(_12277_[0]),
    .SUM(_12278_[0]));
 sky130_fd_sc_hd__ha_1 _24633_ (.A(net3863),
    .B(net3672),
    .COUT(_12279_[0]),
    .SUM(_12280_[0]));
 sky130_fd_sc_hd__ha_1 _24634_ (.A(_11076_),
    .B(net3868),
    .COUT(_12282_[0]),
    .SUM(_12283_[0]));
 sky130_fd_sc_hd__ha_1 _24635_ (.A(_11076_),
    .B(net3868),
    .COUT(_12284_[0]),
    .SUM(_12285_[0]));
 sky130_fd_sc_hd__ha_1 _24636_ (.A(_11076_),
    .B(net3672),
    .COUT(_12286_[0]),
    .SUM(_12287_[0]));
 sky130_fd_sc_hd__ha_1 _24637_ (.A(_11076_),
    .B(_11065_),
    .COUT(_12288_[0]),
    .SUM(_12289_[0]));
 sky130_fd_sc_hd__ha_4 _24638_ (.A(_11622_),
    .B(_11617_),
    .COUT(_12292_[0]),
    .SUM(_12293_[0]));
 sky130_fd_sc_hd__ha_4 _24639_ (.A(_11622_),
    .B(_11617_),
    .COUT(_12294_[0]),
    .SUM(_12295_[0]));
 sky130_fd_sc_hd__ha_4 _24640_ (.A(_11622_),
    .B(_11618_),
    .COUT(_12297_[0]),
    .SUM(_12298_[0]));
 sky130_fd_sc_hd__ha_4 _24641_ (.A(_11622_),
    .B(_11618_),
    .COUT(_12299_[0]),
    .SUM(_12300_[0]));
 sky130_fd_sc_hd__ha_4 _24642_ (.A(_11623_),
    .B(_11617_),
    .COUT(_12302_[0]),
    .SUM(_12303_[0]));
 sky130_fd_sc_hd__ha_4 _24643_ (.A(_11623_),
    .B(_11617_),
    .COUT(_12304_[0]),
    .SUM(_12305_[0]));
 sky130_fd_sc_hd__ha_4 _24644_ (.A(_11623_),
    .B(_11618_),
    .COUT(_12306_[0]),
    .SUM(_12307_[0]));
 sky130_fd_sc_hd__ha_4 _24645_ (.A(_11623_),
    .B(_11618_),
    .COUT(_12308_[0]),
    .SUM(_12309_[0]));
 sky130_fd_sc_hd__ha_1 _24646_ (.A(net3848),
    .B(net3851),
    .COUT(_12311_[0]),
    .SUM(_12312_[0]));
 sky130_fd_sc_hd__ha_1 _24647_ (.A(net3848),
    .B(_11618_),
    .COUT(_12313_[0]),
    .SUM(_12314_[0]));
 sky130_fd_sc_hd__ha_1 _24648_ (.A(net3848),
    .B(_11618_),
    .COUT(_12315_[0]),
    .SUM(_12316_[0]));
 sky130_fd_sc_hd__ha_1 _24649_ (.A(_11628_),
    .B(net3850),
    .COUT(_12318_[0]),
    .SUM(_12319_[0]));
 sky130_fd_sc_hd__ha_1 _24650_ (.A(_11628_),
    .B(net3851),
    .COUT(_12320_[0]),
    .SUM(_12321_[0]));
 sky130_fd_sc_hd__ha_2 _24651_ (.A(_11628_),
    .B(net3665),
    .COUT(_12322_[0]),
    .SUM(_12323_[0]));
 sky130_fd_sc_hd__ha_1 _24652_ (.A(_11628_),
    .B(_11618_),
    .COUT(_12324_[0]),
    .SUM(_12325_[0]));
 sky130_fd_sc_hd__ha_4 _24653_ (.A(_00783_),
    .B(_00776_),
    .COUT(_12328_[0]),
    .SUM(_12329_[0]));
 sky130_fd_sc_hd__ha_4 _24654_ (.A(_00783_),
    .B(_00776_),
    .COUT(_12330_[0]),
    .SUM(_12331_[0]));
 sky130_fd_sc_hd__ha_4 _24655_ (.A(net3829),
    .B(_00777_),
    .COUT(_12333_[0]),
    .SUM(_12334_[0]));
 sky130_fd_sc_hd__ha_4 _24656_ (.A(_00783_),
    .B(_00777_),
    .COUT(_12335_[0]),
    .SUM(_12336_[0]));
 sky130_fd_sc_hd__ha_4 _24657_ (.A(_00784_),
    .B(net3831),
    .COUT(_12338_[0]),
    .SUM(_12339_[0]));
 sky130_fd_sc_hd__ha_4 _24658_ (.A(_00784_),
    .B(_00776_),
    .COUT(_12340_[0]),
    .SUM(_12341_[0]));
 sky130_fd_sc_hd__ha_4 _24659_ (.A(_00784_),
    .B(_00777_),
    .COUT(_12342_[0]),
    .SUM(_12343_[0]));
 sky130_fd_sc_hd__ha_4 _24660_ (.A(_00784_),
    .B(_00777_),
    .COUT(_12344_[0]),
    .SUM(_12345_[0]));
 sky130_fd_sc_hd__ha_1 _24661_ (.A(net3827),
    .B(net3831),
    .COUT(_12347_[0]),
    .SUM(_12348_[0]));
 sky130_fd_sc_hd__ha_1 _24662_ (.A(net3828),
    .B(_00777_),
    .COUT(_12349_[0]),
    .SUM(_12350_[0]));
 sky130_fd_sc_hd__ha_1 _24663_ (.A(net3827),
    .B(_00777_),
    .COUT(_12351_[0]),
    .SUM(_12352_[0]));
 sky130_fd_sc_hd__ha_1 _24664_ (.A(_00798_),
    .B(net3831),
    .COUT(_12354_[0]),
    .SUM(_12355_[0]));
 sky130_fd_sc_hd__ha_1 _24665_ (.A(_00798_),
    .B(net3831),
    .COUT(_12356_[0]),
    .SUM(_12357_[0]));
 sky130_fd_sc_hd__ha_4 _24666_ (.A(_00798_),
    .B(_00777_),
    .COUT(_12358_[0]),
    .SUM(_12359_[0]));
 sky130_fd_sc_hd__ha_1 _24667_ (.A(_00798_),
    .B(_00777_),
    .COUT(_12360_[0]),
    .SUM(_12361_[0]));
 sky130_fd_sc_hd__ha_4 _24668_ (.A(net3799),
    .B(_01342_),
    .COUT(_12364_[0]),
    .SUM(_12365_[0]));
 sky130_fd_sc_hd__ha_4 _24669_ (.A(net3799),
    .B(_01342_),
    .COUT(_12366_[0]),
    .SUM(_12367_[0]));
 sky130_fd_sc_hd__ha_4 _24670_ (.A(net3800),
    .B(_01343_),
    .COUT(_12369_[0]),
    .SUM(_12370_[0]));
 sky130_fd_sc_hd__ha_4 _24671_ (.A(_01349_),
    .B(_01342_),
    .COUT(_12372_[0]),
    .SUM(_12373_[0]));
 sky130_fd_sc_hd__ha_4 _24672_ (.A(_01349_),
    .B(_01342_),
    .COUT(_12374_[0]),
    .SUM(_12375_[0]));
 sky130_fd_sc_hd__ha_1 _24673_ (.A(_01349_),
    .B(_01343_),
    .COUT(_12376_[0]),
    .SUM(_12377_[0]));
 sky130_fd_sc_hd__ha_4 _24674_ (.A(_01349_),
    .B(_01343_),
    .COUT(_12378_[0]),
    .SUM(_12379_[0]));
 sky130_fd_sc_hd__ha_1 _24675_ (.A(net3797),
    .B(net3802),
    .COUT(_12381_[0]),
    .SUM(_12382_[0]));
 sky130_fd_sc_hd__ha_1 _24676_ (.A(net3796),
    .B(net3656),
    .COUT(_12383_[0]),
    .SUM(_12384_[0]));
 sky130_fd_sc_hd__ha_1 _24677_ (.A(net3797),
    .B(_01343_),
    .COUT(_12385_[0]),
    .SUM(_12386_[0]));
 sky130_fd_sc_hd__ha_2 _24678_ (.A(_01354_),
    .B(net3802),
    .COUT(_12388_[0]),
    .SUM(_12389_[0]));
 sky130_fd_sc_hd__ha_1 _24679_ (.A(_01354_),
    .B(net3802),
    .COUT(_12390_[0]),
    .SUM(_12391_[0]));
 sky130_fd_sc_hd__ha_1 _24680_ (.A(net3653),
    .B(net3656),
    .COUT(_12392_[0]),
    .SUM(_12393_[0]));
 sky130_fd_sc_hd__ha_4 _24681_ (.A(_01885_),
    .B(net3778),
    .COUT(_12396_[0]),
    .SUM(_12397_[0]));
 sky130_fd_sc_hd__ha_4 _24682_ (.A(net3777),
    .B(net3778),
    .COUT(_12398_[0]),
    .SUM(_12399_[0]));
 sky130_fd_sc_hd__ha_4 _24683_ (.A(net3777),
    .B(_01882_),
    .COUT(_12401_[0]),
    .SUM(_12402_[0]));
 sky130_fd_sc_hd__ha_4 _24684_ (.A(_01886_),
    .B(net3778),
    .COUT(_12404_[0]),
    .SUM(_12405_[0]));
 sky130_fd_sc_hd__ha_4 _24685_ (.A(_01886_),
    .B(net3778),
    .COUT(_12406_[0]),
    .SUM(_12407_[0]));
 sky130_fd_sc_hd__ha_1 _24686_ (.A(net3650),
    .B(_01882_),
    .COUT(_12408_[0]),
    .SUM(_12409_[0]));
 sky130_fd_sc_hd__ha_4 _24687_ (.A(_01886_),
    .B(_01882_),
    .COUT(_12410_[0]),
    .SUM(_12411_[0]));
 sky130_fd_sc_hd__ha_1 _24688_ (.A(net3771),
    .B(net3779),
    .COUT(_12413_[0]),
    .SUM(_12414_[0]));
 sky130_fd_sc_hd__ha_1 _24689_ (.A(net3773),
    .B(_01882_),
    .COUT(_12415_[0]),
    .SUM(_12416_[0]));
 sky130_fd_sc_hd__ha_1 _24690_ (.A(net3771),
    .B(_01882_),
    .COUT(_12417_[0]),
    .SUM(_12418_[0]));
 sky130_fd_sc_hd__ha_1 _24691_ (.A(_01892_),
    .B(net3779),
    .COUT(_12420_[0]),
    .SUM(_12421_[0]));
 sky130_fd_sc_hd__ha_1 _24692_ (.A(_01892_),
    .B(net3779),
    .COUT(_12422_[0]),
    .SUM(_12423_[0]));
 sky130_fd_sc_hd__ha_1 _24693_ (.A(net3648),
    .B(_01882_),
    .COUT(_12424_[0]),
    .SUM(_12425_[0]));
 sky130_fd_sc_hd__ha_4 _24694_ (.A(_02443_),
    .B(_02437_),
    .COUT(_12428_[0]),
    .SUM(_12429_[0]));
 sky130_fd_sc_hd__ha_4 _24695_ (.A(net3748),
    .B(net3750),
    .COUT(_12430_[0]),
    .SUM(_12431_[0]));
 sky130_fd_sc_hd__ha_4 _24696_ (.A(net3748),
    .B(_02438_),
    .COUT(_12433_[0]),
    .SUM(_12434_[0]));
 sky130_fd_sc_hd__ha_4 _24697_ (.A(_02444_),
    .B(net3751),
    .COUT(_12436_[0]),
    .SUM(_12437_[0]));
 sky130_fd_sc_hd__ha_4 _24698_ (.A(_02444_),
    .B(_02437_),
    .COUT(_12438_[0]),
    .SUM(_12439_[0]));
 sky130_fd_sc_hd__ha_1 _24699_ (.A(_02444_),
    .B(net3643),
    .COUT(_12440_[0]),
    .SUM(_12441_[0]));
 sky130_fd_sc_hd__ha_4 _24700_ (.A(_02444_),
    .B(_02438_),
    .COUT(_12442_[0]),
    .SUM(_12443_[0]));
 sky130_fd_sc_hd__ha_4 _24701_ (.A(_02448_),
    .B(net3751),
    .COUT(_12445_[0]),
    .SUM(_12446_[0]));
 sky130_fd_sc_hd__ha_1 _24702_ (.A(net3746),
    .B(net3643),
    .COUT(_12447_[0]),
    .SUM(_12448_[0]));
 sky130_fd_sc_hd__ha_1 _24703_ (.A(net3746),
    .B(net3643),
    .COUT(_12449_[0]),
    .SUM(_12450_[0]));
 sky130_fd_sc_hd__ha_1 _24704_ (.A(_02449_),
    .B(net3751),
    .COUT(_12452_[0]),
    .SUM(_12453_[0]));
 sky130_fd_sc_hd__ha_2 _24705_ (.A(_02449_),
    .B(net3751),
    .COUT(_12454_[0]),
    .SUM(_12455_[0]));
 sky130_fd_sc_hd__ha_1 _24706_ (.A(_02449_),
    .B(net3643),
    .COUT(_12456_[0]),
    .SUM(_12457_[0]));
 sky130_fd_sc_hd__ha_4 _24707_ (.A(_02986_),
    .B(_02980_),
    .COUT(_12460_[0]),
    .SUM(_12461_[0]));
 sky130_fd_sc_hd__ha_4 _24708_ (.A(_02986_),
    .B(_02980_),
    .COUT(_12462_[0]),
    .SUM(_12463_[0]));
 sky130_fd_sc_hd__ha_4 _24709_ (.A(_02986_),
    .B(_02981_),
    .COUT(_12465_[0]),
    .SUM(_12466_[0]));
 sky130_fd_sc_hd__ha_4 _24710_ (.A(net3639),
    .B(net3727),
    .COUT(_12468_[0]),
    .SUM(_12469_[0]));
 sky130_fd_sc_hd__ha_4 _24711_ (.A(_02987_),
    .B(net3727),
    .COUT(_12470_[0]),
    .SUM(_12471_[0]));
 sky130_fd_sc_hd__ha_1 _24712_ (.A(_02987_),
    .B(_02981_),
    .COUT(_12472_[0]),
    .SUM(_12473_[0]));
 sky130_fd_sc_hd__ha_4 _24713_ (.A(_02987_),
    .B(_02981_),
    .COUT(_12474_[0]),
    .SUM(_12475_[0]));
 sky130_fd_sc_hd__ha_1 _24714_ (.A(net3724),
    .B(net3728),
    .COUT(_12477_[0]),
    .SUM(_12478_[0]));
 sky130_fd_sc_hd__ha_1 _24715_ (.A(net3724),
    .B(_02981_),
    .COUT(_12479_[0]),
    .SUM(_12480_[0]));
 sky130_fd_sc_hd__ha_1 _24716_ (.A(net3724),
    .B(_02981_),
    .COUT(_12481_[0]),
    .SUM(_12482_[0]));
 sky130_fd_sc_hd__ha_1 _24717_ (.A(net3638),
    .B(net3727),
    .COUT(_12484_[0]),
    .SUM(_12485_[0]));
 sky130_fd_sc_hd__ha_1 _24718_ (.A(_02993_),
    .B(net3728),
    .COUT(_12486_[0]),
    .SUM(_12487_[0]));
 sky130_fd_sc_hd__ha_1 _24719_ (.A(net3638),
    .B(_02981_),
    .COUT(_12488_[0]),
    .SUM(_12489_[0]));
 sky130_fd_sc_hd__ha_1 _24720_ (.A(\u0.r0.rcnt_next[0] ),
    .B(_12490_[0]),
    .COUT(_12491_[0]),
    .SUM(\u0.r0.rcnt_next[1] ));
 sky130_fd_sc_hd__ha_1 _24721_ (.A(\u0.r0.rcnt_next[0] ),
    .B(\u0.r0.rcnt[1] ),
    .COUT(_12492_[0]),
    .SUM(_12493_[0]));
 sky130_fd_sc_hd__ha_1 _24722_ (.A(\u0.r0.rcnt[0] ),
    .B(_12490_[0]),
    .COUT(_12494_[0]),
    .SUM(_12495_[0]));
 sky130_fd_sc_hd__ha_1 _24723_ (.A(\u0.r0.rcnt[0] ),
    .B(\u0.r0.rcnt[1] ),
    .COUT(_12496_[0]),
    .SUM(_12497_[0]));
 sky130_fd_sc_hd__ha_1 _24724_ (.A(\u0.r0.rcnt[0] ),
    .B(\u0.r0.rcnt[1] ),
    .COUT(_12498_[0]),
    .SUM(_12499_[0]));
 sky130_fd_sc_hd__dfxtp_1 \dcnt[0]$_SDFFE_PN0P_  (.D(_00405_),
    .Q(\dcnt[0] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 \dcnt[1]$_SDFFE_PN0P_  (.D(_00406_),
    .Q(\dcnt[1] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 \dcnt[2]$_SDFFE_PP0P_  (.D(_00407_),
    .Q(\dcnt[2] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 \dcnt[3]$_SDFFE_PN0P_  (.D(_00408_),
    .Q(\dcnt[3] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 \done$_DFF_P_  (.D(_00160_),
    .Q(net259),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_2 \ld_r$_DFF_P_  (.D(net4236),
    .Q(ld_r),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa00_sr[0]$_DFF_P_  (.D(_00032_),
    .Q(\sa00_sr[0] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa00_sr[1]$_DFF_P_  (.D(_00033_),
    .Q(\sa00_sr[1] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa00_sr[2]$_DFF_P_  (.D(_00034_),
    .Q(\sa00_sr[2] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa00_sr[3]$_DFF_P_  (.D(_00035_),
    .Q(\sa00_sr[3] ),
    .CLK(clknet_3_6_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa00_sr[4]$_DFF_P_  (.D(_00036_),
    .Q(\sa00_sr[4] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa00_sr[5]$_DFF_P_  (.D(_00037_),
    .Q(\sa00_sr[5] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa00_sr[6]$_DFF_P_  (.D(_00038_),
    .Q(\sa00_sr[6] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa00_sr[7]$_DFF_P_  (.D(_00039_),
    .Q(\sa00_sr[7] ),
    .CLK(clknet_3_6_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa01_sr[0]$_DFF_P_  (.D(_00040_),
    .Q(\sa01_sr[0] ),
    .CLK(clknet_3_7_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa01_sr[1]$_DFF_P_  (.D(_00041_),
    .Q(\sa01_sr[1] ),
    .CLK(clknet_3_7_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa01_sr[2]$_DFF_P_  (.D(_00042_),
    .Q(\sa01_sr[2] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa01_sr[3]$_DFF_P_  (.D(_00043_),
    .Q(\sa01_sr[3] ),
    .CLK(clknet_3_7_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa01_sr[4]$_DFF_P_  (.D(_00044_),
    .Q(\sa01_sr[4] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa01_sr[5]$_DFF_P_  (.D(_00045_),
    .Q(\sa01_sr[5] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa01_sr[6]$_DFF_P_  (.D(_00046_),
    .Q(\sa01_sr[6] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa01_sr[7]$_DFF_P_  (.D(_00047_),
    .Q(\sa01_sr[7] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa02_sr[0]$_DFF_P_  (.D(_00048_),
    .Q(\sa02_sr[0] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa02_sr[1]$_DFF_P_  (.D(_00049_),
    .Q(\sa02_sr[1] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa02_sr[2]$_DFF_P_  (.D(_00050_),
    .Q(\sa02_sr[2] ),
    .CLK(clknet_3_5_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa02_sr[3]$_DFF_P_  (.D(net3564),
    .Q(\sa02_sr[3] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa02_sr[4]$_DFF_P_  (.D(_00052_),
    .Q(\sa02_sr[4] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa02_sr[5]$_DFF_P_  (.D(_00053_),
    .Q(\sa02_sr[5] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa02_sr[6]$_DFF_P_  (.D(_00054_),
    .Q(\sa02_sr[6] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa02_sr[7]$_DFF_P_  (.D(_00055_),
    .Q(\sa02_sr[7] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa03_sr[0]$_DFF_P_  (.D(_00056_),
    .Q(\sa03_sr[0] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa03_sr[1]$_DFF_P_  (.D(_00057_),
    .Q(\sa03_sr[1] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa03_sr[2]$_DFF_P_  (.D(_00058_),
    .Q(\sa03_sr[2] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa03_sr[3]$_DFF_P_  (.D(_00059_),
    .Q(\sa03_sr[3] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa03_sr[4]$_DFF_P_  (.D(_00060_),
    .Q(\sa03_sr[4] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa03_sr[5]$_DFF_P_  (.D(_00061_),
    .Q(\sa03_sr[5] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa03_sr[6]$_DFF_P_  (.D(_00062_),
    .Q(\sa03_sr[6] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa03_sr[7]$_DFF_P_  (.D(_00063_),
    .Q(\sa03_sr[7] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_2 \sa10_sr[0]$_DFF_P_  (.D(_00072_),
    .Q(\sa10_sr[0] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa10_sr[1]$_DFF_P_  (.D(_00073_),
    .Q(\sa10_sr[1] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa10_sr[2]$_DFF_P_  (.D(_00074_),
    .Q(\sa10_sr[2] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa10_sr[3]$_DFF_P_  (.D(_00075_),
    .Q(\sa10_sr[3] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa10_sr[4]$_DFF_P_  (.D(_00076_),
    .Q(\sa10_sr[4] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa10_sr[5]$_DFF_P_  (.D(_00077_),
    .Q(\sa10_sr[5] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa10_sr[6]$_DFF_P_  (.D(_00078_),
    .Q(\sa10_sr[6] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa10_sr[7]$_DFF_P_  (.D(_00079_),
    .Q(\sa10_sr[7] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa11_sr[0]$_DFF_P_  (.D(_00080_),
    .Q(\sa11_sr[0] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa11_sr[1]$_DFF_P_  (.D(net3563),
    .Q(\sa11_sr[1] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa11_sr[2]$_DFF_P_  (.D(_00082_),
    .Q(\sa11_sr[2] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa11_sr[3]$_DFF_P_  (.D(_00083_),
    .Q(\sa11_sr[3] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa11_sr[4]$_DFF_P_  (.D(_00084_),
    .Q(\sa11_sr[4] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa11_sr[5]$_DFF_P_  (.D(_00085_),
    .Q(\sa11_sr[5] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa11_sr[6]$_DFF_P_  (.D(_00086_),
    .Q(\sa11_sr[6] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa11_sr[7]$_DFF_P_  (.D(_00087_),
    .Q(\sa11_sr[7] ),
    .CLK(clknet_3_5_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa12_sr[0]$_DFF_P_  (.D(_00088_),
    .Q(\sa12_sr[0] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa12_sr[1]$_DFF_P_  (.D(_00089_),
    .Q(\sa12_sr[1] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa12_sr[2]$_DFF_P_  (.D(_00090_),
    .Q(\sa12_sr[2] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa12_sr[3]$_DFF_P_  (.D(_00091_),
    .Q(\sa12_sr[3] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa12_sr[4]$_DFF_P_  (.D(_00092_),
    .Q(\sa12_sr[4] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa12_sr[5]$_DFF_P_  (.D(_00093_),
    .Q(\sa12_sr[5] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa12_sr[6]$_DFF_P_  (.D(_00094_),
    .Q(\sa12_sr[6] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa12_sr[7]$_DFF_P_  (.D(_00095_),
    .Q(\sa12_sr[7] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa13_sr[0]$_DFF_P_  (.D(_00064_),
    .Q(\sa10_sub[0] ),
    .CLK(clknet_3_2_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa13_sr[1]$_DFF_P_  (.D(_00065_),
    .Q(\sa10_sub[1] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa13_sr[2]$_DFF_P_  (.D(_00066_),
    .Q(\sa10_sub[2] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa13_sr[3]$_DFF_P_  (.D(_00067_),
    .Q(\sa10_sub[3] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa13_sr[4]$_DFF_P_  (.D(_00068_),
    .Q(\sa10_sub[4] ),
    .CLK(clknet_3_2_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa13_sr[5]$_DFF_P_  (.D(_00069_),
    .Q(\sa10_sub[5] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa13_sr[6]$_DFF_P_  (.D(_00070_),
    .Q(\sa10_sub[6] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa13_sr[7]$_DFF_P_  (.D(_00071_),
    .Q(\sa10_sub[7] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa20_sr[0]$_DFF_P_  (.D(_00112_),
    .Q(\sa20_sr[0] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa20_sr[1]$_DFF_P_  (.D(_00113_),
    .Q(\sa20_sr[1] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa20_sr[2]$_DFF_P_  (.D(_00114_),
    .Q(\sa20_sr[2] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa20_sr[3]$_DFF_P_  (.D(_00115_),
    .Q(\sa20_sr[3] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa20_sr[4]$_DFF_P_  (.D(_00116_),
    .Q(\sa20_sr[4] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa20_sr[5]$_DFF_P_  (.D(_00117_),
    .Q(\sa20_sr[5] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa20_sr[6]$_DFF_P_  (.D(net3562),
    .Q(\sa20_sr[6] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa20_sr[7]$_DFF_P_  (.D(_00119_),
    .Q(\sa20_sr[7] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa21_sr[0]$_DFF_P_  (.D(_00120_),
    .Q(\sa21_sr[0] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa21_sr[1]$_DFF_P_  (.D(_00121_),
    .Q(\sa21_sr[1] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa21_sr[2]$_DFF_P_  (.D(_00122_),
    .Q(\sa21_sr[2] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa21_sr[3]$_DFF_P_  (.D(_00123_),
    .Q(\sa21_sr[3] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa21_sr[4]$_DFF_P_  (.D(_00124_),
    .Q(\sa21_sr[4] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa21_sr[5]$_DFF_P_  (.D(_00125_),
    .Q(\sa21_sr[5] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa21_sr[6]$_DFF_P_  (.D(_00126_),
    .Q(\sa21_sr[6] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa21_sr[7]$_DFF_P_  (.D(_00127_),
    .Q(\sa21_sr[7] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa22_sr[0]$_DFF_P_  (.D(_00096_),
    .Q(\sa20_sub[0] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa22_sr[1]$_DFF_P_  (.D(net3561),
    .Q(\sa20_sub[1] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa22_sr[2]$_DFF_P_  (.D(_00098_),
    .Q(\sa20_sub[2] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa22_sr[3]$_DFF_P_  (.D(_00099_),
    .Q(\sa20_sub[3] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa22_sr[4]$_DFF_P_  (.D(_00100_),
    .Q(\sa20_sub[4] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa22_sr[5]$_DFF_P_  (.D(_00101_),
    .Q(\sa20_sub[5] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa22_sr[6]$_DFF_P_  (.D(_00102_),
    .Q(\sa20_sub[6] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa22_sr[7]$_DFF_P_  (.D(_00103_),
    .Q(\sa20_sub[7] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa23_sr[0]$_DFF_P_  (.D(_00104_),
    .Q(\sa21_sub[0] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa23_sr[1]$_DFF_P_  (.D(net3560),
    .Q(\sa21_sub[1] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa23_sr[2]$_DFF_P_  (.D(_00106_),
    .Q(\sa21_sub[2] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa23_sr[3]$_DFF_P_  (.D(_00107_),
    .Q(\sa21_sub[3] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa23_sr[4]$_DFF_P_  (.D(_00108_),
    .Q(\sa21_sub[4] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa23_sr[5]$_DFF_P_  (.D(_00109_),
    .Q(\sa21_sub[5] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa23_sr[6]$_DFF_P_  (.D(_00110_),
    .Q(\sa21_sub[6] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa23_sr[7]$_DFF_P_  (.D(_00111_),
    .Q(\sa21_sub[7] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa30_sr[0]$_DFF_P_  (.D(_00152_),
    .Q(\sa30_sr[0] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa30_sr[1]$_DFF_P_  (.D(_00153_),
    .Q(\sa30_sr[1] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa30_sr[2]$_DFF_P_  (.D(_00154_),
    .Q(\sa30_sr[2] ),
    .CLK(clknet_3_3_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa30_sr[3]$_DFF_P_  (.D(_00155_),
    .Q(\sa30_sr[3] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa30_sr[4]$_DFF_P_  (.D(_00156_),
    .Q(\sa30_sr[4] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa30_sr[5]$_DFF_P_  (.D(_00157_),
    .Q(\sa30_sr[5] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa30_sr[6]$_DFF_P_  (.D(_00158_),
    .Q(\sa30_sr[6] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa30_sr[7]$_DFF_P_  (.D(_00159_),
    .Q(\sa30_sr[7] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa31_sr[0]$_DFF_P_  (.D(_00128_),
    .Q(\sa30_sub[0] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa31_sr[1]$_DFF_P_  (.D(_00129_),
    .Q(\sa30_sub[1] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa31_sr[2]$_DFF_P_  (.D(_00130_),
    .Q(\sa30_sub[2] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa31_sr[3]$_DFF_P_  (.D(_00131_),
    .Q(\sa30_sub[3] ),
    .CLK(clknet_3_5_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa31_sr[4]$_DFF_P_  (.D(_00132_),
    .Q(\sa30_sub[4] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa31_sr[5]$_DFF_P_  (.D(_00133_),
    .Q(\sa30_sub[5] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa31_sr[6]$_DFF_P_  (.D(_00134_),
    .Q(\sa30_sub[6] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa31_sr[7]$_DFF_P_  (.D(_00135_),
    .Q(\sa30_sub[7] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa32_sr[0]$_DFF_P_  (.D(_00136_),
    .Q(\sa31_sub[0] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa32_sr[1]$_DFF_P_  (.D(_00137_),
    .Q(\sa31_sub[1] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa32_sr[2]$_DFF_P_  (.D(_00138_),
    .Q(\sa31_sub[2] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa32_sr[3]$_DFF_P_  (.D(_00139_),
    .Q(\sa31_sub[3] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa32_sr[4]$_DFF_P_  (.D(_00140_),
    .Q(\sa31_sub[4] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa32_sr[5]$_DFF_P_  (.D(_00141_),
    .Q(\sa31_sub[5] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa32_sr[6]$_DFF_P_  (.D(_00142_),
    .Q(\sa31_sub[6] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa32_sr[7]$_DFF_P_  (.D(_00143_),
    .Q(\sa31_sub[7] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa33_sr[0]$_DFF_P_  (.D(_00144_),
    .Q(\sa32_sub[0] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa33_sr[1]$_DFF_P_  (.D(_00145_),
    .Q(\sa32_sub[1] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa33_sr[2]$_DFF_P_  (.D(_00146_),
    .Q(\sa32_sub[2] ),
    .CLK(clknet_3_0_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa33_sr[3]$_DFF_P_  (.D(_00147_),
    .Q(\sa32_sub[3] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa33_sr[4]$_DFF_P_  (.D(_00148_),
    .Q(\sa32_sub[4] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa33_sr[5]$_DFF_P_  (.D(_00149_),
    .Q(\sa32_sub[5] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa33_sr[6]$_DFF_P_  (.D(_00150_),
    .Q(\sa32_sub[6] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__dfxtp_1 \sa33_sr[7]$_DFF_P_  (.D(_00151_),
    .Q(\sa32_sub[7] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[0]$_DFFE_PP_  (.D(net131),
    .DE(net4233),
    .Q(\text_in_r[0] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[100]$_DFFE_PP_  (.D(net132),
    .DE(net4236),
    .Q(\text_in_r[100] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[101]$_DFFE_PP_  (.D(net133),
    .DE(net4236),
    .Q(\text_in_r[101] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[102]$_DFFE_PP_  (.D(net134),
    .DE(net4236),
    .Q(\text_in_r[102] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[103]$_DFFE_PP_  (.D(net135),
    .DE(net4236),
    .Q(\text_in_r[103] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[104]$_DFFE_PP_  (.D(net136),
    .DE(net4240),
    .Q(\text_in_r[104] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[105]$_DFFE_PP_  (.D(net137),
    .DE(net4236),
    .Q(\text_in_r[105] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[106]$_DFFE_PP_  (.D(net138),
    .DE(net4236),
    .Q(\text_in_r[106] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[107]$_DFFE_PP_  (.D(net139),
    .DE(net4236),
    .Q(\text_in_r[107] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[108]$_DFFE_PP_  (.D(net140),
    .DE(net4236),
    .Q(\text_in_r[108] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[109]$_DFFE_PP_  (.D(net141),
    .DE(net4236),
    .Q(\text_in_r[109] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[10]$_DFFE_PP_  (.D(net142),
    .DE(net4234),
    .Q(\text_in_r[10] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[110]$_DFFE_PP_  (.D(net143),
    .DE(net4236),
    .Q(\text_in_r[110] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[111]$_DFFE_PP_  (.D(net144),
    .DE(net4236),
    .Q(\text_in_r[111] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[112]$_DFFE_PP_  (.D(net145),
    .DE(net4237),
    .Q(\text_in_r[112] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[113]$_DFFE_PP_  (.D(net146),
    .DE(net4239),
    .Q(\text_in_r[113] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[114]$_DFFE_PP_  (.D(net147),
    .DE(net4238),
    .Q(\text_in_r[114] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[115]$_DFFE_PP_  (.D(net148),
    .DE(net4238),
    .Q(\text_in_r[115] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[116]$_DFFE_PP_  (.D(net149),
    .DE(net4238),
    .Q(\text_in_r[116] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[117]$_DFFE_PP_  (.D(net150),
    .DE(net4238),
    .Q(\text_in_r[117] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[118]$_DFFE_PP_  (.D(net151),
    .DE(net4238),
    .Q(\text_in_r[118] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[119]$_DFFE_PP_  (.D(net152),
    .DE(net4239),
    .Q(\text_in_r[119] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[11]$_DFFE_PP_  (.D(net153),
    .DE(net4237),
    .Q(\text_in_r[11] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[120]$_DFFE_PP_  (.D(net154),
    .DE(net4240),
    .Q(\text_in_r[120] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[121]$_DFFE_PP_  (.D(net155),
    .DE(net4236),
    .Q(\text_in_r[121] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[122]$_DFFE_PP_  (.D(net156),
    .DE(net4236),
    .Q(\text_in_r[122] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[123]$_DFFE_PP_  (.D(net157),
    .DE(net4236),
    .Q(\text_in_r[123] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[124]$_DFFE_PP_  (.D(net158),
    .DE(net4236),
    .Q(\text_in_r[124] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[125]$_DFFE_PP_  (.D(net159),
    .DE(net4236),
    .Q(\text_in_r[125] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[126]$_DFFE_PP_  (.D(net160),
    .DE(net4236),
    .Q(\text_in_r[126] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[127]$_DFFE_PP_  (.D(net161),
    .DE(net4236),
    .Q(\text_in_r[127] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[12]$_DFFE_PP_  (.D(net162),
    .DE(net4234),
    .Q(\text_in_r[12] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[13]$_DFFE_PP_  (.D(net163),
    .DE(net4237),
    .Q(\text_in_r[13] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[14]$_DFFE_PP_  (.D(net164),
    .DE(net4234),
    .Q(\text_in_r[14] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[15]$_DFFE_PP_  (.D(net165),
    .DE(net4237),
    .Q(\text_in_r[15] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[16]$_DFFE_PP_  (.D(net166),
    .DE(net4233),
    .Q(\text_in_r[16] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[17]$_DFFE_PP_  (.D(net167),
    .DE(net4233),
    .Q(\text_in_r[17] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[18]$_DFFE_PP_  (.D(net168),
    .DE(net4233),
    .Q(\text_in_r[18] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[19]$_DFFE_PP_  (.D(net169),
    .DE(net4233),
    .Q(\text_in_r[19] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[1]$_DFFE_PP_  (.D(net170),
    .DE(net4233),
    .Q(\text_in_r[1] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[20]$_DFFE_PP_  (.D(net171),
    .DE(net4233),
    .Q(\text_in_r[20] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[21]$_DFFE_PP_  (.D(net172),
    .DE(net4233),
    .Q(\text_in_r[21] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[22]$_DFFE_PP_  (.D(net173),
    .DE(net4233),
    .Q(\text_in_r[22] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[23]$_DFFE_PP_  (.D(net174),
    .DE(net4233),
    .Q(\text_in_r[23] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[24]$_DFFE_PP_  (.D(net175),
    .DE(net4233),
    .Q(\text_in_r[24] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[25]$_DFFE_PP_  (.D(net176),
    .DE(net4233),
    .Q(\text_in_r[25] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[26]$_DFFE_PP_  (.D(net177),
    .DE(net4233),
    .Q(\text_in_r[26] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[27]$_DFFE_PP_  (.D(net178),
    .DE(net4233),
    .Q(\text_in_r[27] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[28]$_DFFE_PP_  (.D(net179),
    .DE(net4233),
    .Q(\text_in_r[28] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[29]$_DFFE_PP_  (.D(net180),
    .DE(net4233),
    .Q(\text_in_r[29] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[2]$_DFFE_PP_  (.D(net181),
    .DE(net4233),
    .Q(\text_in_r[2] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[30]$_DFFE_PP_  (.D(net182),
    .DE(net4233),
    .Q(\text_in_r[30] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[31]$_DFFE_PP_  (.D(net183),
    .DE(net4233),
    .Q(\text_in_r[31] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[32]$_DFFE_PP_  (.D(net184),
    .DE(net4232),
    .Q(\text_in_r[32] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[33]$_DFFE_PP_  (.D(net185),
    .DE(net129),
    .Q(\text_in_r[33] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[34]$_DFFE_PP_  (.D(net186),
    .DE(net4232),
    .Q(\text_in_r[34] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[35]$_DFFE_PP_  (.D(net187),
    .DE(net129),
    .Q(\text_in_r[35] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[36]$_DFFE_PP_  (.D(net188),
    .DE(net4232),
    .Q(\text_in_r[36] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[37]$_DFFE_PP_  (.D(net189),
    .DE(net129),
    .Q(\text_in_r[37] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[38]$_DFFE_PP_  (.D(net190),
    .DE(net4232),
    .Q(\text_in_r[38] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[39]$_DFFE_PP_  (.D(net191),
    .DE(net129),
    .Q(\text_in_r[39] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[3]$_DFFE_PP_  (.D(net192),
    .DE(net4233),
    .Q(\text_in_r[3] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[40]$_DFFE_PP_  (.D(net193),
    .DE(net4235),
    .Q(\text_in_r[40] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[41]$_DFFE_PP_  (.D(net194),
    .DE(net4235),
    .Q(\text_in_r[41] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[42]$_DFFE_PP_  (.D(net195),
    .DE(net4235),
    .Q(\text_in_r[42] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[43]$_DFFE_PP_  (.D(net196),
    .DE(net4236),
    .Q(\text_in_r[43] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[44]$_DFFE_PP_  (.D(net197),
    .DE(net4236),
    .Q(\text_in_r[44] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[45]$_DFFE_PP_  (.D(net198),
    .DE(net4236),
    .Q(\text_in_r[45] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[46]$_DFFE_PP_  (.D(net199),
    .DE(net4235),
    .Q(\text_in_r[46] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[47]$_DFFE_PP_  (.D(net200),
    .DE(net4236),
    .Q(\text_in_r[47] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[48]$_DFFE_PP_  (.D(net201),
    .DE(net4232),
    .Q(\text_in_r[48] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[49]$_DFFE_PP_  (.D(net202),
    .DE(net4232),
    .Q(\text_in_r[49] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[4]$_DFFE_PP_  (.D(net203),
    .DE(net4234),
    .Q(\text_in_r[4] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[50]$_DFFE_PP_  (.D(net204),
    .DE(net4232),
    .Q(\text_in_r[50] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[51]$_DFFE_PP_  (.D(net205),
    .DE(net4235),
    .Q(\text_in_r[51] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[52]$_DFFE_PP_  (.D(net206),
    .DE(net4235),
    .Q(\text_in_r[52] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[53]$_DFFE_PP_  (.D(net207),
    .DE(net4235),
    .Q(\text_in_r[53] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[54]$_DFFE_PP_  (.D(net208),
    .DE(net4235),
    .Q(\text_in_r[54] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[55]$_DFFE_PP_  (.D(net209),
    .DE(net4232),
    .Q(\text_in_r[55] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[56]$_DFFE_PP_  (.D(net210),
    .DE(net4232),
    .Q(\text_in_r[56] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[57]$_DFFE_PP_  (.D(net211),
    .DE(net4232),
    .Q(\text_in_r[57] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[58]$_DFFE_PP_  (.D(net212),
    .DE(net4232),
    .Q(\text_in_r[58] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[59]$_DFFE_PP_  (.D(net213),
    .DE(net4232),
    .Q(\text_in_r[59] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[5]$_DFFE_PP_  (.D(net214),
    .DE(net4233),
    .Q(\text_in_r[5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[60]$_DFFE_PP_  (.D(net215),
    .DE(net4232),
    .Q(\text_in_r[60] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[61]$_DFFE_PP_  (.D(net216),
    .DE(net4235),
    .Q(\text_in_r[61] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[62]$_DFFE_PP_  (.D(net217),
    .DE(net4232),
    .Q(\text_in_r[62] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[63]$_DFFE_PP_  (.D(net218),
    .DE(net4232),
    .Q(\text_in_r[63] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[64]$_DFFE_PP_  (.D(net219),
    .DE(net4236),
    .Q(\text_in_r[64] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[65]$_DFFE_PP_  (.D(net220),
    .DE(net4236),
    .Q(\text_in_r[65] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[66]$_DFFE_PP_  (.D(net221),
    .DE(net4236),
    .Q(\text_in_r[66] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[67]$_DFFE_PP_  (.D(net222),
    .DE(net4235),
    .Q(\text_in_r[67] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[68]$_DFFE_PP_  (.D(net223),
    .DE(net4236),
    .Q(\text_in_r[68] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[69]$_DFFE_PP_  (.D(net224),
    .DE(net4236),
    .Q(\text_in_r[69] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[6]$_DFFE_PP_  (.D(net225),
    .DE(net4234),
    .Q(\text_in_r[6] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[70]$_DFFE_PP_  (.D(net226),
    .DE(net4235),
    .Q(\text_in_r[70] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[71]$_DFFE_PP_  (.D(net227),
    .DE(net4235),
    .Q(\text_in_r[71] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[72]$_DFFE_PP_  (.D(net228),
    .DE(net4240),
    .Q(\text_in_r[72] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[73]$_DFFE_PP_  (.D(net229),
    .DE(net4236),
    .Q(\text_in_r[73] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[74]$_DFFE_PP_  (.D(net230),
    .DE(net4237),
    .Q(\text_in_r[74] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[75]$_DFFE_PP_  (.D(net231),
    .DE(net4237),
    .Q(\text_in_r[75] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[76]$_DFFE_PP_  (.D(net232),
    .DE(net4238),
    .Q(\text_in_r[76] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[77]$_DFFE_PP_  (.D(net233),
    .DE(net4239),
    .Q(\text_in_r[77] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[78]$_DFFE_PP_  (.D(net234),
    .DE(net4237),
    .Q(\text_in_r[78] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[79]$_DFFE_PP_  (.D(net235),
    .DE(net4239),
    .Q(\text_in_r[79] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[7]$_DFFE_PP_  (.D(net236),
    .DE(net4234),
    .Q(\text_in_r[7] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[80]$_DFFE_PP_  (.D(net237),
    .DE(net4236),
    .Q(\text_in_r[80] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[81]$_DFFE_PP_  (.D(net238),
    .DE(net4236),
    .Q(\text_in_r[81] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[82]$_DFFE_PP_  (.D(net239),
    .DE(net4236),
    .Q(\text_in_r[82] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[83]$_DFFE_PP_  (.D(net240),
    .DE(net4236),
    .Q(\text_in_r[83] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[84]$_DFFE_PP_  (.D(net241),
    .DE(net4236),
    .Q(\text_in_r[84] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[85]$_DFFE_PP_  (.D(net242),
    .DE(net4236),
    .Q(\text_in_r[85] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[86]$_DFFE_PP_  (.D(net243),
    .DE(net4236),
    .Q(\text_in_r[86] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[87]$_DFFE_PP_  (.D(net244),
    .DE(net4236),
    .Q(\text_in_r[87] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[88]$_DFFE_PP_  (.D(net245),
    .DE(net4236),
    .Q(\text_in_r[88] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[89]$_DFFE_PP_  (.D(net246),
    .DE(net4236),
    .Q(\text_in_r[89] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[8]$_DFFE_PP_  (.D(net247),
    .DE(net4234),
    .Q(\text_in_r[8] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[90]$_DFFE_PP_  (.D(net248),
    .DE(net4236),
    .Q(\text_in_r[90] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[91]$_DFFE_PP_  (.D(net249),
    .DE(net4236),
    .Q(\text_in_r[91] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[92]$_DFFE_PP_  (.D(net250),
    .DE(net4236),
    .Q(\text_in_r[92] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[93]$_DFFE_PP_  (.D(net251),
    .DE(net4236),
    .Q(\text_in_r[93] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[94]$_DFFE_PP_  (.D(net252),
    .DE(net4236),
    .Q(\text_in_r[94] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[95]$_DFFE_PP_  (.D(net253),
    .DE(net4236),
    .Q(\text_in_r[95] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[96]$_DFFE_PP_  (.D(net254),
    .DE(net4236),
    .Q(\text_in_r[96] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[97]$_DFFE_PP_  (.D(net255),
    .DE(net4240),
    .Q(\text_in_r[97] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[98]$_DFFE_PP_  (.D(net256),
    .DE(net4236),
    .Q(\text_in_r[98] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[99]$_DFFE_PP_  (.D(net257),
    .DE(net4236),
    .Q(\text_in_r[99] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \text_in_r[9]$_DFFE_PP_  (.D(net258),
    .DE(net4237),
    .Q(\text_in_r[9] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[0]$_DFF_P_  (.D(_00265_),
    .Q(net260),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[100]$_DFF_P_  (.D(_00165_),
    .Q(net261),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[101]$_DFF_P_  (.D(_00166_),
    .Q(net262),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[102]$_DFF_P_  (.D(_00167_),
    .Q(net263),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[103]$_DFF_P_  (.D(_00168_),
    .Q(net264),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[104]$_DFF_P_  (.D(_00169_),
    .Q(net265),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[105]$_DFF_P_  (.D(_00170_),
    .Q(net266),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[106]$_DFF_P_  (.D(_00171_),
    .Q(net267),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[107]$_DFF_P_  (.D(_00172_),
    .Q(net268),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[108]$_DFF_P_  (.D(_00173_),
    .Q(net269),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[109]$_DFF_P_  (.D(_00174_),
    .Q(net270),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[10]$_DFF_P_  (.D(_00195_),
    .Q(net271),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[110]$_DFF_P_  (.D(_00175_),
    .Q(net272),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[111]$_DFF_P_  (.D(_00176_),
    .Q(net273),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[112]$_DFF_P_  (.D(_00177_),
    .Q(net274),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[113]$_DFF_P_  (.D(_00178_),
    .Q(net275),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[114]$_DFF_P_  (.D(_00179_),
    .Q(net276),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[115]$_DFF_P_  (.D(_00180_),
    .Q(net277),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[116]$_DFF_P_  (.D(_00181_),
    .Q(net278),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[117]$_DFF_P_  (.D(_00182_),
    .Q(net279),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[118]$_DFF_P_  (.D(_00183_),
    .Q(net280),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[119]$_DFF_P_  (.D(_00184_),
    .Q(net281),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[11]$_DFF_P_  (.D(_00196_),
    .Q(net282),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[120]$_DFF_P_  (.D(_00185_),
    .Q(net283),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[121]$_DFF_P_  (.D(_00186_),
    .Q(net284),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[122]$_DFF_P_  (.D(_00187_),
    .Q(net285),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[123]$_DFF_P_  (.D(_00188_),
    .Q(net286),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[124]$_DFF_P_  (.D(_00189_),
    .Q(net287),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[125]$_DFF_P_  (.D(_00190_),
    .Q(net288),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[126]$_DFF_P_  (.D(_00191_),
    .Q(net289),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[127]$_DFF_P_  (.D(_00192_),
    .Q(net290),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[12]$_DFF_P_  (.D(_00197_),
    .Q(net291),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[13]$_DFF_P_  (.D(_00198_),
    .Q(net292),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[14]$_DFF_P_  (.D(_00199_),
    .Q(net293),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[15]$_DFF_P_  (.D(_00200_),
    .Q(net294),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[16]$_DFF_P_  (.D(_00201_),
    .Q(net295),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[17]$_DFF_P_  (.D(_00202_),
    .Q(net296),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[18]$_DFF_P_  (.D(_00203_),
    .Q(net297),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[19]$_DFF_P_  (.D(_00204_),
    .Q(net298),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[1]$_DFF_P_  (.D(_00266_),
    .Q(net299),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[20]$_DFF_P_  (.D(_00205_),
    .Q(net300),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[21]$_DFF_P_  (.D(_00206_),
    .Q(net301),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[22]$_DFF_P_  (.D(_00207_),
    .Q(net302),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[23]$_DFF_P_  (.D(_00208_),
    .Q(net303),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[24]$_DFF_P_  (.D(_00209_),
    .Q(net304),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[25]$_DFF_P_  (.D(_00210_),
    .Q(net305),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[26]$_DFF_P_  (.D(_00211_),
    .Q(net306),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[27]$_DFF_P_  (.D(_00212_),
    .Q(net307),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[28]$_DFF_P_  (.D(_00213_),
    .Q(net308),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[29]$_DFF_P_  (.D(_00214_),
    .Q(net309),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[2]$_DFF_P_  (.D(_00267_),
    .Q(net310),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[30]$_DFF_P_  (.D(_00215_),
    .Q(net311),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[31]$_DFF_P_  (.D(_00216_),
    .Q(net312),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[32]$_DFF_P_  (.D(_00217_),
    .Q(net313),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[33]$_DFF_P_  (.D(_00218_),
    .Q(net314),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[34]$_DFF_P_  (.D(_00219_),
    .Q(net315),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[35]$_DFF_P_  (.D(_00220_),
    .Q(net316),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[36]$_DFF_P_  (.D(_00221_),
    .Q(net317),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[37]$_DFF_P_  (.D(_00222_),
    .Q(net318),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[38]$_DFF_P_  (.D(_00223_),
    .Q(net319),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[39]$_DFF_P_  (.D(_00224_),
    .Q(net320),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[3]$_DFF_P_  (.D(_00268_),
    .Q(net321),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[40]$_DFF_P_  (.D(_00225_),
    .Q(net322),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[41]$_DFF_P_  (.D(_00226_),
    .Q(net323),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[42]$_DFF_P_  (.D(_00227_),
    .Q(net324),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[43]$_DFF_P_  (.D(_00228_),
    .Q(net325),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[44]$_DFF_P_  (.D(_00229_),
    .Q(net326),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[45]$_DFF_P_  (.D(_00230_),
    .Q(net327),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[46]$_DFF_P_  (.D(_00231_),
    .Q(net328),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[47]$_DFF_P_  (.D(_00232_),
    .Q(net329),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[48]$_DFF_P_  (.D(_00233_),
    .Q(net330),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[49]$_DFF_P_  (.D(_00234_),
    .Q(net331),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[4]$_DFF_P_  (.D(_00269_),
    .Q(net332),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[50]$_DFF_P_  (.D(_00235_),
    .Q(net333),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[51]$_DFF_P_  (.D(_00236_),
    .Q(net334),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[52]$_DFF_P_  (.D(_00237_),
    .Q(net335),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[53]$_DFF_P_  (.D(_00238_),
    .Q(net336),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[54]$_DFF_P_  (.D(_00239_),
    .Q(net337),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[55]$_DFF_P_  (.D(_00240_),
    .Q(net338),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[56]$_DFF_P_  (.D(_00241_),
    .Q(net339),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[57]$_DFF_P_  (.D(_00242_),
    .Q(net340),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[58]$_DFF_P_  (.D(_00243_),
    .Q(net341),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[59]$_DFF_P_  (.D(_00244_),
    .Q(net342),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[5]$_DFF_P_  (.D(_00270_),
    .Q(net343),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[60]$_DFF_P_  (.D(_00245_),
    .Q(net344),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[61]$_DFF_P_  (.D(_00246_),
    .Q(net345),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[62]$_DFF_P_  (.D(_00247_),
    .Q(net346),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[63]$_DFF_P_  (.D(_00248_),
    .Q(net347),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[64]$_DFF_P_  (.D(_00249_),
    .Q(net348),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[65]$_DFF_P_  (.D(_00250_),
    .Q(net349),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[66]$_DFF_P_  (.D(_00251_),
    .Q(net350),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[67]$_DFF_P_  (.D(_00252_),
    .Q(net351),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[68]$_DFF_P_  (.D(_00253_),
    .Q(net352),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[69]$_DFF_P_  (.D(_00254_),
    .Q(net353),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[6]$_DFF_P_  (.D(_00271_),
    .Q(net354),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[70]$_DFF_P_  (.D(_00255_),
    .Q(net355),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[71]$_DFF_P_  (.D(_00256_),
    .Q(net356),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[72]$_DFF_P_  (.D(_00257_),
    .Q(net357),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[73]$_DFF_P_  (.D(_00258_),
    .Q(net358),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[74]$_DFF_P_  (.D(_00259_),
    .Q(net359),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[75]$_DFF_P_  (.D(_00260_),
    .Q(net360),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[76]$_DFF_P_  (.D(_00261_),
    .Q(net361),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[77]$_DFF_P_  (.D(_00262_),
    .Q(net362),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[78]$_DFF_P_  (.D(_00263_),
    .Q(net363),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[79]$_DFF_P_  (.D(_00264_),
    .Q(net364),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[7]$_DFF_P_  (.D(_00272_),
    .Q(net365),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[80]$_DFF_P_  (.D(_00273_),
    .Q(net366),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[81]$_DFF_P_  (.D(_00274_),
    .Q(net367),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[82]$_DFF_P_  (.D(_00275_),
    .Q(net368),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[83]$_DFF_P_  (.D(_00276_),
    .Q(net369),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[84]$_DFF_P_  (.D(_00277_),
    .Q(net370),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[85]$_DFF_P_  (.D(_00278_),
    .Q(net371),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[86]$_DFF_P_  (.D(_00279_),
    .Q(net372),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[87]$_DFF_P_  (.D(_00280_),
    .Q(net373),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[88]$_DFF_P_  (.D(_00281_),
    .Q(net374),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[89]$_DFF_P_  (.D(_00282_),
    .Q(net375),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[8]$_DFF_P_  (.D(_00193_),
    .Q(net376),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[90]$_DFF_P_  (.D(_00283_),
    .Q(net377),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[91]$_DFF_P_  (.D(_00284_),
    .Q(net378),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[92]$_DFF_P_  (.D(_00285_),
    .Q(net379),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[93]$_DFF_P_  (.D(_00286_),
    .Q(net380),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[94]$_DFF_P_  (.D(_00287_),
    .Q(net381),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[95]$_DFF_P_  (.D(_00288_),
    .Q(net382),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[96]$_DFF_P_  (.D(_00161_),
    .Q(net383),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[97]$_DFF_P_  (.D(_00162_),
    .Q(net384),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[98]$_DFF_P_  (.D(_00163_),
    .Q(net385),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[99]$_DFF_P_  (.D(_00164_),
    .Q(net386),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__dfxtp_1 \text_out[9]$_DFF_P_  (.D(_00194_),
    .Q(net387),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.r0.out[24]$_SDFF_PP1_  (.D(_00409_),
    .Q(\u0.r0.out[24] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.r0.out[25]$_SDFF_PP0_  (.D(_00410_),
    .Q(\u0.r0.out[25] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.r0.out[26]$_SDFF_PP0_  (.D(_00411_),
    .Q(\u0.r0.out[26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.r0.out[27]$_SDFF_PP0_  (.D(_00412_),
    .Q(\u0.r0.out[27] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.r0.out[28]$_SDFF_PP0_  (.D(_00413_),
    .Q(\u0.r0.out[28] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.r0.out[29]$_SDFF_PP0_  (.D(_00414_),
    .Q(\u0.r0.out[29] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.r0.out[30]$_SDFF_PP0_  (.D(_00415_),
    .Q(\u0.r0.out[30] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.r0.out[31]$_SDFF_PP0_  (.D(_00416_),
    .Q(\u0.r0.out[31] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.r0.rcnt[0]$_SDFF_PP0_  (.D(_00417_),
    .Q(\u0.r0.rcnt[0] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.r0.rcnt[1]$_SDFF_PP0_  (.D(_00418_),
    .Q(\u0.r0.rcnt[1] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.r0.rcnt[2]$_SDFF_PP0_  (.D(_00419_),
    .Q(\u0.r0.rcnt[2] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.r0.rcnt[3]$_SDFF_PP0_  (.D(_00420_),
    .Q(\u0.r0.rcnt[3] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u0.d[0]$_DFF_P_  (.D(_00000_),
    .Q(\u0.subword[24] ),
    .CLK(clknet_3_2_0_clk));
 sky130_fd_sc_hd__dfxtp_2 \u0.u0.d[1]$_DFF_P_  (.D(_00001_),
    .Q(\u0.subword[25] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u0.d[2]$_DFF_P_  (.D(_00002_),
    .Q(\u0.subword[26] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_2 \u0.u0.d[3]$_DFF_P_  (.D(_00003_),
    .Q(\u0.subword[27] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u0.d[4]$_DFF_P_  (.D(_00004_),
    .Q(\u0.subword[28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u0.d[5]$_DFF_P_  (.D(_00005_),
    .Q(\u0.subword[29] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u0.d[6]$_DFF_P_  (.D(_00006_),
    .Q(\u0.subword[30] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u0.d[7]$_DFF_P_  (.D(_00007_),
    .Q(\u0.subword[31] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u1.d[0]$_DFF_P_  (.D(_00008_),
    .Q(\u0.subword[16] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u1.d[1]$_DFF_P_  (.D(_00009_),
    .Q(\u0.subword[17] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u1.d[2]$_DFF_P_  (.D(_00010_),
    .Q(\u0.subword[18] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u1.d[3]$_DFF_P_  (.D(_00011_),
    .Q(\u0.subword[19] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u1.d[4]$_DFF_P_  (.D(_00012_),
    .Q(\u0.subword[20] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u1.d[5]$_DFF_P_  (.D(_00013_),
    .Q(\u0.subword[21] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u1.d[6]$_DFF_P_  (.D(_00014_),
    .Q(\u0.subword[22] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u1.d[7]$_DFF_P_  (.D(_00015_),
    .Q(\u0.subword[23] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u2.d[0]$_DFF_P_  (.D(_00016_),
    .Q(\u0.subword[8] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u2.d[1]$_DFF_P_  (.D(net3567),
    .Q(\u0.subword[9] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u2.d[2]$_DFF_P_  (.D(_00018_),
    .Q(\u0.subword[10] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u2.d[3]$_DFF_P_  (.D(_00019_),
    .Q(\u0.subword[11] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u2.d[4]$_DFF_P_  (.D(_00020_),
    .Q(\u0.subword[12] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u2.d[5]$_DFF_P_  (.D(net3566),
    .Q(\u0.subword[13] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u2.d[6]$_DFF_P_  (.D(_00022_),
    .Q(\u0.subword[14] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u2.d[7]$_DFF_P_  (.D(_00023_),
    .Q(\u0.subword[15] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u3.d[0]$_DFF_P_  (.D(_00024_),
    .Q(\u0.subword[0] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u3.d[1]$_DFF_P_  (.D(_00025_),
    .Q(\u0.subword[1] ),
    .CLK(clknet_3_4_0_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u3.d[2]$_DFF_P_  (.D(_00026_),
    .Q(\u0.subword[2] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u3.d[3]$_DFF_P_  (.D(_00027_),
    .Q(\u0.subword[3] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u3.d[4]$_DFF_P_  (.D(_00028_),
    .Q(\u0.subword[4] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u3.d[5]$_DFF_P_  (.D(net3565),
    .Q(\u0.subword[5] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u3.d[6]$_DFF_P_  (.D(_00030_),
    .Q(\u0.subword[6] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.u3.d[7]$_DFF_P_  (.D(_00031_),
    .Q(\u0.subword[7] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][0]$_DFF_P_  (.D(_00289_),
    .Q(\u0.w[0][0] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][10]$_DFF_P_  (.D(_00290_),
    .Q(\u0.w[0][10] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][11]$_DFF_P_  (.D(_00291_),
    .Q(\u0.w[0][11] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][12]$_DFF_P_  (.D(_00292_),
    .Q(\u0.w[0][12] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][13]$_DFF_P_  (.D(_00293_),
    .Q(\u0.w[0][13] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][14]$_DFF_P_  (.D(_00294_),
    .Q(\u0.w[0][14] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][15]$_DFF_P_  (.D(_00295_),
    .Q(\u0.w[0][15] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][16]$_DFF_P_  (.D(_00296_),
    .Q(\u0.w[0][16] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][17]$_DFF_P_  (.D(_00297_),
    .Q(\u0.w[0][17] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][18]$_DFF_P_  (.D(_00298_),
    .Q(\u0.w[0][18] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][19]$_DFF_P_  (.D(_00299_),
    .Q(\u0.w[0][19] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][1]$_DFF_P_  (.D(_00300_),
    .Q(\u0.w[0][1] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][20]$_DFF_P_  (.D(_00301_),
    .Q(\u0.w[0][20] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][21]$_DFF_P_  (.D(_00302_),
    .Q(\u0.w[0][21] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][22]$_DFF_P_  (.D(_00303_),
    .Q(\u0.w[0][22] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][23]$_DFF_P_  (.D(_00304_),
    .Q(\u0.w[0][23] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][24]$_DFF_P_  (.D(_00305_),
    .Q(\u0.w[0][24] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][25]$_DFF_P_  (.D(_00306_),
    .Q(\u0.w[0][25] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][26]$_DFF_P_  (.D(_00307_),
    .Q(\u0.w[0][26] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][27]$_DFF_P_  (.D(_00308_),
    .Q(\u0.w[0][27] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][28]$_DFF_P_  (.D(_00309_),
    .Q(\u0.w[0][28] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][29]$_DFF_P_  (.D(_00310_),
    .Q(\u0.w[0][29] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][2]$_DFF_P_  (.D(_00311_),
    .Q(\u0.w[0][2] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][30]$_DFF_P_  (.D(_00312_),
    .Q(\u0.w[0][30] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][31]$_DFF_P_  (.D(_00313_),
    .Q(\u0.w[0][31] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][3]$_DFF_P_  (.D(_00314_),
    .Q(\u0.w[0][3] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][4]$_DFF_P_  (.D(_00315_),
    .Q(\u0.w[0][4] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][5]$_DFF_P_  (.D(_00316_),
    .Q(\u0.w[0][5] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][6]$_DFF_P_  (.D(_00317_),
    .Q(\u0.w[0][6] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][7]$_DFF_P_  (.D(_00318_),
    .Q(\u0.w[0][7] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][8]$_DFF_P_  (.D(_00319_),
    .Q(\u0.w[0][8] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[0][9]$_DFF_P_  (.D(_00320_),
    .Q(\u0.w[0][9] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][0]$_DFF_P_  (.D(_00321_),
    .Q(\u0.w[1][0] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][10]$_DFF_P_  (.D(_00322_),
    .Q(\u0.w[1][10] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][11]$_DFF_P_  (.D(_00323_),
    .Q(\u0.w[1][11] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][12]$_DFF_P_  (.D(_00324_),
    .Q(\u0.w[1][12] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][13]$_DFF_P_  (.D(_00325_),
    .Q(\u0.w[1][13] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][14]$_DFF_P_  (.D(_00326_),
    .Q(\u0.w[1][14] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][15]$_DFF_P_  (.D(_00327_),
    .Q(\u0.w[1][15] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][16]$_DFF_P_  (.D(_00328_),
    .Q(\u0.w[1][16] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][17]$_DFF_P_  (.D(_00329_),
    .Q(\u0.w[1][17] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][18]$_DFF_P_  (.D(_00330_),
    .Q(\u0.w[1][18] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][19]$_DFF_P_  (.D(_00331_),
    .Q(\u0.w[1][19] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][1]$_DFF_P_  (.D(_00332_),
    .Q(\u0.w[1][1] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][20]$_DFF_P_  (.D(_00333_),
    .Q(\u0.w[1][20] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][21]$_DFF_P_  (.D(_00334_),
    .Q(\u0.w[1][21] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][22]$_DFF_P_  (.D(_00335_),
    .Q(\u0.w[1][22] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][23]$_DFF_P_  (.D(_00336_),
    .Q(\u0.w[1][23] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][24]$_DFF_P_  (.D(_00337_),
    .Q(\u0.w[1][24] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][25]$_DFF_P_  (.D(_00338_),
    .Q(\u0.w[1][25] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][26]$_DFF_P_  (.D(_00339_),
    .Q(\u0.w[1][26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][27]$_DFF_P_  (.D(_00340_),
    .Q(\u0.w[1][27] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][28]$_DFF_P_  (.D(_00341_),
    .Q(\u0.w[1][28] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][29]$_DFF_P_  (.D(_00342_),
    .Q(\u0.w[1][29] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][2]$_DFF_P_  (.D(_00343_),
    .Q(\u0.w[1][2] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][30]$_DFF_P_  (.D(_00344_),
    .Q(\u0.w[1][30] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][31]$_DFF_P_  (.D(_00345_),
    .Q(\u0.w[1][31] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][3]$_DFF_P_  (.D(_00346_),
    .Q(\u0.w[1][3] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][4]$_DFF_P_  (.D(_00347_),
    .Q(\u0.w[1][4] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][5]$_DFF_P_  (.D(_00348_),
    .Q(\u0.w[1][5] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][6]$_DFF_P_  (.D(_00349_),
    .Q(\u0.w[1][6] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][7]$_DFF_P_  (.D(_00350_),
    .Q(\u0.w[1][7] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][8]$_DFF_P_  (.D(_00351_),
    .Q(\u0.w[1][8] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[1][9]$_DFF_P_  (.D(_00352_),
    .Q(\u0.w[1][9] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][0]$_DFF_P_  (.D(_00353_),
    .Q(\u0.w[2][0] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][10]$_DFF_P_  (.D(_00354_),
    .Q(\u0.w[2][10] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][11]$_DFF_P_  (.D(_00355_),
    .Q(\u0.w[2][11] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][12]$_DFF_P_  (.D(_00356_),
    .Q(\u0.w[2][12] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][13]$_DFF_P_  (.D(_00357_),
    .Q(\u0.w[2][13] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][14]$_DFF_P_  (.D(_00358_),
    .Q(\u0.w[2][14] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][15]$_DFF_P_  (.D(_00359_),
    .Q(\u0.w[2][15] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][16]$_DFF_P_  (.D(_00360_),
    .Q(\u0.w[2][16] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][17]$_DFF_P_  (.D(_00361_),
    .Q(\u0.w[2][17] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][18]$_DFF_P_  (.D(_00362_),
    .Q(\u0.w[2][18] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][19]$_DFF_P_  (.D(_00363_),
    .Q(\u0.w[2][19] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][1]$_DFF_P_  (.D(_00364_),
    .Q(\u0.w[2][1] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][20]$_DFF_P_  (.D(_00365_),
    .Q(\u0.w[2][20] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][21]$_DFF_P_  (.D(_00366_),
    .Q(\u0.w[2][21] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][22]$_DFF_P_  (.D(_00367_),
    .Q(\u0.w[2][22] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][23]$_DFF_P_  (.D(_00368_),
    .Q(\u0.w[2][23] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][24]$_DFF_P_  (.D(_00369_),
    .Q(\u0.w[2][24] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][25]$_DFF_P_  (.D(_00370_),
    .Q(\u0.w[2][25] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][26]$_DFF_P_  (.D(_00371_),
    .Q(\u0.w[2][26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][27]$_DFF_P_  (.D(_00372_),
    .Q(\u0.w[2][27] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][28]$_DFF_P_  (.D(_00373_),
    .Q(\u0.w[2][28] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][29]$_DFF_P_  (.D(_00374_),
    .Q(\u0.w[2][29] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][2]$_DFF_P_  (.D(_00375_),
    .Q(\u0.w[2][2] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][30]$_DFF_P_  (.D(_00376_),
    .Q(\u0.w[2][30] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][31]$_DFF_P_  (.D(_00377_),
    .Q(\u0.w[2][31] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][3]$_DFF_P_  (.D(_00378_),
    .Q(\u0.w[2][3] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][4]$_DFF_P_  (.D(_00379_),
    .Q(\u0.w[2][4] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][5]$_DFF_P_  (.D(_00380_),
    .Q(\u0.w[2][5] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][6]$_DFF_P_  (.D(_00381_),
    .Q(\u0.w[2][6] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][7]$_DFF_P_  (.D(_00382_),
    .Q(\u0.w[2][7] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][8]$_DFF_P_  (.D(_00383_),
    .Q(\u0.w[2][8] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[2][9]$_DFF_P_  (.D(_00384_),
    .Q(\u0.w[2][9] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][0]$_DFF_P_  (.D(_03624_),
    .Q(\u0.tmp_w[0] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][10]$_DFF_P_  (.D(_03704_),
    .Q(\u0.tmp_w[10] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][11]$_DFF_P_  (.D(_03715_),
    .Q(\u0.tmp_w[11] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][12]$_DFF_P_  (.D(_03725_),
    .Q(\u0.tmp_w[12] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][13]$_DFF_P_  (.D(_03735_),
    .Q(\u0.tmp_w[13] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][14]$_DFF_P_  (.D(_03744_),
    .Q(\u0.tmp_w[14] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][15]$_DFF_P_  (.D(_03751_),
    .Q(\u0.tmp_w[15] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][16]$_DFF_P_  (.D(net4106),
    .Q(\u0.tmp_w[16] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][17]$_DFF_P_  (.D(net4104),
    .Q(\u0.tmp_w[17] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][18]$_DFF_P_  (.D(_03618_),
    .Q(\u0.tmp_w[18] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][19]$_DFF_P_  (.D(_03579_),
    .Q(\u0.tmp_w[19] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][1]$_DFF_P_  (.D(net4094),
    .Q(\u0.tmp_w[1] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][20]$_DFF_P_  (.D(_03611_),
    .Q(\u0.tmp_w[20] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][21]$_DFF_P_  (.D(_03602_),
    .Q(\u0.tmp_w[21] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][22]$_DFF_P_  (.D(_03759_),
    .Q(\u0.tmp_w[22] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][23]$_DFF_P_  (.D(_03767_),
    .Q(\u0.tmp_w[23] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][24]$_DFF_P_  (.D(_03772_),
    .Q(\u0.tmp_w[24] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][25]$_DFF_P_  (.D(net4082),
    .Q(\u0.tmp_w[25] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_2 \u0.w[3][26]$_DFF_P_  (.D(net4079),
    .Q(\u0.tmp_w[26] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][27]$_DFF_P_  (.D(_03792_),
    .Q(\u0.tmp_w[27] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][28]$_DFF_P_  (.D(_03801_),
    .Q(\u0.tmp_w[28] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][29]$_DFF_P_  (.D(_03810_),
    .Q(\u0.tmp_w[29] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][2]$_DFF_P_  (.D(_03639_),
    .Q(\u0.tmp_w[2] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][30]$_DFF_P_  (.D(_00398_),
    .Q(\u0.tmp_w[30] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][31]$_DFF_P_  (.D(_03824_),
    .Q(\u0.tmp_w[31] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][3]$_DFF_P_  (.D(_03648_),
    .Q(\u0.tmp_w[3] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][4]$_DFF_P_  (.D(_03658_),
    .Q(\u0.tmp_w[4] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][5]$_DFF_P_  (.D(_03667_),
    .Q(\u0.tmp_w[5] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][6]$_DFF_P_  (.D(_03676_),
    .Q(\u0.tmp_w[6] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][7]$_DFF_P_  (.D(_03685_),
    .Q(\u0.tmp_w[7] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][8]$_DFF_P_  (.D(net4090),
    .Q(\u0.tmp_w[8] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__dfxtp_1 \u0.w[3][9]$_DFF_P_  (.D(_11860_[0]),
    .Q(\u0.tmp_w[9] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5709 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(key[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(key[100]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(key[101]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(key[102]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(key[103]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(key[104]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(key[105]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(key[106]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(key[107]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(key[108]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(key[109]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(key[10]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(key[110]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(key[111]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(key[112]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(key[113]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(key[114]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(key[115]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(key[116]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(key[117]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(key[118]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(key[119]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(key[11]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(key[120]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(key[121]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(key[122]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(key[123]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(key[124]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(key[125]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(key[126]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(key[127]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(key[12]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(key[13]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(key[14]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(key[15]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(key[16]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(key[17]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(key[18]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(key[19]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input40 (.A(key[1]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(key[20]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(key[21]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(key[22]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(key[23]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(key[24]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(key[25]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(key[26]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(key[27]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(key[28]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input50 (.A(key[29]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(key[2]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(key[30]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(key[31]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(key[32]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(key[33]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(key[34]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(key[35]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(key[36]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(key[37]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input60 (.A(key[38]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(key[39]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(key[3]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(key[40]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(key[41]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input65 (.A(key[42]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(key[43]),
    .X(net66));
 sky130_fd_sc_hd__buf_1 input67 (.A(key[44]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input68 (.A(key[45]),
    .X(net68));
 sky130_fd_sc_hd__buf_1 input69 (.A(key[46]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input70 (.A(key[47]),
    .X(net70));
 sky130_fd_sc_hd__buf_1 input71 (.A(key[48]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 input72 (.A(key[49]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input73 (.A(key[4]),
    .X(net73));
 sky130_fd_sc_hd__buf_1 input74 (.A(key[50]),
    .X(net74));
 sky130_fd_sc_hd__buf_1 input75 (.A(key[51]),
    .X(net75));
 sky130_fd_sc_hd__buf_1 input76 (.A(key[52]),
    .X(net76));
 sky130_fd_sc_hd__buf_1 input77 (.A(key[53]),
    .X(net77));
 sky130_fd_sc_hd__buf_1 input78 (.A(key[54]),
    .X(net78));
 sky130_fd_sc_hd__buf_1 input79 (.A(key[55]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input80 (.A(key[56]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 input81 (.A(key[57]),
    .X(net81));
 sky130_fd_sc_hd__buf_1 input82 (.A(key[58]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input83 (.A(key[59]),
    .X(net83));
 sky130_fd_sc_hd__buf_1 input84 (.A(key[5]),
    .X(net84));
 sky130_fd_sc_hd__buf_1 input85 (.A(key[60]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 input86 (.A(key[61]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 input87 (.A(key[62]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 input88 (.A(key[63]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 input89 (.A(key[64]),
    .X(net89));
 sky130_fd_sc_hd__buf_1 input90 (.A(key[65]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 input91 (.A(key[66]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 input92 (.A(key[67]),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input93 (.A(key[68]),
    .X(net93));
 sky130_fd_sc_hd__buf_1 input94 (.A(key[69]),
    .X(net94));
 sky130_fd_sc_hd__buf_1 input95 (.A(key[6]),
    .X(net95));
 sky130_fd_sc_hd__buf_1 input96 (.A(key[70]),
    .X(net96));
 sky130_fd_sc_hd__buf_1 input97 (.A(key[71]),
    .X(net97));
 sky130_fd_sc_hd__buf_1 input98 (.A(key[72]),
    .X(net98));
 sky130_fd_sc_hd__buf_1 input99 (.A(key[73]),
    .X(net99));
 sky130_fd_sc_hd__buf_1 input100 (.A(key[74]),
    .X(net100));
 sky130_fd_sc_hd__buf_1 input101 (.A(key[75]),
    .X(net101));
 sky130_fd_sc_hd__buf_1 input102 (.A(key[76]),
    .X(net102));
 sky130_fd_sc_hd__buf_1 input103 (.A(key[77]),
    .X(net103));
 sky130_fd_sc_hd__buf_1 input104 (.A(key[78]),
    .X(net104));
 sky130_fd_sc_hd__buf_1 input105 (.A(key[79]),
    .X(net105));
 sky130_fd_sc_hd__buf_1 input106 (.A(key[7]),
    .X(net106));
 sky130_fd_sc_hd__buf_1 input107 (.A(key[80]),
    .X(net107));
 sky130_fd_sc_hd__buf_1 input108 (.A(key[81]),
    .X(net108));
 sky130_fd_sc_hd__buf_1 input109 (.A(key[82]),
    .X(net109));
 sky130_fd_sc_hd__buf_1 input110 (.A(key[83]),
    .X(net110));
 sky130_fd_sc_hd__buf_1 input111 (.A(key[84]),
    .X(net111));
 sky130_fd_sc_hd__buf_1 input112 (.A(key[85]),
    .X(net112));
 sky130_fd_sc_hd__buf_1 input113 (.A(key[86]),
    .X(net113));
 sky130_fd_sc_hd__buf_1 input114 (.A(key[87]),
    .X(net114));
 sky130_fd_sc_hd__buf_1 input115 (.A(key[88]),
    .X(net115));
 sky130_fd_sc_hd__buf_1 input116 (.A(key[89]),
    .X(net116));
 sky130_fd_sc_hd__buf_1 input117 (.A(key[8]),
    .X(net117));
 sky130_fd_sc_hd__buf_1 input118 (.A(key[90]),
    .X(net118));
 sky130_fd_sc_hd__buf_1 input119 (.A(key[91]),
    .X(net119));
 sky130_fd_sc_hd__buf_1 input120 (.A(key[92]),
    .X(net120));
 sky130_fd_sc_hd__buf_1 input121 (.A(key[93]),
    .X(net121));
 sky130_fd_sc_hd__buf_1 input122 (.A(key[94]),
    .X(net122));
 sky130_fd_sc_hd__buf_1 input123 (.A(key[95]),
    .X(net123));
 sky130_fd_sc_hd__buf_1 input124 (.A(key[96]),
    .X(net124));
 sky130_fd_sc_hd__buf_1 input125 (.A(key[97]),
    .X(net125));
 sky130_fd_sc_hd__buf_1 input126 (.A(key[98]),
    .X(net126));
 sky130_fd_sc_hd__buf_1 input127 (.A(key[99]),
    .X(net127));
 sky130_fd_sc_hd__buf_1 input128 (.A(key[9]),
    .X(net128));
 sky130_fd_sc_hd__buf_12 input129 (.A(ld),
    .X(net129));
 sky130_fd_sc_hd__buf_1 input130 (.A(rst),
    .X(net130));
 sky130_fd_sc_hd__buf_1 input131 (.A(text_in[0]),
    .X(net131));
 sky130_fd_sc_hd__buf_1 input132 (.A(text_in[100]),
    .X(net132));
 sky130_fd_sc_hd__buf_1 input133 (.A(text_in[101]),
    .X(net133));
 sky130_fd_sc_hd__buf_1 input134 (.A(text_in[102]),
    .X(net134));
 sky130_fd_sc_hd__buf_1 input135 (.A(text_in[103]),
    .X(net135));
 sky130_fd_sc_hd__buf_1 input136 (.A(text_in[104]),
    .X(net136));
 sky130_fd_sc_hd__buf_1 input137 (.A(text_in[105]),
    .X(net137));
 sky130_fd_sc_hd__buf_1 input138 (.A(text_in[106]),
    .X(net138));
 sky130_fd_sc_hd__buf_1 input139 (.A(text_in[107]),
    .X(net139));
 sky130_fd_sc_hd__buf_1 input140 (.A(text_in[108]),
    .X(net140));
 sky130_fd_sc_hd__buf_1 input141 (.A(text_in[109]),
    .X(net141));
 sky130_fd_sc_hd__buf_1 input142 (.A(text_in[10]),
    .X(net142));
 sky130_fd_sc_hd__buf_1 input143 (.A(text_in[110]),
    .X(net143));
 sky130_fd_sc_hd__buf_1 input144 (.A(text_in[111]),
    .X(net144));
 sky130_fd_sc_hd__buf_1 input145 (.A(text_in[112]),
    .X(net145));
 sky130_fd_sc_hd__buf_1 input146 (.A(text_in[113]),
    .X(net146));
 sky130_fd_sc_hd__buf_1 input147 (.A(text_in[114]),
    .X(net147));
 sky130_fd_sc_hd__buf_1 input148 (.A(text_in[115]),
    .X(net148));
 sky130_fd_sc_hd__buf_1 input149 (.A(text_in[116]),
    .X(net149));
 sky130_fd_sc_hd__buf_1 input150 (.A(text_in[117]),
    .X(net150));
 sky130_fd_sc_hd__buf_1 input151 (.A(text_in[118]),
    .X(net151));
 sky130_fd_sc_hd__buf_1 input152 (.A(text_in[119]),
    .X(net152));
 sky130_fd_sc_hd__buf_1 input153 (.A(text_in[11]),
    .X(net153));
 sky130_fd_sc_hd__buf_1 input154 (.A(text_in[120]),
    .X(net154));
 sky130_fd_sc_hd__buf_1 input155 (.A(text_in[121]),
    .X(net155));
 sky130_fd_sc_hd__buf_1 input156 (.A(text_in[122]),
    .X(net156));
 sky130_fd_sc_hd__buf_1 input157 (.A(text_in[123]),
    .X(net157));
 sky130_fd_sc_hd__buf_1 input158 (.A(text_in[124]),
    .X(net158));
 sky130_fd_sc_hd__buf_1 input159 (.A(text_in[125]),
    .X(net159));
 sky130_fd_sc_hd__buf_1 input160 (.A(text_in[126]),
    .X(net160));
 sky130_fd_sc_hd__buf_1 input161 (.A(text_in[127]),
    .X(net161));
 sky130_fd_sc_hd__buf_1 input162 (.A(text_in[12]),
    .X(net162));
 sky130_fd_sc_hd__buf_1 input163 (.A(text_in[13]),
    .X(net163));
 sky130_fd_sc_hd__buf_1 input164 (.A(text_in[14]),
    .X(net164));
 sky130_fd_sc_hd__buf_1 input165 (.A(text_in[15]),
    .X(net165));
 sky130_fd_sc_hd__buf_1 input166 (.A(text_in[16]),
    .X(net166));
 sky130_fd_sc_hd__buf_1 input167 (.A(text_in[17]),
    .X(net167));
 sky130_fd_sc_hd__buf_1 input168 (.A(text_in[18]),
    .X(net168));
 sky130_fd_sc_hd__buf_1 input169 (.A(text_in[19]),
    .X(net169));
 sky130_fd_sc_hd__buf_1 input170 (.A(text_in[1]),
    .X(net170));
 sky130_fd_sc_hd__buf_1 input171 (.A(text_in[20]),
    .X(net171));
 sky130_fd_sc_hd__buf_1 input172 (.A(text_in[21]),
    .X(net172));
 sky130_fd_sc_hd__buf_1 input173 (.A(text_in[22]),
    .X(net173));
 sky130_fd_sc_hd__buf_1 input174 (.A(text_in[23]),
    .X(net174));
 sky130_fd_sc_hd__buf_1 input175 (.A(text_in[24]),
    .X(net175));
 sky130_fd_sc_hd__buf_1 input176 (.A(text_in[25]),
    .X(net176));
 sky130_fd_sc_hd__buf_1 input177 (.A(text_in[26]),
    .X(net177));
 sky130_fd_sc_hd__buf_1 input178 (.A(text_in[27]),
    .X(net178));
 sky130_fd_sc_hd__buf_1 input179 (.A(text_in[28]),
    .X(net179));
 sky130_fd_sc_hd__buf_1 input180 (.A(text_in[29]),
    .X(net180));
 sky130_fd_sc_hd__buf_1 input181 (.A(text_in[2]),
    .X(net181));
 sky130_fd_sc_hd__buf_1 input182 (.A(text_in[30]),
    .X(net182));
 sky130_fd_sc_hd__buf_1 input183 (.A(text_in[31]),
    .X(net183));
 sky130_fd_sc_hd__buf_1 input184 (.A(text_in[32]),
    .X(net184));
 sky130_fd_sc_hd__buf_1 input185 (.A(text_in[33]),
    .X(net185));
 sky130_fd_sc_hd__buf_1 input186 (.A(text_in[34]),
    .X(net186));
 sky130_fd_sc_hd__buf_1 input187 (.A(text_in[35]),
    .X(net187));
 sky130_fd_sc_hd__buf_1 input188 (.A(text_in[36]),
    .X(net188));
 sky130_fd_sc_hd__buf_1 input189 (.A(text_in[37]),
    .X(net189));
 sky130_fd_sc_hd__buf_1 input190 (.A(text_in[38]),
    .X(net190));
 sky130_fd_sc_hd__buf_1 input191 (.A(text_in[39]),
    .X(net191));
 sky130_fd_sc_hd__buf_1 input192 (.A(text_in[3]),
    .X(net192));
 sky130_fd_sc_hd__buf_1 input193 (.A(text_in[40]),
    .X(net193));
 sky130_fd_sc_hd__buf_1 input194 (.A(text_in[41]),
    .X(net194));
 sky130_fd_sc_hd__buf_1 input195 (.A(text_in[42]),
    .X(net195));
 sky130_fd_sc_hd__buf_1 input196 (.A(text_in[43]),
    .X(net196));
 sky130_fd_sc_hd__buf_1 input197 (.A(text_in[44]),
    .X(net197));
 sky130_fd_sc_hd__buf_1 input198 (.A(text_in[45]),
    .X(net198));
 sky130_fd_sc_hd__buf_1 input199 (.A(text_in[46]),
    .X(net199));
 sky130_fd_sc_hd__buf_1 input200 (.A(text_in[47]),
    .X(net200));
 sky130_fd_sc_hd__buf_1 input201 (.A(text_in[48]),
    .X(net201));
 sky130_fd_sc_hd__buf_1 input202 (.A(text_in[49]),
    .X(net202));
 sky130_fd_sc_hd__buf_1 input203 (.A(text_in[4]),
    .X(net203));
 sky130_fd_sc_hd__buf_1 input204 (.A(text_in[50]),
    .X(net204));
 sky130_fd_sc_hd__buf_1 input205 (.A(text_in[51]),
    .X(net205));
 sky130_fd_sc_hd__buf_1 input206 (.A(text_in[52]),
    .X(net206));
 sky130_fd_sc_hd__buf_1 input207 (.A(text_in[53]),
    .X(net207));
 sky130_fd_sc_hd__buf_1 input208 (.A(text_in[54]),
    .X(net208));
 sky130_fd_sc_hd__buf_1 input209 (.A(text_in[55]),
    .X(net209));
 sky130_fd_sc_hd__buf_1 input210 (.A(text_in[56]),
    .X(net210));
 sky130_fd_sc_hd__buf_1 input211 (.A(text_in[57]),
    .X(net211));
 sky130_fd_sc_hd__buf_1 input212 (.A(text_in[58]),
    .X(net212));
 sky130_fd_sc_hd__buf_1 input213 (.A(text_in[59]),
    .X(net213));
 sky130_fd_sc_hd__buf_1 input214 (.A(text_in[5]),
    .X(net214));
 sky130_fd_sc_hd__buf_1 input215 (.A(text_in[60]),
    .X(net215));
 sky130_fd_sc_hd__buf_1 input216 (.A(text_in[61]),
    .X(net216));
 sky130_fd_sc_hd__buf_1 input217 (.A(text_in[62]),
    .X(net217));
 sky130_fd_sc_hd__buf_1 input218 (.A(text_in[63]),
    .X(net218));
 sky130_fd_sc_hd__buf_1 input219 (.A(text_in[64]),
    .X(net219));
 sky130_fd_sc_hd__buf_1 input220 (.A(text_in[65]),
    .X(net220));
 sky130_fd_sc_hd__buf_1 input221 (.A(text_in[66]),
    .X(net221));
 sky130_fd_sc_hd__buf_1 input222 (.A(text_in[67]),
    .X(net222));
 sky130_fd_sc_hd__buf_1 input223 (.A(text_in[68]),
    .X(net223));
 sky130_fd_sc_hd__buf_1 input224 (.A(text_in[69]),
    .X(net224));
 sky130_fd_sc_hd__buf_1 input225 (.A(text_in[6]),
    .X(net225));
 sky130_fd_sc_hd__buf_1 input226 (.A(text_in[70]),
    .X(net226));
 sky130_fd_sc_hd__buf_1 input227 (.A(text_in[71]),
    .X(net227));
 sky130_fd_sc_hd__buf_1 input228 (.A(text_in[72]),
    .X(net228));
 sky130_fd_sc_hd__buf_1 input229 (.A(text_in[73]),
    .X(net229));
 sky130_fd_sc_hd__buf_1 input230 (.A(text_in[74]),
    .X(net230));
 sky130_fd_sc_hd__buf_1 input231 (.A(text_in[75]),
    .X(net231));
 sky130_fd_sc_hd__buf_1 input232 (.A(text_in[76]),
    .X(net232));
 sky130_fd_sc_hd__buf_1 input233 (.A(text_in[77]),
    .X(net233));
 sky130_fd_sc_hd__buf_1 input234 (.A(text_in[78]),
    .X(net234));
 sky130_fd_sc_hd__buf_1 input235 (.A(text_in[79]),
    .X(net235));
 sky130_fd_sc_hd__buf_1 input236 (.A(text_in[7]),
    .X(net236));
 sky130_fd_sc_hd__buf_1 input237 (.A(text_in[80]),
    .X(net237));
 sky130_fd_sc_hd__buf_1 input238 (.A(text_in[81]),
    .X(net238));
 sky130_fd_sc_hd__buf_1 input239 (.A(text_in[82]),
    .X(net239));
 sky130_fd_sc_hd__buf_1 input240 (.A(text_in[83]),
    .X(net240));
 sky130_fd_sc_hd__buf_1 input241 (.A(text_in[84]),
    .X(net241));
 sky130_fd_sc_hd__buf_1 input242 (.A(text_in[85]),
    .X(net242));
 sky130_fd_sc_hd__buf_1 input243 (.A(text_in[86]),
    .X(net243));
 sky130_fd_sc_hd__buf_1 input244 (.A(text_in[87]),
    .X(net244));
 sky130_fd_sc_hd__buf_1 input245 (.A(text_in[88]),
    .X(net245));
 sky130_fd_sc_hd__buf_1 input246 (.A(text_in[89]),
    .X(net246));
 sky130_fd_sc_hd__buf_1 input247 (.A(text_in[8]),
    .X(net247));
 sky130_fd_sc_hd__buf_1 input248 (.A(text_in[90]),
    .X(net248));
 sky130_fd_sc_hd__buf_1 input249 (.A(text_in[91]),
    .X(net249));
 sky130_fd_sc_hd__buf_1 input250 (.A(text_in[92]),
    .X(net250));
 sky130_fd_sc_hd__buf_1 input251 (.A(text_in[93]),
    .X(net251));
 sky130_fd_sc_hd__buf_1 input252 (.A(text_in[94]),
    .X(net252));
 sky130_fd_sc_hd__buf_1 input253 (.A(text_in[95]),
    .X(net253));
 sky130_fd_sc_hd__buf_1 input254 (.A(text_in[96]),
    .X(net254));
 sky130_fd_sc_hd__buf_1 input255 (.A(text_in[97]),
    .X(net255));
 sky130_fd_sc_hd__buf_1 input256 (.A(text_in[98]),
    .X(net256));
 sky130_fd_sc_hd__buf_1 input257 (.A(text_in[99]),
    .X(net257));
 sky130_fd_sc_hd__buf_1 input258 (.A(text_in[9]),
    .X(net258));
 sky130_fd_sc_hd__buf_1 output259 (.A(net259),
    .X(done));
 sky130_fd_sc_hd__buf_1 output260 (.A(net260),
    .X(text_out[0]));
 sky130_fd_sc_hd__buf_1 output261 (.A(net261),
    .X(text_out[100]));
 sky130_fd_sc_hd__buf_1 output262 (.A(net262),
    .X(text_out[101]));
 sky130_fd_sc_hd__buf_1 output263 (.A(net263),
    .X(text_out[102]));
 sky130_fd_sc_hd__clkbuf_2 output264 (.A(net264),
    .X(text_out[103]));
 sky130_fd_sc_hd__buf_1 output265 (.A(net265),
    .X(text_out[104]));
 sky130_fd_sc_hd__buf_1 output266 (.A(net266),
    .X(text_out[105]));
 sky130_fd_sc_hd__buf_1 output267 (.A(net267),
    .X(text_out[106]));
 sky130_fd_sc_hd__buf_1 output268 (.A(net268),
    .X(text_out[107]));
 sky130_fd_sc_hd__buf_1 output269 (.A(net269),
    .X(text_out[108]));
 sky130_fd_sc_hd__buf_1 output270 (.A(net270),
    .X(text_out[109]));
 sky130_fd_sc_hd__buf_1 output271 (.A(net271),
    .X(text_out[10]));
 sky130_fd_sc_hd__buf_1 output272 (.A(net272),
    .X(text_out[110]));
 sky130_fd_sc_hd__buf_1 output273 (.A(net273),
    .X(text_out[111]));
 sky130_fd_sc_hd__buf_1 output274 (.A(net274),
    .X(text_out[112]));
 sky130_fd_sc_hd__buf_1 output275 (.A(net275),
    .X(text_out[113]));
 sky130_fd_sc_hd__buf_1 output276 (.A(net276),
    .X(text_out[114]));
 sky130_fd_sc_hd__buf_1 output277 (.A(net277),
    .X(text_out[115]));
 sky130_fd_sc_hd__buf_1 output278 (.A(net278),
    .X(text_out[116]));
 sky130_fd_sc_hd__buf_1 output279 (.A(net279),
    .X(text_out[117]));
 sky130_fd_sc_hd__buf_1 output280 (.A(net280),
    .X(text_out[118]));
 sky130_fd_sc_hd__buf_1 output281 (.A(net281),
    .X(text_out[119]));
 sky130_fd_sc_hd__buf_1 output282 (.A(net282),
    .X(text_out[11]));
 sky130_fd_sc_hd__buf_1 output283 (.A(net283),
    .X(text_out[120]));
 sky130_fd_sc_hd__buf_1 output284 (.A(net284),
    .X(text_out[121]));
 sky130_fd_sc_hd__buf_1 output285 (.A(net285),
    .X(text_out[122]));
 sky130_fd_sc_hd__buf_1 output286 (.A(net286),
    .X(text_out[123]));
 sky130_fd_sc_hd__buf_1 output287 (.A(net287),
    .X(text_out[124]));
 sky130_fd_sc_hd__buf_1 output288 (.A(net288),
    .X(text_out[125]));
 sky130_fd_sc_hd__buf_1 output289 (.A(net289),
    .X(text_out[126]));
 sky130_fd_sc_hd__buf_1 output290 (.A(net290),
    .X(text_out[127]));
 sky130_fd_sc_hd__buf_1 output291 (.A(net291),
    .X(text_out[12]));
 sky130_fd_sc_hd__buf_1 output292 (.A(net292),
    .X(text_out[13]));
 sky130_fd_sc_hd__buf_1 output293 (.A(net293),
    .X(text_out[14]));
 sky130_fd_sc_hd__buf_1 output294 (.A(net294),
    .X(text_out[15]));
 sky130_fd_sc_hd__buf_1 output295 (.A(net295),
    .X(text_out[16]));
 sky130_fd_sc_hd__buf_1 output296 (.A(net296),
    .X(text_out[17]));
 sky130_fd_sc_hd__buf_1 output297 (.A(net297),
    .X(text_out[18]));
 sky130_fd_sc_hd__buf_1 output298 (.A(net298),
    .X(text_out[19]));
 sky130_fd_sc_hd__buf_1 output299 (.A(net299),
    .X(text_out[1]));
 sky130_fd_sc_hd__buf_1 output300 (.A(net300),
    .X(text_out[20]));
 sky130_fd_sc_hd__buf_1 output301 (.A(net301),
    .X(text_out[21]));
 sky130_fd_sc_hd__buf_1 output302 (.A(net302),
    .X(text_out[22]));
 sky130_fd_sc_hd__buf_1 output303 (.A(net303),
    .X(text_out[23]));
 sky130_fd_sc_hd__buf_1 output304 (.A(net304),
    .X(text_out[24]));
 sky130_fd_sc_hd__buf_1 output305 (.A(net305),
    .X(text_out[25]));
 sky130_fd_sc_hd__buf_1 output306 (.A(net306),
    .X(text_out[26]));
 sky130_fd_sc_hd__buf_1 output307 (.A(net307),
    .X(text_out[27]));
 sky130_fd_sc_hd__buf_1 output308 (.A(net308),
    .X(text_out[28]));
 sky130_fd_sc_hd__buf_1 output309 (.A(net309),
    .X(text_out[29]));
 sky130_fd_sc_hd__buf_1 output310 (.A(net310),
    .X(text_out[2]));
 sky130_fd_sc_hd__buf_1 output311 (.A(net311),
    .X(text_out[30]));
 sky130_fd_sc_hd__buf_1 output312 (.A(net312),
    .X(text_out[31]));
 sky130_fd_sc_hd__buf_1 output313 (.A(net313),
    .X(text_out[32]));
 sky130_fd_sc_hd__buf_1 output314 (.A(net314),
    .X(text_out[33]));
 sky130_fd_sc_hd__buf_1 output315 (.A(net315),
    .X(text_out[34]));
 sky130_fd_sc_hd__buf_1 output316 (.A(net316),
    .X(text_out[35]));
 sky130_fd_sc_hd__buf_1 output317 (.A(net317),
    .X(text_out[36]));
 sky130_fd_sc_hd__buf_1 output318 (.A(net318),
    .X(text_out[37]));
 sky130_fd_sc_hd__buf_1 output319 (.A(net319),
    .X(text_out[38]));
 sky130_fd_sc_hd__buf_1 output320 (.A(net320),
    .X(text_out[39]));
 sky130_fd_sc_hd__buf_1 output321 (.A(net321),
    .X(text_out[3]));
 sky130_fd_sc_hd__buf_1 output322 (.A(net322),
    .X(text_out[40]));
 sky130_fd_sc_hd__buf_1 output323 (.A(net323),
    .X(text_out[41]));
 sky130_fd_sc_hd__buf_1 output324 (.A(net324),
    .X(text_out[42]));
 sky130_fd_sc_hd__buf_1 output325 (.A(net325),
    .X(text_out[43]));
 sky130_fd_sc_hd__buf_1 output326 (.A(net326),
    .X(text_out[44]));
 sky130_fd_sc_hd__buf_1 output327 (.A(net327),
    .X(text_out[45]));
 sky130_fd_sc_hd__buf_1 output328 (.A(net328),
    .X(text_out[46]));
 sky130_fd_sc_hd__buf_1 output329 (.A(net329),
    .X(text_out[47]));
 sky130_fd_sc_hd__buf_1 output330 (.A(net330),
    .X(text_out[48]));
 sky130_fd_sc_hd__buf_1 output331 (.A(net331),
    .X(text_out[49]));
 sky130_fd_sc_hd__buf_1 output332 (.A(net332),
    .X(text_out[4]));
 sky130_fd_sc_hd__buf_1 output333 (.A(net333),
    .X(text_out[50]));
 sky130_fd_sc_hd__buf_1 output334 (.A(net334),
    .X(text_out[51]));
 sky130_fd_sc_hd__buf_1 output335 (.A(net335),
    .X(text_out[52]));
 sky130_fd_sc_hd__buf_1 output336 (.A(net336),
    .X(text_out[53]));
 sky130_fd_sc_hd__buf_1 output337 (.A(net337),
    .X(text_out[54]));
 sky130_fd_sc_hd__buf_1 output338 (.A(net338),
    .X(text_out[55]));
 sky130_fd_sc_hd__buf_1 output339 (.A(net339),
    .X(text_out[56]));
 sky130_fd_sc_hd__buf_1 output340 (.A(net340),
    .X(text_out[57]));
 sky130_fd_sc_hd__buf_1 output341 (.A(net341),
    .X(text_out[58]));
 sky130_fd_sc_hd__buf_1 output342 (.A(net342),
    .X(text_out[59]));
 sky130_fd_sc_hd__buf_1 output343 (.A(net343),
    .X(text_out[5]));
 sky130_fd_sc_hd__buf_1 output344 (.A(net344),
    .X(text_out[60]));
 sky130_fd_sc_hd__buf_1 output345 (.A(net345),
    .X(text_out[61]));
 sky130_fd_sc_hd__buf_1 output346 (.A(net346),
    .X(text_out[62]));
 sky130_fd_sc_hd__buf_1 output347 (.A(net347),
    .X(text_out[63]));
 sky130_fd_sc_hd__buf_1 output348 (.A(net348),
    .X(text_out[64]));
 sky130_fd_sc_hd__buf_1 output349 (.A(net349),
    .X(text_out[65]));
 sky130_fd_sc_hd__buf_1 output350 (.A(net350),
    .X(text_out[66]));
 sky130_fd_sc_hd__buf_1 output351 (.A(net351),
    .X(text_out[67]));
 sky130_fd_sc_hd__buf_1 output352 (.A(net352),
    .X(text_out[68]));
 sky130_fd_sc_hd__buf_1 output353 (.A(net353),
    .X(text_out[69]));
 sky130_fd_sc_hd__buf_1 output354 (.A(net354),
    .X(text_out[6]));
 sky130_fd_sc_hd__buf_1 output355 (.A(net355),
    .X(text_out[70]));
 sky130_fd_sc_hd__buf_1 output356 (.A(net356),
    .X(text_out[71]));
 sky130_fd_sc_hd__buf_1 output357 (.A(net357),
    .X(text_out[72]));
 sky130_fd_sc_hd__buf_1 output358 (.A(net358),
    .X(text_out[73]));
 sky130_fd_sc_hd__buf_1 output359 (.A(net359),
    .X(text_out[74]));
 sky130_fd_sc_hd__buf_1 output360 (.A(net360),
    .X(text_out[75]));
 sky130_fd_sc_hd__buf_1 output361 (.A(net361),
    .X(text_out[76]));
 sky130_fd_sc_hd__buf_1 output362 (.A(net362),
    .X(text_out[77]));
 sky130_fd_sc_hd__buf_1 output363 (.A(net363),
    .X(text_out[78]));
 sky130_fd_sc_hd__buf_1 output364 (.A(net364),
    .X(text_out[79]));
 sky130_fd_sc_hd__buf_1 output365 (.A(net365),
    .X(text_out[7]));
 sky130_fd_sc_hd__buf_1 output366 (.A(net366),
    .X(text_out[80]));
 sky130_fd_sc_hd__buf_1 output367 (.A(net367),
    .X(text_out[81]));
 sky130_fd_sc_hd__buf_1 output368 (.A(net368),
    .X(text_out[82]));
 sky130_fd_sc_hd__buf_1 output369 (.A(net369),
    .X(text_out[83]));
 sky130_fd_sc_hd__buf_1 output370 (.A(net370),
    .X(text_out[84]));
 sky130_fd_sc_hd__buf_1 output371 (.A(net371),
    .X(text_out[85]));
 sky130_fd_sc_hd__buf_1 output372 (.A(net372),
    .X(text_out[86]));
 sky130_fd_sc_hd__buf_1 output373 (.A(net373),
    .X(text_out[87]));
 sky130_fd_sc_hd__buf_1 output374 (.A(net374),
    .X(text_out[88]));
 sky130_fd_sc_hd__buf_1 output375 (.A(net375),
    .X(text_out[89]));
 sky130_fd_sc_hd__buf_1 output376 (.A(net376),
    .X(text_out[8]));
 sky130_fd_sc_hd__buf_1 output377 (.A(net377),
    .X(text_out[90]));
 sky130_fd_sc_hd__buf_1 output378 (.A(net378),
    .X(text_out[91]));
 sky130_fd_sc_hd__buf_1 output379 (.A(net379),
    .X(text_out[92]));
 sky130_fd_sc_hd__buf_1 output380 (.A(net380),
    .X(text_out[93]));
 sky130_fd_sc_hd__buf_1 output381 (.A(net381),
    .X(text_out[94]));
 sky130_fd_sc_hd__buf_1 output382 (.A(net382),
    .X(text_out[95]));
 sky130_fd_sc_hd__buf_1 output383 (.A(net383),
    .X(text_out[96]));
 sky130_fd_sc_hd__buf_1 output384 (.A(net384),
    .X(text_out[97]));
 sky130_fd_sc_hd__buf_1 output385 (.A(net385),
    .X(text_out[98]));
 sky130_fd_sc_hd__buf_1 output386 (.A(net386),
    .X(text_out[99]));
 sky130_fd_sc_hd__buf_1 output387 (.A(net387),
    .X(text_out[9]));
 sky130_fd_sc_hd__buf_12 place3738 (.A(_02480_),
    .X(net3738));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__buf_1 place3793 (.A(net3792),
    .X(net3793));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__buf_12 place3813 (.A(_00830_),
    .X(net3813));
 sky130_fd_sc_hd__buf_8 place3857 (.A(_11122_),
    .X(net3857));
 sky130_fd_sc_hd__buf_1 place3923 (.A(_09406_),
    .X(net3923));
 sky130_fd_sc_hd__buf_8 place3892 (.A(_09998_),
    .X(net3892));
 sky130_fd_sc_hd__buf_1 place3915 (.A(_09412_),
    .X(net3915));
 sky130_fd_sc_hd__buf_1 place4030 (.A(net4029),
    .X(net4030));
 sky130_fd_sc_hd__buf_12 place3961 (.A(_08293_),
    .X(net3961));
 sky130_fd_sc_hd__buf_1 place3975 (.A(net3974),
    .X(net3975));
 sky130_fd_sc_hd__buf_8 place3990 (.A(net3987),
    .X(net3990));
 sky130_fd_sc_hd__buf_12 place4023 (.A(_06541_),
    .X(net4023));
 sky130_fd_sc_hd__buf_12 place4004 (.A(_07174_),
    .X(net4004));
 sky130_fd_sc_hd__buf_12 place4016 (.A(_06590_),
    .X(net4016));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(text_in[0]));
 sky130_fd_sc_hd__buf_1 place3576 (.A(_02542_),
    .X(net3576));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(text_in[114]));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(text_in[114]));
 sky130_fd_sc_hd__buf_12 place4101 (.A(_03617_),
    .X(net4101));
 sky130_fd_sc_hd__buf_1 place3574 (.A(_06081_),
    .X(net3574));
 sky130_fd_sc_hd__buf_12 place4108 (.A(_03578_),
    .X(net4108));
 sky130_fd_sc_hd__buf_1 place4132 (.A(\u0.tmp_w[22] ),
    .X(net4132));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__buf_1 place4125 (.A(_03574_),
    .X(net4125));
 sky130_fd_sc_hd__buf_1 place4114 (.A(_05879_),
    .X(net4114));
 sky130_fd_sc_hd__buf_1 place4136 (.A(\u0.w[2][8] ),
    .X(net4136));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__buf_1 place4137 (.A(\u0.w[2][25] ),
    .X(net4137));
 sky130_fd_sc_hd__buf_1 place4138 (.A(\u0.w[2][20] ),
    .X(net4138));
 sky130_fd_sc_hd__buf_8 place3818 (.A(net3813),
    .X(net3818));
 sky130_fd_sc_hd__buf_1 place3570 (.A(_00563_),
    .X(net3570));
 sky130_fd_sc_hd__buf_1 place3563 (.A(_00081_),
    .X(net3563));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(text_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(text_in[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(text_in[126]));
 sky130_fd_sc_hd__buf_1 place3564 (.A(_00051_),
    .X(net3564));
 sky130_fd_sc_hd__buf_8 place3566 (.A(_00021_),
    .X(net3566));
 sky130_fd_sc_hd__buf_1 place3571 (.A(_08952_),
    .X(net3571));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(text_in[116]));
 sky130_fd_sc_hd__buf_1 place3568 (.A(_01224_),
    .X(net3568));
 sky130_fd_sc_hd__buf_12 place3704 (.A(net3703),
    .X(net3704));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(text_in[102]));
 sky130_fd_sc_hd__buf_8 place3819 (.A(net3813),
    .X(net3819));
 sky130_fd_sc_hd__buf_1 place3565 (.A(_00029_),
    .X(net3565));
 sky130_fd_sc_hd__buf_8 place3795 (.A(net393),
    .X(net3795));
 sky130_fd_sc_hd__buf_6 place3575 (.A(_03225_),
    .X(net3575));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(key[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(key[88]));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(text_in[104]));
 sky130_fd_sc_hd__buf_1 place3577 (.A(_02138_),
    .X(net3577));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(key[87]));
 sky130_fd_sc_hd__buf_1 place3583 (.A(_09591_),
    .X(net3583));
 sky130_fd_sc_hd__buf_1 place3585 (.A(_08911_),
    .X(net3585));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(key[66]));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(key[58]));
 sky130_fd_sc_hd__buf_12 place3863 (.A(_11075_),
    .X(net3863));
 sky130_fd_sc_hd__buf_1 place3586 (.A(_08585_),
    .X(net3586));
 sky130_fd_sc_hd__buf_8 place3925 (.A(_09406_),
    .X(net3925));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(key[65]));
 sky130_fd_sc_hd__buf_1 place3589 (.A(_06643_),
    .X(net3589));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(key[64]));
 sky130_fd_sc_hd__buf_12 place3859 (.A(_11109_),
    .X(net3859));
 sky130_fd_sc_hd__buf_12 place3855 (.A(_11125_),
    .X(net3855));
 sky130_fd_sc_hd__clkbuf_2 place3876 (.A(net3871),
    .X(net3876));
 sky130_fd_sc_hd__buf_12 place3849 (.A(_11622_),
    .X(net3849));
 sky130_fd_sc_hd__buf_12 place3851 (.A(net410),
    .X(net3851));
 sky130_fd_sc_hd__buf_1 place3860 (.A(net3859),
    .X(net3860));
 sky130_fd_sc_hd__buf_8 place3874 (.A(net3873),
    .X(net3874));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(key[60]));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(key[62]));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(key[59]));
 sky130_fd_sc_hd__buf_12 place3848 (.A(_11627_),
    .X(net3848));
 sky130_fd_sc_hd__buf_12 place3934 (.A(net3932),
    .X(net3934));
 sky130_fd_sc_hd__buf_8 place3926 (.A(_09406_),
    .X(net3926));
 sky130_fd_sc_hd__buf_12 place3862 (.A(_11103_),
    .X(net3862));
 sky130_fd_sc_hd__buf_12 place3873 (.A(net3871),
    .X(net3873));
 sky130_fd_sc_hd__buf_12 place3847 (.A(_11639_),
    .X(net3847));
 sky130_fd_sc_hd__buf_1 place3846 (.A(_11639_),
    .X(net3846));
 sky130_fd_sc_hd__buf_12 place3936 (.A(_09363_),
    .X(net3936));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(net3565));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(net3565));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(net3565));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(net3565));
 sky130_fd_sc_hd__buf_1 place3621 (.A(_06767_),
    .X(net3621));
 sky130_fd_sc_hd__buf_4 place3622 (.A(_06540_),
    .X(net3622));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_10040_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_07881_));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net3566));
 sky130_fd_sc_hd__buf_8 place3618 (.A(_08361_),
    .X(net3618));
 sky130_fd_sc_hd__buf_1 place3620 (.A(_07199_),
    .X(net3620));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net3566));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(net3565));
 sky130_fd_sc_hd__buf_1 place3615 (.A(_08902_),
    .X(net3615));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(key[40]));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(key[40]));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(key[48]));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(key[47]));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(key[46]));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net3566));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(net3567));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(key[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(key[28]));
 sky130_fd_sc_hd__buf_1 place3602 (.A(_01991_),
    .X(net3602));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(net3567));
 sky130_fd_sc_hd__buf_1 place3598 (.A(_11978_[0]),
    .X(net3598));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_01033_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(key[110]));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(key[116]));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(key[118]));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(key[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(key[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(key[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(key[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(key[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(key[33]));
 sky130_fd_sc_hd__buf_1 place3601 (.A(_01991_),
    .X(net3601));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(key[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(key[113]));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(key[100]));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(net3567));
 sky130_fd_sc_hd__buf_1 place3616 (.A(_08472_),
    .X(net3616));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_08429_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_08078_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(net3565));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_07457_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_06443_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_06412_));
 sky130_fd_sc_hd__buf_1 place3624 (.A(_06041_),
    .X(net3624));
 sky130_fd_sc_hd__buf_12 place3845 (.A(_11655_),
    .X(net3845));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_00114_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(net3567));
 sky130_fd_sc_hd__buf_12 place3831 (.A(_00776_),
    .X(net3831));
 sky130_fd_sc_hd__buf_4 place3829 (.A(_00783_),
    .X(net3829));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__buf_12 place3821 (.A(_00822_),
    .X(net3821));
 sky130_fd_sc_hd__buf_12 place3950 (.A(_08842_),
    .X(net3950));
 sky130_fd_sc_hd__buf_1 place3949 (.A(_08842_),
    .X(net3949));
 sky130_fd_sc_hd__buf_1 place3812 (.A(net3811),
    .X(net3812));
 sky130_fd_sc_hd__buf_12 place3811 (.A(_00830_),
    .X(net3811));
 sky130_fd_sc_hd__buf_1 place3810 (.A(_00830_),
    .X(net3810));
 sky130_fd_sc_hd__buf_12 place3809 (.A(_00843_),
    .X(net3809));
 sky130_fd_sc_hd__buf_12 place3808 (.A(_00843_),
    .X(net3808));
 sky130_fd_sc_hd__buf_1 place3801 (.A(net3800),
    .X(net3801));
 sky130_fd_sc_hd__buf_12 place3800 (.A(net3799),
    .X(net3800));
 sky130_fd_sc_hd__buf_6 place3942 (.A(_08860_),
    .X(net3942));
 sky130_fd_sc_hd__buf_1 place3822 (.A(net3821),
    .X(net3822));
 sky130_fd_sc_hd__buf_8 place3823 (.A(_00822_),
    .X(net3823));
 sky130_fd_sc_hd__buf_12 place3839 (.A(_11684_),
    .X(net3839));
 sky130_fd_sc_hd__buf_8 place3817 (.A(net3813),
    .X(net3817));
 sky130_fd_sc_hd__buf_1 place3816 (.A(net3813),
    .X(net3816));
 sky130_fd_sc_hd__buf_12 place3796 (.A(_01353_),
    .X(net3796));
 sky130_fd_sc_hd__buf_1 place3815 (.A(net3813),
    .X(net3815));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__buf_12 place3792 (.A(_01367_),
    .X(net3792));
 sky130_fd_sc_hd__buf_8 place3791 (.A(net392),
    .X(net3791));
 sky130_fd_sc_hd__buf_1 place3790 (.A(_01367_),
    .X(net3790));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__buf_12 place3789 (.A(_01373_),
    .X(net3789));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__buf_8 place3787 (.A(_01379_),
    .X(net3787));
 sky130_fd_sc_hd__buf_12 place3786 (.A(_01379_),
    .X(net3786));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__buf_12 place3780 (.A(_01395_),
    .X(net3780));
 sky130_fd_sc_hd__buf_12 place3779 (.A(net3778),
    .X(net3779));
 sky130_fd_sc_hd__buf_12 place3778 (.A(_01881_),
    .X(net3778));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__buf_6 place3770 (.A(_01891_),
    .X(net3770));
 sky130_fd_sc_hd__buf_6 place3776 (.A(net3775),
    .X(net3776));
 sky130_fd_sc_hd__buf_12 place3775 (.A(net3770),
    .X(net3775));
 sky130_fd_sc_hd__buf_1 place3766 (.A(net3765),
    .X(net3766));
 sky130_fd_sc_hd__buf_12 place3762 (.A(_01929_),
    .X(net3762));
 sky130_fd_sc_hd__buf_12 place3774 (.A(net3770),
    .X(net3774));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__buf_1 place3747 (.A(net3746),
    .X(net3747));
 sky130_fd_sc_hd__inv_16 clkload1 (.A(clknet_3_1_0_clk));
 sky130_fd_sc_hd__buf_12 place3737 (.A(_02480_),
    .X(net3737));
 sky130_fd_sc_hd__buf_12 place3736 (.A(_02480_),
    .X(net3736));
 sky130_fd_sc_hd__buf_6 place3754 (.A(_01968_),
    .X(net3754));
 sky130_fd_sc_hd__buf_12 place3724 (.A(_02992_),
    .X(net3724));
 sky130_fd_sc_hd__buf_6 place3753 (.A(_01968_),
    .X(net3753));
 sky130_fd_sc_hd__buf_8 place3740 (.A(_02472_),
    .X(net3740));
 sky130_fd_sc_hd__clkinv_16 clkload3 (.A(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkinv_16 clkload2 (.A(clknet_3_2_0_clk));
 sky130_fd_sc_hd__buf_1 place3726 (.A(_02986_),
    .X(net3726));
 sky130_fd_sc_hd__buf_12 place3734 (.A(_02489_),
    .X(net3734));
 sky130_fd_sc_hd__buf_1 place3731 (.A(_02504_),
    .X(net3731));
 sky130_fd_sc_hd__buf_1 place3730 (.A(_02504_),
    .X(net3730));
 sky130_fd_sc_hd__buf_8 place3719 (.A(_03017_),
    .X(net3719));
 sky130_fd_sc_hd__buf_12 place3720 (.A(_03017_),
    .X(net3720));
 sky130_fd_sc_hd__buf_12 place3712 (.A(_03086_),
    .X(net3712));
 sky130_fd_sc_hd__buf_1 place3711 (.A(_03743_),
    .X(net3711));
 sky130_fd_sc_hd__buf_12 place3716 (.A(_03047_),
    .X(net3716));
 sky130_fd_sc_hd__buf_6 place3760 (.A(_01950_),
    .X(net3760));
 sky130_fd_sc_hd__buf_1 place3713 (.A(_03086_),
    .X(net3713));
 sky130_fd_sc_hd__buf_1 place3735 (.A(net3734),
    .X(net3735));
 sky130_fd_sc_hd__buf_8 place3722 (.A(_03012_),
    .X(net3722));
 sky130_fd_sc_hd__inv_8 clkload4 (.A(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkinv_16 clkload5 (.A(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkinv_16 clkload6 (.A(clknet_3_7_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload8 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__bufinv_16 clkload7 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkinv_4 clkload9 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkinv_4 clkload10 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__buf_1 place3761 (.A(_01950_),
    .X(net3761));
 sky130_fd_sc_hd__inv_8 clkload11 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__inv_8 clkload12 (.A(clknet_leaf_89_clk));
 sky130_fd_sc_hd__buf_1 place3637 (.A(_03179_),
    .X(net3637));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_00022_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_00019_));
 sky130_fd_sc_hd__buf_12 place3635 (.A(_11997_[0]),
    .X(net3635));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_00015_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_00019_));
 sky130_fd_sc_hd__inv_8 clkload13 (.A(clknet_leaf_90_clk));
 sky130_fd_sc_hd__inv_8 clkload14 (.A(clknet_leaf_91_clk));
 sky130_fd_sc_hd__buf_12 place3710 (.A(_05884_),
    .X(net3710));
 sky130_fd_sc_hd__buf_2 rebuffer22 (.A(net408),
    .X(net409));
 sky130_fd_sc_hd__buf_8 place3767 (.A(_01921_),
    .X(net3767));
 sky130_fd_sc_hd__buf_12 place3709 (.A(_05900_),
    .X(net3709));
 sky130_fd_sc_hd__bufinv_16 clkload20 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkinv_8 clkload25 (.A(clknet_leaf_81_clk));
 sky130_fd_sc_hd__buf_1 place3705 (.A(_06035_),
    .X(net3705));
 sky130_fd_sc_hd__clkbuf_8 clkload34 (.A(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkinv_8 clkload32 (.A(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkinv_8 clkload33 (.A(clknet_leaf_78_clk));
 sky130_fd_sc_hd__inv_8 clkload35 (.A(clknet_leaf_80_clk));
 sky130_fd_sc_hd__buf_8 place3700 (.A(_06505_),
    .X(net3700));
 sky130_fd_sc_hd__inv_12 clkload39 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__inv_12 clkload40 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__buf_12 place3690 (.A(_08238_),
    .X(net3690));
 sky130_fd_sc_hd__inv_6 clkload19 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__buf_1 place3794 (.A(net3792),
    .X(net3794));
 sky130_fd_sc_hd__buf_1 place3768 (.A(_01921_),
    .X(net3768));
 sky130_fd_sc_hd__buf_1 place3707 (.A(_05988_),
    .X(net3707));
 sky130_fd_sc_hd__clkinv_8 clkload23 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload30 (.A(clknet_leaf_67_clk));
 sky130_fd_sc_hd__inv_12 clkload29 (.A(clknet_leaf_88_clk));
 sky130_fd_sc_hd__buf_8 place3689 (.A(_08244_),
    .X(net3689));
 sky130_fd_sc_hd__clkinvlp_4 clkload52 (.A(clknet_leaf_28_clk));
 sky130_fd_sc_hd__bufinv_16 clkload54 (.A(clknet_leaf_44_clk));
 sky130_fd_sc_hd__inv_12 clkload58 (.A(clknet_leaf_55_clk));
 sky130_fd_sc_hd__inv_12 clkload57 (.A(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload56 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__buf_1 place3684 (.A(_08812_),
    .X(net3684));
 sky130_fd_sc_hd__clkinv_2 clkload60 (.A(clknet_leaf_57_clk));
 sky130_fd_sc_hd__buf_1 place3657 (.A(_00784_),
    .X(net3657));
 sky130_fd_sc_hd__buf_1 place3646 (.A(_01936_),
    .X(net3646));
 sky130_fd_sc_hd__buf_12 rebuffer16 (.A(_05937_),
    .X(net403));
 sky130_fd_sc_hd__buf_1 rebuffer17 (.A(_05937_),
    .X(net404));
 sky130_fd_sc_hd__buf_1 place3644 (.A(net3643),
    .X(net3644));
 sky130_fd_sc_hd__buf_1 place3663 (.A(_11628_),
    .X(net3663));
 sky130_fd_sc_hd__buf_12 place3649 (.A(_01892_),
    .X(net3649));
 sky130_fd_sc_hd__buf_1 place3664 (.A(_11628_),
    .X(net3664));
 sky130_fd_sc_hd__buf_1 place3647 (.A(_01936_),
    .X(net3647));
 sky130_fd_sc_hd__buf_12 place3643 (.A(_02438_),
    .X(net3643));
 sky130_fd_sc_hd__buf_1 place3659 (.A(_00777_),
    .X(net3659));
 sky130_fd_sc_hd__buf_12 place3640 (.A(_02525_),
    .X(net3640));
 sky130_fd_sc_hd__buf_1 place3641 (.A(_02525_),
    .X(net3641));
 sky130_fd_sc_hd__buf_1 rebuffer20 (.A(net406),
    .X(net407));
 sky130_fd_sc_hd__buf_12 place3642 (.A(_02467_),
    .X(net3642));
 sky130_fd_sc_hd__buf_1 place3655 (.A(_01354_),
    .X(net3655));
 sky130_fd_sc_hd__or2_2 clone12 (.A(_06536_),
    .B(_06534_),
    .X(net399));
 sky130_fd_sc_hd__buf_1 rebuffer5 (.A(_01367_),
    .X(net392));
 sky130_fd_sc_hd__buf_12 place3670 (.A(_11076_),
    .X(net3670));
 sky130_fd_sc_hd__inv_6 clkload63 (.A(clknet_leaf_62_clk));
 sky130_fd_sc_hd__inv_8 clkload62 (.A(clknet_leaf_61_clk));
 sky130_fd_sc_hd__buf_12 place3667 (.A(_11214_),
    .X(net3667));
 sky130_fd_sc_hd__buf_1 place3668 (.A(_11076_),
    .X(net3668));
 sky130_fd_sc_hd__buf_8 place3669 (.A(_11076_),
    .X(net3669));
 sky130_fd_sc_hd__buf_8 place3676 (.A(_09936_),
    .X(net3676));
 sky130_fd_sc_hd__inv_6 clkload18 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkinv_4 clkload59 (.A(clknet_leaf_56_clk));
 sky130_fd_sc_hd__inv_6 clkload17 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__buf_6 place3674 (.A(_10528_),
    .X(net3674));
 sky130_fd_sc_hd__buf_12 place3678 (.A(_09364_),
    .X(net3678));
 sky130_fd_sc_hd__buf_8 place3675 (.A(_10509_),
    .X(net3675));
 sky130_fd_sc_hd__clkinvlp_4 clkload53 (.A(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload55 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkinv_8 clkload22 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__buf_12 place3677 (.A(_09375_),
    .X(net3677));
 sky130_fd_sc_hd__clkinv_8 clkload21 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__buf_1 place3683 (.A(_08812_),
    .X(net3683));
 sky130_fd_sc_hd__inv_4 clkload44 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkinv_8 clkload43 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hd__inv_12 clkload28 (.A(clknet_leaf_87_clk));
 sky130_fd_sc_hd__inv_6 clkload42 (.A(clknet_leaf_30_clk));
 sky130_fd_sc_hd__buf_1 place3687 (.A(_08330_),
    .X(net3687));
 sky130_fd_sc_hd__inv_6 clkload41 (.A(clknet_leaf_29_clk));
 sky130_fd_sc_hd__buf_1 place3691 (.A(_07684_),
    .X(net3691));
 sky130_fd_sc_hd__inv_8 clkload36 (.A(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload38 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__buf_1 place3697 (.A(_07122_),
    .X(net3697));
 sky130_fd_sc_hd__inv_12 clkload27 (.A(clknet_leaf_86_clk));
 sky130_fd_sc_hd__buf_12 place3701 (.A(_06505_),
    .X(net3701));
 sky130_fd_sc_hd__clkinv_8 clkload26 (.A(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkinv_8 clkload37 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkinv_8 clkload31 (.A(clknet_leaf_70_clk));
 sky130_fd_sc_hd__buf_1 place3699 (.A(_06542_),
    .X(net3699));
 sky130_fd_sc_hd__inv_6 clkload24 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__buf_8 place3708 (.A(_05917_),
    .X(net3708));
 sky130_fd_sc_hd__buf_1 place3688 (.A(_08244_),
    .X(net3688));
 sky130_fd_sc_hd__buf_12 place3685 (.A(_08806_),
    .X(net3685));
 sky130_fd_sc_hd__clkinv_1 clkload16 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__inv_6 clkload15 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__buf_1 place3681 (.A(_08858_),
    .X(net3681));
 sky130_fd_sc_hd__buf_1 place3680 (.A(_08931_),
    .X(net3680));
 sky130_fd_sc_hd__inv_12 clkload47 (.A(clknet_leaf_37_clk));
 sky130_fd_sc_hd__inv_8 clkload46 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkinv_8 clkload45 (.A(clknet_leaf_34_clk));
 sky130_fd_sc_hd__buf_1 place3682 (.A(_08818_),
    .X(net3682));
 sky130_fd_sc_hd__buf_1 place3679 (.A(_09016_),
    .X(net3679));
 sky130_fd_sc_hd__inv_16 clkload48 (.A(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload49 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__bufinv_16 clkload51 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__bufinv_16 clkload50 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__inv_6 clkload61 (.A(clknet_leaf_60_clk));
 sky130_fd_sc_hd__buf_1 place3666 (.A(_11291_),
    .X(net3666));
 sky130_fd_sc_hd__buf_12 place3665 (.A(_11618_),
    .X(net3665));
 sky130_fd_sc_hd__inv_6 clkload64 (.A(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload66 (.A(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload65 (.A(clknet_leaf_64_clk));
 sky130_fd_sc_hd__buf_12 place3662 (.A(_11628_),
    .X(net3662));
 sky130_fd_sc_hd__buf_8 place3661 (.A(_11696_),
    .X(net3661));
 sky130_fd_sc_hd__inv_12 clkload69 (.A(clknet_leaf_72_clk));
 sky130_fd_sc_hd__inv_12 clkload68 (.A(clknet_leaf_69_clk));
 sky130_fd_sc_hd__inv_6 clkload67 (.A(clknet_leaf_68_clk));
 sky130_fd_sc_hd__bufinv_16 clkload70 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__bufinv_16 clkload71 (.A(clknet_leaf_40_clk));
 sky130_fd_sc_hd__bufinv_16 clkload72 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__buf_1 place3660 (.A(_11707_),
    .X(net3660));
 sky130_fd_sc_hd__buf_4 rebuffer2 (.A(net388),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_1 clkload77 (.A(clknet_leaf_59_clk));
 sky130_fd_sc_hd__bufinv_16 clkload73 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__bufinv_16 clkload76 (.A(clknet_leaf_53_clk));
 sky130_fd_sc_hd__bufinv_16 clkload75 (.A(clknet_leaf_51_clk));
 sky130_fd_sc_hd__bufinv_16 clkload74 (.A(clknet_leaf_48_clk));
 sky130_fd_sc_hd__buf_1 place3658 (.A(_00784_),
    .X(net3658));
 sky130_fd_sc_hd__buf_1 rebuffer4 (.A(_10550_),
    .X(net391));
 sky130_fd_sc_hd__buf_6 rebuffer3 (.A(_10550_),
    .X(net390));
 sky130_fd_sc_hd__buf_6 clone11 (.A(ld_r),
    .X(net398));
 sky130_fd_sc_hd__and2_2 clone10 (.A(_08265_),
    .B(_08260_),
    .X(net397));
 sky130_fd_sc_hd__buf_1 rebuffer9 (.A(net395),
    .X(net396));
 sky130_fd_sc_hd__buf_8 rebuffer8 (.A(_11931_[0]),
    .X(net395));
 sky130_fd_sc_hd__buf_2 rebuffer7 (.A(_01367_),
    .X(net394));
 sky130_fd_sc_hd__buf_2 rebuffer6 (.A(_01367_),
    .X(net393));
 sky130_fd_sc_hd__buf_1 place3656 (.A(_01343_),
    .X(net3656));
 sky130_fd_sc_hd__buf_6 place3652 (.A(_01354_),
    .X(net3652));
 sky130_fd_sc_hd__buf_1 place3653 (.A(_01354_),
    .X(net3653));
 sky130_fd_sc_hd__buf_4 rebuffer15 (.A(net401),
    .X(net402));
 sky130_fd_sc_hd__buf_4 rebuffer14 (.A(_12227_[0]),
    .X(net401));
 sky130_fd_sc_hd__buf_12 place3650 (.A(_01886_),
    .X(net3650));
 sky130_fd_sc_hd__buf_8 place3651 (.A(_01439_),
    .X(net3651));
 sky130_fd_sc_hd__buf_1 place3654 (.A(_01354_),
    .X(net3654));
 sky130_fd_sc_hd__buf_1 place3648 (.A(_01892_),
    .X(net3648));
 sky130_fd_sc_hd__buf_1 place3645 (.A(_02033_),
    .X(net3645));
 sky130_fd_sc_hd__buf_1 rebuffer18 (.A(_07081_),
    .X(net405));
 sky130_fd_sc_hd__buf_1 place3671 (.A(_11071_),
    .X(net3671));
 sky130_fd_sc_hd__buf_4 rebuffer19 (.A(_07081_),
    .X(net406));
 sky130_fd_sc_hd__buf_12 rebuffer21 (.A(_09928_),
    .X(net408));
 sky130_fd_sc_hd__buf_1 place3638 (.A(_02993_),
    .X(net3638));
 sky130_fd_sc_hd__buf_1 rebuffer23 (.A(_11617_),
    .X(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_00019_));
 sky130_fd_sc_hd__buf_12 place3636 (.A(_11965_[0]),
    .X(net3636));
 sky130_fd_sc_hd__buf_1 place3634 (.A(_12029_[0]),
    .X(net3634));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_00019_));
 sky130_fd_sc_hd__buf_12 place3639 (.A(_02987_),
    .X(net3639));
 sky130_fd_sc_hd__buf_12 place3632 (.A(_12093_[0]),
    .X(net3632));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_00019_));
 sky130_fd_sc_hd__buf_1 place3631 (.A(_12257_[0]),
    .X(net3631));
 sky130_fd_sc_hd__buf_1 place3633 (.A(_12092_[0]),
    .X(net3633));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_00019_));
 sky130_fd_sc_hd__buf_12 place3672 (.A(_11065_),
    .X(net3672));
 sky130_fd_sc_hd__buf_1 place3673 (.A(_10534_),
    .X(net3673));
 sky130_fd_sc_hd__buf_1 place3686 (.A(_08806_),
    .X(net3686));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_00022_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_00022_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_00022_));
 sky130_fd_sc_hd__buf_6 place3630 (.A(_12365_[0]),
    .X(net3630));
 sky130_fd_sc_hd__buf_12 place3629 (.A(_12461_[0]),
    .X(net3629));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_00022_));
 sky130_fd_sc_hd__buf_6 place3628 (.A(_03684_),
    .X(net3628));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_00022_));
 sky130_fd_sc_hd__buf_1 place3627 (.A(_03766_),
    .X(net3627));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_00022_));
 sky130_fd_sc_hd__buf_12 place3626 (.A(_03824_),
    .X(net3626));
 sky130_fd_sc_hd__buf_1 place3692 (.A(_07684_),
    .X(net3692));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_00022_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_00022_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_00022_));
 sky130_fd_sc_hd__buf_12 place3693 (.A(_07684_),
    .X(net3693));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_00099_));
 sky130_fd_sc_hd__buf_1 place3694 (.A(_07684_),
    .X(net3694));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_00119_));
 sky130_fd_sc_hd__buf_1 place3625 (.A(_05600_),
    .X(net3625));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_00956_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net3566));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net3566));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net3566));
 sky130_fd_sc_hd__buf_1 place3613 (.A(_09465_),
    .X(net3613));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net3566));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net3566));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(key[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(key[101]));
 sky130_fd_sc_hd__buf_1 place4047 (.A(_05945_),
    .X(net4047));
 sky130_fd_sc_hd__buf_6 place4040 (.A(_05958_),
    .X(net4040));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__buf_12 place4027 (.A(_06537_),
    .X(net4027));
 sky130_fd_sc_hd__buf_8 place4026 (.A(_06537_),
    .X(net4026));
 sky130_fd_sc_hd__buf_1 place4020 (.A(_06565_),
    .X(net4020));
 sky130_fd_sc_hd__buf_1 place4018 (.A(_06569_),
    .X(net4018));
 sky130_fd_sc_hd__buf_12 place3715 (.A(_03047_),
    .X(net3715));
 sky130_fd_sc_hd__buf_12 place4015 (.A(net407),
    .X(net4015));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__buf_6 place4007 (.A(_07140_),
    .X(net4007));
 sky130_fd_sc_hd__buf_1 place4024 (.A(net4023),
    .X(net4024));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__buf_12 place4019 (.A(_06565_),
    .X(net4019));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__buf_8 place4029 (.A(_06537_),
    .X(net4029));
 sky130_fd_sc_hd__buf_12 place3968 (.A(_08286_),
    .X(net3968));
 sky130_fd_sc_hd__buf_12 place3963 (.A(_08290_),
    .X(net3963));
 sky130_fd_sc_hd__buf_6 place3977 (.A(_08266_),
    .X(net3977));
 sky130_fd_sc_hd__buf_1 place3965 (.A(net3964),
    .X(net3965));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__buf_1 place3898 (.A(_09977_),
    .X(net3898));
 sky130_fd_sc_hd__buf_8 place3897 (.A(_09977_),
    .X(net3897));
 sky130_fd_sc_hd__buf_1 place3889 (.A(_10090_),
    .X(net3889));
 sky130_fd_sc_hd__clkbuf_2 place3884 (.A(net3883),
    .X(net3884));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__buf_12 place3858 (.A(_11109_),
    .X(net3858));
 sky130_fd_sc_hd__buf_12 place3843 (.A(_11655_),
    .X(net3843));
 sky130_fd_sc_hd__buf_8 place3854 (.A(_11140_),
    .X(net3854));
 sky130_fd_sc_hd__buf_1 place3842 (.A(_11655_),
    .X(net3842));
 sky130_fd_sc_hd__buf_8 place3838 (.A(_11684_),
    .X(net3838));
 sky130_fd_sc_hd__buf_1 place3837 (.A(_11684_),
    .X(net3837));
 sky130_fd_sc_hd__buf_12 place3714 (.A(_03075_),
    .X(net3714));
 sky130_fd_sc_hd__buf_12 place3872 (.A(net3871),
    .X(net3872));
 sky130_fd_sc_hd__buf_1 place3844 (.A(net3843),
    .X(net3844));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__buf_8 place3806 (.A(_00855_),
    .X(net3806));
 sky130_fd_sc_hd__buf_12 place3784 (.A(_01384_),
    .X(net3784));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__buf_1 place3783 (.A(_01386_),
    .X(net3783));
 sky130_fd_sc_hd__buf_12 place3777 (.A(_01885_),
    .X(net3777));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__buf_1 place3785 (.A(_01384_),
    .X(net3785));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__buf_1 place3769 (.A(_01910_),
    .X(net3769));
 sky130_fd_sc_hd__buf_1 place3773 (.A(net3771),
    .X(net3773));
 sky130_fd_sc_hd__buf_6 place3759 (.A(_01950_),
    .X(net3759));
 sky130_fd_sc_hd__buf_6 place3758 (.A(_01950_),
    .X(net3758));
 sky130_fd_sc_hd__buf_12 place3757 (.A(_01954_),
    .X(net3757));
 sky130_fd_sc_hd__buf_8 place3756 (.A(_01954_),
    .X(net3756));
 sky130_fd_sc_hd__buf_12 place3748 (.A(_02443_),
    .X(net3748));
 sky130_fd_sc_hd__buf_1 place3750 (.A(_02437_),
    .X(net3750));
 sky130_fd_sc_hd__buf_12 place3751 (.A(_02437_),
    .X(net3751));
 sky130_fd_sc_hd__clkinv_16 clkload0 (.A(clknet_3_0_0_clk));
 sky130_fd_sc_hd__buf_12 place3725 (.A(_02986_),
    .X(net3725));
 sky130_fd_sc_hd__buf_1 place3728 (.A(_02980_),
    .X(net3728));
 sky130_fd_sc_hd__buf_12 place3749 (.A(net3748),
    .X(net3749));
 sky130_fd_sc_hd__buf_1 place3739 (.A(net3738),
    .X(net3739));
 sky130_fd_sc_hd__buf_1 place3718 (.A(net3717),
    .X(net3718));
 sky130_fd_sc_hd__buf_12 place3721 (.A(_03012_),
    .X(net3721));
 sky130_fd_sc_hd__buf_8 place3717 (.A(_03017_),
    .X(net3717));
 sky130_fd_sc_hd__buf_12 place3723 (.A(_03003_),
    .X(net3723));
 sky130_fd_sc_hd__buf_12 place3743 (.A(_02472_),
    .X(net3743));
 sky130_fd_sc_hd__buf_1 place3733 (.A(net3732),
    .X(net3733));
 sky130_fd_sc_hd__buf_12 place3727 (.A(_02980_),
    .X(net3727));
 sky130_fd_sc_hd__buf_12 place3729 (.A(_02504_),
    .X(net3729));
 sky130_fd_sc_hd__buf_6 place3742 (.A(_02472_),
    .X(net3742));
 sky130_fd_sc_hd__buf_12 place3732 (.A(_02489_),
    .X(net3732));
 sky130_fd_sc_hd__buf_8 place3741 (.A(_02472_),
    .X(net3741));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__buf_12 place3746 (.A(_02448_),
    .X(net3746));
 sky130_fd_sc_hd__buf_12 place3745 (.A(_02448_),
    .X(net3745));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__buf_12 place3752 (.A(_01968_),
    .X(net3752));
 sky130_fd_sc_hd__buf_8 place3755 (.A(_01954_),
    .X(net3755));
 sky130_fd_sc_hd__buf_8 place3764 (.A(_01929_),
    .X(net3764));
 sky130_fd_sc_hd__buf_12 place3763 (.A(_01929_),
    .X(net3763));
 sky130_fd_sc_hd__buf_1 place3772 (.A(net3771),
    .X(net3772));
 sky130_fd_sc_hd__buf_12 place3771 (.A(net3770),
    .X(net3771));
 sky130_fd_sc_hd__buf_12 place3765 (.A(_01921_),
    .X(net3765));
 sky130_fd_sc_hd__buf_8 place3782 (.A(_01386_),
    .X(net3782));
 sky130_fd_sc_hd__buf_12 place3781 (.A(_01386_),
    .X(net3781));
 sky130_fd_sc_hd__buf_12 place3788 (.A(_01373_),
    .X(net3788));
 sky130_fd_sc_hd__buf_12 place3798 (.A(_01353_),
    .X(net3798));
 sky130_fd_sc_hd__buf_12 place3797 (.A(_01353_),
    .X(net3797));
 sky130_fd_sc_hd__buf_12 place3802 (.A(_01342_),
    .X(net3802));
 sky130_fd_sc_hd__buf_12 place3799 (.A(_01348_),
    .X(net3799));
 sky130_fd_sc_hd__buf_1 place3814 (.A(net3813),
    .X(net3814));
 sky130_fd_sc_hd__buf_6 place3804 (.A(_00903_),
    .X(net3804));
 sky130_fd_sc_hd__buf_8 place3803 (.A(_00938_),
    .X(net3803));
 sky130_fd_sc_hd__buf_12 place3807 (.A(_00843_),
    .X(net3807));
 sky130_fd_sc_hd__buf_12 place3830 (.A(net3829),
    .X(net3830));
 sky130_fd_sc_hd__buf_1 place3828 (.A(net3827),
    .X(net3828));
 sky130_fd_sc_hd__buf_8 place3805 (.A(_00855_),
    .X(net3805));
 sky130_fd_sc_hd__buf_1 place3825 (.A(_00816_),
    .X(net3825));
 sky130_fd_sc_hd__buf_12 place3833 (.A(_11719_),
    .X(net3833));
 sky130_fd_sc_hd__buf_12 place3841 (.A(_11670_),
    .X(net3841));
 sky130_fd_sc_hd__buf_1 place3826 (.A(_00806_),
    .X(net3826));
 sky130_fd_sc_hd__buf_8 place3836 (.A(_11684_),
    .X(net3836));
 sky130_fd_sc_hd__buf_12 place3827 (.A(_00797_),
    .X(net3827));
 sky130_fd_sc_hd__buf_12 place3835 (.A(_11715_),
    .X(net3835));
 sky130_fd_sc_hd__buf_1 place3832 (.A(_11719_),
    .X(net3832));
 sky130_fd_sc_hd__buf_12 place3834 (.A(_11715_),
    .X(net3834));
 sky130_fd_sc_hd__buf_8 place3840 (.A(_11670_),
    .X(net3840));
 sky130_fd_sc_hd__buf_1 place3850 (.A(_11617_),
    .X(net3850));
 sky130_fd_sc_hd__buf_12 place3852 (.A(_11194_),
    .X(net3852));
 sky130_fd_sc_hd__buf_12 place3866 (.A(net3865),
    .X(net3866));
 sky130_fd_sc_hd__buf_1 place3875 (.A(net3871),
    .X(net3875));
 sky130_fd_sc_hd__buf_1 place3856 (.A(_11122_),
    .X(net3856));
 sky130_fd_sc_hd__buf_6 place3864 (.A(net3863),
    .X(net3864));
 sky130_fd_sc_hd__buf_1 place3853 (.A(_11140_),
    .X(net3853));
 sky130_fd_sc_hd__buf_12 place3861 (.A(_11103_),
    .X(net3861));
 sky130_fd_sc_hd__buf_12 place3868 (.A(net3867),
    .X(net3868));
 sky130_fd_sc_hd__buf_12 place3867 (.A(_11064_),
    .X(net3867));
 sky130_fd_sc_hd__buf_12 place3865 (.A(_11070_),
    .X(net3865));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__buf_1 place3880 (.A(net3879),
    .X(net3880));
 sky130_fd_sc_hd__buf_12 place3869 (.A(_10585_),
    .X(net3869));
 sky130_fd_sc_hd__buf_1 place3909 (.A(net3908),
    .X(net3909));
 sky130_fd_sc_hd__buf_12 place3881 (.A(_10541_),
    .X(net3881));
 sky130_fd_sc_hd__buf_12 place3870 (.A(_10574_),
    .X(net3870));
 sky130_fd_sc_hd__buf_12 place3879 (.A(net390),
    .X(net3879));
 sky130_fd_sc_hd__buf_1 place3924 (.A(_09406_),
    .X(net3924));
 sky130_fd_sc_hd__buf_12 place3906 (.A(net409),
    .X(net3906));
 sky130_fd_sc_hd__buf_12 place3883 (.A(_10507_),
    .X(net3883));
 sky130_fd_sc_hd__buf_12 place3888 (.A(net388),
    .X(net3888));
 sky130_fd_sc_hd__clkbuf_2 place3886 (.A(net3885),
    .X(net3886));
 sky130_fd_sc_hd__buf_12 place3890 (.A(_10073_),
    .X(net3890));
 sky130_fd_sc_hd__buf_12 place3900 (.A(_09972_),
    .X(net3900));
 sky130_fd_sc_hd__buf_8 place3894 (.A(_09998_),
    .X(net3894));
 sky130_fd_sc_hd__buf_12 place3895 (.A(_09990_),
    .X(net3895));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__buf_12 place3899 (.A(_09972_),
    .X(net3899));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__buf_1 place3914 (.A(_09412_),
    .X(net3914));
 sky130_fd_sc_hd__buf_1 place3905 (.A(net409),
    .X(net3905));
 sky130_fd_sc_hd__buf_1 place3922 (.A(_09406_),
    .X(net3922));
 sky130_fd_sc_hd__buf_6 place3910 (.A(_09432_),
    .X(net3910));
 sky130_fd_sc_hd__buf_8 place3951 (.A(_08838_),
    .X(net3951));
 sky130_fd_sc_hd__buf_12 place3933 (.A(net3932),
    .X(net3933));
 sky130_fd_sc_hd__buf_12 place3931 (.A(_09374_),
    .X(net3931));
 sky130_fd_sc_hd__buf_12 place3964 (.A(_08290_),
    .X(net3964));
 sky130_fd_sc_hd__buf_1 place3966 (.A(net3964),
    .X(net3966));
 sky130_fd_sc_hd__buf_1 place3941 (.A(_08860_),
    .X(net3941));
 sky130_fd_sc_hd__buf_1 place3935 (.A(_09363_),
    .X(net3935));
 sky130_fd_sc_hd__buf_1 place3940 (.A(net3939),
    .X(net3940));
 sky130_fd_sc_hd__buf_1 place3954 (.A(_08838_),
    .X(net3954));
 sky130_fd_sc_hd__buf_1 place3953 (.A(net3952),
    .X(net3953));
 sky130_fd_sc_hd__buf_12 place3956 (.A(_08817_),
    .X(net3956));
 sky130_fd_sc_hd__buf_12 place3957 (.A(_08811_),
    .X(net3957));
 sky130_fd_sc_hd__buf_12 place3960 (.A(_08293_),
    .X(net3960));
 sky130_fd_sc_hd__buf_8 place3976 (.A(_08266_),
    .X(net3976));
 sky130_fd_sc_hd__buf_1 place3962 (.A(_08290_),
    .X(net3962));
 sky130_fd_sc_hd__buf_12 place3970 (.A(_08284_),
    .X(net3970));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__buf_8 place3972 (.A(_08279_),
    .X(net3972));
 sky130_fd_sc_hd__buf_12 place3993 (.A(_07718_),
    .X(net3993));
 sky130_fd_sc_hd__buf_1 place4028 (.A(_06537_),
    .X(net4028));
 sky130_fd_sc_hd__buf_12 place3987 (.A(_07728_),
    .X(net3987));
 sky130_fd_sc_hd__buf_1 place3984 (.A(_07791_),
    .X(net3984));
 sky130_fd_sc_hd__buf_1 place4022 (.A(_06541_),
    .X(net4022));
 sky130_fd_sc_hd__buf_4 place4025 (.A(_06541_),
    .X(net4025));
 sky130_fd_sc_hd__buf_8 place3992 (.A(_07718_),
    .X(net3992));
 sky130_fd_sc_hd__buf_1 place3991 (.A(_07718_),
    .X(net3991));
 sky130_fd_sc_hd__buf_12 place4010 (.A(_07099_),
    .X(net4010));
 sky130_fd_sc_hd__buf_1 place4008 (.A(_07140_),
    .X(net4008));
 sky130_fd_sc_hd__buf_1 place4003 (.A(net4001),
    .X(net4003));
 sky130_fd_sc_hd__buf_12 place4000 (.A(_07237_),
    .X(net4000));
 sky130_fd_sc_hd__buf_1 place3998 (.A(_07675_),
    .X(net3998));
 sky130_fd_sc_hd__buf_6 place4051 (.A(net403),
    .X(net4051));
 sky130_fd_sc_hd__buf_12 place4009 (.A(_07131_),
    .X(net4009));
 sky130_fd_sc_hd__buf_1 place4006 (.A(_07140_),
    .X(net4006));
 sky130_fd_sc_hd__buf_12 place4001 (.A(_07190_),
    .X(net4001));
 sky130_fd_sc_hd__buf_12 place4005 (.A(_07163_),
    .X(net4005));
 sky130_fd_sc_hd__buf_12 place4011 (.A(_07099_),
    .X(net4011));
 sky130_fd_sc_hd__buf_1 place4014 (.A(net405),
    .X(net4014));
 sky130_fd_sc_hd__buf_12 place4013 (.A(net4012),
    .X(net4013));
 sky130_fd_sc_hd__buf_12 place4021 (.A(_06541_),
    .X(net4021));
 sky130_fd_sc_hd__buf_12 place4017 (.A(_06569_),
    .X(net4017));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__buf_6 place4046 (.A(_05945_),
    .X(net4046));
 sky130_fd_sc_hd__buf_12 place4033 (.A(_06503_),
    .X(net4033));
 sky130_fd_sc_hd__buf_12 place4120 (.A(net4119),
    .X(net4120));
 sky130_fd_sc_hd__buf_12 place4054 (.A(_05899_),
    .X(net4054));
 sky130_fd_sc_hd__buf_12 place4036 (.A(_06493_),
    .X(net4036));
 sky130_fd_sc_hd__buf_8 place4043 (.A(_05954_),
    .X(net4043));
 sky130_fd_sc_hd__buf_12 place4039 (.A(_05958_),
    .X(net4039));
 sky130_fd_sc_hd__buf_12 place4042 (.A(_05954_),
    .X(net4042));
 sky130_fd_sc_hd__buf_1 place4045 (.A(net4044),
    .X(net4045));
 sky130_fd_sc_hd__buf_12 place4050 (.A(net403),
    .X(net4050));
 sky130_fd_sc_hd__buf_12 place4049 (.A(net403),
    .X(net4049));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__buf_12 place4060 (.A(_03809_),
    .X(net4060));
 sky130_fd_sc_hd__buf_6 place4058 (.A(net4057),
    .X(net4058));
 sky130_fd_sc_hd__buf_1 place3612 (.A(_09517_),
    .X(net3612));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__buf_12 place4119 (.A(_05879_),
    .X(net4119));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(key[102]));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(key[103]));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(key[104]));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(key[106]));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(key[108]));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(key[109]));
 sky130_fd_sc_hd__buf_1 place3608 (.A(_11771_),
    .X(net3608));
 sky130_fd_sc_hd__buf_1 place3610 (.A(_11149_),
    .X(net3610));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(key[111]));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(key[113]));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(key[113]));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(key[113]));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(key[113]));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(key[114]));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(key[116]));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(key[116]));
 sky130_fd_sc_hd__buf_1 place3611 (.A(_10565_),
    .X(net3611));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(key[119]));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(key[116]));
 sky130_fd_sc_hd__buf_1 place3609 (.A(_11771_),
    .X(net3609));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(key[116]));
 sky130_fd_sc_hd__buf_1 place3607 (.A(_01427_),
    .X(net3607));
 sky130_fd_sc_hd__buf_1 place3606 (.A(_01433_),
    .X(net3606));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(key[121]));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(key[122]));
 sky130_fd_sc_hd__buf_1 place3604 (.A(_01493_),
    .X(net3604));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(key[123]));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(key[125]));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(key[125]));
 sky130_fd_sc_hd__buf_1 place3605 (.A(_01456_),
    .X(net3605));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(key[126]));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(key[127]));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(key[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(key[24]));
 sky130_fd_sc_hd__buf_8 place3600 (.A(_03119_),
    .X(net3600));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(key[23]));
 sky130_fd_sc_hd__buf_1 place3599 (.A(_03132_),
    .X(net3599));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(key[39]));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(key[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(key[36]));
 sky130_fd_sc_hd__buf_1 place3596 (.A(_12106_[0]),
    .X(net3596));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(key[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(key[34]));
 sky130_fd_sc_hd__buf_1 place4075 (.A(net4074),
    .X(net4075));
 sky130_fd_sc_hd__buf_8 place3597 (.A(_12102_[0]),
    .X(net3597));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(key[40]));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(key[3]));
 sky130_fd_sc_hd__buf_1 place3603 (.A(_01677_),
    .X(net3603));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(key[40]));
 sky130_fd_sc_hd__buf_1 place3614 (.A(_08983_),
    .X(net3614));
 sky130_fd_sc_hd__buf_1 place3593 (.A(_12299_[0]),
    .X(net3593));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(key[44]));
 sky130_fd_sc_hd__buf_1 place3617 (.A(_08472_),
    .X(net3617));
 sky130_fd_sc_hd__buf_1 place3595 (.A(_12225_[0]),
    .X(net3595));
 sky130_fd_sc_hd__buf_1 place3594 (.A(_12272_[0]),
    .X(net3594));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(key[44]));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(key[40]));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(key[44]));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(key[40]));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(key[41]));
 sky130_fd_sc_hd__buf_1 place3619 (.A(_08342_),
    .X(net3619));
 sky130_fd_sc_hd__buf_1 place3623 (.A(net3622),
    .X(net3623));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(key[44]));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(key[46]));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(key[44]));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(key[44]));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(key[46]));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(key[46]));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(key[46]));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(key[46]));
 sky130_fd_sc_hd__buf_1 place4240 (.A(net129),
    .X(net4240));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(key[46]));
 sky130_fd_sc_hd__buf_1 place3592 (.A(_12378_[0]),
    .X(net3592));
 sky130_fd_sc_hd__buf_1 place3591 (.A(_12433_[0]),
    .X(net3591));
 sky130_fd_sc_hd__buf_1 place4239 (.A(net129),
    .X(net4239));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(key[50]));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(key[51]));
 sky130_fd_sc_hd__buf_1 place4238 (.A(net4237),
    .X(net4238));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(key[53]));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(key[54]));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(key[55]));
 sky130_fd_sc_hd__buf_1 place3590 (.A(_12474_[0]),
    .X(net3590));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(key[56]));
 sky130_fd_sc_hd__buf_1 place3695 (.A(_07676_),
    .X(net3695));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(key[57]));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(key[67]));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(key[68]));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(key[70]));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(key[6]));
 sky130_fd_sc_hd__buf_1 place3587 (.A(_08489_),
    .X(net3587));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(key[78]));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(key[79]));
 sky130_fd_sc_hd__buf_1 place3580 (.A(_11257_),
    .X(net3580));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(key[81]));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(key[72]));
 sky130_fd_sc_hd__buf_8 place3696 (.A(_07668_),
    .X(net3696));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(key[73]));
 sky130_fd_sc_hd__buf_1 place3584 (.A(_09421_),
    .X(net3584));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(key[74]));
 sky130_fd_sc_hd__buf_6 place3588 (.A(_08461_),
    .X(net3588));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(key[75]));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(key[76]));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(key[77]));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(key[82]));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(key[83]));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(key[89]));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(key[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(key[90]));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(key[91]));
 sky130_fd_sc_hd__buf_1 place3581 (.A(_11234_),
    .X(net3581));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(key[94]));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(key[93]));
 sky130_fd_sc_hd__buf_1 place3698 (.A(_07100_),
    .X(net3698));
 sky130_fd_sc_hd__buf_6 place3582 (.A(_10211_),
    .X(net3582));
 sky130_fd_sc_hd__buf_6 place4229 (.A(\sa00_sr[7] ),
    .X(net4229));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(key[95]));
 sky130_fd_sc_hd__buf_12 place3579 (.A(_00889_),
    .X(net3579));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(key[95]));
 sky130_fd_sc_hd__buf_12 place4080 (.A(net4078),
    .X(net4080));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(key[95]));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(key[95]));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(key[95]));
 sky130_fd_sc_hd__buf_1 place3578 (.A(_01067_),
    .X(net3578));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(key[96]));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(key[98]));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(key[99]));
 sky130_fd_sc_hd__buf_8 place3702 (.A(_06505_),
    .X(net3702));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(ld));
 sky130_fd_sc_hd__buf_6 place4088 (.A(_03702_),
    .X(net4088));
 sky130_fd_sc_hd__buf_12 place4079 (.A(net4078),
    .X(net4079));
 sky130_fd_sc_hd__buf_1 place4228 (.A(\sa01_sr[0] ),
    .X(net4228));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(rst));
 sky130_fd_sc_hd__buf_12 place4084 (.A(_03714_),
    .X(net4084));
 sky130_fd_sc_hd__buf_12 place4086 (.A(_03702_),
    .X(net4086));
 sky130_fd_sc_hd__buf_12 place4089 (.A(_11860_[0]),
    .X(net4089));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(text_in[100]));
 sky130_fd_sc_hd__buf_12 place3703 (.A(_06487_),
    .X(net3703));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(text_in[101]));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(text_in[105]));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(text_in[106]));
 sky130_fd_sc_hd__buf_12 place4098 (.A(net4097),
    .X(net4098));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(text_in[107]));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(text_in[109]));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(text_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(text_in[110]));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(text_in[111]));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(text_in[112]));
 sky130_fd_sc_hd__buf_1 place4096 (.A(net4095),
    .X(net4096));
 sky130_fd_sc_hd__buf_12 place4092 (.A(_03647_),
    .X(net4092));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(text_in[113]));
 sky130_fd_sc_hd__buf_1 place4095 (.A(_03630_),
    .X(net4095));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(text_in[114]));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(text_in[114]));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(text_in[114]));
 sky130_fd_sc_hd__buf_12 place4105 (.A(_03592_),
    .X(net4105));
 sky130_fd_sc_hd__buf_8 place4097 (.A(_03624_),
    .X(net4097));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(text_in[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(text_in[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(text_in[21]));
 sky130_fd_sc_hd__buf_12 place4100 (.A(_03617_),
    .X(net4100));
 sky130_fd_sc_hd__buf_12 place4103 (.A(_03610_),
    .X(net4103));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(text_in[13]));
 sky130_fd_sc_hd__buf_8 place4179 (.A(\sa32_sub[7] ),
    .X(net4179));
 sky130_fd_sc_hd__buf_1 place4104 (.A(_03592_),
    .X(net4104));
 sky130_fd_sc_hd__buf_1 place4124 (.A(_03581_),
    .X(net4124));
 sky130_fd_sc_hd__buf_12 place4106 (.A(_03585_),
    .X(net4106));
 sky130_fd_sc_hd__buf_1 place4113 (.A(net4111),
    .X(net4113));
 sky130_fd_sc_hd__buf_1 place4135 (.A(\u0.w[2][9] ),
    .X(net4135));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__buf_1 place4109 (.A(_05970_),
    .X(net4109));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__buf_1 place4133 (.A(\u0.tmp_w[21] ),
    .X(net4133));
 sky130_fd_sc_hd__buf_1 place4131 (.A(\u0.tmp_w[24] ),
    .X(net4131));
 sky130_fd_sc_hd__buf_1 place4140 (.A(\u0.w[2][12] ),
    .X(net4140));
 sky130_fd_sc_hd__buf_1 place4177 (.A(\u0.w[0][11] ),
    .X(net4177));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__buf_1 place4157 (.A(\u0.w[1][0] ),
    .X(net4157));
 sky130_fd_sc_hd__buf_1 place4152 (.A(\u0.w[1][22] ),
    .X(net4152));
 sky130_fd_sc_hd__buf_1 place4141 (.A(\u0.w[2][11] ),
    .X(net4141));
 sky130_fd_sc_hd__buf_1 place4139 (.A(\u0.w[2][17] ),
    .X(net4139));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__buf_1 place4148 (.A(\u0.w[1][27] ),
    .X(net4148));
 sky130_fd_sc_hd__buf_1 place4149 (.A(\u0.w[1][26] ),
    .X(net4149));
 sky130_fd_sc_hd__buf_1 place4153 (.A(\u0.w[1][1] ),
    .X(net4153));
 sky130_fd_sc_hd__buf_1 place4154 (.A(\u0.w[1][17] ),
    .X(net4154));
 sky130_fd_sc_hd__buf_8 place4163 (.A(\u0.w[0][3] ),
    .X(net4163));
 sky130_fd_sc_hd__buf_1 place4162 (.A(\u0.w[0][4] ),
    .X(net4162));
 sky130_fd_sc_hd__buf_1 place4161 (.A(\u0.w[0][5] ),
    .X(net4161));
 sky130_fd_sc_hd__buf_1 place4175 (.A(\u0.w[0][13] ),
    .X(net4175));
 sky130_fd_sc_hd__buf_1 place4164 (.A(\u0.w[0][30] ),
    .X(net4164));
 sky130_fd_sc_hd__buf_12 place4172 (.A(\u0.w[0][21] ),
    .X(net4172));
 sky130_fd_sc_hd__buf_1 place4173 (.A(\u0.w[0][1] ),
    .X(net4173));
 sky130_fd_sc_hd__buf_1 place4188 (.A(\sa30_sub[3] ),
    .X(net4188));
 sky130_fd_sc_hd__buf_1 place4178 (.A(\u0.w[0][0] ),
    .X(net4178));
 sky130_fd_sc_hd__buf_1 place4180 (.A(\sa32_sub[3] ),
    .X(net4180));
 sky130_fd_sc_hd__buf_6 place4182 (.A(\sa31_sub[7] ),
    .X(net4182));
 sky130_fd_sc_hd__buf_1 place4181 (.A(\sa32_sub[1] ),
    .X(net4181));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(text_in[20]));
 sky130_fd_sc_hd__buf_1 place4185 (.A(\sa31_sub[1] ),
    .X(net4185));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(text_in[1]));
 sky130_fd_sc_hd__buf_1 place4194 (.A(\sa21_sub[1] ),
    .X(net4194));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(text_in[19]));
 sky130_fd_sc_hd__buf_6 place4197 (.A(\sa20_sub[5] ),
    .X(net4197));
 sky130_fd_sc_hd__buf_1 place4209 (.A(\sa10_sub[2] ),
    .X(net4209));
 sky130_fd_sc_hd__buf_8 place4227 (.A(\sa01_sr[1] ),
    .X(net4227));
 sky130_fd_sc_hd__buf_1 place4208 (.A(\sa20_sr[5] ),
    .X(net4208));
 sky130_fd_sc_hd__buf_1 place4204 (.A(\sa21_sr[4] ),
    .X(net4204));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__buf_1 place4220 (.A(\sa10_sr[0] ),
    .X(net4220));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(text_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(text_in[16]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__buf_1 place4222 (.A(\sa03_sr[2] ),
    .X(net4222));
 sky130_fd_sc_hd__buf_1 place4218 (.A(\sa10_sr[3] ),
    .X(net4218));
 sky130_fd_sc_hd__buf_1 place3560 (.A(_00105_),
    .X(net3560));
 sky130_fd_sc_hd__buf_1 place4224 (.A(\sa02_sr[2] ),
    .X(net4224));
 sky130_fd_sc_hd__buf_6 place4225 (.A(\sa01_sr[3] ),
    .X(net4225));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__buf_12 place4235 (.A(net129),
    .X(net4235));
 sky130_fd_sc_hd__buf_1 place4231 (.A(net4230),
    .X(net4231));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(text_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(text_in[17]));
 sky130_fd_sc_hd__buf_1 place3820 (.A(net3819),
    .X(net3820));
 sky130_fd_sc_hd__buf_12 place3824 (.A(_00816_),
    .X(net3824));
 sky130_fd_sc_hd__buf_1 place3744 (.A(_02461_),
    .X(net3744));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(text_in[127]));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(text_in[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(text_in[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(text_in[117]));
 sky130_fd_sc_hd__buf_8 place3706 (.A(_06035_),
    .X(net3706));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(text_in[118]));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(text_in[119]));
 sky130_fd_sc_hd__buf_1 place3569 (.A(_05794_),
    .X(net3569));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(text_in[11]));
 sky130_fd_sc_hd__buf_1 place3572 (.A(_07036_),
    .X(net3572));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(text_in[120]));
 sky130_fd_sc_hd__buf_1 place3573 (.A(_06097_),
    .X(net3573));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(text_in[121]));
 sky130_fd_sc_hd__buf_8 place3567 (.A(_00017_),
    .X(net3567));
 sky130_fd_sc_hd__buf_12 place3878 (.A(_10550_),
    .X(net3878));
 sky130_fd_sc_hd__buf_8 place3877 (.A(net391),
    .X(net3877));
 sky130_fd_sc_hd__buf_12 place3871 (.A(_10556_),
    .X(net3871));
 sky130_fd_sc_hd__buf_12 place3891 (.A(_10073_),
    .X(net3891));
 sky130_fd_sc_hd__buf_12 place3893 (.A(_09998_),
    .X(net3893));
 sky130_fd_sc_hd__buf_12 place3885 (.A(_10499_),
    .X(net3885));
 sky130_fd_sc_hd__buf_12 rebuffer1 (.A(_10494_),
    .X(net388));
 sky130_fd_sc_hd__buf_12 place3882 (.A(_10519_),
    .X(net3882));
 sky130_fd_sc_hd__buf_1 place3896 (.A(_09977_),
    .X(net3896));
 sky130_fd_sc_hd__buf_1 place3913 (.A(_09412_),
    .X(net3913));
 sky130_fd_sc_hd__buf_8 place3902 (.A(_09957_),
    .X(net3902));
 sky130_fd_sc_hd__buf_1 place3901 (.A(_09957_),
    .X(net3901));
 sky130_fd_sc_hd__buf_8 place3911 (.A(_09431_),
    .X(net3911));
 sky130_fd_sc_hd__buf_1 place3916 (.A(_09412_),
    .X(net3916));
 sky130_fd_sc_hd__buf_1 place3903 (.A(_09944_),
    .X(net3903));
 sky130_fd_sc_hd__buf_12 place3908 (.A(net3907),
    .X(net3908));
 sky130_fd_sc_hd__buf_12 place3904 (.A(_09935_),
    .X(net3904));
 sky130_fd_sc_hd__buf_12 place3907 (.A(_09922_),
    .X(net3907));
 sky130_fd_sc_hd__buf_12 place3917 (.A(_09412_),
    .X(net3917));
 sky130_fd_sc_hd__buf_12 place3912 (.A(_09431_),
    .X(net3912));
 sky130_fd_sc_hd__buf_1 place3921 (.A(_09406_),
    .X(net3921));
 sky130_fd_sc_hd__buf_6 place3920 (.A(_09406_),
    .X(net3920));
 sky130_fd_sc_hd__buf_6 place3919 (.A(_09406_),
    .X(net3919));
 sky130_fd_sc_hd__buf_1 place3918 (.A(_09406_),
    .X(net3918));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__buf_12 place3930 (.A(_09385_),
    .X(net3930));
 sky130_fd_sc_hd__buf_1 place3928 (.A(_09391_),
    .X(net3928));
 sky130_fd_sc_hd__buf_12 place3927 (.A(_09391_),
    .X(net3927));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__buf_1 place3967 (.A(_08286_),
    .X(net3967));
 sky130_fd_sc_hd__buf_12 place3929 (.A(_09385_),
    .X(net3929));
 sky130_fd_sc_hd__buf_12 place3952 (.A(_08838_),
    .X(net3952));
 sky130_fd_sc_hd__buf_12 place3932 (.A(_09369_),
    .X(net3932));
 sky130_fd_sc_hd__buf_12 place3937 (.A(_08930_),
    .X(net3937));
 sky130_fd_sc_hd__buf_12 place3938 (.A(_08896_),
    .X(net3938));
 sky130_fd_sc_hd__buf_8 place3945 (.A(_08849_),
    .X(net3945));
 sky130_fd_sc_hd__buf_1 place3944 (.A(_08849_),
    .X(net3944));
 sky130_fd_sc_hd__buf_8 place3939 (.A(_08860_),
    .X(net3939));
 sky130_fd_sc_hd__buf_12 place3943 (.A(_08849_),
    .X(net3943));
 sky130_fd_sc_hd__buf_1 place3948 (.A(net3946),
    .X(net3948));
 sky130_fd_sc_hd__buf_6 place3947 (.A(net3946),
    .X(net3947));
 sky130_fd_sc_hd__buf_12 place3946 (.A(_08842_),
    .X(net3946));
 sky130_fd_sc_hd__buf_12 place3955 (.A(_08827_),
    .X(net3955));
 sky130_fd_sc_hd__buf_1 place3959 (.A(net3958),
    .X(net3959));
 sky130_fd_sc_hd__buf_12 place3958 (.A(_08805_),
    .X(net3958));
 sky130_fd_sc_hd__buf_1 place3969 (.A(_08284_),
    .X(net3969));
 sky130_fd_sc_hd__buf_1 place3971 (.A(_08279_),
    .X(net3971));
 sky130_fd_sc_hd__buf_12 place3974 (.A(_08266_),
    .X(net3974));
 sky130_fd_sc_hd__buf_12 place3982 (.A(net3981),
    .X(net3982));
 sky130_fd_sc_hd__buf_12 place3973 (.A(_08266_),
    .X(net3973));
 sky130_fd_sc_hd__buf_1 place3979 (.A(net3978),
    .X(net3979));
 sky130_fd_sc_hd__buf_12 place3978 (.A(_08249_),
    .X(net3978));
 sky130_fd_sc_hd__buf_12 place4012 (.A(_07089_),
    .X(net4012));
 sky130_fd_sc_hd__buf_12 place3989 (.A(net3987),
    .X(net3989));
 sky130_fd_sc_hd__buf_8 place3983 (.A(_07791_),
    .X(net3983));
 sky130_fd_sc_hd__buf_12 place3980 (.A(_08243_),
    .X(net3980));
 sky130_fd_sc_hd__buf_12 place3981 (.A(_08237_),
    .X(net3981));
 sky130_fd_sc_hd__buf_12 place3985 (.A(_07776_),
    .X(net3985));
 sky130_fd_sc_hd__buf_12 place3988 (.A(net3987),
    .X(net3988));
 sky130_fd_sc_hd__buf_12 place3986 (.A(_07740_),
    .X(net3986));
 sky130_fd_sc_hd__buf_1 place4002 (.A(net4001),
    .X(net4002));
 sky130_fd_sc_hd__buf_12 place3997 (.A(_07675_),
    .X(net3997));
 sky130_fd_sc_hd__buf_12 place3996 (.A(_07683_),
    .X(net3996));
 sky130_fd_sc_hd__buf_12 place3994 (.A(_07704_),
    .X(net3994));
 sky130_fd_sc_hd__buf_12 place3995 (.A(_07683_),
    .X(net3995));
 sky130_fd_sc_hd__buf_12 place3999 (.A(_07667_),
    .X(net3999));
 sky130_fd_sc_hd__buf_6 place4041 (.A(_05958_),
    .X(net4041));
 sky130_fd_sc_hd__buf_1 place4034 (.A(net4033),
    .X(net4034));
 sky130_fd_sc_hd__buf_12 place4032 (.A(_06520_),
    .X(net4032));
 sky130_fd_sc_hd__buf_1 place4038 (.A(net4037),
    .X(net4038));
 sky130_fd_sc_hd__buf_12 place4037 (.A(_06486_),
    .X(net4037));
 sky130_fd_sc_hd__clkbuf_2 place4035 (.A(_06493_),
    .X(net4035));
 sky130_fd_sc_hd__buf_12 place4044 (.A(_05945_),
    .X(net4044));
 sky130_fd_sc_hd__buf_8 place4048 (.A(net404),
    .X(net4048));
 sky130_fd_sc_hd__buf_1 place4055 (.A(net4054),
    .X(net4055));
 sky130_fd_sc_hd__buf_12 place4057 (.A(_05883_),
    .X(net4057));
 sky130_fd_sc_hd__buf_12 place4056 (.A(_05890_),
    .X(net4056));
 sky130_fd_sc_hd__buf_6 place4059 (.A(_05883_),
    .X(net4059));
 sky130_fd_sc_hd__buf_1 place4121 (.A(_05879_),
    .X(net4121));
 sky130_fd_sc_hd__buf_1 place4061 (.A(_03734_),
    .X(net4061));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__buf_1 place4070 (.A(_02479_),
    .X(net4070));
 sky130_fd_sc_hd__buf_12 place4117 (.A(_05879_),
    .X(net4117));
 sky130_fd_sc_hd__buf_6 place4207 (.A(\sa20_sr[7] ),
    .X(net4207));
 sky130_fd_sc_hd__buf_1 place4150 (.A(\u0.w[1][25] ),
    .X(net4150));
 sky130_fd_sc_hd__buf_1 place4065 (.A(_03625_),
    .X(net4065));
 sky130_fd_sc_hd__buf_12 place4069 (.A(_03579_),
    .X(net4069));
 sky130_fd_sc_hd__buf_1 place4068 (.A(_03579_),
    .X(net4068));
 sky130_fd_sc_hd__buf_12 place4116 (.A(_05879_),
    .X(net4116));
 sky130_fd_sc_hd__buf_1 place4115 (.A(_05879_),
    .X(net4115));
 sky130_fd_sc_hd__buf_6 place4102 (.A(net4101),
    .X(net4102));
 sky130_fd_sc_hd__buf_12 place4062 (.A(_03724_),
    .X(net4062));
 sky130_fd_sc_hd__buf_8 place4118 (.A(net4117),
    .X(net4118));
 sky130_fd_sc_hd__buf_12 place4063 (.A(_03691_),
    .X(net4063));
 sky130_fd_sc_hd__buf_12 place4066 (.A(_03601_),
    .X(net4066));
 sky130_fd_sc_hd__buf_12 place4076 (.A(net4074),
    .X(net4076));
 sky130_fd_sc_hd__buf_6 place4077 (.A(net4074),
    .X(net4077));
 sky130_fd_sc_hd__buf_12 place4064 (.A(_03648_),
    .X(net4064));
 sky130_fd_sc_hd__buf_6 place4067 (.A(_03579_),
    .X(net4067));
 sky130_fd_sc_hd__buf_1 place4134 (.A(\u0.tmp_w[1] ),
    .X(net4134));
 sky130_fd_sc_hd__buf_1 place4127 (.A(\u0.tmp_w[5] ),
    .X(net4127));
 sky130_fd_sc_hd__buf_1 place4072 (.A(_11650_),
    .X(net4072));
 sky130_fd_sc_hd__buf_6 place4071 (.A(_01371_),
    .X(net4071));
 sky130_fd_sc_hd__buf_12 place4073 (.A(_03800_),
    .X(net4073));
 sky130_fd_sc_hd__buf_12 place4074 (.A(_03791_),
    .X(net4074));
 sky130_fd_sc_hd__buf_12 place4078 (.A(_03783_),
    .X(net4078));
 sky130_fd_sc_hd__buf_1 place4081 (.A(net4078),
    .X(net4081));
 sky130_fd_sc_hd__buf_12 place4087 (.A(_03702_),
    .X(net4087));
 sky130_fd_sc_hd__buf_12 place4082 (.A(_03777_),
    .X(net4082));
 sky130_fd_sc_hd__buf_1 place4099 (.A(_03624_),
    .X(net4099));
 sky130_fd_sc_hd__buf_1 place4085 (.A(net4084),
    .X(net4085));
 sky130_fd_sc_hd__buf_12 place4083 (.A(_03772_),
    .X(net4083));
 sky130_fd_sc_hd__buf_12 place4093 (.A(_03637_),
    .X(net4093));
 sky130_fd_sc_hd__buf_12 place4090 (.A(_03690_),
    .X(net4090));
 sky130_fd_sc_hd__buf_1 place4091 (.A(_03656_),
    .X(net4091));
 sky130_fd_sc_hd__buf_1 place4122 (.A(_05875_),
    .X(net4122));
 sky130_fd_sc_hd__buf_12 place4111 (.A(_05879_),
    .X(net4111));
 sky130_fd_sc_hd__buf_1 place4112 (.A(net4111),
    .X(net4112));
 sky130_fd_sc_hd__buf_1 place4110 (.A(_05885_),
    .X(net4110));
 sky130_fd_sc_hd__buf_12 place4094 (.A(_03630_),
    .X(net4094));
 sky130_fd_sc_hd__buf_12 place4107 (.A(_03578_),
    .X(net4107));
 sky130_fd_sc_hd__buf_1 place4130 (.A(\u0.tmp_w[25] ),
    .X(net4130));
 sky130_fd_sc_hd__buf_1 place4123 (.A(_03587_),
    .X(net4123));
 sky130_fd_sc_hd__buf_1 place4129 (.A(\u0.tmp_w[28] ),
    .X(net4129));
 sky130_fd_sc_hd__buf_1 place4128 (.A(\u0.tmp_w[29] ),
    .X(net4128));
 sky130_fd_sc_hd__buf_1 place4126 (.A(\u0.tmp_w[8] ),
    .X(net4126));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__buf_1 place4142 (.A(\u0.w[1][6] ),
    .X(net4142));
 sky130_fd_sc_hd__buf_1 place4143 (.A(\u0.w[1][5] ),
    .X(net4143));
 sky130_fd_sc_hd__buf_1 place4144 (.A(\u0.w[1][4] ),
    .X(net4144));
 sky130_fd_sc_hd__buf_1 place4145 (.A(\u0.w[1][30] ),
    .X(net4145));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__buf_1 place4146 (.A(\u0.w[1][29] ),
    .X(net4146));
 sky130_fd_sc_hd__buf_1 place4147 (.A(\u0.w[1][28] ),
    .X(net4147));
 sky130_fd_sc_hd__buf_1 place4191 (.A(\sa21_sub[7] ),
    .X(net4191));
 sky130_fd_sc_hd__buf_8 place4151 (.A(\u0.w[1][24] ),
    .X(net4151));
 sky130_fd_sc_hd__buf_1 place4206 (.A(\sa21_sr[0] ),
    .X(net4206));
 sky130_fd_sc_hd__buf_1 place4155 (.A(\u0.w[1][16] ),
    .X(net4155));
 sky130_fd_sc_hd__buf_1 place4156 (.A(\u0.w[1][13] ),
    .X(net4156));
 sky130_fd_sc_hd__buf_1 place4158 (.A(\u0.w[0][9] ),
    .X(net4158));
 sky130_fd_sc_hd__buf_1 place4159 (.A(\u0.w[0][7] ),
    .X(net4159));
 sky130_fd_sc_hd__buf_1 place4160 (.A(\u0.w[0][6] ),
    .X(net4160));
 sky130_fd_sc_hd__buf_1 place4165 (.A(\u0.w[0][29] ),
    .X(net4165));
 sky130_fd_sc_hd__buf_12 place4166 (.A(\u0.w[0][28] ),
    .X(net4166));
 sky130_fd_sc_hd__buf_1 place4167 (.A(\u0.w[0][27] ),
    .X(net4167));
 sky130_fd_sc_hd__buf_1 place4168 (.A(\u0.w[0][26] ),
    .X(net4168));
 sky130_fd_sc_hd__buf_1 place4169 (.A(\u0.w[0][25] ),
    .X(net4169));
 sky130_fd_sc_hd__buf_1 place4170 (.A(\u0.w[0][24] ),
    .X(net4170));
 sky130_fd_sc_hd__buf_1 place4171 (.A(\u0.w[0][22] ),
    .X(net4171));
 sky130_fd_sc_hd__buf_1 place4174 (.A(\u0.w[0][14] ),
    .X(net4174));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__buf_1 place4183 (.A(\sa31_sub[3] ),
    .X(net4183));
 sky130_fd_sc_hd__buf_12 place4176 (.A(\u0.w[0][12] ),
    .X(net4176));
 sky130_fd_sc_hd__buf_1 place4184 (.A(\sa31_sub[2] ),
    .X(net4184));
 sky130_fd_sc_hd__buf_1 place4186 (.A(\sa30_sub[7] ),
    .X(net4186));
 sky130_fd_sc_hd__buf_1 place4187 (.A(\sa30_sub[4] ),
    .X(net4187));
 sky130_fd_sc_hd__clkbuf_2 place4189 (.A(\sa30_sr[7] ),
    .X(net4189));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__buf_1 place4190 (.A(\sa30_sr[4] ),
    .X(net4190));
 sky130_fd_sc_hd__buf_1 place4192 (.A(\sa21_sub[3] ),
    .X(net4192));
 sky130_fd_sc_hd__buf_1 place4193 (.A(\sa21_sub[2] ),
    .X(net4193));
 sky130_fd_sc_hd__buf_1 place4195 (.A(\sa21_sub[0] ),
    .X(net4195));
 sky130_fd_sc_hd__buf_12 place4196 (.A(\sa20_sub[7] ),
    .X(net4196));
 sky130_fd_sc_hd__buf_1 place4200 (.A(\sa20_sub[2] ),
    .X(net4200));
 sky130_fd_sc_hd__buf_1 place4199 (.A(\sa20_sub[3] ),
    .X(net4199));
 sky130_fd_sc_hd__buf_1 place4198 (.A(\sa20_sub[4] ),
    .X(net4198));
 sky130_fd_sc_hd__buf_6 place4201 (.A(\sa20_sub[0] ),
    .X(net4201));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__buf_1 place4202 (.A(\sa21_sr[7] ),
    .X(net4202));
 sky130_fd_sc_hd__buf_1 place4203 (.A(\sa21_sr[5] ),
    .X(net4203));
 sky130_fd_sc_hd__buf_1 place4205 (.A(\sa21_sr[2] ),
    .X(net4205));
 sky130_fd_sc_hd__buf_1 place4210 (.A(\sa10_sub[1] ),
    .X(net4210));
 sky130_fd_sc_hd__buf_8 place4211 (.A(\sa10_sub[0] ),
    .X(net4211));
 sky130_fd_sc_hd__buf_1 place4212 (.A(\sa12_sr[7] ),
    .X(net4212));
 sky130_fd_sc_hd__buf_1 place4214 (.A(\sa11_sr[7] ),
    .X(net4214));
 sky130_fd_sc_hd__buf_12 place4219 (.A(\sa10_sr[2] ),
    .X(net4219));
 sky130_fd_sc_hd__buf_1 place4213 (.A(\sa12_sr[2] ),
    .X(net4213));
 sky130_fd_sc_hd__buf_1 place4216 (.A(\sa10_sr[7] ),
    .X(net4216));
 sky130_fd_sc_hd__buf_1 place4215 (.A(\sa11_sr[0] ),
    .X(net4215));
 sky130_fd_sc_hd__buf_1 place4217 (.A(\sa10_sr[4] ),
    .X(net4217));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__buf_12 place4234 (.A(net129),
    .X(net4234));
 sky130_fd_sc_hd__buf_1 place4221 (.A(\sa03_sr[7] ),
    .X(net4221));
 sky130_fd_sc_hd__buf_12 place4233 (.A(net129),
    .X(net4233));
 sky130_fd_sc_hd__buf_1 place4223 (.A(\sa02_sr[7] ),
    .X(net4223));
 sky130_fd_sc_hd__buf_6 place4226 (.A(\sa01_sr[2] ),
    .X(net4226));
 sky130_fd_sc_hd__buf_12 place4232 (.A(net129),
    .X(net4232));
 sky130_fd_sc_hd__buf_12 place4236 (.A(net4235),
    .X(net4236));
 sky130_fd_sc_hd__clkbuf_16 place4230 (.A(ld_r),
    .X(net4230));
 sky130_fd_sc_hd__buf_12 place4237 (.A(net129),
    .X(net4237));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__buf_1 place4053 (.A(net403),
    .X(net4053));
 sky130_fd_sc_hd__buf_1 place4052 (.A(net403),
    .X(net4052));
 sky130_fd_sc_hd__buf_8 place4031 (.A(_06537_),
    .X(net4031));
 sky130_fd_sc_hd__buf_1 place3562 (.A(_00118_),
    .X(net3562));
 sky130_fd_sc_hd__buf_1 place3561 (.A(_00097_),
    .X(net3561));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(text_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(text_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(text_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(text_in[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(text_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(text_in[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(text_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(text_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(text_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(text_in[38]));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(text_in[39]));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(text_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(text_in[40]));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(text_in[42]));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(text_in[42]));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(text_in[42]));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(text_in[43]));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(text_in[45]));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(text_in[46]));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(text_in[47]));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(text_in[48]));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(text_in[51]));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(text_in[52]));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(text_in[53]));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(text_in[54]));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(text_in[55]));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(text_in[56]));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(text_in[57]));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(text_in[58]));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(text_in[59]));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(text_in[61]));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(text_in[64]));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(text_in[65]));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(text_in[67]));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(text_in[69]));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(text_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(text_in[70]));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(text_in[71]));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(text_in[72]));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(text_in[73]));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(text_in[74]));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(text_in[75]));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(text_in[76]));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(text_in[77]));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(text_in[78]));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(text_in[79]));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(text_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(text_in[81]));
 sky130_fd_sc_hd__diode_2 ANTENNA_263 (.DIODE(text_in[83]));
 sky130_fd_sc_hd__diode_2 ANTENNA_264 (.DIODE(text_in[84]));
 sky130_fd_sc_hd__diode_2 ANTENNA_265 (.DIODE(text_in[85]));
 sky130_fd_sc_hd__diode_2 ANTENNA_266 (.DIODE(text_in[86]));
 sky130_fd_sc_hd__diode_2 ANTENNA_267 (.DIODE(text_in[87]));
 sky130_fd_sc_hd__diode_2 ANTENNA_268 (.DIODE(text_in[89]));
 sky130_fd_sc_hd__diode_2 ANTENNA_269 (.DIODE(text_in[89]));
 sky130_fd_sc_hd__diode_2 ANTENNA_270 (.DIODE(text_in[89]));
 sky130_fd_sc_hd__diode_2 ANTENNA_271 (.DIODE(text_in[89]));
 sky130_fd_sc_hd__diode_2 ANTENNA_272 (.DIODE(text_in[89]));
 sky130_fd_sc_hd__diode_2 ANTENNA_273 (.DIODE(text_in[89]));
 sky130_fd_sc_hd__diode_2 ANTENNA_274 (.DIODE(text_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_275 (.DIODE(text_in[90]));
 sky130_fd_sc_hd__diode_2 ANTENNA_276 (.DIODE(text_in[91]));
 sky130_fd_sc_hd__diode_2 ANTENNA_277 (.DIODE(text_in[92]));
 sky130_fd_sc_hd__diode_2 ANTENNA_278 (.DIODE(text_in[93]));
 sky130_fd_sc_hd__diode_2 ANTENNA_279 (.DIODE(text_in[95]));
 sky130_fd_sc_hd__diode_2 ANTENNA_280 (.DIODE(text_in[96]));
 sky130_fd_sc_hd__diode_2 ANTENNA_281 (.DIODE(text_in[97]));
 sky130_fd_sc_hd__diode_2 ANTENNA_282 (.DIODE(text_in[98]));
 sky130_fd_sc_hd__diode_2 ANTENNA_283 (.DIODE(text_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_284 (.DIODE(net3561));
 sky130_fd_sc_hd__diode_2 ANTENNA_285 (.DIODE(_00096_));
 sky130_fd_sc_hd__diode_2 ANTENNA_286 (.DIODE(key[120]));
 sky130_fd_sc_hd__diode_2 ANTENNA_287 (.DIODE(key[127]));
 sky130_fd_sc_hd__diode_2 ANTENNA_288 (.DIODE(key[127]));
 sky130_fd_sc_hd__diode_2 ANTENNA_289 (.DIODE(key[127]));
 sky130_fd_sc_hd__diode_2 ANTENNA_290 (.DIODE(key[127]));
 sky130_fd_sc_hd__diode_2 ANTENNA_291 (.DIODE(key[127]));
 sky130_fd_sc_hd__diode_2 ANTENNA_292 (.DIODE(key[43]));
 sky130_fd_sc_hd__diode_2 ANTENNA_293 (.DIODE(key[43]));
 sky130_fd_sc_hd__diode_2 ANTENNA_294 (.DIODE(key[43]));
 sky130_fd_sc_hd__diode_2 ANTENNA_295 (.DIODE(key[43]));
 sky130_fd_sc_hd__diode_2 ANTENNA_296 (.DIODE(key[97]));
 sky130_fd_sc_hd__diode_2 ANTENNA_297 (.DIODE(text_in[113]));
 sky130_fd_sc_hd__diode_2 ANTENNA_298 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_299 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_300 (.DIODE(_01621_));
 sky130_fd_sc_hd__diode_2 ANTENNA_301 (.DIODE(net3560));
 sky130_fd_sc_hd__diode_2 ANTENNA_302 (.DIODE(_06575_));
 sky130_fd_sc_hd__diode_2 ANTENNA_303 (.DIODE(_08936_));
 sky130_fd_sc_hd__diode_2 ANTENNA_304 (.DIODE(_09482_));
 sky130_fd_sc_hd__diode_2 ANTENNA_305 (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_306 (.DIODE(key[112]));
 sky130_fd_sc_hd__diode_2 ANTENNA_307 (.DIODE(key[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_308 (.DIODE(key[127]));
 sky130_fd_sc_hd__diode_2 ANTENNA_309 (.DIODE(key[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_310 (.DIODE(key[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_311 (.DIODE(key[42]));
 sky130_fd_sc_hd__diode_2 ANTENNA_312 (.DIODE(key[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_313 (.DIODE(key[71]));
 sky130_fd_sc_hd__diode_2 ANTENNA_314 (.DIODE(key[84]));
 sky130_fd_sc_hd__diode_2 ANTENNA_315 (.DIODE(text_in[103]));
 sky130_fd_sc_hd__diode_2 ANTENNA_316 (.DIODE(text_in[108]));
 sky130_fd_sc_hd__diode_2 ANTENNA_317 (.DIODE(text_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_318 (.DIODE(text_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_319 (.DIODE(text_in[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA_320 (.DIODE(text_in[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA_321 (.DIODE(text_in[49]));
 sky130_fd_sc_hd__diode_2 ANTENNA_322 (.DIODE(text_in[63]));
 sky130_fd_sc_hd__diode_2 ANTENNA_323 (.DIODE(text_in[66]));
 sky130_fd_sc_hd__diode_2 ANTENNA_324 (.DIODE(text_in[82]));
 sky130_fd_sc_hd__diode_2 ANTENNA_325 (.DIODE(text_in[88]));
 sky130_fd_sc_hd__diode_2 ANTENNA_326 (.DIODE(text_in[99]));
 sky130_fd_sc_hd__diode_2 ANTENNA_327 (.DIODE(key[112]));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1367 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1397 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_744 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_673 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_828 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_743 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_798 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_740 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_801 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_806 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_830 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_761 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_799 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_774 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_743 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_774 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_782 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_834 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_842 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_670 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_704 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_771 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_773 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_828 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_747 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_810 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_733 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_747 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_824 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_833 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_507 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_822 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_495 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_674 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_801 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_830 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_460 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_492 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_792 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_504 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_698 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_766 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_806 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_486 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_660 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_782 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_804 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_501 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_761 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_812 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_470 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_540 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_588 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_840 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_507 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_520 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_460 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_537 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_654 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_774 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_828 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_567 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_750 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_758 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_792 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_434 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_443 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_495 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_673 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_807 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_683 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_452 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_516 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_747 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_812 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_490 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_773 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_892 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_922 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_330 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_507 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_860 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_983 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_468 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_552 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_768 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_863 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_975 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_452 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_750 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_858 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_890 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_914 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_932 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_940 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_830 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_852 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_906 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_976 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_504 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_514 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_854 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_867 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_950 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_494 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_890 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1008 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1024 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1032 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_854 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_907 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_952 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_852 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_903 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_498 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_650 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_874 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_914 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_919 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_927 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_949 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_979 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_240 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_470 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_492 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_780 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_842 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_860 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_876 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_960 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_978 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_464 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_507 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_884 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_980 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_996 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_602 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_708 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_720 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_837 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_895 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_914 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_683 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_740 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_829 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_852 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_934 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_970 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_702 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_766 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_774 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_782 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_835 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_933 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_942 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_951 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_998 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1006 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1014 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1022 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_327 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_644 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_730 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_858 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_866 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_891 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_933 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_963 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_979 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_708 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_743 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_882 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_934 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_270 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_330 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_733 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_803 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_884 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_910 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_932 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_823 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_842 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_854 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_918 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1020 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_336 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_364 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_733 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_801 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_987 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_730 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_902 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_944 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_980 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_687 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_764 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_854 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_866 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_923 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_774 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_813 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_895 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_962 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_567 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_711 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_761 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_923 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_996 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_702 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_766 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_774 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_782 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_821 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_906 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_919 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_949 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_963 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_492 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_673 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_870 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_882 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_915 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_920 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_936 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_294 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_771 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_863 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_923 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_462 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_524 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_604 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_966 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_580 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_524 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_696 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_708 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_773 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_834 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_919 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_944 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_966 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_980 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_387 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_674 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_938 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_953 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1011 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_413 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_602 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_638 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_674 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_730 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_955 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1024 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1032 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_798 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_924 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_932 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_996 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_614 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_840 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_906 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_938 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_998 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1006 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_650 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_684 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_726 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_734 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_981 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1035 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1043 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_696 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1010 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_912 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1042 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1050 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_353 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_953 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1039 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_865 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_927 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_990 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_422 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_606 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_866 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1028 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1042 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_392 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_548 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_903 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_951 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_984 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1000 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_297 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_490 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_650 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_792 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_923 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1027 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_272 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_803 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_963 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_324 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_726 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_906 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_976 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1014 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1026 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_270 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_644 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_739 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_747 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_850 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_878 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_906 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_915 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1026 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1039 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_254 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_354 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_761 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_916 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_979 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1066 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1074 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1082 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_554 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_684 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_696 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_750 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_762 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_813 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_906 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_963 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1039 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1047 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_240 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_646 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_660 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_897 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1038 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_280 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_694 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_710 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_768 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_831 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_878 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_913 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_966 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_974 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1023 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1050 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_417 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_847 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_902 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_946 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1148 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1185 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_406 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_514 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_588 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_700 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_792 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_884 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_936 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_992 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1091 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1203 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1219 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1224 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_353 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_702 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_862 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_891 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_982 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_995 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1154 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1183 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1195 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_709 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_744 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_950 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_985 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1043 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1151 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1170 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_53 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_362 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_880 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_985 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1039 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1077 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1118 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1147 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1159 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1253 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_134 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_340 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_567 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_606 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_700 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_760 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_800 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_864 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_992 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1113 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1170 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1198 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1219 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1245 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_542 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_662 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_954 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_968 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1013 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1083 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1117 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1144 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1156 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1204 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1212 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_147 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_884 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_942 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1110 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1118 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1143 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1221 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1248 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_891 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_940 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_954 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_966 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1022 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1088 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1125 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1133 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1186 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1210 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_692 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_932 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_987 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1038 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1054 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1062 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1116 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1158 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1184 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1205 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1239 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_182 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_224 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_362 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_473 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_602 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_835 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1075 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1129 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1155 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1253 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1266 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_82 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_567 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_709 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_979 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_987 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1126 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1147 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1185 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1219 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1227 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1235 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1248 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_56 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_660 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_800 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_888 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_904 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_912 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_957 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_980 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1008 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1024 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1032 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1140 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1148 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1162 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1188 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1246 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1254 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1262 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1270 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1278 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1286 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_267 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_280 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_380 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_404 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_583 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_821 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_864 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_872 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_995 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1004 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1090 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1155 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1220 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1233 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1242 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_54 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_180 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_294 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_426 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_660 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_890 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_933 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_942 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_954 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1008 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1024 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1032 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1133 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1144 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1185 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1253 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1266 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_454 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_588 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_867 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_927 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_932 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_976 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_984 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_998 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1116 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1158 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1174 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1238 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1246 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_800 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_964 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1003 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1034 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1042 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1122 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1130 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1192 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1257 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_87 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_464 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_560 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_828 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_876 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_924 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1053 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1115 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1156 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1180 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_458 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_673 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_890 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1073 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1104 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1121 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1206 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1253 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_397 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_684 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1099 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1235 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_120 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_162 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1010 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1024 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1032 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1086 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1129 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1145 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1215 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1245 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1253 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1101 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1161 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1206 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_164 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_998 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1078 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1124 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1200 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1266 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_747 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1174 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1243 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_45 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_840 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_878 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1083 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1094 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1154 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1159 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1188 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1196 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1264 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1272 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_750 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_996 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1010 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1098 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1173 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1148 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1192 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1214 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1235 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1249 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_823 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_921 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_934 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_994 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1120 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1153 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1216 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1264 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1272 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1280 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1296 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1304 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1312 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_51 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_302 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_831 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_890 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_981 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1063 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1092 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1176 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1185 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1195 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1221 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_460 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_583 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_630 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_694 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_866 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1027 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1114 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1120 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1176 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1215 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1230 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_949 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_973 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1039 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_504 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_674 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1146 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_267 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_346 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_730 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_907 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1092 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1163 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1183 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1221 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_406 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_490 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_711 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_818 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_960 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1092 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1125 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1143 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1185 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_435 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_627 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_803 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_927 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1040 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1113 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1206 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1242 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_384 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_420 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_507 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_900 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_922 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1024 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1137 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1143 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1206 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1242 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1250 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1266 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1052 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1104 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1116 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1156 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1225 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1248 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_711 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_773 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_782 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_921 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1077 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1137 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1145 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1202 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1212 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1260 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1268 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_404 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_794 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_998 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1056 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1120 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1223 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_830 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_866 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1071 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1077 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1095 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1125 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1147 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1221 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_336 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_372 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_512 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_870 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1047 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1104 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1133 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1170 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_240 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_730 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_994 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1070 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1082 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1088 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1219 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1246 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1254 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1262 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1270 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1278 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1286 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_152 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_316 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_413 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_732 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_973 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1122 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1219 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1234 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1242 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_52 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_913 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1000 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1080 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1152 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1249 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1257 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_116 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_670 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_844 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_950 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1086 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1116 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1146 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1218 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1227 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1235 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_74 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_422 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_434 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_963 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1069 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1148 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_30 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_387 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_624 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_692 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1053 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1110 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1118 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1130 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1160 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1213 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1230 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_66 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_74 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_673 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1026 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1034 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1042 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1092 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1130 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1146 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1250 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1266 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_34 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_692 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_704 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_973 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1076 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1121 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1134 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1163 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1227 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1073 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1134 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1148 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1160 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1200 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1216 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1245 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1249 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1257 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_400 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_878 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_886 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1163 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1238 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1246 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_366 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_848 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_890 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_945 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1026 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1034 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1042 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1063 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1124 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1144 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1180 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1192 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1250 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1266 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_504 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_976 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_984 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_996 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1060 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1099 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1159 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1167 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1209 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1223 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_33 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_46 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_70 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_540 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_606 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_702 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_904 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_912 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1126 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1140 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1148 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1238 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1246 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1254 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1262 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1270 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1278 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1286 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_386 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_428 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1120 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1162 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1186 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1249 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_594 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_623 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_831 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_914 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1064 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1134 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1140 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1205 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1251 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1267 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1275 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_54 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_762 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_864 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_922 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_934 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_983 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1155 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1220 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1240 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1248 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_140 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_484 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_520 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_886 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_892 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_923 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_940 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_957 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_967 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_981 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1053 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1070 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1126 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1191 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1216 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1260 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1268 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_814 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1056 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1110 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1118 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1130 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1216 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1240 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1248 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_31 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_80 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_290 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_308 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_727 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_842 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_950 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_970 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1071 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_1101 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1138 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1166 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1212 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_30 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_606 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_829 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_847 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_858 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_966 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_976 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1086 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1094 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1112 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1116 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1130 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1230 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1238 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1246 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_722 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_833 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_951 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_960 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1058 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1129 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1137 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1145 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1186 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1219 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_76 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_812 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_847 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_918 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_932 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_938 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_950 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_968 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_976 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_983 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1050 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1099 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1123 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1163 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1206 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1230 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1238 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1246 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_294 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_918 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_983 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1145 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_83 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_640 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_878 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_890 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_983 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1054 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1116 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1210 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1218 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1226 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1234 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1242 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_41 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_49 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_473 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_891 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_916 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1010 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1026 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1034 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1042 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1091 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1099 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1133 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1161 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_32 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_400 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_614 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_821 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_890 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_914 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_936 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_978 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1039 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1056 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1072 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1173 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_122 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_144 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_650 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_698 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_724 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_800 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_904 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_920 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1186 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1202 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1210 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1218 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1226 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_78 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_383 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_760 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_855 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_954 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_996 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1043 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_122 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_304 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_683 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_906 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_960 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_972 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1070 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1086 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_90 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_576 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_747 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_975 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_987 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1185 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_55 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_473 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_490 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_825 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_830 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_846 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_975 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1099 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1209 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_50 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_462 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_886 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_892 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_916 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_923 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_945 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_979 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_987 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1003 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1173 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1191 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1196 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1205 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1218 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1226 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1234 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1242 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_784 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_837 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_888 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_904 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_912 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_980 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1206 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_761 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_825 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_863 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_944 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_975 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_997 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1009 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1052 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1056 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1087 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1101 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1125 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1160 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_813 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_895 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_953 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1060 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1068 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1144 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1200 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1216 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_380 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_750 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_821 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_934 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_948 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_976 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_984 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_992 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1000 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1043 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1102 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1170 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1185 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_460 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_468 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_775 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_837 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_904 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_914 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_950 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_964 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1084 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1129 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1150 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1186 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1200 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1216 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_327 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_458 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_564 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_696 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_876 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_921 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1038 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1056 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1132 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1155 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1164 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1172 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_440 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_600 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_955 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1034 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1135 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_438 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_582 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_624 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_687 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_696 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_932 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_936 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_970 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_984 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_992 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1027 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1091 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1103 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1150 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_458 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_600 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_825 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1070 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1204 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_350 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_383 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_452 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_683 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_807 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_923 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1042 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1170 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_895 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1015 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1140 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1202 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1210 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1218 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1226 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_932 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1042 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1092 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1104 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1163 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1173 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_413 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_593 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_859 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_904 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_964 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1159 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_606 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_829 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1009 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1087 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1100 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1116 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1219 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1227 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1235 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_653 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_668 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_733 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_817 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_891 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_966 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1073 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_294 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_392 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_627 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_636 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_807 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1003 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1088 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1120 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1215 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1223 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_410 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_474 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_490 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_534 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_580 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_903 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_951 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1071 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1087 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1130 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_387 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_993 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1047 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1061 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1098 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1155 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1206 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1230 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1238 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1246 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_360 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_844 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_904 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1120 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1134 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_374 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_630 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_804 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_895 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_936 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1112 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1120 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1122 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1130 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1136 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1145 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1161 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1215 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1223 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_726 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_826 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_902 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1015 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1069 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1137 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1150 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1197 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_376 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_384 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_398 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_555 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_802 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_858 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_921 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_936 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1043 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1056 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1162 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1189 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_893 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_916 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_966 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1015 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1039 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1080 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1173 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1182 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1206 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_496 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_520 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_570 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_630 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_747 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_370 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_410 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_548 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_945 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1066 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1074 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1088 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1190 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1204 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1212 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_604 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_798 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1043 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1053 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1189 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_840 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_862 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_957 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1101 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1166 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_567 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_802 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_848 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_860 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1044 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1095 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1125 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1190 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_468 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_516 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_662 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1015 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1043 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1069 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_563 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_747 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_936 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_484 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_784 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_831 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_904 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_555 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_630 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_823 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_860 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_892 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_923 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_462 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_484 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_583 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_770 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_833 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_798 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_858 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_891 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_921 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_488 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_804 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_815 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_826 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_833 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_904 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_960 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_520 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_636 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_796 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_804 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_858 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_882 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_775 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_464 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_552 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_570 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_848 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_866 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_942 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_433 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_530 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_784 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_801 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_826 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_830 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_948 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_964 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_486 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_860 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_894 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_927 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_606 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_717 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_828 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_844 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_900 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_458 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_743 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_468 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_530 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_642 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_708 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_514 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_673 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_768 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_501 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_593 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_768 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_700 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_711 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_745 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_812 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_533 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_732 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_747 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_804 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_457 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_709 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_777 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_840 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_614 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_864 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_726 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_773 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_820 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_828 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_683 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_714 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_733 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_814 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_501 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_593 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_657 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_743 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_814 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_758 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_777 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_520 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_683 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_734 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_702 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_774 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_842 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_747 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_678 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_726 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_762 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_727 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_768 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_777 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_831 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_815 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_825 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_787 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_690 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_858 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_756 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_764 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_842 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_850 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_743 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_774 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_724 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_792 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_766 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_815 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_681 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_733 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_673 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1421 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1367 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1397 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_1427 ();
endmodule
