module parameterized_ring_counter (clk,
    enable,
    rst_n,
    count);
 input clk;
 input enable;
 input rst_n;
 output [3:0] count;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;

 INV_X1 _14_ (.A(net1),
    .ZN(_04_));
 BUF_X4 _15_ (.A(enable),
    .Z(_05_));
 MUX2_X1 _16_ (.A(net2),
    .B(net5),
    .S(_05_),
    .Z(_06_));
 OR2_X1 _17_ (.A1(_04_),
    .A2(_06_),
    .ZN(_00_));
 MUX2_X1 _18_ (.A(net3),
    .B(net2),
    .S(_05_),
    .Z(_07_));
 AND2_X1 _19_ (.A1(net1),
    .A2(_07_),
    .ZN(_01_));
 MUX2_X1 _20_ (.A(net4),
    .B(net3),
    .S(_05_),
    .Z(_08_));
 AND2_X1 _21_ (.A1(net1),
    .A2(_08_),
    .ZN(_02_));
 MUX2_X1 _22_ (.A(net5),
    .B(net4),
    .S(_05_),
    .Z(_09_));
 AND2_X1 _23_ (.A1(net1),
    .A2(_09_),
    .ZN(_03_));
 DFF_X1 \counter_reg[0]$_SDFFE_PN1P_  (.D(_00_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net2),
    .QN(_13_));
 DFF_X1 \counter_reg[1]$_SDFFE_PN0P_  (.D(_01_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net3),
    .QN(_12_));
 DFF_X1 \counter_reg[2]$_SDFFE_PN0P_  (.D(_02_),
    .CK(clknet_1_0__leaf_clk),
    .Q(net4),
    .QN(_11_));
 DFF_X1 \counter_reg[3]$_SDFFE_PN0P_  (.D(_03_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net5),
    .QN(_10_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_45 ();
 BUF_X1 input1 (.A(rst_n),
    .Z(net1));
 BUF_X1 output2 (.A(net2),
    .Z(count[0]));
 BUF_X1 output3 (.A(net3),
    .Z(count[1]));
 BUF_X1 output4 (.A(net4),
    .Z(count[2]));
 BUF_X1 output5 (.A(net5),
    .Z(count[3]));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X8 FILLER_0_161 ();
 FILLCELL_X2 FILLER_0_169 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X8 FILLER_1_161 ();
 FILLCELL_X2 FILLER_1_169 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X8 FILLER_2_161 ();
 FILLCELL_X2 FILLER_2_169 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X8 FILLER_3_161 ();
 FILLCELL_X2 FILLER_3_169 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X8 FILLER_4_161 ();
 FILLCELL_X2 FILLER_4_169 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X8 FILLER_5_161 ();
 FILLCELL_X2 FILLER_5_169 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X8 FILLER_6_161 ();
 FILLCELL_X2 FILLER_6_169 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X8 FILLER_7_161 ();
 FILLCELL_X2 FILLER_7_169 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X8 FILLER_8_161 ();
 FILLCELL_X2 FILLER_8_169 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X8 FILLER_9_161 ();
 FILLCELL_X2 FILLER_9_169 ();
 FILLCELL_X1 FILLER_10_30 ();
 FILLCELL_X1 FILLER_10_38 ();
 FILLCELL_X2 FILLER_10_43 ();
 FILLCELL_X32 FILLER_10_62 ();
 FILLCELL_X32 FILLER_10_94 ();
 FILLCELL_X32 FILLER_10_126 ();
 FILLCELL_X8 FILLER_10_158 ();
 FILLCELL_X4 FILLER_10_166 ();
 FILLCELL_X1 FILLER_10_170 ();
 FILLCELL_X1 FILLER_11_4 ();
 FILLCELL_X1 FILLER_11_29 ();
 FILLCELL_X1 FILLER_11_44 ();
 FILLCELL_X8 FILLER_11_62 ();
 FILLCELL_X4 FILLER_11_70 ();
 FILLCELL_X32 FILLER_11_79 ();
 FILLCELL_X32 FILLER_11_111 ();
 FILLCELL_X4 FILLER_11_143 ();
 FILLCELL_X1 FILLER_11_147 ();
 FILLCELL_X2 FILLER_11_151 ();
 FILLCELL_X8 FILLER_11_156 ();
 FILLCELL_X4 FILLER_11_164 ();
 FILLCELL_X2 FILLER_11_168 ();
 FILLCELL_X1 FILLER_11_170 ();
 FILLCELL_X8 FILLER_12_11 ();
 FILLCELL_X4 FILLER_12_19 ();
 FILLCELL_X8 FILLER_12_34 ();
 FILLCELL_X1 FILLER_12_42 ();
 FILLCELL_X32 FILLER_12_47 ();
 FILLCELL_X32 FILLER_12_79 ();
 FILLCELL_X32 FILLER_12_111 ();
 FILLCELL_X16 FILLER_12_143 ();
 FILLCELL_X8 FILLER_12_159 ();
 FILLCELL_X4 FILLER_12_167 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X32 FILLER_13_129 ();
 FILLCELL_X8 FILLER_13_161 ();
 FILLCELL_X2 FILLER_13_169 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X32 FILLER_14_129 ();
 FILLCELL_X8 FILLER_14_161 ();
 FILLCELL_X2 FILLER_14_169 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X8 FILLER_15_161 ();
 FILLCELL_X2 FILLER_15_169 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X32 FILLER_16_129 ();
 FILLCELL_X8 FILLER_16_161 ();
 FILLCELL_X2 FILLER_16_169 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X32 FILLER_17_129 ();
 FILLCELL_X8 FILLER_17_161 ();
 FILLCELL_X2 FILLER_17_169 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X8 FILLER_18_161 ();
 FILLCELL_X2 FILLER_18_169 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X8 FILLER_19_161 ();
 FILLCELL_X2 FILLER_19_169 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X8 FILLER_20_161 ();
 FILLCELL_X2 FILLER_20_169 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X8 FILLER_21_161 ();
 FILLCELL_X2 FILLER_21_169 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X8 FILLER_22_161 ();
 FILLCELL_X2 FILLER_22_169 ();
endmodule
