module parameterized_serdes (clk,
    enable,
    load,
    mode,
    rst_n,
    rx_done,
    serial_in,
    serial_out,
    tx_done,
    parallel_in,
    parallel_out);
 input clk;
 input enable;
 input load;
 input mode;
 input rst_n;
 output rx_done;
 input serial_in;
 output serial_out;
 output tx_done;
 input [7:0] parallel_in;
 output [7:0] parallel_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire \rx_bit_counter[0] ;
 wire \rx_bit_counter[1] ;
 wire \rx_bit_counter[2] ;
 wire \rx_bit_counter[3] ;
 wire \rx_shift_reg[0] ;
 wire \rx_shift_reg[1] ;
 wire \rx_shift_reg[2] ;
 wire \rx_shift_reg[3] ;
 wire \rx_shift_reg[4] ;
 wire \rx_shift_reg[5] ;
 wire \rx_shift_reg[6] ;
 wire \tx_bit_counter[0] ;
 wire \tx_bit_counter[1] ;
 wire \tx_bit_counter[2] ;
 wire \tx_bit_counter[3] ;
 wire \tx_shift_reg[0] ;
 wire \tx_shift_reg[1] ;
 wire \tx_shift_reg[2] ;
 wire \tx_shift_reg[3] ;
 wire \tx_shift_reg[4] ;
 wire \tx_shift_reg[5] ;
 wire \tx_shift_reg[6] ;
 wire \tx_shift_reg[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;

 CLKBUF_X2 _167_ (.A(rst_n),
    .Z(_122_));
 BUF_X2 _168_ (.A(_122_),
    .Z(_123_));
 BUF_X2 _169_ (.A(_123_),
    .Z(_124_));
 BUF_X2 _170_ (.A(net19),
    .Z(_125_));
 BUF_X4 _171_ (.A(load),
    .Z(_126_));
 BUF_X4 _172_ (.A(_163_),
    .Z(_127_));
 AOI21_X4 _173_ (.A(\rx_bit_counter[3] ),
    .B1(\rx_bit_counter[2] ),
    .B2(_127_),
    .ZN(_128_));
 BUF_X4 _174_ (.A(enable),
    .Z(_129_));
 NAND2_X2 _175_ (.A1(_129_),
    .A2(net1),
    .ZN(_130_));
 NOR4_X4 _176_ (.A1(_125_),
    .A2(_126_),
    .A3(_128_),
    .A4(_130_),
    .ZN(_131_));
 MUX2_X1 _177_ (.A(net16),
    .B(\rx_shift_reg[4] ),
    .S(_131_),
    .Z(_132_));
 AND2_X1 _178_ (.A1(_124_),
    .A2(_132_),
    .ZN(_003_));
 MUX2_X1 _179_ (.A(net17),
    .B(\rx_shift_reg[5] ),
    .S(_131_),
    .Z(_036_));
 AND2_X1 _180_ (.A1(_124_),
    .A2(_036_),
    .ZN(_004_));
 MUX2_X1 _181_ (.A(net18),
    .B(\rx_shift_reg[6] ),
    .S(_131_),
    .Z(_037_));
 AND2_X1 _182_ (.A1(_124_),
    .A2(_037_),
    .ZN(_005_));
 INV_X2 _183_ (.A(_123_),
    .ZN(_038_));
 INV_X1 _184_ (.A(\rx_bit_counter[0] ),
    .ZN(_039_));
 NAND2_X1 _185_ (.A1(\rx_bit_counter[2] ),
    .A2(_127_),
    .ZN(_040_));
 INV_X2 _186_ (.A(_126_),
    .ZN(_041_));
 AOI21_X4 _187_ (.A(_130_),
    .B1(_041_),
    .B2(_125_),
    .ZN(_042_));
 NOR2_X2 _188_ (.A1(_126_),
    .A2(\rx_bit_counter[3] ),
    .ZN(_043_));
 NAND4_X1 _189_ (.A1(_039_),
    .A2(_040_),
    .A3(_042_),
    .A4(_043_),
    .ZN(_044_));
 AND2_X1 _190_ (.A1(_129_),
    .A2(net1),
    .ZN(_045_));
 INV_X1 _191_ (.A(_125_),
    .ZN(_046_));
 OAI21_X2 _192_ (.A(_045_),
    .B1(_126_),
    .B2(_046_),
    .ZN(_047_));
 NAND2_X1 _193_ (.A1(\rx_bit_counter[0] ),
    .A2(_047_),
    .ZN(_048_));
 AOI21_X1 _194_ (.A(_038_),
    .B1(_044_),
    .B2(_048_),
    .ZN(_006_));
 NAND2_X1 _195_ (.A1(\rx_bit_counter[1] ),
    .A2(_047_),
    .ZN(_049_));
 NAND4_X1 _196_ (.A1(_164_),
    .A2(_040_),
    .A3(_042_),
    .A4(_043_),
    .ZN(_050_));
 AOI21_X1 _197_ (.A(_038_),
    .B1(_049_),
    .B2(_050_),
    .ZN(_007_));
 NOR3_X1 _198_ (.A1(_126_),
    .A2(\rx_bit_counter[3] ),
    .A3(_127_),
    .ZN(_051_));
 OAI21_X1 _199_ (.A(\rx_bit_counter[2] ),
    .B1(_047_),
    .B2(_051_),
    .ZN(_052_));
 INV_X1 _200_ (.A(\rx_bit_counter[2] ),
    .ZN(_053_));
 NAND4_X1 _201_ (.A1(_053_),
    .A2(_127_),
    .A3(_042_),
    .A4(_043_),
    .ZN(_054_));
 AOI21_X1 _202_ (.A(_038_),
    .B1(_052_),
    .B2(_054_),
    .ZN(_008_));
 NAND3_X1 _203_ (.A1(\rx_bit_counter[0] ),
    .A2(\rx_bit_counter[1] ),
    .A3(_043_),
    .ZN(_055_));
 OR4_X1 _204_ (.A1(_053_),
    .A2(_127_),
    .A3(_047_),
    .A4(_055_),
    .ZN(_056_));
 NAND2_X1 _205_ (.A1(\rx_bit_counter[3] ),
    .A2(_047_),
    .ZN(_057_));
 AOI21_X1 _206_ (.A(_038_),
    .B1(_056_),
    .B2(_057_),
    .ZN(_009_));
 NAND2_X1 _207_ (.A1(_125_),
    .A2(_130_),
    .ZN(_058_));
 AOI21_X1 _208_ (.A(_126_),
    .B1(_002_),
    .B2(_128_),
    .ZN(_059_));
 NAND2_X1 _209_ (.A1(_045_),
    .A2(_059_),
    .ZN(_060_));
 AOI21_X1 _210_ (.A(_038_),
    .B1(_058_),
    .B2(_060_),
    .ZN(_010_));
 AND3_X1 _211_ (.A1(_041_),
    .A2(net10),
    .A3(_122_),
    .ZN(_061_));
 AND2_X1 _212_ (.A1(\rx_shift_reg[0] ),
    .A2(_123_),
    .ZN(_062_));
 NAND2_X1 _213_ (.A1(_041_),
    .A2(_002_),
    .ZN(_063_));
 OAI21_X4 _214_ (.A(_042_),
    .B1(_063_),
    .B2(_128_),
    .ZN(_064_));
 MUX2_X1 _215_ (.A(_061_),
    .B(_062_),
    .S(_064_),
    .Z(_011_));
 AND3_X1 _216_ (.A1(_041_),
    .A2(\rx_shift_reg[0] ),
    .A3(_122_),
    .ZN(_065_));
 AND2_X1 _217_ (.A1(\rx_shift_reg[1] ),
    .A2(_123_),
    .ZN(_066_));
 MUX2_X1 _218_ (.A(_065_),
    .B(_066_),
    .S(_064_),
    .Z(_012_));
 AND3_X1 _219_ (.A1(_041_),
    .A2(\rx_shift_reg[1] ),
    .A3(_122_),
    .ZN(_067_));
 AND2_X1 _220_ (.A1(\rx_shift_reg[2] ),
    .A2(_123_),
    .ZN(_068_));
 MUX2_X1 _221_ (.A(_067_),
    .B(_068_),
    .S(_064_),
    .Z(_013_));
 AND3_X1 _222_ (.A1(_041_),
    .A2(\rx_shift_reg[2] ),
    .A3(_122_),
    .ZN(_069_));
 AND2_X1 _223_ (.A1(\rx_shift_reg[3] ),
    .A2(_123_),
    .ZN(_070_));
 MUX2_X1 _224_ (.A(_069_),
    .B(_070_),
    .S(_064_),
    .Z(_014_));
 AND3_X1 _225_ (.A1(_041_),
    .A2(\rx_shift_reg[3] ),
    .A3(_122_),
    .ZN(_071_));
 AND2_X1 _226_ (.A1(\rx_shift_reg[4] ),
    .A2(_123_),
    .ZN(_072_));
 MUX2_X1 _227_ (.A(_071_),
    .B(_072_),
    .S(_064_),
    .Z(_015_));
 AND3_X1 _228_ (.A1(_041_),
    .A2(\rx_shift_reg[4] ),
    .A3(_122_),
    .ZN(_073_));
 AND2_X1 _229_ (.A1(\rx_shift_reg[5] ),
    .A2(_123_),
    .ZN(_074_));
 MUX2_X1 _230_ (.A(_073_),
    .B(_074_),
    .S(_064_),
    .Z(_016_));
 AND3_X1 _231_ (.A1(_041_),
    .A2(\rx_shift_reg[5] ),
    .A3(_122_),
    .ZN(_075_));
 AND2_X1 _232_ (.A1(\rx_shift_reg[6] ),
    .A2(_123_),
    .ZN(_076_));
 MUX2_X1 _233_ (.A(_075_),
    .B(_076_),
    .S(_064_),
    .Z(_017_));
 INV_X1 _234_ (.A(net1),
    .ZN(_077_));
 INV_X1 _235_ (.A(net21),
    .ZN(_078_));
 CLKBUF_X2 _236_ (.A(\tx_bit_counter[2] ),
    .Z(_079_));
 AOI211_X2 _237_ (.A(_126_),
    .B(\tx_bit_counter[3] ),
    .C1(_079_),
    .C2(_165_),
    .ZN(_080_));
 AND4_X1 _238_ (.A1(_129_),
    .A2(_077_),
    .A3(_078_),
    .A4(_080_),
    .ZN(_081_));
 OAI211_X2 _239_ (.A(_129_),
    .B(_077_),
    .C1(_126_),
    .C2(_078_),
    .ZN(_082_));
 BUF_X1 _240_ (.A(\tx_bit_counter[0] ),
    .Z(_083_));
 MUX2_X1 _241_ (.A(_081_),
    .B(_082_),
    .S(_083_),
    .Z(_084_));
 AND2_X1 _242_ (.A1(_124_),
    .A2(_084_),
    .ZN(_018_));
 BUF_X2 _243_ (.A(\tx_bit_counter[1] ),
    .Z(_085_));
 AOI22_X1 _244_ (.A1(_085_),
    .A2(_082_),
    .B1(_081_),
    .B2(_166_),
    .ZN(_086_));
 NOR2_X1 _245_ (.A1(_038_),
    .A2(_086_),
    .ZN(_019_));
 NAND2_X1 _246_ (.A1(_079_),
    .A2(_082_),
    .ZN(_087_));
 XNOR2_X1 _247_ (.A(_165_),
    .B(_000_),
    .ZN(_088_));
 NAND2_X1 _248_ (.A1(_080_),
    .A2(_088_),
    .ZN(_089_));
 OR2_X1 _249_ (.A1(_082_),
    .A2(_089_),
    .ZN(_090_));
 AOI21_X1 _250_ (.A(_038_),
    .B1(_087_),
    .B2(_090_),
    .ZN(_020_));
 BUF_X2 _251_ (.A(_123_),
    .Z(_091_));
 NAND3_X1 _252_ (.A1(_079_),
    .A2(_083_),
    .A3(_085_),
    .ZN(_092_));
 XOR2_X1 _253_ (.A(_001_),
    .B(_092_),
    .Z(_093_));
 NAND3_X1 _254_ (.A1(_091_),
    .A2(_081_),
    .A3(_093_),
    .ZN(_094_));
 NAND3_X1 _255_ (.A1(\tx_bit_counter[3] ),
    .A2(_091_),
    .A3(_082_),
    .ZN(_095_));
 NAND2_X1 _256_ (.A1(_094_),
    .A2(_095_),
    .ZN(_021_));
 NAND3_X4 _257_ (.A1(_129_),
    .A2(_077_),
    .A3(_126_),
    .ZN(_096_));
 NAND2_X1 _258_ (.A1(_091_),
    .A2(_096_),
    .ZN(_097_));
 INV_X1 _259_ (.A(_129_),
    .ZN(_098_));
 AOI21_X1 _260_ (.A(\tx_bit_counter[3] ),
    .B1(_079_),
    .B2(_165_),
    .ZN(_099_));
 OR3_X1 _261_ (.A1(_098_),
    .A2(net1),
    .A3(_099_),
    .ZN(_100_));
 AOI21_X1 _262_ (.A(_097_),
    .B1(_100_),
    .B2(_078_),
    .ZN(_022_));
 MUX2_X1 _263_ (.A(net2),
    .B(\tx_shift_reg[0] ),
    .S(_096_),
    .Z(_101_));
 AND2_X1 _264_ (.A1(_124_),
    .A2(_101_),
    .ZN(_023_));
 MUX2_X1 _265_ (.A(net3),
    .B(\tx_shift_reg[1] ),
    .S(_096_),
    .Z(_102_));
 AND2_X1 _266_ (.A1(_124_),
    .A2(_102_),
    .ZN(_024_));
 MUX2_X1 _267_ (.A(net4),
    .B(\tx_shift_reg[2] ),
    .S(_096_),
    .Z(_103_));
 AND2_X1 _268_ (.A1(_124_),
    .A2(_103_),
    .ZN(_025_));
 MUX2_X1 _269_ (.A(net5),
    .B(\tx_shift_reg[3] ),
    .S(_096_),
    .Z(_104_));
 AND2_X1 _270_ (.A1(_124_),
    .A2(_104_),
    .ZN(_026_));
 MUX2_X1 _271_ (.A(net6),
    .B(\tx_shift_reg[4] ),
    .S(_096_),
    .Z(_105_));
 AND2_X1 _272_ (.A1(_124_),
    .A2(_105_),
    .ZN(_027_));
 MUX2_X1 _273_ (.A(net7),
    .B(\tx_shift_reg[5] ),
    .S(_096_),
    .Z(_106_));
 AND2_X1 _274_ (.A1(_124_),
    .A2(_106_),
    .ZN(_028_));
 MUX2_X1 _275_ (.A(net8),
    .B(\tx_shift_reg[6] ),
    .S(_096_),
    .Z(_107_));
 AND2_X1 _276_ (.A1(_091_),
    .A2(_107_),
    .ZN(_029_));
 MUX2_X1 _277_ (.A(net9),
    .B(\tx_shift_reg[7] ),
    .S(_096_),
    .Z(_108_));
 AND2_X1 _278_ (.A1(_091_),
    .A2(_108_),
    .ZN(_030_));
 MUX2_X1 _279_ (.A(net11),
    .B(net10),
    .S(_131_),
    .Z(_109_));
 AND2_X1 _280_ (.A1(_091_),
    .A2(_109_),
    .ZN(_031_));
 MUX2_X1 _281_ (.A(net12),
    .B(\rx_shift_reg[0] ),
    .S(_131_),
    .Z(_110_));
 AND2_X1 _282_ (.A1(_091_),
    .A2(_110_),
    .ZN(_032_));
 MUX2_X1 _283_ (.A(net13),
    .B(\rx_shift_reg[1] ),
    .S(_131_),
    .Z(_111_));
 AND2_X1 _284_ (.A1(_091_),
    .A2(_111_),
    .ZN(_033_));
 MUX2_X1 _285_ (.A(net14),
    .B(\rx_shift_reg[2] ),
    .S(_131_),
    .Z(_112_));
 AND2_X1 _286_ (.A1(_091_),
    .A2(_112_),
    .ZN(_034_));
 MUX2_X1 _287_ (.A(net15),
    .B(\rx_shift_reg[3] ),
    .S(_131_),
    .Z(_113_));
 AND2_X1 _288_ (.A1(_091_),
    .A2(_113_),
    .ZN(_035_));
 INV_X1 _289_ (.A(\tx_bit_counter[3] ),
    .ZN(_114_));
 MUX2_X1 _290_ (.A(\tx_shift_reg[7] ),
    .B(\tx_shift_reg[5] ),
    .S(_085_),
    .Z(_115_));
 MUX2_X1 _291_ (.A(\tx_shift_reg[6] ),
    .B(\tx_shift_reg[4] ),
    .S(_085_),
    .Z(_116_));
 MUX2_X1 _292_ (.A(_115_),
    .B(_116_),
    .S(_083_),
    .Z(_117_));
 MUX2_X1 _293_ (.A(\tx_shift_reg[3] ),
    .B(\tx_shift_reg[1] ),
    .S(_085_),
    .Z(_118_));
 MUX2_X1 _294_ (.A(\tx_shift_reg[2] ),
    .B(\tx_shift_reg[0] ),
    .S(_085_),
    .Z(_119_));
 MUX2_X1 _295_ (.A(_118_),
    .B(_119_),
    .S(_083_),
    .Z(_120_));
 MUX2_X1 _296_ (.A(_117_),
    .B(_120_),
    .S(_079_),
    .Z(_121_));
 AND3_X1 _297_ (.A1(_114_),
    .A2(_001_),
    .A3(_121_),
    .ZN(net20));
 HA_X1 _298_ (.A(\rx_bit_counter[0] ),
    .B(\rx_bit_counter[1] ),
    .CO(_163_),
    .S(_164_));
 HA_X1 _299_ (.A(\tx_bit_counter[0] ),
    .B(\tx_bit_counter[1] ),
    .CO(_165_),
    .S(_166_));
 DFF_X1 \parallel_out[0]$_SDFFE_PN0P_  (.D(_031_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net11),
    .QN(_162_));
 DFF_X1 \parallel_out[1]$_SDFFE_PN0P_  (.D(_032_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net12),
    .QN(_161_));
 DFF_X1 \parallel_out[2]$_SDFFE_PN0P_  (.D(_033_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net13),
    .QN(_160_));
 DFF_X1 \parallel_out[3]$_SDFFE_PN0P_  (.D(_034_),
    .CK(clknet_2_0__leaf_clk),
    .Q(net14),
    .QN(_159_));
 DFF_X1 \parallel_out[4]$_SDFFE_PN0P_  (.D(_035_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net15),
    .QN(_158_));
 DFF_X1 \parallel_out[5]$_SDFFE_PN0P_  (.D(_003_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net16),
    .QN(_157_));
 DFF_X1 \parallel_out[6]$_SDFFE_PN0P_  (.D(_004_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net17),
    .QN(_156_));
 DFF_X1 \parallel_out[7]$_SDFFE_PN0P_  (.D(_005_),
    .CK(clknet_2_2__leaf_clk),
    .Q(net18),
    .QN(_155_));
 DFF_X1 \rx_bit_counter[0]$_SDFFE_PN0P_  (.D(_006_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\rx_bit_counter[0] ),
    .QN(_154_));
 DFF_X1 \rx_bit_counter[1]$_SDFFE_PN0P_  (.D(_007_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\rx_bit_counter[1] ),
    .QN(_153_));
 DFF_X2 \rx_bit_counter[2]$_SDFFE_PN0P_  (.D(_008_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\rx_bit_counter[2] ),
    .QN(_152_));
 DFF_X2 \rx_bit_counter[3]$_SDFFE_PN0P_  (.D(_009_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\rx_bit_counter[3] ),
    .QN(_151_));
 DFF_X1 \rx_done$_SDFFE_PN0P_  (.D(_010_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net19),
    .QN(_002_));
 DFF_X1 \rx_shift_reg[0]$_SDFFE_PN0P_  (.D(_011_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\rx_shift_reg[0] ),
    .QN(_150_));
 DFF_X1 \rx_shift_reg[1]$_SDFFE_PN0P_  (.D(_012_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\rx_shift_reg[1] ),
    .QN(_149_));
 DFF_X1 \rx_shift_reg[2]$_SDFFE_PN0P_  (.D(_013_),
    .CK(clknet_2_0__leaf_clk),
    .Q(\rx_shift_reg[2] ),
    .QN(_148_));
 DFF_X1 \rx_shift_reg[3]$_SDFFE_PN0P_  (.D(_014_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\rx_shift_reg[3] ),
    .QN(_147_));
 DFF_X1 \rx_shift_reg[4]$_SDFFE_PN0P_  (.D(_015_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\rx_shift_reg[4] ),
    .QN(_146_));
 DFF_X1 \rx_shift_reg[5]$_SDFFE_PN0P_  (.D(_016_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\rx_shift_reg[5] ),
    .QN(_145_));
 DFF_X1 \rx_shift_reg[6]$_SDFFE_PN0P_  (.D(_017_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\rx_shift_reg[6] ),
    .QN(_144_));
 DFF_X1 \tx_bit_counter[0]$_SDFFE_PN0P_  (.D(_018_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\tx_bit_counter[0] ),
    .QN(_143_));
 DFF_X1 \tx_bit_counter[1]$_SDFFE_PN0P_  (.D(_019_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\tx_bit_counter[1] ),
    .QN(_142_));
 DFF_X1 \tx_bit_counter[2]$_SDFFE_PN0P_  (.D(_020_),
    .CK(clknet_2_1__leaf_clk),
    .Q(\tx_bit_counter[2] ),
    .QN(_000_));
 DFF_X2 \tx_bit_counter[3]$_SDFFE_PN0P_  (.D(_021_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\tx_bit_counter[3] ),
    .QN(_001_));
 DFF_X1 \tx_done_reg$_SDFFE_PN0P_  (.D(_022_),
    .CK(clknet_2_1__leaf_clk),
    .Q(net21),
    .QN(_141_));
 DFF_X1 \tx_shift_reg[0]$_SDFFE_PN0P_  (.D(_023_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\tx_shift_reg[0] ),
    .QN(_140_));
 DFF_X1 \tx_shift_reg[1]$_SDFFE_PN0P_  (.D(_024_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\tx_shift_reg[1] ),
    .QN(_139_));
 DFF_X1 \tx_shift_reg[2]$_SDFFE_PN0P_  (.D(_025_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\tx_shift_reg[2] ),
    .QN(_138_));
 DFF_X1 \tx_shift_reg[3]$_SDFFE_PN0P_  (.D(_026_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\tx_shift_reg[3] ),
    .QN(_137_));
 DFF_X1 \tx_shift_reg[4]$_SDFFE_PN0P_  (.D(_027_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\tx_shift_reg[4] ),
    .QN(_136_));
 DFF_X1 \tx_shift_reg[5]$_SDFFE_PN0P_  (.D(_028_),
    .CK(clknet_2_2__leaf_clk),
    .Q(\tx_shift_reg[5] ),
    .QN(_135_));
 DFF_X1 \tx_shift_reg[6]$_SDFFE_PN0P_  (.D(_029_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\tx_shift_reg[6] ),
    .QN(_134_));
 DFF_X1 \tx_shift_reg[7]$_SDFFE_PN0P_  (.D(_030_),
    .CK(clknet_2_3__leaf_clk),
    .Q(\tx_shift_reg[7] ),
    .QN(_133_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_49 ();
 BUF_X1 input1 (.A(mode),
    .Z(net1));
 BUF_X1 input2 (.A(parallel_in[0]),
    .Z(net2));
 BUF_X1 input3 (.A(parallel_in[1]),
    .Z(net3));
 BUF_X1 input4 (.A(parallel_in[2]),
    .Z(net4));
 BUF_X1 input5 (.A(parallel_in[3]),
    .Z(net5));
 BUF_X1 input6 (.A(parallel_in[4]),
    .Z(net6));
 BUF_X1 input7 (.A(parallel_in[5]),
    .Z(net7));
 BUF_X1 input8 (.A(parallel_in[6]),
    .Z(net8));
 BUF_X1 input9 (.A(parallel_in[7]),
    .Z(net9));
 BUF_X1 input10 (.A(serial_in),
    .Z(net10));
 BUF_X1 output11 (.A(net11),
    .Z(parallel_out[0]));
 BUF_X1 output12 (.A(net12),
    .Z(parallel_out[1]));
 BUF_X1 output13 (.A(net13),
    .Z(parallel_out[2]));
 BUF_X1 output14 (.A(net14),
    .Z(parallel_out[3]));
 BUF_X1 output15 (.A(net15),
    .Z(parallel_out[4]));
 BUF_X1 output16 (.A(net16),
    .Z(parallel_out[5]));
 BUF_X1 output17 (.A(net17),
    .Z(parallel_out[6]));
 BUF_X1 output18 (.A(net18),
    .Z(parallel_out[7]));
 BUF_X1 output19 (.A(net19),
    .Z(rx_done));
 BUF_X1 output20 (.A(net20),
    .Z(serial_out));
 BUF_X1 output21 (.A(net21),
    .Z(tx_done));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_0__leaf_clk));
 CLKBUF_X3 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_1__leaf_clk));
 CLKBUF_X3 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_2__leaf_clk));
 CLKBUF_X3 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_2_3__leaf_clk));
 INV_X2 clkload0 (.A(clknet_2_0__leaf_clk));
 INV_X2 clkload1 (.A(clknet_2_1__leaf_clk));
 CLKBUF_X1 clkload2 (.A(clknet_2_2__leaf_clk));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X16 FILLER_0_33 ();
 FILLCELL_X8 FILLER_0_49 ();
 FILLCELL_X2 FILLER_0_57 ();
 FILLCELL_X4 FILLER_0_68 ();
 FILLCELL_X2 FILLER_0_72 ();
 FILLCELL_X1 FILLER_0_74 ();
 FILLCELL_X16 FILLER_0_78 ();
 FILLCELL_X4 FILLER_0_94 ();
 FILLCELL_X1 FILLER_0_101 ();
 FILLCELL_X16 FILLER_0_105 ();
 FILLCELL_X8 FILLER_0_121 ();
 FILLCELL_X4 FILLER_0_129 ();
 FILLCELL_X4 FILLER_0_136 ();
 FILLCELL_X2 FILLER_0_140 ();
 FILLCELL_X32 FILLER_0_145 ();
 FILLCELL_X8 FILLER_0_177 ();
 FILLCELL_X4 FILLER_0_185 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X8 FILLER_1_33 ();
 FILLCELL_X2 FILLER_1_41 ();
 FILLCELL_X16 FILLER_1_101 ();
 FILLCELL_X8 FILLER_1_117 ();
 FILLCELL_X16 FILLER_1_166 ();
 FILLCELL_X4 FILLER_1_182 ();
 FILLCELL_X2 FILLER_1_186 ();
 FILLCELL_X1 FILLER_1_188 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X8 FILLER_2_33 ();
 FILLCELL_X2 FILLER_2_41 ();
 FILLCELL_X1 FILLER_2_43 ();
 FILLCELL_X2 FILLER_2_61 ();
 FILLCELL_X4 FILLER_2_67 ();
 FILLCELL_X2 FILLER_2_71 ();
 FILLCELL_X16 FILLER_2_112 ();
 FILLCELL_X4 FILLER_2_128 ();
 FILLCELL_X1 FILLER_2_132 ();
 FILLCELL_X4 FILLER_2_137 ();
 FILLCELL_X1 FILLER_2_141 ();
 FILLCELL_X32 FILLER_2_153 ();
 FILLCELL_X4 FILLER_2_185 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X16 FILLER_3_33 ();
 FILLCELL_X8 FILLER_3_49 ();
 FILLCELL_X16 FILLER_3_68 ();
 FILLCELL_X8 FILLER_3_84 ();
 FILLCELL_X2 FILLER_3_96 ();
 FILLCELL_X1 FILLER_3_102 ();
 FILLCELL_X8 FILLER_3_110 ();
 FILLCELL_X2 FILLER_3_122 ();
 FILLCELL_X1 FILLER_3_124 ();
 FILLCELL_X32 FILLER_3_142 ();
 FILLCELL_X8 FILLER_3_174 ();
 FILLCELL_X4 FILLER_3_182 ();
 FILLCELL_X2 FILLER_3_186 ();
 FILLCELL_X1 FILLER_3_188 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X4 FILLER_4_65 ();
 FILLCELL_X16 FILLER_4_81 ();
 FILLCELL_X8 FILLER_4_97 ();
 FILLCELL_X4 FILLER_4_105 ();
 FILLCELL_X2 FILLER_4_109 ();
 FILLCELL_X1 FILLER_4_111 ();
 FILLCELL_X32 FILLER_4_138 ();
 FILLCELL_X16 FILLER_4_170 ();
 FILLCELL_X2 FILLER_4_186 ();
 FILLCELL_X1 FILLER_4_188 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X16 FILLER_5_33 ();
 FILLCELL_X4 FILLER_5_49 ();
 FILLCELL_X1 FILLER_5_53 ();
 FILLCELL_X16 FILLER_5_87 ();
 FILLCELL_X8 FILLER_5_103 ();
 FILLCELL_X2 FILLER_5_111 ();
 FILLCELL_X32 FILLER_5_132 ();
 FILLCELL_X16 FILLER_5_164 ();
 FILLCELL_X8 FILLER_5_180 ();
 FILLCELL_X1 FILLER_5_188 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X16 FILLER_6_33 ();
 FILLCELL_X8 FILLER_6_49 ();
 FILLCELL_X4 FILLER_6_57 ();
 FILLCELL_X2 FILLER_6_61 ();
 FILLCELL_X1 FILLER_6_63 ();
 FILLCELL_X8 FILLER_6_85 ();
 FILLCELL_X4 FILLER_6_93 ();
 FILLCELL_X1 FILLER_6_97 ();
 FILLCELL_X8 FILLER_6_103 ();
 FILLCELL_X2 FILLER_6_111 ();
 FILLCELL_X4 FILLER_6_118 ();
 FILLCELL_X2 FILLER_6_122 ();
 FILLCELL_X2 FILLER_6_128 ();
 FILLCELL_X4 FILLER_6_154 ();
 FILLCELL_X2 FILLER_6_158 ();
 FILLCELL_X8 FILLER_6_181 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X1 FILLER_7_65 ();
 FILLCELL_X2 FILLER_7_83 ();
 FILLCELL_X4 FILLER_7_96 ();
 FILLCELL_X1 FILLER_7_100 ();
 FILLCELL_X8 FILLER_7_108 ();
 FILLCELL_X4 FILLER_7_116 ();
 FILLCELL_X2 FILLER_7_120 ();
 FILLCELL_X4 FILLER_7_129 ();
 FILLCELL_X2 FILLER_7_133 ();
 FILLCELL_X1 FILLER_7_135 ();
 FILLCELL_X32 FILLER_7_144 ();
 FILLCELL_X8 FILLER_7_176 ();
 FILLCELL_X4 FILLER_7_184 ();
 FILLCELL_X1 FILLER_7_188 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X4 FILLER_8_33 ();
 FILLCELL_X2 FILLER_8_37 ();
 FILLCELL_X1 FILLER_8_39 ();
 FILLCELL_X4 FILLER_8_44 ();
 FILLCELL_X1 FILLER_8_48 ();
 FILLCELL_X4 FILLER_8_67 ();
 FILLCELL_X1 FILLER_8_71 ();
 FILLCELL_X8 FILLER_8_75 ();
 FILLCELL_X1 FILLER_8_117 ();
 FILLCELL_X32 FILLER_8_122 ();
 FILLCELL_X16 FILLER_8_154 ();
 FILLCELL_X8 FILLER_8_170 ();
 FILLCELL_X2 FILLER_8_178 ();
 FILLCELL_X4 FILLER_8_183 ();
 FILLCELL_X2 FILLER_8_187 ();
 FILLCELL_X16 FILLER_9_1 ();
 FILLCELL_X8 FILLER_9_17 ();
 FILLCELL_X2 FILLER_9_42 ();
 FILLCELL_X1 FILLER_9_44 ();
 FILLCELL_X2 FILLER_9_58 ();
 FILLCELL_X32 FILLER_9_63 ();
 FILLCELL_X2 FILLER_9_95 ();
 FILLCELL_X1 FILLER_9_97 ();
 FILLCELL_X16 FILLER_9_101 ();
 FILLCELL_X2 FILLER_9_117 ();
 FILLCELL_X1 FILLER_9_119 ();
 FILLCELL_X4 FILLER_9_124 ();
 FILLCELL_X2 FILLER_9_128 ();
 FILLCELL_X1 FILLER_9_130 ();
 FILLCELL_X8 FILLER_9_152 ();
 FILLCELL_X4 FILLER_9_160 ();
 FILLCELL_X8 FILLER_9_181 ();
 FILLCELL_X16 FILLER_10_1 ();
 FILLCELL_X4 FILLER_10_17 ();
 FILLCELL_X2 FILLER_10_21 ();
 FILLCELL_X4 FILLER_10_26 ();
 FILLCELL_X2 FILLER_10_30 ();
 FILLCELL_X2 FILLER_10_48 ();
 FILLCELL_X32 FILLER_10_63 ();
 FILLCELL_X32 FILLER_10_95 ();
 FILLCELL_X4 FILLER_10_127 ();
 FILLCELL_X1 FILLER_10_131 ();
 FILLCELL_X2 FILLER_10_170 ();
 FILLCELL_X1 FILLER_10_172 ();
 FILLCELL_X8 FILLER_10_177 ();
 FILLCELL_X4 FILLER_10_185 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X2 FILLER_11_33 ();
 FILLCELL_X1 FILLER_11_35 ();
 FILLCELL_X8 FILLER_11_47 ();
 FILLCELL_X4 FILLER_11_55 ();
 FILLCELL_X2 FILLER_11_59 ();
 FILLCELL_X1 FILLER_11_61 ();
 FILLCELL_X16 FILLER_11_67 ();
 FILLCELL_X8 FILLER_11_83 ();
 FILLCELL_X4 FILLER_11_91 ();
 FILLCELL_X32 FILLER_11_100 ();
 FILLCELL_X1 FILLER_11_132 ();
 FILLCELL_X8 FILLER_11_137 ();
 FILLCELL_X4 FILLER_11_145 ();
 FILLCELL_X2 FILLER_11_149 ();
 FILLCELL_X4 FILLER_11_158 ();
 FILLCELL_X1 FILLER_11_162 ();
 FILLCELL_X8 FILLER_11_177 ();
 FILLCELL_X4 FILLER_11_185 ();
 FILLCELL_X8 FILLER_12_1 ();
 FILLCELL_X4 FILLER_12_9 ();
 FILLCELL_X2 FILLER_12_13 ();
 FILLCELL_X1 FILLER_12_15 ();
 FILLCELL_X16 FILLER_12_48 ();
 FILLCELL_X8 FILLER_12_64 ();
 FILLCELL_X4 FILLER_12_72 ();
 FILLCELL_X1 FILLER_12_76 ();
 FILLCELL_X2 FILLER_12_79 ();
 FILLCELL_X16 FILLER_12_105 ();
 FILLCELL_X8 FILLER_12_121 ();
 FILLCELL_X2 FILLER_12_129 ();
 FILLCELL_X1 FILLER_12_131 ();
 FILLCELL_X8 FILLER_12_136 ();
 FILLCELL_X1 FILLER_12_151 ();
 FILLCELL_X4 FILLER_12_166 ();
 FILLCELL_X4 FILLER_12_176 ();
 FILLCELL_X2 FILLER_12_180 ();
 FILLCELL_X1 FILLER_12_182 ();
 FILLCELL_X2 FILLER_12_186 ();
 FILLCELL_X1 FILLER_12_188 ();
 FILLCELL_X1 FILLER_13_8 ();
 FILLCELL_X1 FILLER_13_40 ();
 FILLCELL_X8 FILLER_13_45 ();
 FILLCELL_X1 FILLER_13_53 ();
 FILLCELL_X8 FILLER_13_62 ();
 FILLCELL_X4 FILLER_13_70 ();
 FILLCELL_X2 FILLER_13_74 ();
 FILLCELL_X1 FILLER_13_76 ();
 FILLCELL_X4 FILLER_13_107 ();
 FILLCELL_X2 FILLER_13_111 ();
 FILLCELL_X1 FILLER_13_113 ();
 FILLCELL_X8 FILLER_13_118 ();
 FILLCELL_X16 FILLER_13_136 ();
 FILLCELL_X4 FILLER_13_159 ();
 FILLCELL_X16 FILLER_13_166 ();
 FILLCELL_X4 FILLER_13_182 ();
 FILLCELL_X2 FILLER_13_186 ();
 FILLCELL_X1 FILLER_13_188 ();
 FILLCELL_X8 FILLER_14_1 ();
 FILLCELL_X2 FILLER_14_16 ();
 FILLCELL_X1 FILLER_14_18 ();
 FILLCELL_X1 FILLER_14_22 ();
 FILLCELL_X2 FILLER_14_47 ();
 FILLCELL_X1 FILLER_14_49 ();
 FILLCELL_X8 FILLER_14_57 ();
 FILLCELL_X4 FILLER_14_65 ();
 FILLCELL_X2 FILLER_14_69 ();
 FILLCELL_X1 FILLER_14_71 ();
 FILLCELL_X1 FILLER_14_107 ();
 FILLCELL_X1 FILLER_14_112 ();
 FILLCELL_X1 FILLER_14_116 ();
 FILLCELL_X2 FILLER_14_148 ();
 FILLCELL_X32 FILLER_14_157 ();
 FILLCELL_X16 FILLER_15_1 ();
 FILLCELL_X8 FILLER_15_17 ();
 FILLCELL_X1 FILLER_15_51 ();
 FILLCELL_X16 FILLER_15_56 ();
 FILLCELL_X8 FILLER_15_72 ();
 FILLCELL_X8 FILLER_15_89 ();
 FILLCELL_X1 FILLER_15_97 ();
 FILLCELL_X8 FILLER_15_101 ();
 FILLCELL_X4 FILLER_15_109 ();
 FILLCELL_X16 FILLER_15_128 ();
 FILLCELL_X8 FILLER_15_144 ();
 FILLCELL_X2 FILLER_15_152 ();
 FILLCELL_X1 FILLER_15_154 ();
 FILLCELL_X2 FILLER_15_179 ();
 FILLCELL_X4 FILLER_15_184 ();
 FILLCELL_X1 FILLER_15_188 ();
 FILLCELL_X8 FILLER_16_1 ();
 FILLCELL_X4 FILLER_16_9 ();
 FILLCELL_X4 FILLER_16_30 ();
 FILLCELL_X1 FILLER_16_34 ();
 FILLCELL_X4 FILLER_16_45 ();
 FILLCELL_X2 FILLER_16_66 ();
 FILLCELL_X8 FILLER_16_85 ();
 FILLCELL_X2 FILLER_16_93 ();
 FILLCELL_X1 FILLER_16_95 ();
 FILLCELL_X16 FILLER_16_131 ();
 FILLCELL_X8 FILLER_16_147 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X8 FILLER_17_97 ();
 FILLCELL_X2 FILLER_17_105 ();
 FILLCELL_X1 FILLER_17_107 ();
 FILLCELL_X16 FILLER_17_125 ();
 FILLCELL_X8 FILLER_17_141 ();
 FILLCELL_X4 FILLER_17_149 ();
 FILLCELL_X2 FILLER_17_153 ();
 FILLCELL_X4 FILLER_17_162 ();
 FILLCELL_X2 FILLER_17_174 ();
 FILLCELL_X2 FILLER_17_183 ();
 FILLCELL_X1 FILLER_17_185 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X8 FILLER_18_129 ();
 FILLCELL_X4 FILLER_18_137 ();
 FILLCELL_X4 FILLER_18_145 ();
 FILLCELL_X8 FILLER_18_159 ();
 FILLCELL_X2 FILLER_18_167 ();
 FILLCELL_X1 FILLER_18_169 ();
 FILLCELL_X8 FILLER_18_180 ();
 FILLCELL_X1 FILLER_18_188 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X8 FILLER_19_129 ();
 FILLCELL_X8 FILLER_19_154 ();
 FILLCELL_X2 FILLER_19_162 ();
 FILLCELL_X1 FILLER_19_164 ();
 FILLCELL_X16 FILLER_19_169 ();
 FILLCELL_X4 FILLER_19_185 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X2 FILLER_20_161 ();
 FILLCELL_X1 FILLER_20_163 ();
 FILLCELL_X8 FILLER_20_181 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X16 FILLER_21_161 ();
 FILLCELL_X8 FILLER_21_177 ();
 FILLCELL_X4 FILLER_21_185 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X16 FILLER_22_161 ();
 FILLCELL_X8 FILLER_22_177 ();
 FILLCELL_X4 FILLER_22_185 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X16 FILLER_23_161 ();
 FILLCELL_X8 FILLER_23_177 ();
 FILLCELL_X4 FILLER_23_185 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X16 FILLER_24_65 ();
 FILLCELL_X2 FILLER_24_81 ();
 FILLCELL_X1 FILLER_24_83 ();
 FILLCELL_X32 FILLER_24_87 ();
 FILLCELL_X32 FILLER_24_119 ();
 FILLCELL_X32 FILLER_24_151 ();
 FILLCELL_X4 FILLER_24_183 ();
 FILLCELL_X2 FILLER_24_187 ();
endmodule
