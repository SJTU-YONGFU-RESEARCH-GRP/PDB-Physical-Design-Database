module async_fifo (almost_empty,
    almost_full,
    empty,
    full,
    pointer_wraparound_flag,
    rd_clk,
    rd_en,
    rd_rst_n,
    sync_error_flag,
    wr_clk,
    wr_en,
    wr_rst_n,
    rd_count,
    rd_data,
    wr_count,
    wr_data);
 output almost_empty;
 output almost_full;
 output empty;
 output full;
 output pointer_wraparound_flag;
 input rd_clk;
 input rd_en;
 input rd_rst_n;
 output sync_error_flag;
 input wr_clk;
 input wr_en;
 input wr_rst_n;
 output [4:0] rd_count;
 output [7:0] rd_data;
 output [4:0] wr_count;
 input [7:0] wr_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire \mem[0][0] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[10][0] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[11][0] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[12][0] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[13][0] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[14][0] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[15][0] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[1][0] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[2][0] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[3][0] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[4][0] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[5][0] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[6][0] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[7][0] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[8][0] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[9][0] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \rd_ptr_bin[0] ;
 wire \rd_ptr_bin[1] ;
 wire \rd_ptr_bin[2] ;
 wire \rd_ptr_bin[3] ;
 wire \rd_ptr_bin[4] ;
 wire \rd_ptr_gray[0] ;
 wire \rd_ptr_gray[1] ;
 wire \rd_ptr_gray[2] ;
 wire \rd_ptr_gray[3] ;
 wire \rd_ptr_gray_sync1[0] ;
 wire \rd_ptr_gray_sync1[1] ;
 wire \rd_ptr_gray_sync1[2] ;
 wire \rd_ptr_gray_sync1[3] ;
 wire \rd_ptr_gray_sync1[4] ;
 wire \rd_ptr_gray_sync2[0] ;
 wire \rd_ptr_gray_sync2[1] ;
 wire \rd_ptr_gray_sync2[2] ;
 wire \rd_ptr_gray_sync2[3] ;
 wire \rd_ptr_gray_sync2[4] ;
 wire \rd_ptr_sync[0] ;
 wire \rd_ptr_sync[1] ;
 wire \rd_ptr_sync[2] ;
 wire \rd_ptr_sync[3] ;
 wire \rd_ptr_sync[4] ;
 wire \wr_ptr_bin[0] ;
 wire \wr_ptr_bin[1] ;
 wire \wr_ptr_bin[2] ;
 wire \wr_ptr_bin[3] ;
 wire \wr_ptr_bin[4] ;
 wire \wr_ptr_gray[0] ;
 wire \wr_ptr_gray[1] ;
 wire \wr_ptr_gray[2] ;
 wire \wr_ptr_gray[3] ;
 wire \wr_ptr_gray_sync1[0] ;
 wire \wr_ptr_gray_sync1[1] ;
 wire \wr_ptr_gray_sync1[2] ;
 wire \wr_ptr_gray_sync1[3] ;
 wire \wr_ptr_gray_sync1[4] ;
 wire \wr_ptr_gray_sync2[0] ;
 wire \wr_ptr_gray_sync2[1] ;
 wire \wr_ptr_gray_sync2[2] ;
 wire \wr_ptr_gray_sync2[3] ;
 wire \wr_ptr_gray_sync2[4] ;
 wire \wr_ptr_sync[0] ;
 wire \wr_ptr_sync[1] ;
 wire \wr_ptr_sync[2] ;
 wire \wr_ptr_sync[3] ;
 wire \wr_ptr_sync[4] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;

 sky130_fd_sc_hd__inv_1 _338_ (.A(_306_),
    .Y(net20));
 sky130_fd_sc_hd__nand2_1 _339_ (.A(_299_),
    .B(_301_),
    .Y(_057_));
 sky130_fd_sc_hd__nand3_1 _340_ (.A(_296_),
    .B(_304_),
    .C(_306_),
    .Y(_058_));
 sky130_fd_sc_hd__nor2_1 _341_ (.A(_057_),
    .B(_058_),
    .Y(_000_));
 sky130_fd_sc_hd__a21o_1 _342_ (.A1(_304_),
    .A2(_290_),
    .B1(_303_),
    .X(_059_));
 sky130_fd_sc_hd__a21oi_1 _343_ (.A1(_296_),
    .A2(_059_),
    .B1(_295_),
    .Y(_060_));
 sky130_fd_sc_hd__xnor2_1 _344_ (.A(_299_),
    .B(_060_),
    .Y(net24));
 sky130_fd_sc_hd__xor2_1 _345_ (.A(_304_),
    .B(_290_),
    .X(net22));
 sky130_fd_sc_hd__nor2b_1 _346_ (.A(_308_),
    .B_N(_301_),
    .Y(_061_));
 sky130_fd_sc_hd__o21a_1 _347_ (.A1(_300_),
    .A2(_061_),
    .B1(_304_),
    .X(_062_));
 sky130_fd_sc_hd__o21ai_0 _348_ (.A1(_303_),
    .A2(_062_),
    .B1(_296_),
    .Y(_063_));
 sky130_fd_sc_hd__or3_1 _349_ (.A(_296_),
    .B(_303_),
    .C(_062_),
    .X(_064_));
 sky130_fd_sc_hd__and2_0 _350_ (.A(_063_),
    .B(_064_),
    .X(net23));
 sky130_fd_sc_hd__inv_1 _351_ (.A(_313_),
    .Y(net34));
 sky130_fd_sc_hd__inv_1 _352_ (.A(_319_),
    .Y(_065_));
 sky130_fd_sc_hd__nor2b_1 _353_ (.A(_314_),
    .B_N(_310_),
    .Y(_066_));
 sky130_fd_sc_hd__o21ai_0 _354_ (.A1(_316_),
    .A2(_066_),
    .B1(_320_),
    .Y(_067_));
 sky130_fd_sc_hd__a21boi_0 _355_ (.A1(_065_),
    .A2(_067_),
    .B1_N(_324_),
    .Y(_068_));
 sky130_fd_sc_hd__nor3b_1 _356_ (.A(_324_),
    .B(_319_),
    .C_N(_067_),
    .Y(_069_));
 sky130_fd_sc_hd__nor2_1 _357_ (.A(_068_),
    .B(_069_),
    .Y(net37));
 sky130_fd_sc_hd__a21o_1 _358_ (.A1(_320_),
    .A2(_293_),
    .B1(_319_),
    .X(_070_));
 sky130_fd_sc_hd__a21oi_1 _359_ (.A1(_324_),
    .A2(_070_),
    .B1(_323_),
    .Y(_071_));
 sky130_fd_sc_hd__xor2_1 _360_ (.A(_328_),
    .B(_071_),
    .X(_072_));
 sky130_fd_sc_hd__inv_1 _361_ (.A(_072_),
    .Y(net38));
 sky130_fd_sc_hd__nor4_1 _362_ (.A(\rd_ptr_sync[1] ),
    .B(\rd_ptr_sync[0] ),
    .C(\rd_ptr_sync[3] ),
    .D(\rd_ptr_sync[2] ),
    .Y(_073_));
 sky130_fd_sc_hd__clkbuf_4 _363_ (.A(\wr_ptr_bin[3] ),
    .X(_074_));
 sky130_fd_sc_hd__clkbuf_4 _364_ (.A(\wr_ptr_bin[2] ),
    .X(_075_));
 sky130_fd_sc_hd__or2_0 _365_ (.A(_074_),
    .B(_075_),
    .X(_076_));
 sky130_fd_sc_hd__buf_4 _366_ (.A(_076_),
    .X(_077_));
 sky130_fd_sc_hd__nand2_1 _367_ (.A(\wr_ptr_bin[4] ),
    .B(_330_),
    .Y(_078_));
 sky130_fd_sc_hd__nor3_1 _368_ (.A(_073_),
    .B(_077_),
    .C(_078_),
    .Y(_010_));
 sky130_fd_sc_hd__nand3_1 _369_ (.A(_310_),
    .B(_324_),
    .C(_320_),
    .Y(_079_));
 sky130_fd_sc_hd__nor3_1 _370_ (.A(net34),
    .B(_328_),
    .C(_079_),
    .Y(_001_));
 sky130_fd_sc_hd__inv_1 _371_ (.A(_075_),
    .Y(_321_));
 sky130_fd_sc_hd__nand2_4 _372_ (.A(_074_),
    .B(_321_),
    .Y(_080_));
 sky130_fd_sc_hd__nor2b_1 _373_ (.A(net18),
    .B_N(net13),
    .Y(_081_));
 sky130_fd_sc_hd__buf_6 _374_ (.A(_081_),
    .X(_082_));
 sky130_fd_sc_hd__nand2_8 _375_ (.A(_331_),
    .B(_082_),
    .Y(_083_));
 sky130_fd_sc_hd__nor2_4 _376_ (.A(_080_),
    .B(_083_),
    .Y(_012_));
 sky130_fd_sc_hd__nand2_4 _377_ (.A(_333_),
    .B(_082_),
    .Y(_084_));
 sky130_fd_sc_hd__nor2_4 _378_ (.A(_080_),
    .B(_084_),
    .Y(_026_));
 sky130_fd_sc_hd__nand2_8 _379_ (.A(_330_),
    .B(_082_),
    .Y(_085_));
 sky130_fd_sc_hd__nor2_4 _380_ (.A(_080_),
    .B(_085_),
    .Y(_025_));
 sky130_fd_sc_hd__inv_1 _381_ (.A(_074_),
    .Y(_325_));
 sky130_fd_sc_hd__nand2_4 _382_ (.A(_325_),
    .B(_075_),
    .Y(_086_));
 sky130_fd_sc_hd__nand2_8 _383_ (.A(_335_),
    .B(_082_),
    .Y(_087_));
 sky130_fd_sc_hd__nor2_4 _384_ (.A(_086_),
    .B(_087_),
    .Y(_024_));
 sky130_fd_sc_hd__nand2_4 _385_ (.A(_074_),
    .B(_075_),
    .Y(_088_));
 sky130_fd_sc_hd__nor2_4 _386_ (.A(_087_),
    .B(_088_),
    .Y(_017_));
 sky130_fd_sc_hd__nor2_4 _387_ (.A(_083_),
    .B(_086_),
    .Y(_023_));
 sky130_fd_sc_hd__nor2_4 _388_ (.A(_083_),
    .B(_088_),
    .Y(_016_));
 sky130_fd_sc_hd__nor2_4 _389_ (.A(_084_),
    .B(_086_),
    .Y(_022_));
 sky130_fd_sc_hd__buf_4 _390_ (.A(\rd_ptr_bin[2] ),
    .X(_089_));
 sky130_fd_sc_hd__inv_1 _391_ (.A(_089_),
    .Y(_302_));
 sky130_fd_sc_hd__buf_2 _392_ (.A(\rd_ptr_bin[3] ),
    .X(_090_));
 sky130_fd_sc_hd__inv_1 _393_ (.A(_090_),
    .Y(_294_));
 sky130_fd_sc_hd__nor2_4 _394_ (.A(_085_),
    .B(_086_),
    .Y(_021_));
 sky130_fd_sc_hd__nor2_4 _395_ (.A(_077_),
    .B(_087_),
    .Y(_020_));
 sky130_fd_sc_hd__nor2_4 _396_ (.A(_077_),
    .B(_083_),
    .Y(_019_));
 sky130_fd_sc_hd__nor2_4 _397_ (.A(_077_),
    .B(_084_),
    .Y(_018_));
 sky130_fd_sc_hd__nor2_4 _398_ (.A(_077_),
    .B(_085_),
    .Y(_011_));
 sky130_fd_sc_hd__nor2_4 _399_ (.A(_084_),
    .B(_088_),
    .Y(_015_));
 sky130_fd_sc_hd__nor2_4 _400_ (.A(_085_),
    .B(_088_),
    .Y(_014_));
 sky130_fd_sc_hd__xor2_1 _401_ (.A(\wr_ptr_gray_sync2[4] ),
    .B(\wr_ptr_gray_sync2[3] ),
    .X(_005_));
 sky130_fd_sc_hd__xnor2_1 _402_ (.A(\wr_ptr_gray_sync2[2] ),
    .B(_005_),
    .Y(_091_));
 sky130_fd_sc_hd__inv_1 _403_ (.A(_091_),
    .Y(_004_));
 sky130_fd_sc_hd__xnor2_1 _404_ (.A(\wr_ptr_gray_sync2[1] ),
    .B(_091_),
    .Y(_003_));
 sky130_fd_sc_hd__xor2_1 _405_ (.A(\wr_ptr_gray_sync2[0] ),
    .B(_003_),
    .X(_002_));
 sky130_fd_sc_hd__xor2_1 _406_ (.A(\rd_ptr_gray_sync2[4] ),
    .B(\rd_ptr_gray_sync2[3] ),
    .X(_009_));
 sky130_fd_sc_hd__xnor2_1 _407_ (.A(\rd_ptr_gray_sync2[2] ),
    .B(_009_),
    .Y(_092_));
 sky130_fd_sc_hd__inv_1 _408_ (.A(_092_),
    .Y(_008_));
 sky130_fd_sc_hd__xnor2_1 _409_ (.A(\rd_ptr_gray_sync2[1] ),
    .B(_092_),
    .Y(_007_));
 sky130_fd_sc_hd__xor2_1 _410_ (.A(\rd_ptr_gray_sync2[0] ),
    .B(_007_),
    .X(_006_));
 sky130_fd_sc_hd__nor2_4 _411_ (.A(_080_),
    .B(_087_),
    .Y(_013_));
 sky130_fd_sc_hd__buf_2 _412_ (.A(\rd_ptr_bin[1] ),
    .X(_093_));
 sky130_fd_sc_hd__buf_4 _413_ (.A(_093_),
    .X(_094_));
 sky130_fd_sc_hd__inv_1 _414_ (.A(_094_),
    .Y(_288_));
 sky130_fd_sc_hd__clkbuf_4 _415_ (.A(\rd_ptr_bin[0] ),
    .X(_095_));
 sky130_fd_sc_hd__inv_1 _416_ (.A(_095_),
    .Y(_029_));
 sky130_fd_sc_hd__inv_1 _417_ (.A(\rd_ptr_sync[0] ),
    .Y(_311_));
 sky130_fd_sc_hd__inv_1 _418_ (.A(\rd_ptr_sync[1] ),
    .Y(_291_));
 sky130_fd_sc_hd__inv_1 _419_ (.A(\rd_ptr_sync[2] ),
    .Y(_318_));
 sky130_fd_sc_hd__inv_1 _420_ (.A(\rd_ptr_sync[3] ),
    .Y(_322_));
 sky130_fd_sc_hd__clkinvlp_4 _421_ (.A(\wr_ptr_bin[0] ),
    .Y(_027_));
 sky130_fd_sc_hd__inv_1 _422_ (.A(\wr_ptr_sync[4] ),
    .Y(_297_));
 sky130_fd_sc_hd__inv_1 _423_ (.A(_308_),
    .Y(_289_));
 sky130_fd_sc_hd__inv_1 _424_ (.A(\wr_ptr_sync[0] ),
    .Y(_307_));
 sky130_fd_sc_hd__inv_1 _425_ (.A(_314_),
    .Y(_292_));
 sky130_fd_sc_hd__inv_1 _426_ (.A(\wr_ptr_bin[4] ),
    .Y(_326_));
 sky130_fd_sc_hd__inv_1 _427_ (.A(\wr_ptr_bin[1] ),
    .Y(_317_));
 sky130_fd_sc_hd__nand2b_1 _428_ (.A_N(net17),
    .B(net2),
    .Y(_096_));
 sky130_fd_sc_hd__buf_2 _429_ (.A(_096_),
    .X(_097_));
 sky130_fd_sc_hd__buf_2 _430_ (.A(_097_),
    .X(_098_));
 sky130_fd_sc_hd__nand2_1 _431_ (.A(net25),
    .B(_098_),
    .Y(_099_));
 sky130_fd_sc_hd__nor2b_1 _432_ (.A(_089_),
    .B_N(_095_),
    .Y(_100_));
 sky130_fd_sc_hd__buf_2 _433_ (.A(_100_),
    .X(_101_));
 sky130_fd_sc_hd__clkbuf_4 _434_ (.A(_101_),
    .X(_102_));
 sky130_fd_sc_hd__buf_4 _435_ (.A(_094_),
    .X(_103_));
 sky130_fd_sc_hd__mux2i_1 _436_ (.A0(\mem[9][0] ),
    .A1(\mem[11][0] ),
    .S(_103_),
    .Y(_104_));
 sky130_fd_sc_hd__nand2_1 _437_ (.A(_102_),
    .B(_104_),
    .Y(_105_));
 sky130_fd_sc_hd__and2_0 _438_ (.A(_095_),
    .B(_089_),
    .X(_106_));
 sky130_fd_sc_hd__buf_2 _439_ (.A(_106_),
    .X(_107_));
 sky130_fd_sc_hd__buf_6 _440_ (.A(_107_),
    .X(_108_));
 sky130_fd_sc_hd__buf_6 _441_ (.A(_093_),
    .X(_109_));
 sky130_fd_sc_hd__mux2i_1 _442_ (.A0(\mem[13][0] ),
    .A1(\mem[15][0] ),
    .S(_109_),
    .Y(_110_));
 sky130_fd_sc_hd__nor2b_1 _443_ (.A(_095_),
    .B_N(_089_),
    .Y(_111_));
 sky130_fd_sc_hd__buf_2 _444_ (.A(_111_),
    .X(_112_));
 sky130_fd_sc_hd__clkbuf_4 _445_ (.A(_112_),
    .X(_113_));
 sky130_fd_sc_hd__buf_6 _446_ (.A(_093_),
    .X(_114_));
 sky130_fd_sc_hd__mux2i_2 _447_ (.A0(\mem[12][0] ),
    .A1(\mem[14][0] ),
    .S(_114_),
    .Y(_115_));
 sky130_fd_sc_hd__a22oi_2 _448_ (.A1(_108_),
    .A2(_110_),
    .B1(_113_),
    .B2(_115_),
    .Y(_116_));
 sky130_fd_sc_hd__nor2_4 _449_ (.A(_294_),
    .B(_097_),
    .Y(_117_));
 sky130_fd_sc_hd__nor2_4 _450_ (.A(_095_),
    .B(_089_),
    .Y(_118_));
 sky130_fd_sc_hd__clkbuf_4 _451_ (.A(_118_),
    .X(_119_));
 sky130_fd_sc_hd__mux2i_1 _452_ (.A0(\mem[8][0] ),
    .A1(\mem[10][0] ),
    .S(_103_),
    .Y(_120_));
 sky130_fd_sc_hd__nand2_1 _453_ (.A(_119_),
    .B(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__nand4_1 _454_ (.A(_105_),
    .B(_116_),
    .C(_117_),
    .D(_121_),
    .Y(_122_));
 sky130_fd_sc_hd__mux2i_1 _455_ (.A0(\mem[5][0] ),
    .A1(\mem[7][0] ),
    .S(_114_),
    .Y(_123_));
 sky130_fd_sc_hd__buf_6 _456_ (.A(_094_),
    .X(_124_));
 sky130_fd_sc_hd__mux2i_1 _457_ (.A0(\mem[1][0] ),
    .A1(\mem[3][0] ),
    .S(_124_),
    .Y(_125_));
 sky130_fd_sc_hd__a22oi_1 _458_ (.A1(_108_),
    .A2(_123_),
    .B1(_125_),
    .B2(_102_),
    .Y(_126_));
 sky130_fd_sc_hd__nor2_4 _459_ (.A(_090_),
    .B(_097_),
    .Y(_127_));
 sky130_fd_sc_hd__mux2i_1 _460_ (.A0(\mem[4][0] ),
    .A1(\mem[6][0] ),
    .S(_114_),
    .Y(_128_));
 sky130_fd_sc_hd__buf_6 _461_ (.A(_094_),
    .X(_129_));
 sky130_fd_sc_hd__mux2i_1 _462_ (.A0(\mem[0][0] ),
    .A1(\mem[2][0] ),
    .S(_129_),
    .Y(_130_));
 sky130_fd_sc_hd__a22oi_1 _463_ (.A1(_113_),
    .A2(_128_),
    .B1(_130_),
    .B2(_119_),
    .Y(_131_));
 sky130_fd_sc_hd__nand3_1 _464_ (.A(_126_),
    .B(_127_),
    .C(_131_),
    .Y(_132_));
 sky130_fd_sc_hd__nand3_1 _465_ (.A(_099_),
    .B(_122_),
    .C(_132_),
    .Y(_031_));
 sky130_fd_sc_hd__nand2_1 _466_ (.A(net26),
    .B(_098_),
    .Y(_133_));
 sky130_fd_sc_hd__mux2i_1 _467_ (.A0(\mem[9][1] ),
    .A1(\mem[11][1] ),
    .S(_103_),
    .Y(_134_));
 sky130_fd_sc_hd__nand2_1 _468_ (.A(_102_),
    .B(_134_),
    .Y(_135_));
 sky130_fd_sc_hd__mux2i_1 _469_ (.A0(\mem[13][1] ),
    .A1(\mem[15][1] ),
    .S(_109_),
    .Y(_136_));
 sky130_fd_sc_hd__buf_6 _470_ (.A(_093_),
    .X(_137_));
 sky130_fd_sc_hd__mux2i_2 _471_ (.A0(\mem[12][1] ),
    .A1(\mem[14][1] ),
    .S(_137_),
    .Y(_138_));
 sky130_fd_sc_hd__a22oi_2 _472_ (.A1(_108_),
    .A2(_136_),
    .B1(_138_),
    .B2(_113_),
    .Y(_139_));
 sky130_fd_sc_hd__mux2i_1 _473_ (.A0(\mem[8][1] ),
    .A1(\mem[10][1] ),
    .S(_124_),
    .Y(_140_));
 sky130_fd_sc_hd__nand2_1 _474_ (.A(_119_),
    .B(_140_),
    .Y(_141_));
 sky130_fd_sc_hd__nand4_1 _475_ (.A(_117_),
    .B(_135_),
    .C(_139_),
    .D(_141_),
    .Y(_142_));
 sky130_fd_sc_hd__mux2i_1 _476_ (.A0(\mem[0][1] ),
    .A1(\mem[2][1] ),
    .S(_114_),
    .Y(_143_));
 sky130_fd_sc_hd__mux2i_1 _477_ (.A0(\mem[1][1] ),
    .A1(\mem[3][1] ),
    .S(_124_),
    .Y(_144_));
 sky130_fd_sc_hd__a22oi_1 _478_ (.A1(_118_),
    .A2(_143_),
    .B1(_144_),
    .B2(_102_),
    .Y(_145_));
 sky130_fd_sc_hd__mux2i_2 _479_ (.A0(\mem[4][1] ),
    .A1(\mem[6][1] ),
    .S(_109_),
    .Y(_146_));
 sky130_fd_sc_hd__mux2i_1 _480_ (.A0(\mem[5][1] ),
    .A1(\mem[7][1] ),
    .S(_129_),
    .Y(_147_));
 sky130_fd_sc_hd__a22oi_1 _481_ (.A1(_113_),
    .A2(_146_),
    .B1(_147_),
    .B2(_108_),
    .Y(_148_));
 sky130_fd_sc_hd__nand3_1 _482_ (.A(_127_),
    .B(_145_),
    .C(_148_),
    .Y(_149_));
 sky130_fd_sc_hd__nand3_1 _483_ (.A(_133_),
    .B(_142_),
    .C(_149_),
    .Y(_032_));
 sky130_fd_sc_hd__nand2_1 _484_ (.A(net27),
    .B(_098_),
    .Y(_150_));
 sky130_fd_sc_hd__mux2i_1 _485_ (.A0(\mem[9][2] ),
    .A1(\mem[11][2] ),
    .S(_103_),
    .Y(_151_));
 sky130_fd_sc_hd__nand2_1 _486_ (.A(_102_),
    .B(_151_),
    .Y(_152_));
 sky130_fd_sc_hd__mux2i_1 _487_ (.A0(\mem[13][2] ),
    .A1(\mem[15][2] ),
    .S(_109_),
    .Y(_153_));
 sky130_fd_sc_hd__mux2i_2 _488_ (.A0(\mem[12][2] ),
    .A1(\mem[14][2] ),
    .S(_137_),
    .Y(_154_));
 sky130_fd_sc_hd__a22oi_2 _489_ (.A1(_107_),
    .A2(_153_),
    .B1(_154_),
    .B2(_113_),
    .Y(_155_));
 sky130_fd_sc_hd__mux2i_1 _490_ (.A0(\mem[8][2] ),
    .A1(\mem[10][2] ),
    .S(_124_),
    .Y(_156_));
 sky130_fd_sc_hd__nand2_1 _491_ (.A(_119_),
    .B(_156_),
    .Y(_157_));
 sky130_fd_sc_hd__nand4_1 _492_ (.A(_117_),
    .B(_152_),
    .C(_155_),
    .D(_157_),
    .Y(_158_));
 sky130_fd_sc_hd__mux2i_1 _493_ (.A0(\mem[5][2] ),
    .A1(\mem[7][2] ),
    .S(_114_),
    .Y(_159_));
 sky130_fd_sc_hd__mux2i_1 _494_ (.A0(\mem[1][2] ),
    .A1(\mem[3][2] ),
    .S(_124_),
    .Y(_160_));
 sky130_fd_sc_hd__a22oi_1 _495_ (.A1(_108_),
    .A2(_159_),
    .B1(_160_),
    .B2(_101_),
    .Y(_161_));
 sky130_fd_sc_hd__mux2i_2 _496_ (.A0(\mem[4][2] ),
    .A1(\mem[6][2] ),
    .S(_109_),
    .Y(_162_));
 sky130_fd_sc_hd__mux2i_1 _497_ (.A0(\mem[0][2] ),
    .A1(\mem[2][2] ),
    .S(_129_),
    .Y(_163_));
 sky130_fd_sc_hd__a22oi_2 _498_ (.A1(_112_),
    .A2(_162_),
    .B1(_163_),
    .B2(_119_),
    .Y(_164_));
 sky130_fd_sc_hd__nand3_1 _499_ (.A(_127_),
    .B(_161_),
    .C(_164_),
    .Y(_165_));
 sky130_fd_sc_hd__nand3_1 _500_ (.A(_150_),
    .B(_158_),
    .C(_165_),
    .Y(_033_));
 sky130_fd_sc_hd__nand2_1 _501_ (.A(net28),
    .B(_098_),
    .Y(_166_));
 sky130_fd_sc_hd__mux2i_1 _502_ (.A0(\mem[9][3] ),
    .A1(\mem[11][3] ),
    .S(_103_),
    .Y(_167_));
 sky130_fd_sc_hd__nand2_1 _503_ (.A(_102_),
    .B(_167_),
    .Y(_168_));
 sky130_fd_sc_hd__mux2i_1 _504_ (.A0(\mem[13][3] ),
    .A1(\mem[15][3] ),
    .S(_094_),
    .Y(_169_));
 sky130_fd_sc_hd__mux2i_1 _505_ (.A0(\mem[12][3] ),
    .A1(\mem[14][3] ),
    .S(_137_),
    .Y(_170_));
 sky130_fd_sc_hd__a22oi_1 _506_ (.A1(_107_),
    .A2(_169_),
    .B1(_170_),
    .B2(_113_),
    .Y(_171_));
 sky130_fd_sc_hd__mux2i_1 _507_ (.A0(\mem[8][3] ),
    .A1(\mem[10][3] ),
    .S(_124_),
    .Y(_172_));
 sky130_fd_sc_hd__nand2_1 _508_ (.A(_119_),
    .B(_172_),
    .Y(_173_));
 sky130_fd_sc_hd__nand4_1 _509_ (.A(_117_),
    .B(_168_),
    .C(_171_),
    .D(_173_),
    .Y(_174_));
 sky130_fd_sc_hd__mux2i_1 _510_ (.A0(\mem[5][3] ),
    .A1(\mem[7][3] ),
    .S(_114_),
    .Y(_175_));
 sky130_fd_sc_hd__mux2i_1 _511_ (.A0(\mem[1][3] ),
    .A1(\mem[3][3] ),
    .S(_129_),
    .Y(_176_));
 sky130_fd_sc_hd__a22oi_1 _512_ (.A1(_108_),
    .A2(_175_),
    .B1(_176_),
    .B2(_101_),
    .Y(_177_));
 sky130_fd_sc_hd__mux2i_1 _513_ (.A0(\mem[4][3] ),
    .A1(\mem[6][3] ),
    .S(_109_),
    .Y(_178_));
 sky130_fd_sc_hd__mux2i_1 _514_ (.A0(\mem[0][3] ),
    .A1(\mem[2][3] ),
    .S(_129_),
    .Y(_179_));
 sky130_fd_sc_hd__a22oi_2 _515_ (.A1(_112_),
    .A2(_178_),
    .B1(_179_),
    .B2(_118_),
    .Y(_180_));
 sky130_fd_sc_hd__nand3_1 _516_ (.A(_127_),
    .B(_177_),
    .C(_180_),
    .Y(_181_));
 sky130_fd_sc_hd__nand3_1 _517_ (.A(_166_),
    .B(_174_),
    .C(_181_),
    .Y(_034_));
 sky130_fd_sc_hd__nand2_1 _518_ (.A(net29),
    .B(_098_),
    .Y(_182_));
 sky130_fd_sc_hd__mux2i_1 _519_ (.A0(\mem[9][4] ),
    .A1(\mem[11][4] ),
    .S(_103_),
    .Y(_183_));
 sky130_fd_sc_hd__nand2_1 _520_ (.A(_102_),
    .B(_183_),
    .Y(_184_));
 sky130_fd_sc_hd__mux2i_2 _521_ (.A0(\mem[13][4] ),
    .A1(\mem[15][4] ),
    .S(_094_),
    .Y(_185_));
 sky130_fd_sc_hd__mux2i_1 _522_ (.A0(\mem[12][4] ),
    .A1(\mem[14][4] ),
    .S(_137_),
    .Y(_186_));
 sky130_fd_sc_hd__a22oi_2 _523_ (.A1(_107_),
    .A2(_185_),
    .B1(_186_),
    .B2(_113_),
    .Y(_187_));
 sky130_fd_sc_hd__mux2i_1 _524_ (.A0(\mem[8][4] ),
    .A1(\mem[10][4] ),
    .S(_124_),
    .Y(_188_));
 sky130_fd_sc_hd__nand2_1 _525_ (.A(_119_),
    .B(_188_),
    .Y(_189_));
 sky130_fd_sc_hd__nand4_1 _526_ (.A(_117_),
    .B(_184_),
    .C(_187_),
    .D(_189_),
    .Y(_190_));
 sky130_fd_sc_hd__mux2i_1 _527_ (.A0(\mem[5][4] ),
    .A1(\mem[7][4] ),
    .S(_114_),
    .Y(_191_));
 sky130_fd_sc_hd__mux2i_1 _528_ (.A0(\mem[1][4] ),
    .A1(\mem[3][4] ),
    .S(_129_),
    .Y(_192_));
 sky130_fd_sc_hd__a22oi_1 _529_ (.A1(_108_),
    .A2(_191_),
    .B1(_192_),
    .B2(_101_),
    .Y(_193_));
 sky130_fd_sc_hd__mux2i_1 _530_ (.A0(\mem[4][4] ),
    .A1(\mem[6][4] ),
    .S(_109_),
    .Y(_194_));
 sky130_fd_sc_hd__mux2i_1 _531_ (.A0(\mem[0][4] ),
    .A1(\mem[2][4] ),
    .S(_129_),
    .Y(_195_));
 sky130_fd_sc_hd__a22oi_2 _532_ (.A1(_112_),
    .A2(_194_),
    .B1(_195_),
    .B2(_118_),
    .Y(_196_));
 sky130_fd_sc_hd__nand3_1 _533_ (.A(_127_),
    .B(_193_),
    .C(_196_),
    .Y(_197_));
 sky130_fd_sc_hd__nand3_1 _534_ (.A(_182_),
    .B(_190_),
    .C(_197_),
    .Y(_035_));
 sky130_fd_sc_hd__nand2_1 _535_ (.A(net30),
    .B(_098_),
    .Y(_198_));
 sky130_fd_sc_hd__mux2i_1 _536_ (.A0(\mem[9][5] ),
    .A1(\mem[11][5] ),
    .S(_103_),
    .Y(_199_));
 sky130_fd_sc_hd__nand2_1 _537_ (.A(_102_),
    .B(_199_),
    .Y(_200_));
 sky130_fd_sc_hd__mux2i_1 _538_ (.A0(\mem[13][5] ),
    .A1(\mem[15][5] ),
    .S(_094_),
    .Y(_201_));
 sky130_fd_sc_hd__mux2i_1 _539_ (.A0(\mem[12][5] ),
    .A1(\mem[14][5] ),
    .S(_137_),
    .Y(_202_));
 sky130_fd_sc_hd__a22oi_2 _540_ (.A1(_107_),
    .A2(_201_),
    .B1(_202_),
    .B2(_113_),
    .Y(_203_));
 sky130_fd_sc_hd__mux2i_1 _541_ (.A0(\mem[8][5] ),
    .A1(\mem[10][5] ),
    .S(_124_),
    .Y(_204_));
 sky130_fd_sc_hd__nand2_1 _542_ (.A(_119_),
    .B(_204_),
    .Y(_205_));
 sky130_fd_sc_hd__nand4_1 _543_ (.A(_117_),
    .B(_200_),
    .C(_203_),
    .D(_205_),
    .Y(_206_));
 sky130_fd_sc_hd__mux2i_1 _544_ (.A0(\mem[0][5] ),
    .A1(\mem[2][5] ),
    .S(_114_),
    .Y(_207_));
 sky130_fd_sc_hd__mux2i_1 _545_ (.A0(\mem[1][5] ),
    .A1(\mem[3][5] ),
    .S(_129_),
    .Y(_208_));
 sky130_fd_sc_hd__a22oi_1 _546_ (.A1(_118_),
    .A2(_207_),
    .B1(_208_),
    .B2(_101_),
    .Y(_209_));
 sky130_fd_sc_hd__mux2i_2 _547_ (.A0(\mem[4][5] ),
    .A1(\mem[6][5] ),
    .S(_109_),
    .Y(_210_));
 sky130_fd_sc_hd__mux2i_1 _548_ (.A0(\mem[5][5] ),
    .A1(\mem[7][5] ),
    .S(_137_),
    .Y(_211_));
 sky130_fd_sc_hd__a22oi_1 _549_ (.A1(_112_),
    .A2(_210_),
    .B1(_211_),
    .B2(_108_),
    .Y(_212_));
 sky130_fd_sc_hd__nand3_1 _550_ (.A(_127_),
    .B(_209_),
    .C(_212_),
    .Y(_213_));
 sky130_fd_sc_hd__nand3_1 _551_ (.A(_198_),
    .B(_206_),
    .C(_213_),
    .Y(_036_));
 sky130_fd_sc_hd__nand2_1 _552_ (.A(net31),
    .B(_098_),
    .Y(_214_));
 sky130_fd_sc_hd__mux2i_1 _553_ (.A0(\mem[9][6] ),
    .A1(\mem[11][6] ),
    .S(_103_),
    .Y(_215_));
 sky130_fd_sc_hd__nand2_1 _554_ (.A(_102_),
    .B(_215_),
    .Y(_216_));
 sky130_fd_sc_hd__mux2i_1 _555_ (.A0(\mem[13][6] ),
    .A1(\mem[15][6] ),
    .S(_094_),
    .Y(_217_));
 sky130_fd_sc_hd__mux2i_1 _556_ (.A0(\mem[12][6] ),
    .A1(\mem[14][6] ),
    .S(_137_),
    .Y(_218_));
 sky130_fd_sc_hd__a22oi_1 _557_ (.A1(_107_),
    .A2(_217_),
    .B1(_218_),
    .B2(_113_),
    .Y(_219_));
 sky130_fd_sc_hd__mux2i_1 _558_ (.A0(\mem[8][6] ),
    .A1(\mem[10][6] ),
    .S(_124_),
    .Y(_220_));
 sky130_fd_sc_hd__nand2_1 _559_ (.A(_119_),
    .B(_220_),
    .Y(_221_));
 sky130_fd_sc_hd__nand4_1 _560_ (.A(_117_),
    .B(_216_),
    .C(_219_),
    .D(_221_),
    .Y(_222_));
 sky130_fd_sc_hd__mux2i_1 _561_ (.A0(\mem[0][6] ),
    .A1(\mem[2][6] ),
    .S(_114_),
    .Y(_223_));
 sky130_fd_sc_hd__mux2i_1 _562_ (.A0(\mem[1][6] ),
    .A1(\mem[3][6] ),
    .S(_129_),
    .Y(_224_));
 sky130_fd_sc_hd__a22oi_1 _563_ (.A1(_118_),
    .A2(_223_),
    .B1(_224_),
    .B2(_101_),
    .Y(_225_));
 sky130_fd_sc_hd__mux2i_2 _564_ (.A0(\mem[4][6] ),
    .A1(\mem[6][6] ),
    .S(_109_),
    .Y(_226_));
 sky130_fd_sc_hd__mux2i_1 _565_ (.A0(\mem[5][6] ),
    .A1(\mem[7][6] ),
    .S(_137_),
    .Y(_227_));
 sky130_fd_sc_hd__a22oi_1 _566_ (.A1(_112_),
    .A2(_226_),
    .B1(_227_),
    .B2(_108_),
    .Y(_228_));
 sky130_fd_sc_hd__nand3_1 _567_ (.A(_127_),
    .B(_225_),
    .C(_228_),
    .Y(_229_));
 sky130_fd_sc_hd__nand3_1 _568_ (.A(_214_),
    .B(_222_),
    .C(_229_),
    .Y(_037_));
 sky130_fd_sc_hd__nand2_1 _569_ (.A(net32),
    .B(_098_),
    .Y(_230_));
 sky130_fd_sc_hd__mux2i_1 _570_ (.A0(\mem[9][7] ),
    .A1(\mem[11][7] ),
    .S(_103_),
    .Y(_231_));
 sky130_fd_sc_hd__nand2_1 _571_ (.A(_102_),
    .B(_231_),
    .Y(_232_));
 sky130_fd_sc_hd__mux2i_1 _572_ (.A0(\mem[13][7] ),
    .A1(\mem[15][7] ),
    .S(_094_),
    .Y(_233_));
 sky130_fd_sc_hd__mux2i_2 _573_ (.A0(\mem[12][7] ),
    .A1(\mem[14][7] ),
    .S(_137_),
    .Y(_234_));
 sky130_fd_sc_hd__a22oi_2 _574_ (.A1(_107_),
    .A2(_233_),
    .B1(_234_),
    .B2(_113_),
    .Y(_235_));
 sky130_fd_sc_hd__mux2i_1 _575_ (.A0(\mem[8][7] ),
    .A1(\mem[10][7] ),
    .S(_124_),
    .Y(_236_));
 sky130_fd_sc_hd__nand2_1 _576_ (.A(_119_),
    .B(_236_),
    .Y(_237_));
 sky130_fd_sc_hd__nand4_1 _577_ (.A(_117_),
    .B(_232_),
    .C(_235_),
    .D(_237_),
    .Y(_238_));
 sky130_fd_sc_hd__mux2i_1 _578_ (.A0(\mem[5][7] ),
    .A1(\mem[7][7] ),
    .S(_114_),
    .Y(_239_));
 sky130_fd_sc_hd__mux2i_1 _579_ (.A0(\mem[1][7] ),
    .A1(\mem[3][7] ),
    .S(_129_),
    .Y(_240_));
 sky130_fd_sc_hd__a22oi_1 _580_ (.A1(_108_),
    .A2(_239_),
    .B1(_240_),
    .B2(_101_),
    .Y(_241_));
 sky130_fd_sc_hd__mux2i_1 _581_ (.A0(\mem[4][7] ),
    .A1(\mem[6][7] ),
    .S(_109_),
    .Y(_242_));
 sky130_fd_sc_hd__mux2i_1 _582_ (.A0(\mem[0][7] ),
    .A1(\mem[2][7] ),
    .S(_137_),
    .Y(_243_));
 sky130_fd_sc_hd__a22oi_1 _583_ (.A1(_112_),
    .A2(_242_),
    .B1(_243_),
    .B2(_118_),
    .Y(_244_));
 sky130_fd_sc_hd__nand3_1 _584_ (.A(_127_),
    .B(_241_),
    .C(_244_),
    .Y(_245_));
 sky130_fd_sc_hd__nand3_1 _585_ (.A(_230_),
    .B(_238_),
    .C(_245_),
    .Y(_038_));
 sky130_fd_sc_hd__nor2b_1 _586_ (.A(net17),
    .B_N(net2),
    .Y(_246_));
 sky130_fd_sc_hd__clkbuf_2 _587_ (.A(_246_),
    .X(_247_));
 sky130_fd_sc_hd__xnor2_1 _588_ (.A(_029_),
    .B(_247_),
    .Y(_039_));
 sky130_fd_sc_hd__nand2_1 _589_ (.A(_030_),
    .B(_247_),
    .Y(_248_));
 sky130_fd_sc_hd__o21ai_0 _590_ (.A1(_288_),
    .A2(_247_),
    .B1(_248_),
    .Y(_040_));
 sky130_fd_sc_hd__nand2_1 _591_ (.A(_329_),
    .B(_247_),
    .Y(_249_));
 sky130_fd_sc_hd__xnor2_1 _592_ (.A(_089_),
    .B(_249_),
    .Y(_041_));
 sky130_fd_sc_hd__nand4_1 _593_ (.A(_095_),
    .B(_103_),
    .C(_089_),
    .D(_247_),
    .Y(_250_));
 sky130_fd_sc_hd__xnor2_1 _594_ (.A(_090_),
    .B(_250_),
    .Y(_042_));
 sky130_fd_sc_hd__xor2_1 _595_ (.A(_095_),
    .B(_030_),
    .X(_251_));
 sky130_fd_sc_hd__nand2_1 _596_ (.A(\rd_ptr_gray[0] ),
    .B(_098_),
    .Y(_252_));
 sky130_fd_sc_hd__o21ai_0 _597_ (.A1(_097_),
    .A2(_251_),
    .B1(_252_),
    .Y(_043_));
 sky130_fd_sc_hd__xnor2_1 _598_ (.A(_329_),
    .B(_030_),
    .Y(_253_));
 sky130_fd_sc_hd__xnor2_1 _599_ (.A(_302_),
    .B(_253_),
    .Y(_254_));
 sky130_fd_sc_hd__nand2_1 _600_ (.A(\rd_ptr_gray[1] ),
    .B(_098_),
    .Y(_255_));
 sky130_fd_sc_hd__o21ai_0 _601_ (.A1(_097_),
    .A2(_254_),
    .B1(_255_),
    .Y(_044_));
 sky130_fd_sc_hd__xnor2_1 _602_ (.A(_090_),
    .B(_329_),
    .Y(_256_));
 sky130_fd_sc_hd__o21ai_0 _603_ (.A1(_029_),
    .A2(_288_),
    .B1(_089_),
    .Y(_257_));
 sky130_fd_sc_hd__xnor2_1 _604_ (.A(_256_),
    .B(_257_),
    .Y(_258_));
 sky130_fd_sc_hd__nand2_1 _605_ (.A(\rd_ptr_gray[2] ),
    .B(_097_),
    .Y(_259_));
 sky130_fd_sc_hd__o21ai_0 _606_ (.A1(_097_),
    .A2(_258_),
    .B1(_259_),
    .Y(_045_));
 sky130_fd_sc_hd__a31oi_1 _607_ (.A1(_095_),
    .A2(_094_),
    .A3(_089_),
    .B1(_090_),
    .Y(_260_));
 sky130_fd_sc_hd__nand4b_1 _608_ (.A_N(_329_),
    .B(_090_),
    .C(_093_),
    .D(_095_),
    .Y(_261_));
 sky130_fd_sc_hd__a21bo_1 _609_ (.A1(_095_),
    .A2(_093_),
    .B1_N(_329_),
    .X(_262_));
 sky130_fd_sc_hd__a21oi_1 _610_ (.A1(_261_),
    .A2(_262_),
    .B1(_302_),
    .Y(_263_));
 sky130_fd_sc_hd__o21ai_0 _611_ (.A1(_260_),
    .A2(_263_),
    .B1(\rd_ptr_bin[4] ),
    .Y(_264_));
 sky130_fd_sc_hd__or3_1 _612_ (.A(\rd_ptr_bin[4] ),
    .B(_260_),
    .C(_263_),
    .X(_265_));
 sky130_fd_sc_hd__nor2_1 _613_ (.A(\rd_ptr_gray[3] ),
    .B(_247_),
    .Y(_266_));
 sky130_fd_sc_hd__a31oi_1 _614_ (.A1(_247_),
    .A2(_264_),
    .A3(_265_),
    .B1(_266_),
    .Y(_046_));
 sky130_fd_sc_hd__nand3_1 _615_ (.A(_089_),
    .B(_329_),
    .C(_117_),
    .Y(_267_));
 sky130_fd_sc_hd__xnor2_1 _616_ (.A(\rd_ptr_bin[4] ),
    .B(_267_),
    .Y(_047_));
 sky130_fd_sc_hd__xnor2_1 _617_ (.A(_027_),
    .B(_082_),
    .Y(_048_));
 sky130_fd_sc_hd__nand2_1 _618_ (.A(_028_),
    .B(_082_),
    .Y(_268_));
 sky130_fd_sc_hd__o21ai_0 _619_ (.A1(_317_),
    .A2(_082_),
    .B1(_268_),
    .Y(_049_));
 sky130_fd_sc_hd__xnor2_1 _620_ (.A(_075_),
    .B(_087_),
    .Y(_050_));
 sky130_fd_sc_hd__and2_0 _621_ (.A(\wr_ptr_bin[1] ),
    .B(\wr_ptr_bin[0] ),
    .X(_269_));
 sky130_fd_sc_hd__nand3_1 _622_ (.A(_075_),
    .B(_082_),
    .C(_269_),
    .Y(_270_));
 sky130_fd_sc_hd__xnor2_1 _623_ (.A(_074_),
    .B(_270_),
    .Y(_051_));
 sky130_fd_sc_hd__nand2b_2 _624_ (.A_N(net18),
    .B(net13),
    .Y(_271_));
 sky130_fd_sc_hd__xor2_1 _625_ (.A(\wr_ptr_bin[0] ),
    .B(_028_),
    .X(_272_));
 sky130_fd_sc_hd__nand2_1 _626_ (.A(\wr_ptr_gray[0] ),
    .B(_271_),
    .Y(_273_));
 sky130_fd_sc_hd__o21ai_0 _627_ (.A1(_271_),
    .A2(_272_),
    .B1(_273_),
    .Y(_052_));
 sky130_fd_sc_hd__xnor2_1 _628_ (.A(_335_),
    .B(_028_),
    .Y(_274_));
 sky130_fd_sc_hd__xnor2_1 _629_ (.A(_321_),
    .B(_274_),
    .Y(_275_));
 sky130_fd_sc_hd__nand2_1 _630_ (.A(\wr_ptr_gray[1] ),
    .B(_271_),
    .Y(_276_));
 sky130_fd_sc_hd__o21ai_0 _631_ (.A1(_271_),
    .A2(_275_),
    .B1(_276_),
    .Y(_053_));
 sky130_fd_sc_hd__xnor2_1 _632_ (.A(_074_),
    .B(_335_),
    .Y(_277_));
 sky130_fd_sc_hd__o21ai_0 _633_ (.A1(_317_),
    .A2(_027_),
    .B1(_075_),
    .Y(_278_));
 sky130_fd_sc_hd__xnor2_1 _634_ (.A(_277_),
    .B(_278_),
    .Y(_279_));
 sky130_fd_sc_hd__nand2_1 _635_ (.A(\wr_ptr_gray[2] ),
    .B(_271_),
    .Y(_280_));
 sky130_fd_sc_hd__o21ai_0 _636_ (.A1(_271_),
    .A2(_279_),
    .B1(_280_),
    .Y(_054_));
 sky130_fd_sc_hd__a21boi_0 _637_ (.A1(_075_),
    .A2(_335_),
    .B1_N(_074_),
    .Y(_281_));
 sky130_fd_sc_hd__nand4_1 _638_ (.A(_074_),
    .B(_075_),
    .C(\wr_ptr_bin[1] ),
    .D(\wr_ptr_bin[0] ),
    .Y(_282_));
 sky130_fd_sc_hd__o221ai_2 _639_ (.A1(_269_),
    .A2(_281_),
    .B1(_282_),
    .B2(_335_),
    .C1(_077_),
    .Y(_283_));
 sky130_fd_sc_hd__xnor2_1 _640_ (.A(_326_),
    .B(_283_),
    .Y(_284_));
 sky130_fd_sc_hd__nand2_1 _641_ (.A(\wr_ptr_gray[3] ),
    .B(_271_),
    .Y(_285_));
 sky130_fd_sc_hd__o21ai_0 _642_ (.A1(_271_),
    .A2(_284_),
    .B1(_285_),
    .Y(_055_));
 sky130_fd_sc_hd__xnor2_1 _643_ (.A(_326_),
    .B(_017_),
    .Y(_056_));
 sky130_fd_sc_hd__nor2b_1 _644_ (.A(_306_),
    .B_N(net21),
    .Y(_286_));
 sky130_fd_sc_hd__a2111oi_0 _645_ (.A1(_063_),
    .A2(_064_),
    .B1(_286_),
    .C1(net22),
    .D1(net24),
    .Y(net15));
 sky130_fd_sc_hd__xor2_1 _646_ (.A(_320_),
    .B(_293_),
    .X(net36));
 sky130_fd_sc_hd__nand2_1 _647_ (.A(net35),
    .B(net36),
    .Y(_287_));
 sky130_fd_sc_hd__o31ai_1 _648_ (.A1(_068_),
    .A2(_069_),
    .A3(_287_),
    .B1(_072_),
    .Y(net16));
 sky130_fd_sc_hd__fa_1 _649_ (.A(_288_),
    .B(\wr_ptr_sync[1] ),
    .CIN(_289_),
    .COUT(_290_),
    .SUM(net21));
 sky130_fd_sc_hd__fa_1 _650_ (.A(_291_),
    .B(\wr_ptr_bin[1] ),
    .CIN(_292_),
    .COUT(_293_),
    .SUM(net35));
 sky130_fd_sc_hd__ha_1 _651_ (.A(_294_),
    .B(\wr_ptr_sync[3] ),
    .COUT(_295_),
    .SUM(_296_));
 sky130_fd_sc_hd__ha_1 _652_ (.A(\rd_ptr_bin[4] ),
    .B(_297_),
    .COUT(_298_),
    .SUM(_299_));
 sky130_fd_sc_hd__ha_1 _653_ (.A(_288_),
    .B(\wr_ptr_sync[1] ),
    .COUT(_300_),
    .SUM(_301_));
 sky130_fd_sc_hd__ha_1 _654_ (.A(_302_),
    .B(\wr_ptr_sync[2] ),
    .COUT(_303_),
    .SUM(_304_));
 sky130_fd_sc_hd__ha_1 _655_ (.A(_029_),
    .B(\wr_ptr_sync[0] ),
    .COUT(_305_),
    .SUM(_306_));
 sky130_fd_sc_hd__ha_1 _656_ (.A(\rd_ptr_bin[0] ),
    .B(_307_),
    .COUT(_308_),
    .SUM(_309_));
 sky130_fd_sc_hd__ha_1 _657_ (.A(_311_),
    .B(\wr_ptr_bin[0] ),
    .COUT(_312_),
    .SUM(_313_));
 sky130_fd_sc_hd__ha_1 _658_ (.A(\rd_ptr_sync[0] ),
    .B(_027_),
    .COUT(_314_),
    .SUM(_315_));
 sky130_fd_sc_hd__ha_1 _659_ (.A(_291_),
    .B(\wr_ptr_bin[1] ),
    .COUT(_316_),
    .SUM(_310_));
 sky130_fd_sc_hd__ha_1 _660_ (.A(_318_),
    .B(\wr_ptr_bin[2] ),
    .COUT(_319_),
    .SUM(_320_));
 sky130_fd_sc_hd__ha_1 _661_ (.A(_322_),
    .B(\wr_ptr_bin[3] ),
    .COUT(_323_),
    .SUM(_324_));
 sky130_fd_sc_hd__ha_1 _662_ (.A(\rd_ptr_sync[4] ),
    .B(_326_),
    .COUT(_327_),
    .SUM(_328_));
 sky130_fd_sc_hd__ha_2 _663_ (.A(\rd_ptr_bin[0] ),
    .B(\rd_ptr_bin[1] ),
    .COUT(_329_),
    .SUM(_030_));
 sky130_fd_sc_hd__ha_2 _664_ (.A(_027_),
    .B(_317_),
    .COUT(_330_),
    .SUM(_028_));
 sky130_fd_sc_hd__ha_1 _665_ (.A(_027_),
    .B(\wr_ptr_bin[1] ),
    .COUT(_331_),
    .SUM(_332_));
 sky130_fd_sc_hd__ha_1 _666_ (.A(\wr_ptr_bin[0] ),
    .B(_317_),
    .COUT(_333_),
    .SUM(_334_));
 sky130_fd_sc_hd__ha_2 _667_ (.A(\wr_ptr_bin[0] ),
    .B(\wr_ptr_bin[1] ),
    .COUT(_335_),
    .SUM(_336_));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__dfstp_1 \empty_reg$_DFF_PN1_  (.D(_000_),
    .Q(net17),
    .SET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \full_reg$_DFF_PN0_  (.D(_001_),
    .Q(net18),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][0]$_DFFE_PP_  (.D(net5),
    .DE(_011_),
    .Q(\mem[0][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][1]$_DFFE_PP_  (.D(net6),
    .DE(_011_),
    .Q(\mem[0][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][2]$_DFFE_PP_  (.D(net7),
    .DE(_011_),
    .Q(\mem[0][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][3]$_DFFE_PP_  (.D(net8),
    .DE(_011_),
    .Q(\mem[0][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][4]$_DFFE_PP_  (.D(net9),
    .DE(_011_),
    .Q(\mem[0][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][5]$_DFFE_PP_  (.D(net10),
    .DE(_011_),
    .Q(\mem[0][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][6]$_DFFE_PP_  (.D(net11),
    .DE(_011_),
    .Q(\mem[0][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[0][7]$_DFFE_PP_  (.D(net12),
    .DE(_011_),
    .Q(\mem[0][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][0]$_DFFE_PP_  (.D(net5),
    .DE(_012_),
    .Q(\mem[10][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][1]$_DFFE_PP_  (.D(net6),
    .DE(_012_),
    .Q(\mem[10][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][2]$_DFFE_PP_  (.D(net7),
    .DE(_012_),
    .Q(\mem[10][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][3]$_DFFE_PP_  (.D(net8),
    .DE(_012_),
    .Q(\mem[10][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][4]$_DFFE_PP_  (.D(net9),
    .DE(_012_),
    .Q(\mem[10][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][5]$_DFFE_PP_  (.D(net10),
    .DE(_012_),
    .Q(\mem[10][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][6]$_DFFE_PP_  (.D(net11),
    .DE(_012_),
    .Q(\mem[10][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[10][7]$_DFFE_PP_  (.D(net12),
    .DE(_012_),
    .Q(\mem[10][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][0]$_DFFE_PP_  (.D(net5),
    .DE(_013_),
    .Q(\mem[11][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][1]$_DFFE_PP_  (.D(net6),
    .DE(_013_),
    .Q(\mem[11][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][2]$_DFFE_PP_  (.D(net7),
    .DE(_013_),
    .Q(\mem[11][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][3]$_DFFE_PP_  (.D(net8),
    .DE(_013_),
    .Q(\mem[11][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][4]$_DFFE_PP_  (.D(net9),
    .DE(_013_),
    .Q(\mem[11][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][5]$_DFFE_PP_  (.D(net10),
    .DE(_013_),
    .Q(\mem[11][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][6]$_DFFE_PP_  (.D(net11),
    .DE(_013_),
    .Q(\mem[11][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[11][7]$_DFFE_PP_  (.D(net12),
    .DE(_013_),
    .Q(\mem[11][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][0]$_DFFE_PP_  (.D(net5),
    .DE(_014_),
    .Q(\mem[12][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][1]$_DFFE_PP_  (.D(net6),
    .DE(_014_),
    .Q(\mem[12][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][2]$_DFFE_PP_  (.D(net7),
    .DE(_014_),
    .Q(\mem[12][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][3]$_DFFE_PP_  (.D(net8),
    .DE(_014_),
    .Q(\mem[12][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][4]$_DFFE_PP_  (.D(net9),
    .DE(_014_),
    .Q(\mem[12][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][5]$_DFFE_PP_  (.D(net10),
    .DE(_014_),
    .Q(\mem[12][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][6]$_DFFE_PP_  (.D(net11),
    .DE(_014_),
    .Q(\mem[12][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[12][7]$_DFFE_PP_  (.D(net12),
    .DE(_014_),
    .Q(\mem[12][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][0]$_DFFE_PP_  (.D(net5),
    .DE(_015_),
    .Q(\mem[13][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][1]$_DFFE_PP_  (.D(net6),
    .DE(_015_),
    .Q(\mem[13][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][2]$_DFFE_PP_  (.D(net7),
    .DE(_015_),
    .Q(\mem[13][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][3]$_DFFE_PP_  (.D(net8),
    .DE(_015_),
    .Q(\mem[13][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][4]$_DFFE_PP_  (.D(net9),
    .DE(_015_),
    .Q(\mem[13][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][5]$_DFFE_PP_  (.D(net10),
    .DE(_015_),
    .Q(\mem[13][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][6]$_DFFE_PP_  (.D(net11),
    .DE(_015_),
    .Q(\mem[13][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[13][7]$_DFFE_PP_  (.D(net12),
    .DE(_015_),
    .Q(\mem[13][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][0]$_DFFE_PP_  (.D(net5),
    .DE(_016_),
    .Q(\mem[14][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][1]$_DFFE_PP_  (.D(net6),
    .DE(_016_),
    .Q(\mem[14][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][2]$_DFFE_PP_  (.D(net7),
    .DE(_016_),
    .Q(\mem[14][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][3]$_DFFE_PP_  (.D(net8),
    .DE(_016_),
    .Q(\mem[14][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][4]$_DFFE_PP_  (.D(net9),
    .DE(_016_),
    .Q(\mem[14][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][5]$_DFFE_PP_  (.D(net10),
    .DE(_016_),
    .Q(\mem[14][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][6]$_DFFE_PP_  (.D(net11),
    .DE(_016_),
    .Q(\mem[14][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[14][7]$_DFFE_PP_  (.D(net12),
    .DE(_016_),
    .Q(\mem[14][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][0]$_DFFE_PP_  (.D(net5),
    .DE(_017_),
    .Q(\mem[15][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][1]$_DFFE_PP_  (.D(net6),
    .DE(_017_),
    .Q(\mem[15][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][2]$_DFFE_PP_  (.D(net7),
    .DE(_017_),
    .Q(\mem[15][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][3]$_DFFE_PP_  (.D(net8),
    .DE(_017_),
    .Q(\mem[15][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][4]$_DFFE_PP_  (.D(net9),
    .DE(_017_),
    .Q(\mem[15][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][5]$_DFFE_PP_  (.D(net10),
    .DE(_017_),
    .Q(\mem[15][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][6]$_DFFE_PP_  (.D(net11),
    .DE(_017_),
    .Q(\mem[15][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[15][7]$_DFFE_PP_  (.D(net12),
    .DE(_017_),
    .Q(\mem[15][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][0]$_DFFE_PP_  (.D(net5),
    .DE(_018_),
    .Q(\mem[1][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][1]$_DFFE_PP_  (.D(net6),
    .DE(_018_),
    .Q(\mem[1][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][2]$_DFFE_PP_  (.D(net7),
    .DE(_018_),
    .Q(\mem[1][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][3]$_DFFE_PP_  (.D(net8),
    .DE(_018_),
    .Q(\mem[1][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][4]$_DFFE_PP_  (.D(net9),
    .DE(_018_),
    .Q(\mem[1][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][5]$_DFFE_PP_  (.D(net10),
    .DE(_018_),
    .Q(\mem[1][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][6]$_DFFE_PP_  (.D(net11),
    .DE(_018_),
    .Q(\mem[1][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[1][7]$_DFFE_PP_  (.D(net12),
    .DE(_018_),
    .Q(\mem[1][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][0]$_DFFE_PP_  (.D(net5),
    .DE(_019_),
    .Q(\mem[2][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][1]$_DFFE_PP_  (.D(net6),
    .DE(_019_),
    .Q(\mem[2][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][2]$_DFFE_PP_  (.D(net7),
    .DE(_019_),
    .Q(\mem[2][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][3]$_DFFE_PP_  (.D(net8),
    .DE(_019_),
    .Q(\mem[2][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][4]$_DFFE_PP_  (.D(net9),
    .DE(_019_),
    .Q(\mem[2][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][5]$_DFFE_PP_  (.D(net10),
    .DE(_019_),
    .Q(\mem[2][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][6]$_DFFE_PP_  (.D(net11),
    .DE(_019_),
    .Q(\mem[2][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[2][7]$_DFFE_PP_  (.D(net12),
    .DE(_019_),
    .Q(\mem[2][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][0]$_DFFE_PP_  (.D(net5),
    .DE(_020_),
    .Q(\mem[3][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][1]$_DFFE_PP_  (.D(net6),
    .DE(_020_),
    .Q(\mem[3][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][2]$_DFFE_PP_  (.D(net7),
    .DE(_020_),
    .Q(\mem[3][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][3]$_DFFE_PP_  (.D(net8),
    .DE(_020_),
    .Q(\mem[3][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][4]$_DFFE_PP_  (.D(net9),
    .DE(_020_),
    .Q(\mem[3][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][5]$_DFFE_PP_  (.D(net10),
    .DE(_020_),
    .Q(\mem[3][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][6]$_DFFE_PP_  (.D(net11),
    .DE(_020_),
    .Q(\mem[3][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[3][7]$_DFFE_PP_  (.D(net12),
    .DE(_020_),
    .Q(\mem[3][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][0]$_DFFE_PP_  (.D(net5),
    .DE(_021_),
    .Q(\mem[4][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][1]$_DFFE_PP_  (.D(net6),
    .DE(_021_),
    .Q(\mem[4][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][2]$_DFFE_PP_  (.D(net7),
    .DE(_021_),
    .Q(\mem[4][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][3]$_DFFE_PP_  (.D(net8),
    .DE(_021_),
    .Q(\mem[4][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][4]$_DFFE_PP_  (.D(net9),
    .DE(_021_),
    .Q(\mem[4][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][5]$_DFFE_PP_  (.D(net10),
    .DE(_021_),
    .Q(\mem[4][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][6]$_DFFE_PP_  (.D(net11),
    .DE(_021_),
    .Q(\mem[4][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[4][7]$_DFFE_PP_  (.D(net12),
    .DE(_021_),
    .Q(\mem[4][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][0]$_DFFE_PP_  (.D(net5),
    .DE(_022_),
    .Q(\mem[5][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][1]$_DFFE_PP_  (.D(net6),
    .DE(_022_),
    .Q(\mem[5][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][2]$_DFFE_PP_  (.D(net7),
    .DE(_022_),
    .Q(\mem[5][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][3]$_DFFE_PP_  (.D(net8),
    .DE(_022_),
    .Q(\mem[5][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][4]$_DFFE_PP_  (.D(net9),
    .DE(_022_),
    .Q(\mem[5][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][5]$_DFFE_PP_  (.D(net10),
    .DE(_022_),
    .Q(\mem[5][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][6]$_DFFE_PP_  (.D(net11),
    .DE(_022_),
    .Q(\mem[5][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[5][7]$_DFFE_PP_  (.D(net12),
    .DE(_022_),
    .Q(\mem[5][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][0]$_DFFE_PP_  (.D(net5),
    .DE(_023_),
    .Q(\mem[6][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][1]$_DFFE_PP_  (.D(net6),
    .DE(_023_),
    .Q(\mem[6][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][2]$_DFFE_PP_  (.D(net7),
    .DE(_023_),
    .Q(\mem[6][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][3]$_DFFE_PP_  (.D(net8),
    .DE(_023_),
    .Q(\mem[6][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][4]$_DFFE_PP_  (.D(net9),
    .DE(_023_),
    .Q(\mem[6][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][5]$_DFFE_PP_  (.D(net10),
    .DE(_023_),
    .Q(\mem[6][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][6]$_DFFE_PP_  (.D(net11),
    .DE(_023_),
    .Q(\mem[6][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[6][7]$_DFFE_PP_  (.D(net12),
    .DE(_023_),
    .Q(\mem[6][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][0]$_DFFE_PP_  (.D(net5),
    .DE(_024_),
    .Q(\mem[7][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][1]$_DFFE_PP_  (.D(net6),
    .DE(_024_),
    .Q(\mem[7][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][2]$_DFFE_PP_  (.D(net7),
    .DE(_024_),
    .Q(\mem[7][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][3]$_DFFE_PP_  (.D(net8),
    .DE(_024_),
    .Q(\mem[7][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][4]$_DFFE_PP_  (.D(net9),
    .DE(_024_),
    .Q(\mem[7][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][5]$_DFFE_PP_  (.D(net10),
    .DE(_024_),
    .Q(\mem[7][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][6]$_DFFE_PP_  (.D(net11),
    .DE(_024_),
    .Q(\mem[7][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[7][7]$_DFFE_PP_  (.D(net12),
    .DE(_024_),
    .Q(\mem[7][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][0]$_DFFE_PP_  (.D(net5),
    .DE(_025_),
    .Q(\mem[8][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][1]$_DFFE_PP_  (.D(net6),
    .DE(_025_),
    .Q(\mem[8][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][2]$_DFFE_PP_  (.D(net7),
    .DE(_025_),
    .Q(\mem[8][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][3]$_DFFE_PP_  (.D(net8),
    .DE(_025_),
    .Q(\mem[8][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][4]$_DFFE_PP_  (.D(net9),
    .DE(_025_),
    .Q(\mem[8][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][5]$_DFFE_PP_  (.D(net10),
    .DE(_025_),
    .Q(\mem[8][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][6]$_DFFE_PP_  (.D(net11),
    .DE(_025_),
    .Q(\mem[8][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[8][7]$_DFFE_PP_  (.D(net12),
    .DE(_025_),
    .Q(\mem[8][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][0]$_DFFE_PP_  (.D(net5),
    .DE(_026_),
    .Q(\mem[9][0] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][1]$_DFFE_PP_  (.D(net6),
    .DE(_026_),
    .Q(\mem[9][1] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][2]$_DFFE_PP_  (.D(net7),
    .DE(_026_),
    .Q(\mem[9][2] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][3]$_DFFE_PP_  (.D(net8),
    .DE(_026_),
    .Q(\mem[9][3] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][4]$_DFFE_PP_  (.D(net9),
    .DE(_026_),
    .Q(\mem[9][4] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][5]$_DFFE_PP_  (.D(net10),
    .DE(_026_),
    .Q(\mem[9][5] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][6]$_DFFE_PP_  (.D(net11),
    .DE(_026_),
    .Q(\mem[9][6] ),
    .CLK(net4));
 sky130_fd_sc_hd__edfxtp_1 \mem[9][7]$_DFFE_PP_  (.D(net12),
    .DE(_026_),
    .Q(\mem[9][7] ),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \pointer_wraparound_error$_DFF_PN0_  (.D(_010_),
    .Q(net19),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[0]$_DFFE_PN0P_  (.D(_031_),
    .Q(net25),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[1]$_DFFE_PN0P_  (.D(_032_),
    .Q(net26),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[2]$_DFFE_PN0P_  (.D(_033_),
    .Q(net27),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[3]$_DFFE_PN0P_  (.D(_034_),
    .Q(net28),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[4]$_DFFE_PN0P_  (.D(_035_),
    .Q(net29),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[5]$_DFFE_PN0P_  (.D(_036_),
    .Q(net30),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[6]$_DFFE_PN0P_  (.D(_037_),
    .Q(net31),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_data_reg[7]$_DFFE_PN0P_  (.D(_038_),
    .Q(net32),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_bin[0]$_DFFE_PN0P_  (.D(_039_),
    .Q(\rd_ptr_bin[0] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_bin[1]$_DFFE_PN0P_  (.D(_040_),
    .Q(\rd_ptr_bin[1] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_bin[2]$_DFFE_PN0P_  (.D(_041_),
    .Q(\rd_ptr_bin[2] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_bin[3]$_DFFE_PN0P_  (.D(_042_),
    .Q(\rd_ptr_bin[3] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray[0]$_DFFE_PN0P_  (.D(_043_),
    .Q(\rd_ptr_gray[0] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray[1]$_DFFE_PN0P_  (.D(_044_),
    .Q(\rd_ptr_gray[1] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray[2]$_DFFE_PN0P_  (.D(_045_),
    .Q(\rd_ptr_gray[2] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray[3]$_DFFE_PN0P_  (.D(_046_),
    .Q(\rd_ptr_gray[3] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_4 \rd_ptr_gray[4]$_DFFE_PN0P_  (.D(_047_),
    .Q(\rd_ptr_bin[4] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync1[0]$_DFF_PN0_  (.D(\rd_ptr_gray[0] ),
    .Q(\rd_ptr_gray_sync1[0] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync1[1]$_DFF_PN0_  (.D(\rd_ptr_gray[1] ),
    .Q(\rd_ptr_gray_sync1[1] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync1[2]$_DFF_PN0_  (.D(\rd_ptr_gray[2] ),
    .Q(\rd_ptr_gray_sync1[2] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync1[3]$_DFF_PN0_  (.D(\rd_ptr_gray[3] ),
    .Q(\rd_ptr_gray_sync1[3] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync1[4]$_DFF_PN0_  (.D(\rd_ptr_bin[4] ),
    .Q(\rd_ptr_gray_sync1[4] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync2[0]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[0] ),
    .Q(\rd_ptr_gray_sync2[0] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync2[1]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[1] ),
    .Q(\rd_ptr_gray_sync2[1] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync2[2]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[2] ),
    .Q(\rd_ptr_gray_sync2[2] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync2[3]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[3] ),
    .Q(\rd_ptr_gray_sync2[3] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_gray_sync2[4]$_DFF_PN0_  (.D(\rd_ptr_gray_sync1[4] ),
    .Q(\rd_ptr_gray_sync2[4] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_sync[0]$_DFF_PN0_  (.D(_006_),
    .Q(\rd_ptr_sync[0] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_sync[1]$_DFF_PN0_  (.D(_007_),
    .Q(\rd_ptr_sync[1] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_sync[2]$_DFF_PN0_  (.D(_008_),
    .Q(\rd_ptr_sync[2] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_sync[3]$_DFF_PN0_  (.D(_009_),
    .Q(\rd_ptr_sync[3] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \rd_ptr_sync[4]$_DFF_PN0_  (.D(\rd_ptr_gray_sync2[4] ),
    .Q(\rd_ptr_sync[4] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \sync_error$_DFF_PN0_  (.D(net39),
    .Q(net33),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_4 \wr_ptr_bin[0]$_DFFE_PN0P_  (.D(_048_),
    .Q(\wr_ptr_bin[0] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_4 \wr_ptr_bin[1]$_DFFE_PN0P_  (.D(_049_),
    .Q(\wr_ptr_bin[1] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_bin[2]$_DFFE_PN0P_  (.D(_050_),
    .Q(\wr_ptr_bin[2] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_bin[3]$_DFFE_PN0P_  (.D(_051_),
    .Q(\wr_ptr_bin[3] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray[0]$_DFFE_PN0P_  (.D(_052_),
    .Q(\wr_ptr_gray[0] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray[1]$_DFFE_PN0P_  (.D(_053_),
    .Q(\wr_ptr_gray[1] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray[2]$_DFFE_PN0P_  (.D(_054_),
    .Q(\wr_ptr_gray[2] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray[3]$_DFFE_PN0P_  (.D(_055_),
    .Q(\wr_ptr_gray[3] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray[4]$_DFFE_PN0P_  (.D(_056_),
    .Q(\wr_ptr_bin[4] ),
    .RESET_B(net14),
    .CLK(net4));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync1[0]$_DFF_PN0_  (.D(\wr_ptr_gray[0] ),
    .Q(\wr_ptr_gray_sync1[0] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync1[1]$_DFF_PN0_  (.D(\wr_ptr_gray[1] ),
    .Q(\wr_ptr_gray_sync1[1] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync1[2]$_DFF_PN0_  (.D(\wr_ptr_gray[2] ),
    .Q(\wr_ptr_gray_sync1[2] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync1[3]$_DFF_PN0_  (.D(\wr_ptr_gray[3] ),
    .Q(\wr_ptr_gray_sync1[3] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync1[4]$_DFF_PN0_  (.D(\wr_ptr_bin[4] ),
    .Q(\wr_ptr_gray_sync1[4] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync2[0]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[0] ),
    .Q(\wr_ptr_gray_sync2[0] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync2[1]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[1] ),
    .Q(\wr_ptr_gray_sync2[1] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync2[2]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[2] ),
    .Q(\wr_ptr_gray_sync2[2] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync2[3]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[3] ),
    .Q(\wr_ptr_gray_sync2[3] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_gray_sync2[4]$_DFF_PN0_  (.D(\wr_ptr_gray_sync1[4] ),
    .Q(\wr_ptr_gray_sync2[4] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_sync[0]$_DFF_PN0_  (.D(_002_),
    .Q(\wr_ptr_sync[0] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_sync[1]$_DFF_PN0_  (.D(_003_),
    .Q(\wr_ptr_sync[1] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_sync[2]$_DFF_PN0_  (.D(_004_),
    .Q(\wr_ptr_sync[2] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_sync[3]$_DFF_PN0_  (.D(_005_),
    .Q(\wr_ptr_sync[3] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__dfrtp_1 \wr_ptr_sync[4]$_DFF_PN0_  (.D(\wr_ptr_gray_sync2[4] ),
    .Q(\wr_ptr_sync[4] ),
    .RESET_B(net3),
    .CLK(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_329 ();
 sky130_fd_sc_hd__buf_8 input1 (.A(rd_clk),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(rd_en),
    .X(net2));
 sky130_fd_sc_hd__buf_12 input3 (.A(rd_rst_n),
    .X(net3));
 sky130_fd_sc_hd__buf_16 input4 (.A(wr_clk),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(wr_data[0]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input6 (.A(wr_data[1]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input7 (.A(wr_data[2]),
    .X(net7));
 sky130_fd_sc_hd__buf_6 input8 (.A(wr_data[3]),
    .X(net8));
 sky130_fd_sc_hd__buf_6 input9 (.A(wr_data[4]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_8 input10 (.A(wr_data[5]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_8 input11 (.A(wr_data[6]),
    .X(net11));
 sky130_fd_sc_hd__buf_6 input12 (.A(wr_data[7]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(wr_en),
    .X(net13));
 sky130_fd_sc_hd__buf_16 input14 (.A(wr_rst_n),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 output15 (.A(net15),
    .X(almost_empty));
 sky130_fd_sc_hd__clkbuf_1 output16 (.A(net16),
    .X(almost_full));
 sky130_fd_sc_hd__clkbuf_1 output17 (.A(net17),
    .X(empty));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net18),
    .X(full));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net19),
    .X(pointer_wraparound_flag));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net20),
    .X(rd_count[0]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net21),
    .X(rd_count[1]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net22),
    .X(rd_count[2]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net23),
    .X(rd_count[3]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net24),
    .X(rd_count[4]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net25),
    .X(rd_data[0]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net26),
    .X(rd_data[1]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net27),
    .X(rd_data[2]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net28),
    .X(rd_data[3]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net29),
    .X(rd_data[4]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net30),
    .X(rd_data[5]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net31),
    .X(rd_data[6]));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(net32),
    .X(rd_data[7]));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net33),
    .X(sync_error_flag));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net34),
    .X(wr_count[0]));
 sky130_fd_sc_hd__clkbuf_1 output35 (.A(net35),
    .X(wr_count[1]));
 sky130_fd_sc_hd__clkbuf_1 output36 (.A(net36),
    .X(wr_count[2]));
 sky130_fd_sc_hd__clkbuf_1 output37 (.A(net37),
    .X(wr_count[3]));
 sky130_fd_sc_hd__clkbuf_1 output38 (.A(net38),
    .X(wr_count[4]));
 sky130_fd_sc_hd__conb_1 \sync_error$_DFF_PN0__39  (.HI(net39));
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_226 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_234 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_210 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_261 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_242 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_224 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_164 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_92 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_100 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_140 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_195 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_336 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_78 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_102 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_67 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_67 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_75 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_162 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_48 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_64 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_72 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_291 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_212 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_20 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_103 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_11 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_192 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_231 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_244 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_252 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_345 ();
endmodule
