module pulse_width_detector (clk,
    pulse_detected,
    rst,
    signal_in,
    threshold);
 input clk;
 output pulse_detected;
 input rst;
 input signal_in;
 input [7:0] threshold;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire signal_prev;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire net12;

 INV_X4 _089_ (.A(net1),
    .ZN(_000_));
 INV_X1 _090_ (.A(net3),
    .ZN(_084_));
 BUF_X4 _091_ (.A(net2),
    .Z(_013_));
 NOR2_X2 _092_ (.A1(_013_),
    .A2(signal_prev),
    .ZN(_014_));
 NAND2_X1 _093_ (.A1(\counter[0] ),
    .A2(_014_),
    .ZN(_015_));
 NAND2_X2 _094_ (.A1(_013_),
    .A2(signal_prev),
    .ZN(_016_));
 AND3_X1 _095_ (.A1(\counter[3] ),
    .A2(\counter[2] ),
    .A3(_087_),
    .ZN(_017_));
 BUF_X2 _096_ (.A(\counter[4] ),
    .Z(_018_));
 AND4_X1 _097_ (.A1(\counter[5] ),
    .A2(_018_),
    .A3(\counter[6] ),
    .A4(\counter[7] ),
    .ZN(_019_));
 AND2_X1 _098_ (.A1(_017_),
    .A2(_019_),
    .ZN(_020_));
 XOR2_X1 _099_ (.A(\counter[0] ),
    .B(_020_),
    .Z(_021_));
 OAI21_X1 _100_ (.A(_015_),
    .B1(_016_),
    .B2(_021_),
    .ZN(_001_));
 MUX2_X1 _101_ (.A(_088_),
    .B(\counter[1] ),
    .S(_020_),
    .Z(_022_));
 AND2_X1 _102_ (.A1(_013_),
    .A2(signal_prev),
    .ZN(_023_));
 AOI22_X1 _103_ (.A1(\counter[1] ),
    .A2(_014_),
    .B1(_022_),
    .B2(_023_),
    .ZN(_024_));
 INV_X1 _104_ (.A(_024_),
    .ZN(_002_));
 XOR2_X2 _105_ (.A(_013_),
    .B(signal_prev),
    .Z(_025_));
 NAND3_X1 _106_ (.A1(_013_),
    .A2(\counter[2] ),
    .A3(_087_),
    .ZN(_026_));
 NOR2_X1 _107_ (.A1(_020_),
    .A2(_026_),
    .ZN(_027_));
 AOI21_X1 _108_ (.A(\counter[2] ),
    .B1(_087_),
    .B2(_013_),
    .ZN(_028_));
 NOR3_X1 _109_ (.A1(_025_),
    .A2(_027_),
    .A3(_028_),
    .ZN(_003_));
 NAND3_X1 _110_ (.A1(\counter[2] ),
    .A2(\counter[0] ),
    .A3(\counter[1] ),
    .ZN(_029_));
 NAND2_X1 _111_ (.A1(_013_),
    .A2(\counter[3] ),
    .ZN(_030_));
 AOI211_X2 _112_ (.A(_029_),
    .B(_030_),
    .C1(_017_),
    .C2(_019_),
    .ZN(_031_));
 INV_X1 _113_ (.A(\counter[3] ),
    .ZN(_032_));
 AOI21_X1 _114_ (.A(_016_),
    .B1(_029_),
    .B2(_032_),
    .ZN(_033_));
 AOI21_X1 _115_ (.A(_033_),
    .B1(_014_),
    .B2(\counter[3] ),
    .ZN(_034_));
 NOR2_X1 _116_ (.A1(_031_),
    .A2(_034_),
    .ZN(_004_));
 NAND2_X1 _117_ (.A1(_018_),
    .A2(_014_),
    .ZN(_035_));
 OR2_X1 _118_ (.A1(_018_),
    .A2(_017_),
    .ZN(_036_));
 NAND2_X1 _119_ (.A1(_018_),
    .A2(_017_),
    .ZN(_037_));
 OAI21_X1 _120_ (.A(_036_),
    .B1(_037_),
    .B2(_019_),
    .ZN(_038_));
 OAI21_X1 _121_ (.A(_035_),
    .B1(_038_),
    .B2(_016_),
    .ZN(_005_));
 NAND2_X1 _122_ (.A1(_018_),
    .A2(_031_),
    .ZN(_039_));
 XOR2_X1 _123_ (.A(\counter[5] ),
    .B(_039_),
    .Z(_040_));
 NOR2_X1 _124_ (.A1(_025_),
    .A2(_040_),
    .ZN(_006_));
 NAND2_X1 _125_ (.A1(\counter[6] ),
    .A2(_014_),
    .ZN(_041_));
 NAND3_X1 _126_ (.A1(\counter[5] ),
    .A2(_018_),
    .A3(_017_),
    .ZN(_042_));
 NOR2_X1 _127_ (.A1(\counter[7] ),
    .A2(_042_),
    .ZN(_043_));
 MUX2_X1 _128_ (.A(_042_),
    .B(_043_),
    .S(\counter[6] ),
    .Z(_044_));
 OAI21_X1 _129_ (.A(_041_),
    .B1(_044_),
    .B2(_016_),
    .ZN(_007_));
 NAND4_X1 _130_ (.A1(\counter[5] ),
    .A2(_018_),
    .A3(\counter[6] ),
    .A4(_031_),
    .ZN(_045_));
 XOR2_X1 _131_ (.A(\counter[7] ),
    .B(_045_),
    .Z(_046_));
 NOR2_X1 _132_ (.A1(_025_),
    .A2(_046_),
    .ZN(_008_));
 INV_X1 _133_ (.A(net11),
    .ZN(_047_));
 NAND4_X1 _134_ (.A1(_065_),
    .A2(_068_),
    .A3(_071_),
    .A4(_074_),
    .ZN(_048_));
 NAND4_X1 _135_ (.A1(_077_),
    .A2(_080_),
    .A3(_083_),
    .A4(_086_),
    .ZN(_049_));
 OAI21_X1 _136_ (.A(_047_),
    .B1(_048_),
    .B2(_049_),
    .ZN(_050_));
 AOI22_X1 _137_ (.A1(net11),
    .A2(_014_),
    .B1(_050_),
    .B2(_023_),
    .ZN(_051_));
 INV_X1 _138_ (.A(_082_),
    .ZN(_052_));
 INV_X1 _139_ (.A(_083_),
    .ZN(_053_));
 OAI21_X1 _140_ (.A(_052_),
    .B1(_085_),
    .B2(_053_),
    .ZN(_054_));
 NAND3_X1 _141_ (.A1(_077_),
    .A2(_080_),
    .A3(_054_),
    .ZN(_055_));
 AOI21_X1 _142_ (.A(_076_),
    .B1(_079_),
    .B2(_077_),
    .ZN(_056_));
 AOI21_X1 _143_ (.A(_048_),
    .B1(_055_),
    .B2(_056_),
    .ZN(_057_));
 INV_X1 _144_ (.A(_065_),
    .ZN(_058_));
 NAND3_X1 _145_ (.A1(_073_),
    .A2(_068_),
    .A3(_071_),
    .ZN(_059_));
 AOI21_X1 _146_ (.A(_067_),
    .B1(_070_),
    .B2(_068_),
    .ZN(_010_));
 AOI21_X1 _147_ (.A(_058_),
    .B1(_059_),
    .B2(_010_),
    .ZN(_011_));
 OR3_X1 _148_ (.A1(_064_),
    .A2(_016_),
    .A3(_011_),
    .ZN(_012_));
 OAI21_X1 _149_ (.A(_051_),
    .B1(_057_),
    .B2(_012_),
    .ZN(_009_));
 HA_X1 _150_ (.A(_063_),
    .B(net10),
    .CO(_064_),
    .S(_065_));
 HA_X1 _151_ (.A(_066_),
    .B(net9),
    .CO(_067_),
    .S(_068_));
 HA_X1 _152_ (.A(_069_),
    .B(net8),
    .CO(_070_),
    .S(_071_));
 HA_X1 _153_ (.A(_072_),
    .B(net7),
    .CO(_073_),
    .S(_074_));
 HA_X1 _154_ (.A(_075_),
    .B(net6),
    .CO(_076_),
    .S(_077_));
 HA_X1 _155_ (.A(_078_),
    .B(net5),
    .CO(_079_),
    .S(_080_));
 HA_X1 _156_ (.A(_081_),
    .B(net4),
    .CO(_082_),
    .S(_083_));
 HA_X1 _157_ (.A(\counter[0] ),
    .B(_084_),
    .CO(_085_),
    .S(_086_));
 HA_X1 _158_ (.A(\counter[0] ),
    .B(\counter[1] ),
    .CO(_087_),
    .S(_088_));
 DFFR_X2 \counter[0]$_DFFE_PP0P_  (.D(_001_),
    .RN(_000_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\counter[0] ),
    .QN(_062_));
 DFFR_X1 \counter[1]$_DFFE_PP0P_  (.D(_002_),
    .RN(_000_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[1] ),
    .QN(_081_));
 DFFR_X1 \counter[2]$_DFFE_PP0P_  (.D(_003_),
    .RN(_000_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[2] ),
    .QN(_078_));
 DFFR_X1 \counter[3]$_DFFE_PP0P_  (.D(_004_),
    .RN(_000_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[3] ),
    .QN(_075_));
 DFFR_X1 \counter[4]$_DFFE_PP0P_  (.D(_005_),
    .RN(_000_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[4] ),
    .QN(_072_));
 DFFR_X1 \counter[5]$_DFFE_PP0P_  (.D(_006_),
    .RN(_000_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\counter[5] ),
    .QN(_069_));
 DFFR_X1 \counter[6]$_DFFE_PP0P_  (.D(_007_),
    .RN(_000_),
    .CK(clknet_1_1__leaf_clk),
    .Q(\counter[6] ),
    .QN(_066_));
 DFFR_X1 \counter[7]$_DFFE_PP0P_  (.D(_008_),
    .RN(_000_),
    .CK(clknet_1_0__leaf_clk),
    .Q(\counter[7] ),
    .QN(_063_));
 DFFR_X1 \pulse_detected$_DFFE_PP0P_  (.D(_009_),
    .RN(_000_),
    .CK(clknet_1_1__leaf_clk),
    .Q(net11),
    .QN(_061_));
 DFFR_X2 \signal_prev$_DFF_PP0_  (.D(net2),
    .RN(_000_),
    .CK(clknet_1_0__leaf_clk),
    .Q(signal_prev),
    .QN(_060_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_51 ();
 BUF_X1 input1 (.A(net12),
    .Z(net1));
 BUF_X1 input2 (.A(signal_in),
    .Z(net2));
 BUF_X1 input3 (.A(threshold[0]),
    .Z(net3));
 BUF_X1 input4 (.A(threshold[1]),
    .Z(net4));
 BUF_X1 input5 (.A(threshold[2]),
    .Z(net5));
 BUF_X1 input6 (.A(threshold[3]),
    .Z(net6));
 BUF_X1 input7 (.A(threshold[4]),
    .Z(net7));
 BUF_X1 input8 (.A(threshold[5]),
    .Z(net8));
 BUF_X1 input9 (.A(threshold[6]),
    .Z(net9));
 BUF_X1 input10 (.A(threshold[7]),
    .Z(net10));
 BUF_X1 output11 (.A(net11),
    .Z(pulse_detected));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_0__leaf_clk));
 CLKBUF_X3 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_1_1__leaf_clk));
 INV_X1 clkload0 (.A(clknet_1_0__leaf_clk));
 CLKBUF_X1 hold1 (.A(rst),
    .Z(net12));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X1 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_136 ();
 FILLCELL_X16 FILLER_0_168 ();
 FILLCELL_X8 FILLER_0_184 ();
 FILLCELL_X4 FILLER_0_192 ();
 FILLCELL_X2 FILLER_0_196 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X4 FILLER_1_193 ();
 FILLCELL_X1 FILLER_1_197 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X4 FILLER_2_129 ();
 FILLCELL_X2 FILLER_2_133 ();
 FILLCELL_X32 FILLER_2_137 ();
 FILLCELL_X16 FILLER_2_169 ();
 FILLCELL_X8 FILLER_2_185 ();
 FILLCELL_X4 FILLER_2_193 ();
 FILLCELL_X1 FILLER_2_197 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X4 FILLER_3_193 ();
 FILLCELL_X1 FILLER_3_197 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X4 FILLER_4_193 ();
 FILLCELL_X1 FILLER_4_197 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X4 FILLER_5_193 ();
 FILLCELL_X1 FILLER_5_197 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X4 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_155 ();
 FILLCELL_X8 FILLER_6_187 ();
 FILLCELL_X2 FILLER_6_195 ();
 FILLCELL_X1 FILLER_6_197 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X8 FILLER_7_65 ();
 FILLCELL_X4 FILLER_7_73 ();
 FILLCELL_X4 FILLER_7_99 ();
 FILLCELL_X1 FILLER_7_103 ();
 FILLCELL_X2 FILLER_7_107 ();
 FILLCELL_X16 FILLER_7_131 ();
 FILLCELL_X2 FILLER_7_147 ();
 FILLCELL_X32 FILLER_7_155 ();
 FILLCELL_X8 FILLER_7_187 ();
 FILLCELL_X2 FILLER_7_195 ();
 FILLCELL_X1 FILLER_7_197 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X16 FILLER_8_65 ();
 FILLCELL_X8 FILLER_8_81 ();
 FILLCELL_X4 FILLER_8_89 ();
 FILLCELL_X2 FILLER_8_93 ();
 FILLCELL_X1 FILLER_8_95 ();
 FILLCELL_X2 FILLER_8_124 ();
 FILLCELL_X2 FILLER_8_130 ();
 FILLCELL_X4 FILLER_8_152 ();
 FILLCELL_X2 FILLER_8_161 ();
 FILLCELL_X2 FILLER_8_167 ();
 FILLCELL_X1 FILLER_8_169 ();
 FILLCELL_X2 FILLER_8_184 ();
 FILLCELL_X8 FILLER_8_189 ();
 FILLCELL_X1 FILLER_8_197 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X2 FILLER_9_97 ();
 FILLCELL_X4 FILLER_9_103 ();
 FILLCELL_X1 FILLER_9_107 ();
 FILLCELL_X32 FILLER_9_116 ();
 FILLCELL_X8 FILLER_9_148 ();
 FILLCELL_X4 FILLER_9_156 ();
 FILLCELL_X1 FILLER_9_175 ();
 FILLCELL_X2 FILLER_9_186 ();
 FILLCELL_X1 FILLER_9_188 ();
 FILLCELL_X4 FILLER_9_192 ();
 FILLCELL_X2 FILLER_9_196 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X8 FILLER_10_65 ();
 FILLCELL_X4 FILLER_10_73 ();
 FILLCELL_X1 FILLER_10_77 ();
 FILLCELL_X16 FILLER_10_85 ();
 FILLCELL_X2 FILLER_10_101 ();
 FILLCELL_X1 FILLER_10_103 ();
 FILLCELL_X1 FILLER_10_109 ();
 FILLCELL_X2 FILLER_10_117 ();
 FILLCELL_X2 FILLER_10_144 ();
 FILLCELL_X1 FILLER_10_146 ();
 FILLCELL_X8 FILLER_10_171 ();
 FILLCELL_X4 FILLER_10_179 ();
 FILLCELL_X1 FILLER_10_183 ();
 FILLCELL_X8 FILLER_10_187 ();
 FILLCELL_X2 FILLER_10_195 ();
 FILLCELL_X1 FILLER_10_197 ();
 FILLCELL_X8 FILLER_11_1 ();
 FILLCELL_X1 FILLER_11_9 ();
 FILLCELL_X32 FILLER_11_13 ();
 FILLCELL_X16 FILLER_11_45 ();
 FILLCELL_X8 FILLER_11_61 ();
 FILLCELL_X2 FILLER_11_69 ();
 FILLCELL_X1 FILLER_11_71 ();
 FILLCELL_X2 FILLER_11_108 ();
 FILLCELL_X1 FILLER_11_110 ();
 FILLCELL_X1 FILLER_11_118 ();
 FILLCELL_X1 FILLER_11_122 ();
 FILLCELL_X4 FILLER_11_133 ();
 FILLCELL_X1 FILLER_11_137 ();
 FILLCELL_X32 FILLER_11_143 ();
 FILLCELL_X16 FILLER_11_175 ();
 FILLCELL_X4 FILLER_11_191 ();
 FILLCELL_X2 FILLER_11_195 ();
 FILLCELL_X1 FILLER_11_197 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X16 FILLER_12_97 ();
 FILLCELL_X4 FILLER_12_113 ();
 FILLCELL_X32 FILLER_12_130 ();
 FILLCELL_X32 FILLER_12_162 ();
 FILLCELL_X4 FILLER_12_194 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X8 FILLER_13_65 ();
 FILLCELL_X4 FILLER_13_73 ();
 FILLCELL_X2 FILLER_13_77 ();
 FILLCELL_X1 FILLER_13_79 ();
 FILLCELL_X16 FILLER_13_87 ();
 FILLCELL_X8 FILLER_13_103 ();
 FILLCELL_X32 FILLER_13_116 ();
 FILLCELL_X32 FILLER_13_148 ();
 FILLCELL_X16 FILLER_13_180 ();
 FILLCELL_X2 FILLER_13_196 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X16 FILLER_14_97 ();
 FILLCELL_X4 FILLER_14_113 ();
 FILLCELL_X2 FILLER_14_117 ();
 FILLCELL_X1 FILLER_14_119 ();
 FILLCELL_X8 FILLER_14_123 ();
 FILLCELL_X4 FILLER_14_131 ();
 FILLCELL_X2 FILLER_14_135 ();
 FILLCELL_X1 FILLER_14_140 ();
 FILLCELL_X32 FILLER_14_147 ();
 FILLCELL_X16 FILLER_14_179 ();
 FILLCELL_X2 FILLER_14_195 ();
 FILLCELL_X1 FILLER_14_197 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X2 FILLER_15_97 ();
 FILLCELL_X1 FILLER_15_99 ();
 FILLCELL_X4 FILLER_15_103 ();
 FILLCELL_X4 FILLER_15_113 ();
 FILLCELL_X2 FILLER_15_117 ();
 FILLCELL_X2 FILLER_15_170 ();
 FILLCELL_X1 FILLER_15_175 ();
 FILLCELL_X1 FILLER_15_183 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X16 FILLER_16_65 ();
 FILLCELL_X2 FILLER_16_81 ();
 FILLCELL_X4 FILLER_16_103 ();
 FILLCELL_X2 FILLER_16_107 ();
 FILLCELL_X4 FILLER_16_112 ();
 FILLCELL_X2 FILLER_16_116 ();
 FILLCELL_X1 FILLER_16_118 ();
 FILLCELL_X4 FILLER_16_135 ();
 FILLCELL_X1 FILLER_16_139 ();
 FILLCELL_X2 FILLER_16_174 ();
 FILLCELL_X2 FILLER_16_196 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X8 FILLER_17_97 ();
 FILLCELL_X2 FILLER_17_105 ();
 FILLCELL_X32 FILLER_17_127 ();
 FILLCELL_X16 FILLER_17_159 ();
 FILLCELL_X1 FILLER_17_175 ();
 FILLCELL_X2 FILLER_17_196 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X32 FILLER_18_129 ();
 FILLCELL_X8 FILLER_18_161 ();
 FILLCELL_X4 FILLER_18_169 ();
 FILLCELL_X2 FILLER_18_173 ();
 FILLCELL_X1 FILLER_18_175 ();
 FILLCELL_X2 FILLER_18_186 ();
 FILLCELL_X1 FILLER_18_188 ();
 FILLCELL_X4 FILLER_18_192 ();
 FILLCELL_X2 FILLER_18_196 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X32 FILLER_19_97 ();
 FILLCELL_X32 FILLER_19_129 ();
 FILLCELL_X32 FILLER_19_161 ();
 FILLCELL_X4 FILLER_19_193 ();
 FILLCELL_X1 FILLER_19_197 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X32 FILLER_20_97 ();
 FILLCELL_X32 FILLER_20_129 ();
 FILLCELL_X32 FILLER_20_161 ();
 FILLCELL_X4 FILLER_20_193 ();
 FILLCELL_X1 FILLER_20_197 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X32 FILLER_21_97 ();
 FILLCELL_X32 FILLER_21_129 ();
 FILLCELL_X32 FILLER_21_161 ();
 FILLCELL_X4 FILLER_21_193 ();
 FILLCELL_X1 FILLER_21_197 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X32 FILLER_22_97 ();
 FILLCELL_X32 FILLER_22_129 ();
 FILLCELL_X32 FILLER_22_161 ();
 FILLCELL_X4 FILLER_22_193 ();
 FILLCELL_X1 FILLER_22_197 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X4 FILLER_23_193 ();
 FILLCELL_X1 FILLER_23_197 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X32 FILLER_24_129 ();
 FILLCELL_X32 FILLER_24_161 ();
 FILLCELL_X4 FILLER_24_193 ();
 FILLCELL_X1 FILLER_24_197 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X32 FILLER_25_129 ();
 FILLCELL_X32 FILLER_25_161 ();
 FILLCELL_X4 FILLER_25_193 ();
 FILLCELL_X1 FILLER_25_197 ();
endmodule
