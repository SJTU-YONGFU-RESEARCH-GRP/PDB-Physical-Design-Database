module radix4_booth_multiplier (clk,
    done,
    rst_n,
    start,
    multiplicand,
    multiplier,
    product);
 input clk;
 output done;
 input rst_n;
 input start;
 input [7:0] multiplicand;
 input [7:0] multiplier;
 output [15:0] product;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire \a_reg[0] ;
 wire \a_reg[1] ;
 wire \a_reg[2] ;
 wire \a_reg[3] ;
 wire \a_reg[4] ;
 wire \a_reg[5] ;
 wire \a_reg[6] ;
 wire \a_reg[7] ;
 wire \b_reg[0] ;
 wire \b_reg[1] ;
 wire \b_reg[2] ;
 wire \b_reg[3] ;
 wire \b_reg[4] ;
 wire \b_reg[5] ;
 wire \b_reg[6] ;
 wire \b_reg[7] ;
 wire \next_state[0] ;
 wire \next_state[1] ;
 wire \state[0] ;
 wire \state[1] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net36;

 sky130_fd_sc_hd__clkbuf_4 _414_ (.A(\b_reg[0] ),
    .X(_033_));
 sky130_fd_sc_hd__nand2_1 _415_ (.A(_033_),
    .B(\a_reg[6] ),
    .Y(_129_));
 sky130_fd_sc_hd__clkbuf_4 _416_ (.A(\b_reg[1] ),
    .X(_034_));
 sky130_fd_sc_hd__buf_2 _417_ (.A(\a_reg[5] ),
    .X(_035_));
 sky130_fd_sc_hd__nand2_1 _418_ (.A(_034_),
    .B(_035_),
    .Y(_128_));
 sky130_fd_sc_hd__buf_2 _419_ (.A(\a_reg[4] ),
    .X(_036_));
 sky130_fd_sc_hd__nand2_1 _420_ (.A(\b_reg[2] ),
    .B(_036_),
    .Y(_127_));
 sky130_fd_sc_hd__and2_0 _421_ (.A(_034_),
    .B(_036_),
    .X(_141_));
 sky130_fd_sc_hd__and2_0 _422_ (.A(\b_reg[2] ),
    .B(\a_reg[3] ),
    .X(_140_));
 sky130_fd_sc_hd__and2_0 _423_ (.A(\a_reg[3] ),
    .B(\b_reg[3] ),
    .X(_134_));
 sky130_fd_sc_hd__buf_2 _424_ (.A(\a_reg[2] ),
    .X(_037_));
 sky130_fd_sc_hd__and2_0 _425_ (.A(\b_reg[4] ),
    .B(_037_),
    .X(_133_));
 sky130_fd_sc_hd__buf_2 _426_ (.A(\a_reg[1] ),
    .X(_038_));
 sky130_fd_sc_hd__and2_0 _427_ (.A(\b_reg[5] ),
    .B(_038_),
    .X(_132_));
 sky130_fd_sc_hd__and2_0 _428_ (.A(_034_),
    .B(\a_reg[3] ),
    .X(_159_));
 sky130_fd_sc_hd__and2_0 _429_ (.A(\b_reg[2] ),
    .B(_037_),
    .X(_158_));
 sky130_fd_sc_hd__and2_0 _430_ (.A(\a_reg[0] ),
    .B(\b_reg[6] ),
    .X(_326_));
 sky130_fd_sc_hd__nand2_1 _431_ (.A(_033_),
    .B(\a_reg[3] ),
    .Y(_174_));
 sky130_fd_sc_hd__and2_0 _432_ (.A(\b_reg[3] ),
    .B(_038_),
    .X(_329_));
 sky130_fd_sc_hd__and2_0 _433_ (.A(\b_reg[4] ),
    .B(\a_reg[0] ),
    .X(_328_));
 sky130_fd_sc_hd__nand2_1 _434_ (.A(_033_),
    .B(_037_),
    .Y(_182_));
 sky130_fd_sc_hd__and2_0 _435_ (.A(\b_reg[3] ),
    .B(\a_reg[0] ),
    .X(_177_));
 sky130_fd_sc_hd__and2_0 _436_ (.A(_033_),
    .B(_038_),
    .X(_404_));
 sky130_fd_sc_hd__and2_0 _437_ (.A(_034_),
    .B(\a_reg[0] ),
    .X(_405_));
 sky130_fd_sc_hd__nand2_1 _438_ (.A(\a_reg[6] ),
    .B(_034_),
    .Y(_192_));
 sky130_fd_sc_hd__nand2_1 _439_ (.A(_035_),
    .B(\b_reg[2] ),
    .Y(_196_));
 sky130_fd_sc_hd__nand2_1 _440_ (.A(_036_),
    .B(\b_reg[3] ),
    .Y(_198_));
 sky130_fd_sc_hd__nand2_1 _441_ (.A(\a_reg[3] ),
    .B(\b_reg[4] ),
    .Y(_197_));
 sky130_fd_sc_hd__nand2b_1 _442_ (.A_N(\a_reg[0] ),
    .B(\b_reg[7] ),
    .Y(_203_));
 sky130_fd_sc_hd__inv_1 _443_ (.A(_215_),
    .Y(_211_));
 sky130_fd_sc_hd__and2_0 _444_ (.A(\a_reg[6] ),
    .B(\b_reg[2] ),
    .X(_348_));
 sky130_fd_sc_hd__nand2_1 _445_ (.A(_035_),
    .B(\b_reg[3] ),
    .Y(_218_));
 sky130_fd_sc_hd__nand2_1 _446_ (.A(_036_),
    .B(\b_reg[4] ),
    .Y(_217_));
 sky130_fd_sc_hd__nand2_1 _447_ (.A(\a_reg[3] ),
    .B(\b_reg[5] ),
    .Y(_216_));
 sky130_fd_sc_hd__and2_0 _448_ (.A(_037_),
    .B(\b_reg[6] ),
    .X(_353_));
 sky130_fd_sc_hd__inv_2 _449_ (.A(\b_reg[7] ),
    .Y(_191_));
 sky130_fd_sc_hd__nor2_1 _450_ (.A(_038_),
    .B(_191_),
    .Y(_352_));
 sky130_fd_sc_hd__clkbuf_4 _451_ (.A(\a_reg[7] ),
    .X(_039_));
 sky130_fd_sc_hd__and2_0 _452_ (.A(\b_reg[2] ),
    .B(_039_),
    .X(_358_));
 sky130_fd_sc_hd__a31oi_2 _453_ (.A1(_033_),
    .A2(_034_),
    .A3(_039_),
    .B1(_350_),
    .Y(_239_));
 sky130_fd_sc_hd__nand2_1 _454_ (.A(\a_reg[6] ),
    .B(\b_reg[3] ),
    .Y(_235_));
 sky130_fd_sc_hd__nand2_1 _455_ (.A(_035_),
    .B(\b_reg[4] ),
    .Y(_236_));
 sky130_fd_sc_hd__nand2_1 _456_ (.A(_036_),
    .B(\b_reg[5] ),
    .Y(_234_));
 sky130_fd_sc_hd__and2_0 _457_ (.A(\a_reg[3] ),
    .B(\b_reg[6] ),
    .X(_362_));
 sky130_fd_sc_hd__nor2_1 _458_ (.A(_037_),
    .B(_191_),
    .Y(_361_));
 sky130_fd_sc_hd__a31oi_4 _459_ (.A1(_033_),
    .A2(_034_),
    .A3(_039_),
    .B1(_359_),
    .Y(_259_));
 sky130_fd_sc_hd__and2_1 _460_ (.A(\b_reg[3] ),
    .B(_039_),
    .X(_253_));
 sky130_fd_sc_hd__and2_0 _461_ (.A(\a_reg[6] ),
    .B(\b_reg[4] ),
    .X(_254_));
 sky130_fd_sc_hd__and2_0 _462_ (.A(_035_),
    .B(\b_reg[5] ),
    .X(_255_));
 sky130_fd_sc_hd__and2_0 _463_ (.A(_036_),
    .B(\b_reg[6] ),
    .X(_366_));
 sky130_fd_sc_hd__nor2_1 _464_ (.A(\a_reg[3] ),
    .B(_191_),
    .Y(_367_));
 sky130_fd_sc_hd__inv_1 _465_ (.A(_342_),
    .Y(_186_));
 sky130_fd_sc_hd__and2_1 _466_ (.A(\b_reg[4] ),
    .B(_039_),
    .X(_274_));
 sky130_fd_sc_hd__and2_0 _467_ (.A(\a_reg[6] ),
    .B(\b_reg[5] ),
    .X(_273_));
 sky130_fd_sc_hd__and2_0 _468_ (.A(_035_),
    .B(\b_reg[6] ),
    .X(_372_));
 sky130_fd_sc_hd__nor2_1 _469_ (.A(_036_),
    .B(_191_),
    .Y(_373_));
 sky130_fd_sc_hd__and2_0 _470_ (.A(\b_reg[5] ),
    .B(_039_),
    .X(_290_));
 sky130_fd_sc_hd__and2_0 _471_ (.A(\a_reg[6] ),
    .B(\b_reg[6] ),
    .X(_379_));
 sky130_fd_sc_hd__nor2_1 _472_ (.A(_035_),
    .B(_191_),
    .Y(_380_));
 sky130_fd_sc_hd__and2_0 _473_ (.A(\b_reg[6] ),
    .B(_039_),
    .X(_389_));
 sky130_fd_sc_hd__nor2_1 _474_ (.A(\a_reg[6] ),
    .B(_191_),
    .Y(_388_));
 sky130_fd_sc_hd__nand2_1 _475_ (.A(\b_reg[5] ),
    .B(\a_reg[0] ),
    .Y(_145_));
 sky130_fd_sc_hd__nand2_1 _476_ (.A(\b_reg[2] ),
    .B(_038_),
    .Y(_172_));
 sky130_fd_sc_hd__nand2_1 _477_ (.A(\b_reg[2] ),
    .B(\a_reg[0] ),
    .Y(_181_));
 sky130_fd_sc_hd__nand2_1 _478_ (.A(\b_reg[4] ),
    .B(_038_),
    .Y(_146_));
 sky130_fd_sc_hd__inv_1 _479_ (.A(_330_),
    .Y(_163_));
 sky130_fd_sc_hd__nand2_1 _480_ (.A(_034_),
    .B(_037_),
    .Y(_173_));
 sky130_fd_sc_hd__nand2_1 _481_ (.A(_037_),
    .B(\b_reg[5] ),
    .Y(_204_));
 sky130_fd_sc_hd__nand2_1 _482_ (.A(\b_reg[3] ),
    .B(_037_),
    .Y(_147_));
 sky130_fd_sc_hd__nand2_1 _483_ (.A(_034_),
    .B(_038_),
    .Y(_183_));
 sky130_fd_sc_hd__nand2_1 _484_ (.A(_033_),
    .B(_039_),
    .Y(_193_));
 sky130_fd_sc_hd__nand2_1 _485_ (.A(_038_),
    .B(\b_reg[6] ),
    .Y(_205_));
 sky130_fd_sc_hd__inv_1 _486_ (.A(_144_),
    .Y(_156_));
 sky130_fd_sc_hd__inv_1 _487_ (.A(_154_),
    .Y(_332_));
 sky130_fd_sc_hd__inv_1 _488_ (.A(_161_),
    .Y(_168_));
 sky130_fd_sc_hd__inv_1 _489_ (.A(_247_),
    .Y(_248_));
 sky130_fd_sc_hd__inv_1 _490_ (.A(_257_),
    .Y(_258_));
 sky130_fd_sc_hd__inv_1 _491_ (.A(_266_),
    .Y(_267_));
 sky130_fd_sc_hd__inv_1 _492_ (.A(_276_),
    .Y(_277_));
 sky130_fd_sc_hd__inv_1 _493_ (.A(_283_),
    .Y(_284_));
 sky130_fd_sc_hd__inv_1 _494_ (.A(_292_),
    .Y(_293_));
 sky130_fd_sc_hd__inv_1 _495_ (.A(_299_),
    .Y(_300_));
 sky130_fd_sc_hd__inv_1 _496_ (.A(_309_),
    .Y(_310_));
 sky130_fd_sc_hd__inv_1 _497_ (.A(_319_),
    .Y(_320_));
 sky130_fd_sc_hd__inv_1 _498_ (.A(_143_),
    .Y(_137_));
 sky130_fd_sc_hd__inv_1 _499_ (.A(_153_),
    .Y(_212_));
 sky130_fd_sc_hd__inv_1 _500_ (.A(_169_),
    .Y(_162_));
 sky130_fd_sc_hd__inv_1 _501_ (.A(_246_),
    .Y(_270_));
 sky130_fd_sc_hd__inv_1 _502_ (.A(_265_),
    .Y(_287_));
 sky130_fd_sc_hd__inv_1 _503_ (.A(_282_),
    .Y(_303_));
 sky130_fd_sc_hd__inv_1 _504_ (.A(_298_),
    .Y(_313_));
 sky130_fd_sc_hd__inv_1 _505_ (.A(_308_),
    .Y(_323_));
 sky130_fd_sc_hd__inv_1 _506_ (.A(_171_),
    .Y(_167_));
 sky130_fd_sc_hd__inv_1 _507_ (.A(_164_),
    .Y(_331_));
 sky130_fd_sc_hd__inv_1 _508_ (.A(_175_),
    .Y(_176_));
 sky130_fd_sc_hd__inv_1 _509_ (.A(_165_),
    .Y(_338_));
 sky130_fd_sc_hd__inv_1 _510_ (.A(_207_),
    .Y(_343_));
 sky130_fd_sc_hd__inv_1 _511_ (.A(_214_),
    .Y(_345_));
 sky130_fd_sc_hd__inv_1 _512_ (.A(_228_),
    .Y(_229_));
 sky130_fd_sc_hd__inv_1 _513_ (.A(_213_),
    .Y(_355_));
 sky130_fd_sc_hd__inv_1 _514_ (.A(_251_),
    .Y(_368_));
 sky130_fd_sc_hd__inv_1 _515_ (.A(_271_),
    .Y(_374_));
 sky130_fd_sc_hd__inv_1 _516_ (.A(_295_),
    .Y(_378_));
 sky130_fd_sc_hd__inv_1 _517_ (.A(_305_),
    .Y(_381_));
 sky130_fd_sc_hd__inv_1 _518_ (.A(_315_),
    .Y(_390_));
 sky130_fd_sc_hd__inv_1 _519_ (.A(_314_),
    .Y(_398_));
 sky130_fd_sc_hd__and2_0 _520_ (.A(_033_),
    .B(_035_),
    .X(_142_));
 sky130_fd_sc_hd__and2_0 _521_ (.A(_033_),
    .B(_036_),
    .X(_160_));
 sky130_fd_sc_hd__inv_1 _522_ (.A(_139_),
    .Y(_152_));
 sky130_fd_sc_hd__inv_1 _523_ (.A(_148_),
    .Y(_327_));
 sky130_fd_sc_hd__inv_1 _524_ (.A(_184_),
    .Y(_178_));
 sky130_fd_sc_hd__inv_1 _525_ (.A(_209_),
    .Y(_230_));
 sky130_fd_sc_hd__xor2_1 _526_ (.A(\b_reg[0] ),
    .B(\b_reg[1] ),
    .X(_040_));
 sky130_fd_sc_hd__and2_0 _527_ (.A(_039_),
    .B(_040_),
    .X(_349_));
 sky130_fd_sc_hd__inv_1 _528_ (.A(_219_),
    .Y(_244_));
 sky130_fd_sc_hd__inv_1 _529_ (.A(_252_),
    .Y(_363_));
 sky130_fd_sc_hd__inv_1 _530_ (.A(_237_),
    .Y(_264_));
 sky130_fd_sc_hd__inv_1 _531_ (.A(_272_),
    .Y(_369_));
 sky130_fd_sc_hd__inv_1 _532_ (.A(_289_),
    .Y(_375_));
 sky130_fd_sc_hd__inv_1 _533_ (.A(_288_),
    .Y(_382_));
 sky130_fd_sc_hd__inv_1 _534_ (.A(_294_),
    .Y(_385_));
 sky130_fd_sc_hd__inv_1 _535_ (.A(_304_),
    .Y(_391_));
 sky130_fd_sc_hd__nor2_1 _536_ (.A(_039_),
    .B(_191_),
    .Y(_394_));
 sky130_fd_sc_hd__inv_1 _537_ (.A(_325_),
    .Y(_399_));
 sky130_fd_sc_hd__inv_1 _538_ (.A(_185_),
    .Y(_408_));
 sky130_fd_sc_hd__inv_1 _539_ (.A(_334_),
    .Y(_188_));
 sky130_fd_sc_hd__inv_1 _540_ (.A(_344_),
    .Y(_208_));
 sky130_fd_sc_hd__inv_1 _541_ (.A(_351_),
    .Y(_221_));
 sky130_fd_sc_hd__clkinvlp_4 _542_ (.A(_360_),
    .Y(_240_));
 sky130_fd_sc_hd__inv_1 _543_ (.A(_354_),
    .Y(_224_));
 sky130_fd_sc_hd__inv_1 _544_ (.A(_335_),
    .Y(_187_));
 sky130_fd_sc_hd__nand2b_2 _545_ (.A_N(\state[0] ),
    .B(net18),
    .Y(_041_));
 sky130_fd_sc_hd__nor2_8 _546_ (.A(\state[1] ),
    .B(_041_),
    .Y(_042_));
 sky130_fd_sc_hd__buf_4 _547_ (.A(_042_),
    .X(\next_state[0] ));
 sky130_fd_sc_hd__mux2_1 _548_ (.A0(\a_reg[0] ),
    .A1(net2),
    .S(\next_state[0] ),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _549_ (.A0(_038_),
    .A1(net3),
    .S(\next_state[0] ),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _550_ (.A0(_037_),
    .A1(net4),
    .S(\next_state[0] ),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _551_ (.A0(\a_reg[3] ),
    .A1(net5),
    .S(\next_state[0] ),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _552_ (.A0(_036_),
    .A1(net6),
    .S(\next_state[0] ),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _553_ (.A0(_035_),
    .A1(net7),
    .S(\next_state[0] ),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _554_ (.A0(\a_reg[6] ),
    .A1(net8),
    .S(\next_state[0] ),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _555_ (.A0(\a_reg[7] ),
    .A1(net9),
    .S(_042_),
    .X(_007_));
 sky130_fd_sc_hd__mux2_1 _556_ (.A0(\b_reg[0] ),
    .A1(net10),
    .S(_042_),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _557_ (.A0(_034_),
    .A1(net11),
    .S(_042_),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _558_ (.A0(\b_reg[2] ),
    .A1(net12),
    .S(_042_),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _559_ (.A0(\b_reg[3] ),
    .A1(net13),
    .S(_042_),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _560_ (.A0(\b_reg[4] ),
    .A1(net14),
    .S(_042_),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _561_ (.A0(\b_reg[5] ),
    .A1(net15),
    .S(_042_),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _562_ (.A0(\b_reg[6] ),
    .A1(net16),
    .S(_042_),
    .X(_014_));
 sky130_fd_sc_hd__nand2_1 _563_ (.A(net17),
    .B(\next_state[0] ),
    .Y(_043_));
 sky130_fd_sc_hd__o21ai_0 _564_ (.A1(_191_),
    .A2(\next_state[0] ),
    .B1(_043_),
    .Y(_015_));
 sky130_fd_sc_hd__inv_1 _565_ (.A(\state[1] ),
    .Y(_044_));
 sky130_fd_sc_hd__nand2_1 _566_ (.A(net19),
    .B(_041_),
    .Y(_045_));
 sky130_fd_sc_hd__o21ai_0 _567_ (.A1(_044_),
    .A2(\state[0] ),
    .B1(_045_),
    .Y(_016_));
 sky130_fd_sc_hd__nand2_2 _568_ (.A(_044_),
    .B(\state[0] ),
    .Y(_046_));
 sky130_fd_sc_hd__clkbuf_4 _569_ (.A(_046_),
    .X(_047_));
 sky130_fd_sc_hd__nand2_1 _570_ (.A(net20),
    .B(_047_),
    .Y(_048_));
 sky130_fd_sc_hd__inv_1 _571_ (.A(_046_),
    .Y(_049_));
 sky130_fd_sc_hd__clkbuf_4 _572_ (.A(_049_),
    .X(\next_state[1] ));
 sky130_fd_sc_hd__nand3_1 _573_ (.A(_033_),
    .B(\a_reg[0] ),
    .C(\next_state[1] ),
    .Y(_050_));
 sky130_fd_sc_hd__nand2_1 _574_ (.A(_048_),
    .B(_050_),
    .Y(_017_));
 sky130_fd_sc_hd__buf_2 _575_ (.A(_046_),
    .X(_051_));
 sky130_fd_sc_hd__a211oi_1 _576_ (.A1(_337_),
    .A2(_342_),
    .B1(_336_),
    .C1(_346_),
    .Y(_052_));
 sky130_fd_sc_hd__o21ai_0 _577_ (.A1(_347_),
    .A2(_346_),
    .B1(_357_),
    .Y(_053_));
 sky130_fd_sc_hd__o21bai_1 _578_ (.A1(_052_),
    .A2(_053_),
    .B1_N(_356_),
    .Y(_054_));
 sky130_fd_sc_hd__a21oi_1 _579_ (.A1(_365_),
    .A2(_054_),
    .B1(_364_),
    .Y(_055_));
 sky130_fd_sc_hd__xor2_1 _580_ (.A(_371_),
    .B(_055_),
    .X(_056_));
 sky130_fd_sc_hd__nand2_1 _581_ (.A(net21),
    .B(_051_),
    .Y(_057_));
 sky130_fd_sc_hd__o21ai_0 _582_ (.A1(_051_),
    .A2(_056_),
    .B1(_057_),
    .Y(_018_));
 sky130_fd_sc_hd__clkbuf_2 _583_ (.A(_377_),
    .X(_058_));
 sky130_fd_sc_hd__nor2b_1 _584_ (.A(_189_),
    .B_N(_347_),
    .Y(_059_));
 sky130_fd_sc_hd__o21a_1 _585_ (.A1(_357_),
    .A2(_356_),
    .B1(_365_),
    .X(_060_));
 sky130_fd_sc_hd__o31a_1 _586_ (.A1(_346_),
    .A2(_356_),
    .A3(_059_),
    .B1(_060_),
    .X(_061_));
 sky130_fd_sc_hd__o21a_1 _587_ (.A1(_364_),
    .A2(_061_),
    .B1(_371_),
    .X(_062_));
 sky130_fd_sc_hd__nor3_1 _588_ (.A(_058_),
    .B(_370_),
    .C(_062_),
    .Y(_063_));
 sky130_fd_sc_hd__o21a_1 _589_ (.A1(_370_),
    .A2(_062_),
    .B1(_058_),
    .X(_064_));
 sky130_fd_sc_hd__nand2_1 _590_ (.A(net22),
    .B(_047_),
    .Y(_065_));
 sky130_fd_sc_hd__o31ai_1 _591_ (.A1(_046_),
    .A2(_063_),
    .A3(_064_),
    .B1(_065_),
    .Y(_019_));
 sky130_fd_sc_hd__clkbuf_2 _592_ (.A(_384_),
    .X(_066_));
 sky130_fd_sc_hd__and3_1 _593_ (.A(_365_),
    .B(_371_),
    .C(_058_),
    .X(_067_));
 sky130_fd_sc_hd__a21oi_1 _594_ (.A1(_058_),
    .A2(_370_),
    .B1(_376_),
    .Y(_068_));
 sky130_fd_sc_hd__nand3_1 _595_ (.A(_371_),
    .B(_058_),
    .C(_364_),
    .Y(_069_));
 sky130_fd_sc_hd__nand2_1 _596_ (.A(_068_),
    .B(_069_),
    .Y(_070_));
 sky130_fd_sc_hd__a21oi_1 _597_ (.A1(_054_),
    .A2(_067_),
    .B1(_070_),
    .Y(_071_));
 sky130_fd_sc_hd__xor2_1 _598_ (.A(_066_),
    .B(_071_),
    .X(_072_));
 sky130_fd_sc_hd__nand2_1 _599_ (.A(net23),
    .B(_051_),
    .Y(_073_));
 sky130_fd_sc_hd__o21ai_0 _600_ (.A1(_051_),
    .A2(_072_),
    .B1(_073_),
    .Y(_020_));
 sky130_fd_sc_hd__o2111ai_1 _601_ (.A1(_364_),
    .A2(_061_),
    .B1(_371_),
    .C1(_058_),
    .D1(_066_),
    .Y(_074_));
 sky130_fd_sc_hd__nor2b_1 _602_ (.A(_068_),
    .B_N(_066_),
    .Y(_075_));
 sky130_fd_sc_hd__nor2_1 _603_ (.A(_383_),
    .B(_075_),
    .Y(_076_));
 sky130_fd_sc_hd__a211o_1 _604_ (.A1(_074_),
    .A2(_076_),
    .B1(_393_),
    .C1(_046_),
    .X(_077_));
 sky130_fd_sc_hd__nand4_1 _605_ (.A(_393_),
    .B(\next_state[1] ),
    .C(_074_),
    .D(_076_),
    .Y(_078_));
 sky130_fd_sc_hd__nand2_1 _606_ (.A(net24),
    .B(_047_),
    .Y(_079_));
 sky130_fd_sc_hd__nand3_1 _607_ (.A(_077_),
    .B(_078_),
    .C(_079_),
    .Y(_021_));
 sky130_fd_sc_hd__nor2_1 _608_ (.A(net25),
    .B(_049_),
    .Y(_080_));
 sky130_fd_sc_hd__nand4_1 _609_ (.A(_371_),
    .B(_058_),
    .C(_066_),
    .D(_393_),
    .Y(_081_));
 sky130_fd_sc_hd__nand2_1 _610_ (.A(_401_),
    .B(_081_),
    .Y(_082_));
 sky130_fd_sc_hd__nand2_1 _611_ (.A(_066_),
    .B(_393_),
    .Y(_083_));
 sky130_fd_sc_hd__a21oi_1 _612_ (.A1(_393_),
    .A2(_383_),
    .B1(_392_),
    .Y(_084_));
 sky130_fd_sc_hd__o21ai_1 _613_ (.A1(_068_),
    .A2(_083_),
    .B1(_084_),
    .Y(_085_));
 sky130_fd_sc_hd__mux2i_1 _614_ (.A0(_082_),
    .A1(_401_),
    .S(_085_),
    .Y(_086_));
 sky130_fd_sc_hd__nor2_1 _615_ (.A(_046_),
    .B(_086_),
    .Y(_087_));
 sky130_fd_sc_hd__nor2_1 _616_ (.A(_401_),
    .B(_081_),
    .Y(_088_));
 sky130_fd_sc_hd__inv_1 _617_ (.A(_401_),
    .Y(_089_));
 sky130_fd_sc_hd__nor2_1 _618_ (.A(_089_),
    .B(_085_),
    .Y(_090_));
 sky130_fd_sc_hd__mux2i_1 _619_ (.A0(_088_),
    .A1(_090_),
    .S(_055_),
    .Y(_091_));
 sky130_fd_sc_hd__o22ai_1 _620_ (.A1(_080_),
    .A2(_087_),
    .B1(_091_),
    .B2(_047_),
    .Y(_022_));
 sky130_fd_sc_hd__nand4_1 _621_ (.A(_058_),
    .B(_066_),
    .C(_393_),
    .D(_401_),
    .Y(_092_));
 sky130_fd_sc_hd__nor2_1 _622_ (.A(_371_),
    .B(_370_),
    .Y(_093_));
 sky130_fd_sc_hd__nor2_1 _623_ (.A(_092_),
    .B(_093_),
    .Y(_094_));
 sky130_fd_sc_hd__o31ai_1 _624_ (.A1(_364_),
    .A2(_370_),
    .A3(_061_),
    .B1(_094_),
    .Y(_095_));
 sky130_fd_sc_hd__a21o_1 _625_ (.A1(_066_),
    .A2(_376_),
    .B1(_383_),
    .X(_096_));
 sky130_fd_sc_hd__nand3_1 _626_ (.A(_393_),
    .B(_401_),
    .C(_096_),
    .Y(_097_));
 sky130_fd_sc_hd__a21oi_1 _627_ (.A1(_401_),
    .A2(_392_),
    .B1(_400_),
    .Y(_098_));
 sky130_fd_sc_hd__xor2_1 _628_ (.A(_318_),
    .B(_397_),
    .X(_099_));
 sky130_fd_sc_hd__xnor2_1 _629_ (.A(_321_),
    .B(_324_),
    .Y(_100_));
 sky130_fd_sc_hd__xnor2_1 _630_ (.A(_099_),
    .B(_100_),
    .Y(_101_));
 sky130_fd_sc_hd__xnor2_1 _631_ (.A(_395_),
    .B(_387_),
    .Y(_102_));
 sky130_fd_sc_hd__xnor2_1 _632_ (.A(_101_),
    .B(_102_),
    .Y(_103_));
 sky130_fd_sc_hd__a31o_1 _633_ (.A1(_095_),
    .A2(_097_),
    .A3(_098_),
    .B1(_103_),
    .X(_104_));
 sky130_fd_sc_hd__nand4_1 _634_ (.A(_103_),
    .B(_095_),
    .C(_097_),
    .D(_098_),
    .Y(_105_));
 sky130_fd_sc_hd__nor2_1 _635_ (.A(net26),
    .B(\next_state[1] ),
    .Y(_106_));
 sky130_fd_sc_hd__a31oi_1 _636_ (.A1(\next_state[1] ),
    .A2(_104_),
    .A3(_105_),
    .B1(_106_),
    .Y(_023_));
 sky130_fd_sc_hd__nand2_1 _637_ (.A(_407_),
    .B(\next_state[1] ),
    .Y(_107_));
 sky130_fd_sc_hd__nand2_1 _638_ (.A(net27),
    .B(_047_),
    .Y(_108_));
 sky130_fd_sc_hd__nand2_1 _639_ (.A(_107_),
    .B(_108_),
    .Y(_024_));
 sky130_fd_sc_hd__nand2_1 _640_ (.A(_410_),
    .B(\next_state[1] ),
    .Y(_109_));
 sky130_fd_sc_hd__nand2_1 _641_ (.A(net28),
    .B(_047_),
    .Y(_110_));
 sky130_fd_sc_hd__nand2_1 _642_ (.A(_109_),
    .B(_110_),
    .Y(_025_));
 sky130_fd_sc_hd__nand2_1 _643_ (.A(_412_),
    .B(\next_state[1] ),
    .Y(_111_));
 sky130_fd_sc_hd__nand2_1 _644_ (.A(net29),
    .B(_047_),
    .Y(_112_));
 sky130_fd_sc_hd__nand2_1 _645_ (.A(_111_),
    .B(_112_),
    .Y(_026_));
 sky130_fd_sc_hd__nand2_1 _646_ (.A(_413_),
    .B(\next_state[1] ),
    .Y(_113_));
 sky130_fd_sc_hd__nand2_1 _647_ (.A(net30),
    .B(_047_),
    .Y(_114_));
 sky130_fd_sc_hd__nand2_1 _648_ (.A(_113_),
    .B(_114_),
    .Y(_027_));
 sky130_fd_sc_hd__nand2_1 _649_ (.A(_403_),
    .B(\next_state[1] ),
    .Y(_115_));
 sky130_fd_sc_hd__nand2_1 _650_ (.A(net31),
    .B(_047_),
    .Y(_116_));
 sky130_fd_sc_hd__nand2_1 _651_ (.A(_115_),
    .B(_116_),
    .Y(_028_));
 sky130_fd_sc_hd__nand2_1 _652_ (.A(net32),
    .B(_051_),
    .Y(_117_));
 sky130_fd_sc_hd__o21ai_0 _653_ (.A1(_190_),
    .A2(_047_),
    .B1(_117_),
    .Y(_029_));
 sky130_fd_sc_hd__xor2_1 _654_ (.A(_347_),
    .B(_189_),
    .X(_118_));
 sky130_fd_sc_hd__nand2_1 _655_ (.A(net33),
    .B(_051_),
    .Y(_119_));
 sky130_fd_sc_hd__o21ai_0 _656_ (.A1(_051_),
    .A2(_118_),
    .B1(_119_),
    .Y(_030_));
 sky130_fd_sc_hd__a21o_1 _657_ (.A1(_337_),
    .A2(_342_),
    .B1(_336_),
    .X(_120_));
 sky130_fd_sc_hd__a21oi_1 _658_ (.A1(_347_),
    .A2(_120_),
    .B1(_346_),
    .Y(_121_));
 sky130_fd_sc_hd__xor2_1 _659_ (.A(_357_),
    .B(_121_),
    .X(_122_));
 sky130_fd_sc_hd__nand2_1 _660_ (.A(net34),
    .B(_051_),
    .Y(_123_));
 sky130_fd_sc_hd__o21ai_0 _661_ (.A1(_051_),
    .A2(_122_),
    .B1(_123_),
    .Y(_031_));
 sky130_fd_sc_hd__o21ai_0 _662_ (.A1(_346_),
    .A2(_059_),
    .B1(_357_),
    .Y(_124_));
 sky130_fd_sc_hd__nor2_1 _663_ (.A(_365_),
    .B(_356_),
    .Y(_125_));
 sky130_fd_sc_hd__a211oi_1 _664_ (.A1(_124_),
    .A2(_125_),
    .B1(_061_),
    .C1(_046_),
    .Y(_126_));
 sky130_fd_sc_hd__a21o_1 _665_ (.A1(net35),
    .A2(_051_),
    .B1(_126_),
    .X(_032_));
 sky130_fd_sc_hd__fa_1 _666_ (.A(_127_),
    .B(_128_),
    .CIN(_129_),
    .COUT(_130_),
    .SUM(_131_));
 sky130_fd_sc_hd__fa_1 _667_ (.A(_132_),
    .B(_133_),
    .CIN(_134_),
    .COUT(_135_),
    .SUM(_136_));
 sky130_fd_sc_hd__fa_1 _668_ (.A(_136_),
    .B(_137_),
    .CIN(_131_),
    .COUT(_138_),
    .SUM(_139_));
 sky130_fd_sc_hd__fa_1 _669_ (.A(_140_),
    .B(_141_),
    .CIN(_142_),
    .COUT(_143_),
    .SUM(_144_));
 sky130_fd_sc_hd__fa_1 _670_ (.A(_145_),
    .B(_146_),
    .CIN(_147_),
    .COUT(_148_),
    .SUM(_149_));
 sky130_fd_sc_hd__fa_1 _671_ (.A(_150_),
    .B(_151_),
    .CIN(_152_),
    .COUT(_153_),
    .SUM(_154_));
 sky130_fd_sc_hd__fa_1 _672_ (.A(_149_),
    .B(_155_),
    .CIN(_156_),
    .COUT(_151_),
    .SUM(_157_));
 sky130_fd_sc_hd__fa_1 _673_ (.A(_158_),
    .B(_159_),
    .CIN(_160_),
    .COUT(_155_),
    .SUM(_161_));
 sky130_fd_sc_hd__fa_1 _674_ (.A(_162_),
    .B(_163_),
    .CIN(_157_),
    .COUT(_164_),
    .SUM(_165_));
 sky130_fd_sc_hd__fa_1 _675_ (.A(_166_),
    .B(_167_),
    .CIN(_168_),
    .COUT(_169_),
    .SUM(_170_));
 sky130_fd_sc_hd__fa_1 _676_ (.A(_172_),
    .B(_173_),
    .CIN(_174_),
    .COUT(_171_),
    .SUM(_175_));
 sky130_fd_sc_hd__fa_1 _677_ (.A(_176_),
    .B(_177_),
    .CIN(_178_),
    .COUT(_179_),
    .SUM(_180_));
 sky130_fd_sc_hd__fa_1 _678_ (.A(_181_),
    .B(_182_),
    .CIN(_183_),
    .COUT(_184_),
    .SUM(_185_));
 sky130_fd_sc_hd__fa_1 _679_ (.A(_186_),
    .B(_187_),
    .CIN(_188_),
    .COUT(_189_),
    .SUM(_190_));
 sky130_fd_sc_hd__fa_1 _680_ (.A(_191_),
    .B(_192_),
    .CIN(_193_),
    .COUT(_194_),
    .SUM(_195_));
 sky130_fd_sc_hd__fa_1 _681_ (.A(_196_),
    .B(_197_),
    .CIN(_198_),
    .COUT(_199_),
    .SUM(_200_));
 sky130_fd_sc_hd__fa_1 _682_ (.A(_195_),
    .B(_200_),
    .CIN(_130_),
    .COUT(_201_),
    .SUM(_202_));
 sky130_fd_sc_hd__fa_1 _683_ (.A(_203_),
    .B(_204_),
    .CIN(_205_),
    .COUT(_206_),
    .SUM(_207_));
 sky130_fd_sc_hd__fa_1 _684_ (.A(_208_),
    .B(_202_),
    .CIN(_138_),
    .COUT(_209_),
    .SUM(_210_));
 sky130_fd_sc_hd__fa_1 _685_ (.A(_211_),
    .B(_210_),
    .CIN(_212_),
    .COUT(_213_),
    .SUM(_214_));
 sky130_fd_sc_hd__fa_1 _686_ (.A(_216_),
    .B(_217_),
    .CIN(_218_),
    .COUT(_219_),
    .SUM(_220_));
 sky130_fd_sc_hd__fa_1 _687_ (.A(_220_),
    .B(_221_),
    .CIN(_194_),
    .COUT(_222_),
    .SUM(_223_));
 sky130_fd_sc_hd__fa_1 _688_ (.A(_224_),
    .B(_199_),
    .CIN(_206_),
    .COUT(_225_),
    .SUM(_226_));
 sky130_fd_sc_hd__fa_1 _689_ (.A(_223_),
    .B(_201_),
    .CIN(_226_),
    .COUT(_227_),
    .SUM(_228_));
 sky130_fd_sc_hd__fa_1 _690_ (.A(_229_),
    .B(_230_),
    .CIN(_231_),
    .COUT(_232_),
    .SUM(_233_));
 sky130_fd_sc_hd__fa_1 _691_ (.A(_234_),
    .B(_235_),
    .CIN(_236_),
    .COUT(_237_),
    .SUM(_238_));
 sky130_fd_sc_hd__fa_1 _692_ (.A(_238_),
    .B(_239_),
    .CIN(_240_),
    .COUT(_241_),
    .SUM(_242_));
 sky130_fd_sc_hd__fa_1 _693_ (.A(_243_),
    .B(_244_),
    .CIN(_245_),
    .COUT(_246_),
    .SUM(_247_));
 sky130_fd_sc_hd__fa_1 _694_ (.A(_242_),
    .B(_248_),
    .CIN(_222_),
    .COUT(_249_),
    .SUM(_250_));
 sky130_fd_sc_hd__fa_1 _695_ (.A(_227_),
    .B(_225_),
    .CIN(_250_),
    .COUT(_251_),
    .SUM(_252_));
 sky130_fd_sc_hd__fa_1 _696_ (.A(_253_),
    .B(_254_),
    .CIN(_255_),
    .COUT(_256_),
    .SUM(_257_));
 sky130_fd_sc_hd__fa_1 _697_ (.A(_258_),
    .B(_259_),
    .CIN(_240_),
    .COUT(_260_),
    .SUM(_261_));
 sky130_fd_sc_hd__fa_1 _698_ (.A(_262_),
    .B(_263_),
    .CIN(_264_),
    .COUT(_265_),
    .SUM(_266_));
 sky130_fd_sc_hd__fa_1 _699_ (.A(_267_),
    .B(_241_),
    .CIN(_261_),
    .COUT(_268_),
    .SUM(_269_));
 sky130_fd_sc_hd__fa_1 _700_ (.A(_269_),
    .B(_270_),
    .CIN(_249_),
    .COUT(_271_),
    .SUM(_272_));
 sky130_fd_sc_hd__fa_1 _701_ (.A(_273_),
    .B(_274_),
    .CIN(_253_),
    .COUT(_275_),
    .SUM(_276_));
 sky130_fd_sc_hd__fa_1 _702_ (.A(_277_),
    .B(_259_),
    .CIN(_240_),
    .COUT(_278_),
    .SUM(_279_));
 sky130_fd_sc_hd__fa_1 _703_ (.A(_256_),
    .B(_280_),
    .CIN(_281_),
    .COUT(_282_),
    .SUM(_283_));
 sky130_fd_sc_hd__fa_1 _704_ (.A(_260_),
    .B(_279_),
    .CIN(_284_),
    .COUT(_285_),
    .SUM(_286_));
 sky130_fd_sc_hd__fa_1 _705_ (.A(_286_),
    .B(_268_),
    .CIN(_287_),
    .COUT(_288_),
    .SUM(_289_));
 sky130_fd_sc_hd__fa_2 _706_ (.A(_274_),
    .B(_253_),
    .CIN(_290_),
    .COUT(_291_),
    .SUM(_292_));
 sky130_fd_sc_hd__fa_4 _707_ (.A(_259_),
    .B(_240_),
    .CIN(_293_),
    .COUT(_294_),
    .SUM(_295_));
 sky130_fd_sc_hd__fa_1 _708_ (.A(_275_),
    .B(_296_),
    .CIN(_297_),
    .COUT(_298_),
    .SUM(_299_));
 sky130_fd_sc_hd__fa_1 _709_ (.A(_295_),
    .B(_278_),
    .CIN(_300_),
    .COUT(_301_),
    .SUM(_302_));
 sky130_fd_sc_hd__fa_1 _710_ (.A(_285_),
    .B(_302_),
    .CIN(_303_),
    .COUT(_304_),
    .SUM(_305_));
 sky130_fd_sc_hd__fa_1 _711_ (.A(_306_),
    .B(_307_),
    .CIN(_291_),
    .COUT(_308_),
    .SUM(_309_));
 sky130_fd_sc_hd__fa_1 _712_ (.A(_295_),
    .B(_294_),
    .CIN(_310_),
    .COUT(_311_),
    .SUM(_312_));
 sky130_fd_sc_hd__fa_1 _713_ (.A(_313_),
    .B(_301_),
    .CIN(_312_),
    .COUT(_314_),
    .SUM(_315_));
 sky130_fd_sc_hd__fa_1 _714_ (.A(_291_),
    .B(_316_),
    .CIN(_317_),
    .COUT(_318_),
    .SUM(_319_));
 sky130_fd_sc_hd__fa_1 _715_ (.A(_295_),
    .B(_294_),
    .CIN(_320_),
    .COUT(_321_),
    .SUM(_322_));
 sky130_fd_sc_hd__fa_1 _716_ (.A(_311_),
    .B(_323_),
    .CIN(_322_),
    .COUT(_324_),
    .SUM(_325_));
 sky130_fd_sc_hd__ha_1 _717_ (.A(_326_),
    .B(_327_),
    .COUT(_215_),
    .SUM(_150_));
 sky130_fd_sc_hd__ha_1 _718_ (.A(_328_),
    .B(_329_),
    .COUT(_330_),
    .SUM(_166_));
 sky130_fd_sc_hd__ha_1 _719_ (.A(_331_),
    .B(_332_),
    .COUT(_333_),
    .SUM(_334_));
 sky130_fd_sc_hd__ha_1 _720_ (.A(_335_),
    .B(_334_),
    .COUT(_336_),
    .SUM(_337_));
 sky130_fd_sc_hd__ha_1 _721_ (.A(_338_),
    .B(_339_),
    .COUT(_335_),
    .SUM(_340_));
 sky130_fd_sc_hd__ha_1 _722_ (.A(_170_),
    .B(_179_),
    .COUT(_339_),
    .SUM(_341_));
 sky130_fd_sc_hd__ha_1 _723_ (.A(_343_),
    .B(_135_),
    .COUT(_231_),
    .SUM(_344_));
 sky130_fd_sc_hd__ha_1 _724_ (.A(_345_),
    .B(_333_),
    .COUT(_346_),
    .SUM(_347_));
 sky130_fd_sc_hd__ha_1 _725_ (.A(_348_),
    .B(_349_),
    .COUT(_350_),
    .SUM(_351_));
 sky130_fd_sc_hd__ha_1 _726_ (.A(_352_),
    .B(_353_),
    .COUT(_245_),
    .SUM(_354_));
 sky130_fd_sc_hd__ha_1 _727_ (.A(_355_),
    .B(_233_),
    .COUT(_356_),
    .SUM(_357_));
 sky130_fd_sc_hd__ha_1 _728_ (.A(_358_),
    .B(_349_),
    .COUT(_359_),
    .SUM(_360_));
 sky130_fd_sc_hd__ha_1 _729_ (.A(_361_),
    .B(_362_),
    .COUT(_262_),
    .SUM(_243_));
 sky130_fd_sc_hd__ha_1 _730_ (.A(_232_),
    .B(_363_),
    .COUT(_364_),
    .SUM(_365_));
 sky130_fd_sc_hd__ha_1 _731_ (.A(_366_),
    .B(_367_),
    .COUT(_281_),
    .SUM(_263_));
 sky130_fd_sc_hd__ha_2 _732_ (.A(_368_),
    .B(_369_),
    .COUT(_370_),
    .SUM(_371_));
 sky130_fd_sc_hd__ha_1 _733_ (.A(_372_),
    .B(_373_),
    .COUT(_296_),
    .SUM(_280_));
 sky130_fd_sc_hd__ha_1 _734_ (.A(_374_),
    .B(_375_),
    .COUT(_376_),
    .SUM(_377_));
 sky130_fd_sc_hd__ha_1 _735_ (.A(_379_),
    .B(_380_),
    .COUT(_307_),
    .SUM(_297_));
 sky130_fd_sc_hd__ha_1 _736_ (.A(_381_),
    .B(_382_),
    .COUT(_383_),
    .SUM(_384_));
 sky130_fd_sc_hd__ha_1 _737_ (.A(_378_),
    .B(_385_),
    .COUT(_386_),
    .SUM(_387_));
 sky130_fd_sc_hd__ha_1 _738_ (.A(_388_),
    .B(_389_),
    .COUT(_317_),
    .SUM(_306_));
 sky130_fd_sc_hd__ha_1 _739_ (.A(_390_),
    .B(_391_),
    .COUT(_392_),
    .SUM(_393_));
 sky130_fd_sc_hd__ha_1 _740_ (.A(_389_),
    .B(_394_),
    .COUT(_395_),
    .SUM(_316_));
 sky130_fd_sc_hd__ha_1 _741_ (.A(_291_),
    .B(_316_),
    .COUT(_396_),
    .SUM(_397_));
 sky130_fd_sc_hd__ha_2 _742_ (.A(_398_),
    .B(_399_),
    .COUT(_400_),
    .SUM(_401_));
 sky130_fd_sc_hd__ha_1 _743_ (.A(_340_),
    .B(_402_),
    .COUT(_342_),
    .SUM(_403_));
 sky130_fd_sc_hd__ha_1 _744_ (.A(_404_),
    .B(_405_),
    .COUT(_406_),
    .SUM(_407_));
 sky130_fd_sc_hd__ha_1 _745_ (.A(_406_),
    .B(_408_),
    .COUT(_409_),
    .SUM(_410_));
 sky130_fd_sc_hd__ha_1 _746_ (.A(_180_),
    .B(_409_),
    .COUT(_411_),
    .SUM(_412_));
 sky130_fd_sc_hd__ha_1 _747_ (.A(_341_),
    .B(_411_),
    .COUT(_402_),
    .SUM(_413_));
 sky130_fd_sc_hd__dfrtp_4 \a_reg[0]$_DFFE_PN0P_  (.D(_000_),
    .Q(\a_reg[0] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \a_reg[1]$_DFFE_PN0P_  (.D(_001_),
    .Q(\a_reg[1] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \a_reg[2]$_DFFE_PN0P_  (.D(_002_),
    .Q(\a_reg[2] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \a_reg[3]$_DFFE_PN0P_  (.D(_003_),
    .Q(\a_reg[3] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \a_reg[4]$_DFFE_PN0P_  (.D(_004_),
    .Q(\a_reg[4] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \a_reg[5]$_DFFE_PN0P_  (.D(_005_),
    .Q(\a_reg[5] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \a_reg[6]$_DFFE_PN0P_  (.D(_006_),
    .Q(\a_reg[6] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \a_reg[7]$_DFFE_PN0P_  (.D(_007_),
    .Q(\a_reg[7] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \b_reg[0]$_DFFE_PN0P_  (.D(_008_),
    .Q(\b_reg[0] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \b_reg[1]$_DFFE_PN0P_  (.D(_009_),
    .Q(\b_reg[1] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \b_reg[2]$_DFFE_PN0P_  (.D(_010_),
    .Q(\b_reg[2] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \b_reg[3]$_DFFE_PN0P_  (.D(_011_),
    .Q(\b_reg[3] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \b_reg[4]$_DFFE_PN0P_  (.D(_012_),
    .Q(\b_reg[4] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_4 \b_reg[5]$_DFFE_PN0P_  (.D(_013_),
    .Q(\b_reg[5] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \b_reg[6]$_DFFE_PN0P_  (.D(_014_),
    .Q(\b_reg[6] ),
    .RESET_B(net1),
    .CLK(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \b_reg[7]$_DFFE_PN0P_  (.D(_015_),
    .Q(\b_reg[7] ),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \done$_DFFE_PN0P_  (.D(_016_),
    .Q(net19),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[0]$_DFFE_PN0N_  (.D(_017_),
    .Q(net20),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[10]$_DFFE_PN0N_  (.D(_018_),
    .Q(net21),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[11]$_DFFE_PN0N_  (.D(_019_),
    .Q(net22),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[12]$_DFFE_PN0N_  (.D(_020_),
    .Q(net23),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[13]$_DFFE_PN0N_  (.D(_021_),
    .Q(net24),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[14]$_DFFE_PN0N_  (.D(_022_),
    .Q(net25),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[15]$_DFFE_PN0N_  (.D(_023_),
    .Q(net26),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[1]$_DFFE_PN0N_  (.D(_024_),
    .Q(net27),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[2]$_DFFE_PN0N_  (.D(_025_),
    .Q(net28),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[3]$_DFFE_PN0N_  (.D(_026_),
    .Q(net29),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[4]$_DFFE_PN0N_  (.D(_027_),
    .Q(net30),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[5]$_DFFE_PN0N_  (.D(_028_),
    .Q(net31),
    .RESET_B(net1),
    .CLK(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[6]$_DFFE_PN0N_  (.D(_029_),
    .Q(net32),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[7]$_DFFE_PN0N_  (.D(_030_),
    .Q(net33),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[8]$_DFFE_PN0N_  (.D(_031_),
    .Q(net34),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \product[9]$_DFFE_PN0N_  (.D(_032_),
    .Q(net35),
    .RESET_B(net1),
    .CLK(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__dfrtp_1 \state[0]$_DFF_PN0_  (.D(\next_state[0] ),
    .Q(\state[0] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__dfrtp_2 \state[1]$_DFF_PN0_  (.D(\next_state[1] ),
    .Q(\state[1] ),
    .RESET_B(net1),
    .CLK(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__buf_12 hold1 (.A(net36),
    .X(net1));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_76 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(multiplicand[0]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(multiplicand[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(multiplicand[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(multiplicand[3]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(multiplicand[4]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(multiplicand[5]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(multiplicand[6]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(multiplicand[7]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(multiplier[0]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(multiplier[1]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(multiplier[2]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(multiplier[3]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(multiplier[4]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(multiplier[5]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(multiplier[6]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(multiplier[7]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(start),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 output18 (.A(net19),
    .X(done));
 sky130_fd_sc_hd__clkbuf_1 output19 (.A(net20),
    .X(product[0]));
 sky130_fd_sc_hd__clkbuf_1 output20 (.A(net21),
    .X(product[10]));
 sky130_fd_sc_hd__clkbuf_1 output21 (.A(net22),
    .X(product[11]));
 sky130_fd_sc_hd__clkbuf_1 output22 (.A(net23),
    .X(product[12]));
 sky130_fd_sc_hd__clkbuf_1 output23 (.A(net24),
    .X(product[13]));
 sky130_fd_sc_hd__clkbuf_1 output24 (.A(net25),
    .X(product[14]));
 sky130_fd_sc_hd__clkbuf_1 output25 (.A(net26),
    .X(product[15]));
 sky130_fd_sc_hd__clkbuf_1 output26 (.A(net27),
    .X(product[1]));
 sky130_fd_sc_hd__clkbuf_1 output27 (.A(net28),
    .X(product[2]));
 sky130_fd_sc_hd__clkbuf_1 output28 (.A(net29),
    .X(product[3]));
 sky130_fd_sc_hd__clkbuf_1 output29 (.A(net30),
    .X(product[4]));
 sky130_fd_sc_hd__clkbuf_1 output30 (.A(net31),
    .X(product[5]));
 sky130_fd_sc_hd__clkbuf_1 output31 (.A(net32),
    .X(product[6]));
 sky130_fd_sc_hd__clkbuf_1 output32 (.A(net33),
    .X(product[7]));
 sky130_fd_sc_hd__clkbuf_1 output33 (.A(net34),
    .X(product[8]));
 sky130_fd_sc_hd__clkbuf_1 output34 (.A(net35),
    .X(product[9]));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload0 (.A(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload1 (.A(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload2 (.A(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(rst_n),
    .X(net36));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_68 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_6 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_65 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_75 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_102 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_158 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_25 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_37 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_49 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_108 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_73 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_29 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_113 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_163 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_58 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_50 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_62 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_72 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_12 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_59 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_98 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_64 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_142 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_106 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_150 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_88 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_170 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_96 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_108 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_147 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_158 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_44 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_60 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_68 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_80 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_171 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_76 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_173 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_87 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_104 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_174 ();
endmodule
