module parameterized_barrel_rotator (direction,
    data_in,
    data_out,
    rotate_amount);
 input direction;
 input [31:0] data_in;
 output [31:0] data_out;
 input [4:0] rotate_amount;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire net78;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net101;
 wire net73;
 wire net74;
 wire net75;
 wire net79;
 wire net84;
 wire net89;
 wire net99;
 wire net100;
 wire net66;
 wire net67;
 wire net80;
 wire net81;
 wire net91;
 wire net94;
 wire net102;
 wire net103;

 BUF_X32 _0573_ (.A(rotate_amount[0]),
    .Z(_0546_));
 INV_X32 _0574_ (.A(_0546_),
    .ZN(_0547_));
 BUF_X32 _0575_ (.A(_0547_),
    .Z(_0548_));
 BUF_X32 _0576_ (.A(_0548_),
    .Z(_0549_));
 BUF_X32 _0577_ (.A(_0549_),
    .Z(_0550_));
 BUF_X1 rebuffer15 (.A(_0559_),
    .Z(net78));
 CLKBUF_X3 _0579_ (.A(rotate_amount[1]),
    .Z(_0551_));
 INV_X1 _0580_ (.A(_0551_),
    .ZN(_0570_));
 BUF_X8 _0581_ (.A(rotate_amount[2]),
    .Z(_0552_));
 INV_X4 _0582_ (.A(_0552_),
    .ZN(_0553_));
 BUF_X4 _0583_ (.A(_0571_),
    .Z(_0554_));
 INV_X4 _0584_ (.A(_0554_),
    .ZN(_0555_));
 BUF_X8 _0585_ (.A(_0555_),
    .Z(_0556_));
 BUF_X4 _0586_ (.A(direction),
    .Z(_0557_));
 BUF_X16 _0587_ (.A(_0557_),
    .Z(_0558_));
 AOI21_X4 _0588_ (.A(_0553_),
    .B1(_0558_),
    .B2(_0556_),
    .ZN(_0559_));
 BUF_X4 _0589_ (.A(_0559_),
    .Z(_0560_));
 INV_X8 _0590_ (.A(_0557_),
    .ZN(_0561_));
 NOR3_X4 _0591_ (.A1(_0554_),
    .A2(_0552_),
    .A3(_0561_),
    .ZN(_0562_));
 BUF_X4 _0592_ (.A(_0562_),
    .Z(_0563_));
 CLKBUF_X3 _0593_ (.A(rotate_amount[4]),
    .Z(_0564_));
 CLKBUF_X3 _0594_ (.A(rotate_amount[3]),
    .Z(_0565_));
 BUF_X8 _0595_ (.A(_0546_),
    .Z(_0566_));
 OR4_X2 _0596_ (.A1(_0564_),
    .A2(_0565_),
    .A3(_0551_),
    .A4(_0566_),
    .ZN(_0567_));
 BUF_X32 _0597_ (.A(_0558_),
    .Z(_0568_));
 BUF_X4 _0598_ (.A(_0552_),
    .Z(_0000_));
 OR2_X1 _0599_ (.A1(_0568_),
    .A2(_0000_),
    .ZN(_0001_));
 BUF_X4 _0600_ (.A(_0554_),
    .Z(_0002_));
 BUF_X8 _0601_ (.A(_0572_),
    .Z(_0003_));
 INV_X4 _0602_ (.A(_0003_),
    .ZN(_0004_));
 BUF_X8 _0603_ (.A(_0004_),
    .Z(_0005_));
 AOI211_X2 _0604_ (.A(_0567_),
    .B(_0001_),
    .C1(_0002_),
    .C2(_0005_),
    .ZN(_0006_));
 NOR3_X4 _0605_ (.A1(_0560_),
    .A2(_0563_),
    .A3(_0006_),
    .ZN(_0007_));
 BUF_X8 _0606_ (.A(_0566_),
    .Z(_0008_));
 MUX2_X2 _0607_ (.A(net14),
    .B(net15),
    .S(_0008_),
    .Z(_0009_));
 MUX2_X1 _0608_ (.A(net16),
    .B(net17),
    .S(_0566_),
    .Z(_0010_));
 BUF_X16 _0609_ (.A(_0003_),
    .Z(_0011_));
 OAI21_X2 _0610_ (.A(_0011_),
    .B1(_0547_),
    .B2(_0558_),
    .ZN(_0012_));
 BUF_X4 _0611_ (.A(_0012_),
    .Z(_0013_));
 NAND3_X2 _0612_ (.A1(_0561_),
    .A2(_0566_),
    .A3(_0004_),
    .ZN(_0014_));
 BUF_X8 _0613_ (.A(_0014_),
    .Z(_0015_));
 NAND2_X4 _0614_ (.A1(_0013_),
    .A2(_0015_),
    .ZN(_0016_));
 MUX2_X1 _0615_ (.A(_0009_),
    .B(_0010_),
    .S(_0016_),
    .Z(_0017_));
 BUF_X1 _0616_ (.A(data_in[30]),
    .Z(_0018_));
 BUF_X16 _0617_ (.A(_0003_),
    .Z(_0019_));
 BUF_X16 _0618_ (.A(_0019_),
    .Z(_0020_));
 MUX2_X1 _0619_ (.A(net18),
    .B(_0018_),
    .S(_0020_),
    .Z(_0021_));
 CLKBUF_X2 _0620_ (.A(data_in[31]),
    .Z(_0022_));
 XNOR2_X2 _0621_ (.A(_0011_),
    .B(_0558_),
    .ZN(_0023_));
 BUF_X4 _0622_ (.A(_0023_),
    .Z(_0024_));
 MUX2_X1 _0623_ (.A(net19),
    .B(_0022_),
    .S(_0024_),
    .Z(_0025_));
 BUF_X8 _0624_ (.A(_0566_),
    .Z(_0026_));
 BUF_X4 _0625_ (.A(_0026_),
    .Z(_0027_));
 BUF_X4 _0626_ (.A(_0027_),
    .Z(_0028_));
 MUX2_X2 _0627_ (.A(_0021_),
    .B(_0025_),
    .S(_0028_),
    .Z(_0029_));
 OAI21_X4 _0628_ (.A(_0552_),
    .B1(_0554_),
    .B2(_0561_),
    .ZN(_0030_));
 NAND3_X4 _0629_ (.A1(_0558_),
    .A2(_0553_),
    .A3(_0555_),
    .ZN(_0031_));
 NAND2_X2 _0630_ (.A1(_0030_),
    .A2(_0031_),
    .ZN(_0032_));
 BUF_X4 _0631_ (.A(_0032_),
    .Z(_0033_));
 AOI22_X2 _0632_ (.A1(_0007_),
    .A2(_0017_),
    .B1(_0029_),
    .B2(_0033_),
    .ZN(_0034_));
 BUF_X1 _0633_ (.A(data_in[16]),
    .Z(_0035_));
 MUX2_X1 _0634_ (.A(_0035_),
    .B(net7),
    .S(_0016_),
    .Z(_0036_));
 NOR3_X4 _0635_ (.A1(_0028_),
    .A2(_0560_),
    .A3(_0563_),
    .ZN(_0037_));
 BUF_X4 _0636_ (.A(_0548_),
    .Z(_0038_));
 NOR3_X4 _0637_ (.A1(_0038_),
    .A2(net78),
    .A3(_0562_),
    .ZN(_0039_));
 BUF_X32 _0638_ (.A(_0011_),
    .Z(_0040_));
 BUF_X16 _0639_ (.A(_0040_),
    .Z(_0041_));
 NAND2_X1 _0640_ (.A1(_0041_),
    .A2(net8),
    .ZN(_0042_));
 BUF_X8 _0641_ (.A(_0561_),
    .Z(_0043_));
 BUF_X4 _0642_ (.A(_0043_),
    .Z(_0044_));
 AOI21_X2 _0643_ (.A(_0042_),
    .B1(_0027_),
    .B2(_0044_),
    .ZN(_0045_));
 INV_X1 _0644_ (.A(net6),
    .ZN(_0046_));
 BUF_X4 _0645_ (.A(_0043_),
    .Z(_0047_));
 AOI211_X2 _0646_ (.A(_0020_),
    .B(_0046_),
    .C1(_0047_),
    .C2(_0026_),
    .ZN(_0048_));
 BUF_X8 _0647_ (.A(_0568_),
    .Z(_0049_));
 INV_X1 _0648_ (.A(net8),
    .ZN(_0050_));
 NOR4_X2 _0649_ (.A1(_0049_),
    .A2(_0549_),
    .A3(_0041_),
    .A4(_0050_),
    .ZN(_0051_));
 NOR4_X2 _0650_ (.A1(_0049_),
    .A2(_0038_),
    .A3(_0005_),
    .A4(_0046_),
    .ZN(_0052_));
 OR4_X2 _0651_ (.A1(_0045_),
    .A2(_0048_),
    .A3(_0051_),
    .A4(_0052_),
    .ZN(_0053_));
 MUX2_X1 _0652_ (.A(net12),
    .B(net13),
    .S(_0008_),
    .Z(_0054_));
 AOI21_X1 _0653_ (.A(_0054_),
    .B1(_0015_),
    .B2(net81),
    .ZN(_0055_));
 INV_X1 _0654_ (.A(net10),
    .ZN(_0056_));
 INV_X1 _0655_ (.A(net11),
    .ZN(_0057_));
 MUX2_X1 _0656_ (.A(_0056_),
    .B(_0057_),
    .S(_0027_),
    .Z(_0058_));
 AOI21_X4 _0657_ (.A(_0004_),
    .B1(_0008_),
    .B2(_0561_),
    .ZN(_0059_));
 NOR3_X4 _0658_ (.A1(net91),
    .A2(net1),
    .A3(_0568_),
    .ZN(_0060_));
 NOR2_X2 _0659_ (.A1(_0059_),
    .A2(_0060_),
    .ZN(_0061_));
 AOI21_X1 _0660_ (.A(_0055_),
    .B1(_0058_),
    .B2(_0061_),
    .ZN(_0062_));
 AOI222_X2 _0661_ (.A1(_0036_),
    .A2(_0037_),
    .B1(_0053_),
    .B2(_0039_),
    .C1(_0033_),
    .C2(_0062_),
    .ZN(_0063_));
 NOR2_X2 _0662_ (.A1(_0551_),
    .A2(_0011_),
    .ZN(_0064_));
 OAI221_X2 _0663_ (.A(_0561_),
    .B1(net101),
    .B2(_0554_),
    .C1(_0064_),
    .C2(_0552_),
    .ZN(_0065_));
 NOR2_X1 _0664_ (.A1(_0552_),
    .A2(_0554_),
    .ZN(_0066_));
 OAI211_X2 _0665_ (.A(_0561_),
    .B(_0551_),
    .C1(_0019_),
    .C2(_0066_),
    .ZN(_0067_));
 NAND2_X1 _0666_ (.A1(_0561_),
    .A2(_0566_),
    .ZN(_0068_));
 NOR2_X1 _0667_ (.A1(_0551_),
    .A2(_0566_),
    .ZN(_0069_));
 NAND3_X1 _0668_ (.A1(_0568_),
    .A2(_0553_),
    .A3(_0069_),
    .ZN(_0070_));
 NAND4_X4 _0669_ (.A1(_0065_),
    .A2(_0067_),
    .A3(_0068_),
    .A4(_0070_),
    .ZN(_0071_));
 XOR2_X2 _0670_ (.A(_0565_),
    .B(_0071_),
    .Z(_0072_));
 BUF_X8 _0671_ (.A(_0072_),
    .Z(_0073_));
 BUF_X8 _0672_ (.A(_0073_),
    .Z(_0074_));
 MUX2_X1 _0673_ (.A(_0034_),
    .B(_0063_),
    .S(_0074_),
    .Z(_0075_));
 BUF_X16 _0674_ (.A(_0568_),
    .Z(_0076_));
 NOR3_X2 _0675_ (.A1(_0000_),
    .A2(_0556_),
    .A3(_0069_),
    .ZN(_0077_));
 NAND2_X2 _0676_ (.A1(_0568_),
    .A2(_0002_),
    .ZN(_0078_));
 OR2_X1 _0677_ (.A1(_0565_),
    .A2(_0552_),
    .ZN(_0079_));
 OAI22_X4 _0678_ (.A1(_0076_),
    .A2(_0077_),
    .B1(_0078_),
    .B2(_0079_),
    .ZN(_0080_));
 XOR2_X2 _0679_ (.A(_0564_),
    .B(_0080_),
    .Z(_0081_));
 BUF_X4 _0680_ (.A(_0081_),
    .Z(_0082_));
 CLKBUF_X2 _0681_ (.A(data_in[11]),
    .Z(_0083_));
 AND2_X1 _0682_ (.A1(_0019_),
    .A2(_0083_),
    .ZN(_0084_));
 OAI21_X1 _0683_ (.A(_0084_),
    .B1(net1),
    .B2(_0568_),
    .ZN(_0085_));
 CLKBUF_X2 _0684_ (.A(data_in[9]),
    .Z(_0086_));
 OAI211_X2 _0685_ (.A(_0005_),
    .B(_0086_),
    .C1(_0568_),
    .C2(net1),
    .ZN(_0087_));
 NAND4_X1 _0686_ (.A1(_0043_),
    .A2(_0008_),
    .A3(_0005_),
    .A4(_0083_),
    .ZN(_0088_));
 NAND2_X1 _0687_ (.A1(_0011_),
    .A2(_0086_),
    .ZN(_0089_));
 OR3_X1 _0688_ (.A1(_0568_),
    .A2(_0548_),
    .A3(_0089_),
    .ZN(_0090_));
 AND4_X4 _0689_ (.A1(_0085_),
    .A2(_0087_),
    .A3(_0088_),
    .A4(_0090_),
    .ZN(_0091_));
 NAND2_X1 _0690_ (.A1(net91),
    .A2(net5),
    .ZN(_0092_));
 AOI21_X2 _0691_ (.A(_0092_),
    .B1(_0008_),
    .B2(_0043_),
    .ZN(_0093_));
 INV_X1 _0692_ (.A(net3),
    .ZN(_0094_));
 AOI211_X2 _0693_ (.A(_0003_),
    .B(_0094_),
    .C1(_0561_),
    .C2(_0566_),
    .ZN(_0095_));
 INV_X1 _0694_ (.A(net5),
    .ZN(_0096_));
 NOR4_X2 _0695_ (.A1(_0558_),
    .A2(_0548_),
    .A3(net101),
    .A4(_0096_),
    .ZN(_0097_));
 NOR4_X2 _0696_ (.A1(_0558_),
    .A2(_0548_),
    .A3(_0004_),
    .A4(_0094_),
    .ZN(_0098_));
 NOR4_X4 _0697_ (.A1(_0093_),
    .A2(_0095_),
    .A3(_0097_),
    .A4(_0098_),
    .ZN(_0099_));
 AOI21_X4 _0698_ (.A(net65),
    .B1(_0030_),
    .B2(_0031_),
    .ZN(_0100_));
 AOI22_X1 _0699_ (.A1(_0039_),
    .A2(_0091_),
    .B1(net60),
    .B2(_0100_),
    .ZN(_0101_));
 BUF_X1 _0700_ (.A(data_in[10]),
    .Z(_0102_));
 AND2_X1 _0701_ (.A1(_0020_),
    .A2(_0102_),
    .ZN(_0103_));
 BUF_X4 _0702_ (.A(_0038_),
    .Z(_0104_));
 OAI21_X1 _0703_ (.A(_0103_),
    .B1(_0104_),
    .B2(_0049_),
    .ZN(_0105_));
 BUF_X4 _0704_ (.A(_0005_),
    .Z(_0106_));
 OAI211_X2 _0705_ (.A(_0106_),
    .B(net24),
    .C1(_0049_),
    .C2(_0104_),
    .ZN(_0107_));
 BUF_X4 _0706_ (.A(_0026_),
    .Z(_0108_));
 NAND4_X1 _0707_ (.A1(_0044_),
    .A2(_0108_),
    .A3(_0106_),
    .A4(_0102_),
    .ZN(_0109_));
 NAND2_X4 _0708_ (.A1(_0040_),
    .A2(net24),
    .ZN(_0110_));
 OR3_X4 _0709_ (.A1(_0076_),
    .A2(_0038_),
    .A3(_0110_),
    .ZN(_0111_));
 AND4_X2 _0710_ (.A1(_0105_),
    .A2(_0107_),
    .A3(_0109_),
    .A4(_0111_),
    .ZN(_0112_));
 BUF_X4 _0711_ (.A(_0020_),
    .Z(_0113_));
 NAND2_X2 _0712_ (.A1(_0113_),
    .A2(net4),
    .ZN(_0114_));
 AOI21_X4 _0713_ (.A(_0114_),
    .B1(_0028_),
    .B2(_0044_),
    .ZN(_0115_));
 INV_X2 _0714_ (.A(net2),
    .ZN(_0116_));
 AOI211_X2 _0715_ (.A(_0041_),
    .B(_0116_),
    .C1(_0047_),
    .C2(_0108_),
    .ZN(_0117_));
 BUF_X4 _0716_ (.A(_0049_),
    .Z(_0118_));
 INV_X2 _0717_ (.A(net4),
    .ZN(_0119_));
 NOR4_X4 _0718_ (.A1(_0113_),
    .A2(_0104_),
    .A3(_0118_),
    .A4(_0119_),
    .ZN(_0120_));
 NOR4_X4 _0719_ (.A1(_0106_),
    .A2(_0104_),
    .A3(_0118_),
    .A4(_0116_),
    .ZN(_0121_));
 NOR4_X4 _0720_ (.A1(_0115_),
    .A2(_0117_),
    .A3(_0120_),
    .A4(_0121_),
    .ZN(_0122_));
 CLKBUF_X3 _0721_ (.A(_0030_),
    .Z(_0123_));
 CLKBUF_X3 _0722_ (.A(_0031_),
    .Z(_0124_));
 AOI21_X2 _0723_ (.A(_0028_),
    .B1(_0123_),
    .B2(_0124_),
    .ZN(_0125_));
 AOI22_X1 _0724_ (.A1(_0037_),
    .A2(_0112_),
    .B1(_0122_),
    .B2(_0125_),
    .ZN(_0126_));
 NAND2_X1 _0725_ (.A1(_0101_),
    .A2(_0126_),
    .ZN(_0127_));
 NAND3_X4 _0726_ (.A1(_0027_),
    .A2(_0030_),
    .A3(_0031_),
    .ZN(_0128_));
 AND2_X1 _0727_ (.A1(_0040_),
    .A2(net21),
    .ZN(_0129_));
 OAI21_X1 _0728_ (.A(_0129_),
    .B1(net63),
    .B2(_0076_),
    .ZN(_0130_));
 OAI211_X2 _0729_ (.A(_0005_),
    .B(net9),
    .C1(_0076_),
    .C2(_0038_),
    .ZN(_0131_));
 NAND4_X2 _0730_ (.A1(_0047_),
    .A2(_0026_),
    .A3(_0005_),
    .A4(net21),
    .ZN(_0132_));
 AND2_X1 _0731_ (.A1(_0040_),
    .A2(net9),
    .ZN(_0133_));
 NAND3_X1 _0732_ (.A1(_0047_),
    .A2(_0026_),
    .A3(_0133_),
    .ZN(_0134_));
 AND4_X2 _0733_ (.A1(_0130_),
    .A2(_0131_),
    .A3(_0132_),
    .A4(_0134_),
    .ZN(_0135_));
 AND2_X1 _0734_ (.A1(net101),
    .A2(net23),
    .ZN(_0136_));
 OAI21_X1 _0735_ (.A(_0136_),
    .B1(_0104_),
    .B2(_0049_),
    .ZN(_0137_));
 BUF_X1 _0736_ (.A(data_in[5]),
    .Z(_0138_));
 OAI211_X2 _0737_ (.A(_0106_),
    .B(_0138_),
    .C1(_0049_),
    .C2(_0549_),
    .ZN(_0139_));
 NAND4_X1 _0738_ (.A1(_0047_),
    .A2(_0108_),
    .A3(_0005_),
    .A4(net23),
    .ZN(_0140_));
 NAND2_X4 _0739_ (.A1(_0040_),
    .A2(_0138_),
    .ZN(_0141_));
 OR3_X4 _0740_ (.A1(_0076_),
    .A2(_0038_),
    .A3(_0141_),
    .ZN(_0142_));
 AND4_X4 _0741_ (.A1(_0137_),
    .A2(_0139_),
    .A3(_0140_),
    .A4(_0142_),
    .ZN(_0143_));
 OAI21_X4 _0742_ (.A(_0108_),
    .B1(_0559_),
    .B2(_0562_),
    .ZN(_0144_));
 OAI22_X2 _0743_ (.A1(_0128_),
    .A2(_0135_),
    .B1(_0143_),
    .B2(_0144_),
    .ZN(_0145_));
 CLKBUF_X2 _0744_ (.A(data_in[0]),
    .Z(_0146_));
 MUX2_X1 _0745_ (.A(_0146_),
    .B(net20),
    .S(_0020_),
    .Z(_0147_));
 NOR3_X1 _0746_ (.A1(_0560_),
    .A2(_0563_),
    .A3(_0147_),
    .ZN(_0148_));
 AND2_X1 _0747_ (.A1(_0019_),
    .A2(net22),
    .ZN(_0149_));
 OAI21_X2 _0748_ (.A(_0149_),
    .B1(_0549_),
    .B2(_0049_),
    .ZN(_0150_));
 CLKBUF_X2 _0749_ (.A(data_in[4]),
    .Z(_0151_));
 OAI211_X2 _0750_ (.A(_0106_),
    .B(_0151_),
    .C1(_0049_),
    .C2(_0549_),
    .ZN(_0152_));
 NAND4_X2 _0751_ (.A1(_0047_),
    .A2(_0108_),
    .A3(_0005_),
    .A4(net22),
    .ZN(_0153_));
 NAND2_X4 _0752_ (.A1(_0040_),
    .A2(_0151_),
    .ZN(_0154_));
 OR3_X4 _0753_ (.A1(_0076_),
    .A2(net1),
    .A3(_0154_),
    .ZN(_0155_));
 AND4_X4 _0754_ (.A1(_0150_),
    .A2(_0152_),
    .A3(_0153_),
    .A4(_0155_),
    .ZN(_0156_));
 AOI211_X2 _0755_ (.A(_0028_),
    .B(_0148_),
    .C1(_0156_),
    .C2(_0032_),
    .ZN(_0157_));
 NOR2_X1 _0756_ (.A1(_0145_),
    .A2(_0157_),
    .ZN(_0158_));
 MUX2_X1 _0757_ (.A(_0127_),
    .B(_0158_),
    .S(_0074_),
    .Z(_0159_));
 NOR4_X4 _0758_ (.A1(_0564_),
    .A2(_0565_),
    .A3(_0551_),
    .A4(_0546_),
    .ZN(_0160_));
 NOR2_X2 _0759_ (.A1(_0558_),
    .A2(_0552_),
    .ZN(_0161_));
 OAI211_X4 _0760_ (.A(_0160_),
    .B(_0161_),
    .C1(_0556_),
    .C2(net91),
    .ZN(_0162_));
 NAND2_X4 _0761_ (.A1(_0162_),
    .A2(_0082_),
    .ZN(_0163_));
 OAI22_X1 _0762_ (.A1(_0075_),
    .A2(_0082_),
    .B1(_0159_),
    .B2(_0163_),
    .ZN(net25));
 XNOR2_X2 _0763_ (.A(_0565_),
    .B(_0071_),
    .ZN(_0164_));
 BUF_X4 _0764_ (.A(_0164_),
    .Z(_0165_));
 BUF_X4 _0765_ (.A(_0165_),
    .Z(_0166_));
 NAND3_X2 _0766_ (.A1(_0033_),
    .A2(_0016_),
    .A3(_0009_),
    .ZN(_0167_));
 NAND3_X1 _0767_ (.A1(net81),
    .A2(_0015_),
    .A3(_0054_),
    .ZN(_0168_));
 MUX2_X1 _0768_ (.A(_0050_),
    .B(_0057_),
    .S(_0023_),
    .Z(_0169_));
 MUX2_X1 _0769_ (.A(net7),
    .B(net10),
    .S(_0040_),
    .Z(_0170_));
 INV_X1 _0770_ (.A(_0170_),
    .ZN(_0171_));
 MUX2_X1 _0771_ (.A(_0169_),
    .B(_0171_),
    .S(_0104_),
    .Z(_0172_));
 NOR2_X1 _0772_ (.A1(_0559_),
    .A2(_0562_),
    .ZN(_0173_));
 BUF_X4 _0773_ (.A(_0173_),
    .Z(_0174_));
 MUX2_X1 _0774_ (.A(_0168_),
    .B(_0172_),
    .S(_0174_),
    .Z(_0175_));
 BUF_X4 _0775_ (.A(_0006_),
    .Z(_0176_));
 OAI211_X2 _0776_ (.A(_0166_),
    .B(_0167_),
    .C1(_0175_),
    .C2(_0176_),
    .ZN(_0177_));
 CLKBUF_X3 _0777_ (.A(_0027_),
    .Z(_0178_));
 MUX2_X1 _0778_ (.A(_0102_),
    .B(net2),
    .S(_0020_),
    .Z(_0179_));
 NOR3_X1 _0779_ (.A1(_0560_),
    .A2(_0563_),
    .A3(_0179_),
    .ZN(_0180_));
 NAND2_X1 _0780_ (.A1(_0020_),
    .A2(_0035_),
    .ZN(_0181_));
 OAI21_X1 _0781_ (.A(_0181_),
    .B1(_0119_),
    .B2(_0020_),
    .ZN(_0182_));
 AOI21_X1 _0782_ (.A(_0182_),
    .B1(_0124_),
    .B2(_0123_),
    .ZN(_0183_));
 OR3_X1 _0783_ (.A1(_0178_),
    .A2(_0180_),
    .A3(_0183_),
    .ZN(_0184_));
 MUX2_X1 _0784_ (.A(_0083_),
    .B(net3),
    .S(_0024_),
    .Z(_0185_));
 MUX2_X1 _0785_ (.A(net5),
    .B(net6),
    .S(_0023_),
    .Z(_0186_));
 AOI22_X2 _0786_ (.A1(_0039_),
    .A2(_0185_),
    .B1(_0186_),
    .B2(_0100_),
    .ZN(_0187_));
 AOI21_X2 _0787_ (.A(_0176_),
    .B1(_0184_),
    .B2(_0187_),
    .ZN(_0188_));
 OAI211_X2 _0788_ (.A(_0082_),
    .B(_0177_),
    .C1(_0188_),
    .C2(_0166_),
    .ZN(_0189_));
 BUF_X4 _0789_ (.A(_0174_),
    .Z(_0190_));
 NOR3_X2 _0790_ (.A1(_0059_),
    .A2(_0060_),
    .A3(_0010_),
    .ZN(_0191_));
 AND2_X1 _0791_ (.A1(_0566_),
    .A2(net19),
    .ZN(_0192_));
 AOI221_X2 _0792_ (.A(_0192_),
    .B1(_0014_),
    .B2(_0012_),
    .C1(_0038_),
    .C2(net18),
    .ZN(_0193_));
 OAI21_X1 _0793_ (.A(_0190_),
    .B1(_0191_),
    .B2(_0193_),
    .ZN(_0194_));
 OR2_X1 _0794_ (.A1(_0551_),
    .A2(_0546_),
    .ZN(_0195_));
 OR3_X1 _0795_ (.A1(_0564_),
    .A2(_0565_),
    .A3(_0552_),
    .ZN(_0196_));
 NOR2_X1 _0796_ (.A1(_0558_),
    .A2(net101),
    .ZN(_0197_));
 AOI211_X2 _0797_ (.A(_0195_),
    .B(_0196_),
    .C1(_0197_),
    .C2(_0002_),
    .ZN(_0198_));
 AND2_X1 _0798_ (.A1(_0551_),
    .A2(_0554_),
    .ZN(_0199_));
 MUX2_X1 _0799_ (.A(_0556_),
    .B(_0199_),
    .S(_0553_),
    .Z(_0200_));
 NAND2_X1 _0800_ (.A1(_0564_),
    .A2(_0565_),
    .ZN(_0201_));
 OR2_X1 _0801_ (.A1(_0566_),
    .A2(net101),
    .ZN(_0202_));
 NOR3_X2 _0802_ (.A1(_0568_),
    .A2(_0201_),
    .A3(_0202_),
    .ZN(_0203_));
 AOI21_X4 _0803_ (.A(_0198_),
    .B1(_0200_),
    .B2(_0203_),
    .ZN(_0204_));
 XOR2_X2 _0804_ (.A(_0557_),
    .B(_0003_),
    .Z(_0205_));
 NAND3_X1 _0805_ (.A1(_0108_),
    .A2(_0022_),
    .A3(_0205_),
    .ZN(_0206_));
 NAND3_X1 _0806_ (.A1(net63),
    .A2(_0106_),
    .A3(_0018_),
    .ZN(_0207_));
 NAND2_X1 _0807_ (.A1(_0206_),
    .A2(_0207_),
    .ZN(_0208_));
 OAI21_X1 _0808_ (.A(_0162_),
    .B1(_0208_),
    .B2(_0190_),
    .ZN(_0209_));
 MUX2_X1 _0809_ (.A(net9),
    .B(_0022_),
    .S(_0205_),
    .Z(_0210_));
 MUX2_X1 _0810_ (.A(_0018_),
    .B(_0146_),
    .S(_0019_),
    .Z(_0211_));
 MUX2_X1 _0811_ (.A(_0210_),
    .B(_0211_),
    .S(_0038_),
    .Z(_0212_));
 OAI21_X1 _0812_ (.A(_0204_),
    .B1(_0212_),
    .B2(_0190_),
    .ZN(_0213_));
 OAI22_X2 _0813_ (.A1(_0204_),
    .A2(_0209_),
    .B1(_0213_),
    .B2(net79),
    .ZN(_0214_));
 AOI21_X1 _0814_ (.A(_0141_),
    .B1(_0108_),
    .B2(_0047_),
    .ZN(_0215_));
 INV_X1 _0815_ (.A(net21),
    .ZN(_0216_));
 AOI211_X2 _0816_ (.A(net91),
    .B(_0216_),
    .C1(_0043_),
    .C2(_0008_),
    .ZN(_0217_));
 INV_X1 _0817_ (.A(_0138_),
    .ZN(_0218_));
 NOR4_X2 _0818_ (.A1(_0076_),
    .A2(net1),
    .A3(_0040_),
    .A4(_0218_),
    .ZN(_0219_));
 NAND2_X1 _0819_ (.A1(_0040_),
    .A2(net21),
    .ZN(_0220_));
 NOR3_X2 _0820_ (.A1(_0076_),
    .A2(_0038_),
    .A3(_0220_),
    .ZN(_0221_));
 OR4_X4 _0821_ (.A1(_0215_),
    .A2(_0217_),
    .A3(_0219_),
    .A4(_0221_),
    .ZN(_0222_));
 AOI21_X1 _0822_ (.A(_0089_),
    .B1(_0026_),
    .B2(_0047_),
    .ZN(_0223_));
 INV_X1 _0823_ (.A(net23),
    .ZN(_0224_));
 AOI211_X2 _0824_ (.A(net91),
    .B(_0224_),
    .C1(_0561_),
    .C2(_0008_),
    .ZN(_0225_));
 AND4_X1 _0825_ (.A1(_0043_),
    .A2(_0008_),
    .A3(_0004_),
    .A4(_0086_),
    .ZN(_0226_));
 AND3_X1 _0826_ (.A1(_0043_),
    .A2(_0008_),
    .A3(_0136_),
    .ZN(_0227_));
 OR4_X4 _0827_ (.A1(_0223_),
    .A2(_0225_),
    .A3(_0226_),
    .A4(_0227_),
    .ZN(_0228_));
 OAI22_X2 _0828_ (.A1(_0128_),
    .A2(_0222_),
    .B1(_0228_),
    .B2(_0144_),
    .ZN(_0229_));
 AOI21_X2 _0829_ (.A(_0110_),
    .B1(_0027_),
    .B2(_0044_),
    .ZN(_0230_));
 INV_X1 _0830_ (.A(net22),
    .ZN(_0231_));
 AOI211_X2 _0831_ (.A(_0040_),
    .B(_0231_),
    .C1(_0043_),
    .C2(_0026_),
    .ZN(_0232_));
 INV_X1 _0832_ (.A(net24),
    .ZN(_0233_));
 NOR4_X2 _0833_ (.A1(_0049_),
    .A2(_0038_),
    .A3(_0020_),
    .A4(_0233_),
    .ZN(_0234_));
 AND3_X1 _0834_ (.A1(_0047_),
    .A2(_0026_),
    .A3(_0149_),
    .ZN(_0235_));
 NOR4_X4 _0835_ (.A1(_0235_),
    .A2(_0232_),
    .A3(_0234_),
    .A4(_0230_),
    .ZN(_0236_));
 INV_X1 _0836_ (.A(net20),
    .ZN(_0237_));
 NOR3_X2 _0837_ (.A1(_0237_),
    .A2(_0059_),
    .A3(_0060_),
    .ZN(_0238_));
 INV_X1 _0838_ (.A(_0151_),
    .ZN(_0239_));
 AOI21_X2 _0839_ (.A(_0239_),
    .B1(_0013_),
    .B2(_0015_),
    .ZN(_0240_));
 NOR2_X2 _0840_ (.A1(_0238_),
    .A2(_0240_),
    .ZN(_0241_));
 AOI221_X2 _0841_ (.A(_0229_),
    .B1(net74),
    .B2(_0125_),
    .C1(_0037_),
    .C2(_0241_),
    .ZN(_0242_));
 NOR2_X4 _0842_ (.A1(net75),
    .A2(_0176_),
    .ZN(_0243_));
 AOI22_X2 _0843_ (.A1(_0194_),
    .A2(_0214_),
    .B1(_0242_),
    .B2(_0243_),
    .ZN(_0244_));
 OAI21_X1 _0844_ (.A(_0189_),
    .B1(_0244_),
    .B2(_0082_),
    .ZN(net26));
 NOR2_X4 _0845_ (.A1(_0026_),
    .A2(_0041_),
    .ZN(_0245_));
 NAND2_X1 _0846_ (.A1(_0044_),
    .A2(_0245_),
    .ZN(_0246_));
 NAND2_X1 _0847_ (.A1(_0551_),
    .A2(_0002_),
    .ZN(_0247_));
 MUX2_X1 _0848_ (.A(_0002_),
    .B(_0247_),
    .S(_0553_),
    .Z(_0248_));
 OR2_X1 _0849_ (.A1(_0076_),
    .A2(_0020_),
    .ZN(_0249_));
 NOR2_X1 _0850_ (.A1(_0556_),
    .A2(_0249_),
    .ZN(_0250_));
 OAI33_X1 _0851_ (.A1(_0246_),
    .A2(_0201_),
    .A3(_0248_),
    .B1(_0250_),
    .B2(_0195_),
    .B3(_0196_),
    .ZN(_0251_));
 BUF_X4 _0852_ (.A(net57),
    .Z(_0252_));
 MUX2_X1 _0853_ (.A(net17),
    .B(net19),
    .S(_0041_),
    .Z(_0253_));
 AND3_X1 _0854_ (.A1(_0123_),
    .A2(_0124_),
    .A3(_0253_),
    .ZN(_0254_));
 AOI21_X1 _0855_ (.A(_0133_),
    .B1(_0022_),
    .B2(_0106_),
    .ZN(_0255_));
 AOI21_X1 _0856_ (.A(_0255_),
    .B1(_0124_),
    .B2(_0123_),
    .ZN(_0256_));
 OAI21_X1 _0857_ (.A(net64),
    .B1(_0254_),
    .B2(_0256_),
    .ZN(_0257_));
 MUX2_X1 _0858_ (.A(_0146_),
    .B(net20),
    .S(net73),
    .Z(_0258_));
 NAND4_X1 _0859_ (.A1(_0118_),
    .A2(_0000_),
    .A3(_0556_),
    .A4(_0021_),
    .ZN(_0259_));
 NAND4_X1 _0860_ (.A1(_0118_),
    .A2(_0553_),
    .A3(_0002_),
    .A4(_0021_),
    .ZN(_0260_));
 MUX2_X1 _0861_ (.A(_0018_),
    .B(net18),
    .S(_0041_),
    .Z(_0261_));
 NAND2_X1 _0862_ (.A1(_0161_),
    .A2(_0261_),
    .ZN(_0262_));
 NAND3_X1 _0863_ (.A1(_0259_),
    .A2(_0260_),
    .A3(_0262_),
    .ZN(_0263_));
 AOI22_X2 _0864_ (.A1(_0100_),
    .A2(_0258_),
    .B1(_0263_),
    .B2(_0178_),
    .ZN(_0264_));
 AOI21_X2 _0865_ (.A(net89),
    .B1(_0257_),
    .B2(_0264_),
    .ZN(_0265_));
 NAND4_X4 _0866_ (.A1(_0152_),
    .A2(_0150_),
    .A3(_0153_),
    .A4(_0155_),
    .ZN(_0266_));
 NAND3_X4 _0867_ (.A1(_0104_),
    .A2(_0030_),
    .A3(_0031_),
    .ZN(_0267_));
 OAI22_X4 _0868_ (.A1(_0128_),
    .A2(net103),
    .B1(_0222_),
    .B2(_0267_),
    .ZN(_0268_));
 OAI21_X4 _0869_ (.A(net63),
    .B1(net80),
    .B2(_0562_),
    .ZN(_0269_));
 NOR2_X2 _0870_ (.A1(_0269_),
    .A2(_0228_),
    .ZN(_0270_));
 NAND4_X2 _0871_ (.A1(_0105_),
    .A2(_0107_),
    .A3(_0109_),
    .A4(_0111_),
    .ZN(_0271_));
 NOR2_X2 _0872_ (.A1(_0144_),
    .A2(_0271_),
    .ZN(_0272_));
 NOR4_X4 _0873_ (.A1(_0268_),
    .A2(_0176_),
    .A3(_0270_),
    .A4(_0272_),
    .ZN(_0273_));
 BUF_X4 _0874_ (.A(_0164_),
    .Z(_0274_));
 AOI211_X2 _0875_ (.A(_0252_),
    .B(_0265_),
    .C1(_0273_),
    .C2(_0274_),
    .ZN(_0275_));
 XNOR2_X2 _0876_ (.A(_0564_),
    .B(_0080_),
    .ZN(_0276_));
 CLKBUF_X3 _0877_ (.A(_0276_),
    .Z(_0277_));
 NAND2_X1 _0878_ (.A1(_0178_),
    .A2(_0263_),
    .ZN(_0278_));
 NAND2_X1 _0879_ (.A1(_0106_),
    .A2(_0022_),
    .ZN(_0279_));
 AOI21_X1 _0880_ (.A(_0279_),
    .B1(_0124_),
    .B2(_0123_),
    .ZN(_0280_));
 OAI21_X1 _0881_ (.A(net64),
    .B1(_0254_),
    .B2(_0280_),
    .ZN(_0281_));
 AOI21_X1 _0882_ (.A(_0274_),
    .B1(_0278_),
    .B2(_0281_),
    .ZN(_0282_));
 NAND4_X4 _0883_ (.A1(_0044_),
    .A2(_0553_),
    .A3(_0556_),
    .A4(_0160_),
    .ZN(_0283_));
 NAND2_X1 _0884_ (.A1(_0252_),
    .A2(_0283_),
    .ZN(_0284_));
 OAI21_X1 _0885_ (.A(_0277_),
    .B1(_0282_),
    .B2(_0284_),
    .ZN(_0285_));
 MUX2_X1 _0886_ (.A(net13),
    .B(net14),
    .S(_0026_),
    .Z(_0286_));
 OR3_X1 _0887_ (.A1(_0059_),
    .A2(_0060_),
    .A3(_0286_),
    .ZN(_0287_));
 NAND2_X1 _0888_ (.A1(net62),
    .A2(net15),
    .ZN(_0288_));
 INV_X1 _0889_ (.A(net16),
    .ZN(_0289_));
 OAI221_X2 _0890_ (.A(_0288_),
    .B1(_0060_),
    .B2(_0059_),
    .C1(_0550_),
    .C2(_0289_),
    .ZN(_0290_));
 NAND3_X2 _0891_ (.A1(_0033_),
    .A2(_0287_),
    .A3(_0290_),
    .ZN(_0291_));
 MUX2_X1 _0892_ (.A(_0050_),
    .B(_0056_),
    .S(_0108_),
    .Z(_0292_));
 AND2_X1 _0893_ (.A1(_0008_),
    .A2(net12),
    .ZN(_0293_));
 AOI21_X1 _0894_ (.A(_0293_),
    .B1(net11),
    .B2(_0549_),
    .ZN(_0294_));
 MUX2_X1 _0895_ (.A(_0292_),
    .B(_0294_),
    .S(_0016_),
    .Z(_0295_));
 NAND3_X2 _0896_ (.A1(_0030_),
    .A2(_0031_),
    .A3(_0162_),
    .ZN(_0296_));
 OAI211_X2 _0897_ (.A(_0274_),
    .B(_0291_),
    .C1(net94),
    .C2(_0296_),
    .ZN(_0297_));
 NAND2_X1 _0898_ (.A1(net62),
    .A2(_0113_),
    .ZN(_0298_));
 NOR3_X1 _0899_ (.A1(_0094_),
    .A2(_0560_),
    .A3(_0563_),
    .ZN(_0299_));
 AOI21_X1 _0900_ (.A(_0046_),
    .B1(_0123_),
    .B2(_0124_),
    .ZN(_0300_));
 NOR3_X1 _0901_ (.A1(_0298_),
    .A2(_0299_),
    .A3(_0300_),
    .ZN(_0301_));
 NAND2_X1 _0902_ (.A1(_0000_),
    .A2(_0035_),
    .ZN(_0302_));
 AOI21_X2 _0903_ (.A(_0302_),
    .B1(_0556_),
    .B2(_0076_),
    .ZN(_0303_));
 AOI211_X2 _0904_ (.A(_0552_),
    .B(_0116_),
    .C1(_0556_),
    .C2(_0558_),
    .ZN(_0304_));
 INV_X1 _0905_ (.A(_0035_),
    .ZN(_0305_));
 NOR4_X2 _0906_ (.A1(_0043_),
    .A2(_0000_),
    .A3(_0002_),
    .A4(_0305_),
    .ZN(_0306_));
 NOR4_X2 _0907_ (.A1(_0043_),
    .A2(_0553_),
    .A3(_0002_),
    .A4(_0116_),
    .ZN(_0307_));
 NOR4_X4 _0908_ (.A1(_0303_),
    .A2(_0304_),
    .A3(_0306_),
    .A4(_0307_),
    .ZN(_0308_));
 NOR2_X1 _0909_ (.A1(_0104_),
    .A2(_0024_),
    .ZN(_0309_));
 AND2_X1 _0910_ (.A1(_0308_),
    .A2(_0309_),
    .ZN(_0310_));
 OAI21_X2 _0911_ (.A(_0249_),
    .B1(_0078_),
    .B2(_0106_),
    .ZN(_0311_));
 INV_X1 _0912_ (.A(net7),
    .ZN(_0312_));
 MUX2_X1 _0913_ (.A(_0119_),
    .B(_0312_),
    .S(_0000_),
    .Z(_0313_));
 NAND3_X1 _0914_ (.A1(_0178_),
    .A2(_0311_),
    .A3(_0313_),
    .ZN(_0314_));
 MUX2_X1 _0915_ (.A(net7),
    .B(net4),
    .S(_0000_),
    .Z(_0315_));
 NAND4_X1 _0916_ (.A1(_0118_),
    .A2(_0178_),
    .A3(_0556_),
    .A4(_0113_),
    .ZN(_0316_));
 OAI21_X1 _0917_ (.A(_0314_),
    .B1(_0315_),
    .B2(_0316_),
    .ZN(_0317_));
 AOI21_X1 _0918_ (.A(_0096_),
    .B1(_0030_),
    .B2(_0031_),
    .ZN(_0318_));
 AOI211_X2 _0919_ (.A(_0202_),
    .B(_0318_),
    .C1(_0083_),
    .C2(_0174_),
    .ZN(_0319_));
 NOR4_X2 _0920_ (.A1(_0301_),
    .A2(_0310_),
    .A3(_0317_),
    .A4(_0319_),
    .ZN(_0320_));
 OAI21_X1 _0921_ (.A(_0297_),
    .B1(_0320_),
    .B2(_0166_),
    .ZN(_0321_));
 CLKBUF_X3 _0922_ (.A(_0277_),
    .Z(_0322_));
 OAI22_X1 _0923_ (.A1(_0275_),
    .A2(_0285_),
    .B1(_0321_),
    .B2(_0322_),
    .ZN(net27));
 INV_X1 _0924_ (.A(_0009_),
    .ZN(_0323_));
 OAI22_X1 _0925_ (.A1(_0190_),
    .A2(_0323_),
    .B1(_0058_),
    .B2(_0296_),
    .ZN(_0324_));
 MUX2_X1 _0926_ (.A(_0010_),
    .B(_0054_),
    .S(_0174_),
    .Z(_0325_));
 NOR2_X1 _0927_ (.A1(_0176_),
    .A2(_0061_),
    .ZN(_0326_));
 AOI22_X1 _0928_ (.A1(_0061_),
    .A2(_0324_),
    .B1(_0325_),
    .B2(_0326_),
    .ZN(_0327_));
 AOI22_X2 _0929_ (.A1(_0039_),
    .A2(net60),
    .B1(_0037_),
    .B2(_0122_),
    .ZN(_0328_));
 OAI221_X2 _0930_ (.A(_0328_),
    .B1(_0269_),
    .B2(_0036_),
    .C1(_0053_),
    .C2(_0144_),
    .ZN(_0329_));
 MUX2_X1 _0931_ (.A(_0327_),
    .B(_0329_),
    .S(_0074_),
    .Z(_0330_));
 NAND2_X4 _0932_ (.A1(_0276_),
    .A2(_0204_),
    .ZN(_0331_));
 CLKBUF_X3 _0933_ (.A(_0331_),
    .Z(_0332_));
 NOR2_X1 _0934_ (.A1(_0027_),
    .A2(_0147_),
    .ZN(_0333_));
 AOI21_X1 _0935_ (.A(_0333_),
    .B1(_0124_),
    .B2(_0123_),
    .ZN(_0334_));
 NAND4_X2 _0936_ (.A1(_0130_),
    .A2(_0131_),
    .A3(_0132_),
    .A4(_0134_),
    .ZN(_0335_));
 OAI21_X1 _0937_ (.A(_0334_),
    .B1(_0335_),
    .B2(net64),
    .ZN(_0336_));
 NAND2_X1 _0938_ (.A1(_0007_),
    .A2(_0029_),
    .ZN(_0337_));
 AOI21_X1 _0939_ (.A(_0165_),
    .B1(_0336_),
    .B2(_0337_),
    .ZN(_0338_));
 MUX2_X1 _0940_ (.A(_0271_),
    .B(_0266_),
    .S(_0174_),
    .Z(_0339_));
 NAND4_X1 _0941_ (.A1(_0085_),
    .A2(_0087_),
    .A3(_0088_),
    .A4(_0090_),
    .ZN(_0340_));
 NAND4_X2 _0942_ (.A1(_0137_),
    .A2(_0139_),
    .A3(_0140_),
    .A4(_0142_),
    .ZN(_0341_));
 MUX2_X1 _0943_ (.A(_0340_),
    .B(_0341_),
    .S(_0174_),
    .Z(_0342_));
 MUX2_X1 _0944_ (.A(_0339_),
    .B(_0342_),
    .S(_0178_),
    .Z(_0343_));
 AOI21_X1 _0945_ (.A(_0338_),
    .B1(_0343_),
    .B2(_0243_),
    .ZN(_0344_));
 OAI22_X1 _0946_ (.A1(_0322_),
    .A2(_0330_),
    .B1(_0332_),
    .B2(_0344_),
    .ZN(net28));
 AND3_X1 _0947_ (.A1(_0013_),
    .A2(_0015_),
    .A3(_0294_),
    .ZN(_0345_));
 AOI21_X2 _0948_ (.A(_0286_),
    .B1(_0015_),
    .B2(net81),
    .ZN(_0346_));
 NOR3_X2 _0949_ (.A1(_0033_),
    .A2(_0345_),
    .A3(_0346_),
    .ZN(_0347_));
 MUX2_X1 _0950_ (.A(net15),
    .B(net17),
    .S(_0041_),
    .Z(_0348_));
 MUX2_X1 _0951_ (.A(net16),
    .B(net18),
    .S(_0024_),
    .Z(_0349_));
 MUX2_X1 _0952_ (.A(_0348_),
    .B(_0349_),
    .S(_0028_),
    .Z(_0350_));
 AND2_X4 _0953_ (.A1(_0033_),
    .A2(_0350_),
    .ZN(_0351_));
 NOR3_X4 _0954_ (.A1(_0351_),
    .A2(_0347_),
    .A3(net99),
    .ZN(_0352_));
 AOI21_X1 _0955_ (.A(_0181_),
    .B1(_0028_),
    .B2(_0044_),
    .ZN(_0353_));
 AOI211_X2 _0956_ (.A(_0113_),
    .B(_0119_),
    .C1(_0044_),
    .C2(_0027_),
    .ZN(_0354_));
 NOR4_X2 _0957_ (.A1(_0118_),
    .A2(net62),
    .A3(_0113_),
    .A4(_0305_),
    .ZN(_0355_));
 NOR3_X1 _0958_ (.A1(_0118_),
    .A2(net65),
    .A3(_0114_),
    .ZN(_0356_));
 NOR4_X2 _0959_ (.A1(_0353_),
    .A2(_0354_),
    .A3(_0355_),
    .A4(_0356_),
    .ZN(_0357_));
 NAND2_X1 _0960_ (.A1(_0113_),
    .A2(net10),
    .ZN(_0358_));
 AOI21_X1 _0961_ (.A(_0358_),
    .B1(_0028_),
    .B2(_0044_),
    .ZN(_0359_));
 AOI211_X2 _0962_ (.A(_0041_),
    .B(_0312_),
    .C1(_0044_),
    .C2(_0027_),
    .ZN(_0360_));
 NOR4_X2 _0963_ (.A1(_0118_),
    .A2(net65),
    .A3(_0113_),
    .A4(_0056_),
    .ZN(_0361_));
 NOR4_X2 _0964_ (.A1(_0118_),
    .A2(net65),
    .A3(_0106_),
    .A4(_0312_),
    .ZN(_0362_));
 NOR4_X2 _0965_ (.A1(_0359_),
    .A2(_0360_),
    .A3(_0361_),
    .A4(_0362_),
    .ZN(_0363_));
 AOI22_X2 _0966_ (.A1(_0039_),
    .A2(_0357_),
    .B1(_0363_),
    .B2(_0100_),
    .ZN(_0364_));
 NOR4_X2 _0967_ (.A1(_0045_),
    .A2(_0048_),
    .A3(_0051_),
    .A4(_0052_),
    .ZN(_0365_));
 AOI22_X2 _0968_ (.A1(_0037_),
    .A2(net61),
    .B1(_0125_),
    .B2(_0365_),
    .ZN(_0366_));
 AOI21_X1 _0969_ (.A(_0165_),
    .B1(_0364_),
    .B2(_0366_),
    .ZN(_0367_));
 NAND4_X1 _0970_ (.A1(_0138_),
    .A2(_0123_),
    .A3(_0124_),
    .A4(_0245_),
    .ZN(_0368_));
 NAND2_X1 _0971_ (.A1(_0086_),
    .A2(_0245_),
    .ZN(_0369_));
 OAI221_X2 _0972_ (.A(_0368_),
    .B1(_0236_),
    .B2(_0128_),
    .C1(_0190_),
    .C2(_0369_),
    .ZN(_0370_));
 NAND3_X1 _0973_ (.A1(net23),
    .A2(_0030_),
    .A3(_0031_),
    .ZN(_0371_));
 OAI21_X1 _0974_ (.A(_0083_),
    .B1(_0560_),
    .B2(_0563_),
    .ZN(_0372_));
 AOI21_X2 _0975_ (.A(_0298_),
    .B1(_0371_),
    .B2(_0372_),
    .ZN(_0373_));
 NAND3_X1 _0976_ (.A1(_0102_),
    .A2(net81),
    .A3(_0015_),
    .ZN(_0374_));
 OAI21_X1 _0977_ (.A(net2),
    .B1(_0059_),
    .B2(_0060_),
    .ZN(_0375_));
 AOI21_X2 _0978_ (.A(_0144_),
    .B1(_0374_),
    .B2(_0375_),
    .ZN(_0376_));
 NOR4_X2 _0979_ (.A1(_0073_),
    .A2(_0370_),
    .A3(_0373_),
    .A4(_0376_),
    .ZN(_0377_));
 MUX2_X1 _0980_ (.A(_0146_),
    .B(_0018_),
    .S(net66),
    .Z(_0378_));
 MUX2_X1 _0981_ (.A(net20),
    .B(_0151_),
    .S(_0024_),
    .Z(_0379_));
 AOI22_X1 _0982_ (.A1(_0039_),
    .A2(_0378_),
    .B1(_0379_),
    .B2(_0100_),
    .ZN(_0380_));
 INV_X1 _0983_ (.A(net9),
    .ZN(_0381_));
 OAI221_X2 _0984_ (.A(_0220_),
    .B1(_0563_),
    .B2(_0560_),
    .C1(_0113_),
    .C2(_0381_),
    .ZN(_0382_));
 MUX2_X1 _0985_ (.A(net19),
    .B(_0022_),
    .S(_0041_),
    .Z(_0383_));
 OAI211_X2 _0986_ (.A(_0550_),
    .B(_0382_),
    .C1(_0383_),
    .C2(_0033_),
    .ZN(_0384_));
 AND3_X4 _0987_ (.A1(_0073_),
    .A2(_0380_),
    .A3(_0384_),
    .ZN(_0385_));
 OAI33_X1 _0988_ (.A1(_0352_),
    .A2(_0277_),
    .A3(_0367_),
    .B1(_0377_),
    .B2(_0385_),
    .B3(_0331_),
    .ZN(_0386_));
 AND2_X1 _0989_ (.A1(_0386_),
    .A2(_0162_),
    .ZN(net29));
 NOR3_X1 _0990_ (.A1(_0059_),
    .A2(_0060_),
    .A3(_0054_),
    .ZN(_0387_));
 AOI21_X1 _0991_ (.A(_0009_),
    .B1(_0014_),
    .B2(_0012_),
    .ZN(_0388_));
 OAI33_X1 _0992_ (.A1(_0193_),
    .A2(_0191_),
    .A3(_0174_),
    .B1(_0387_),
    .B2(_0388_),
    .B3(_0296_),
    .ZN(_0389_));
 NOR2_X1 _0993_ (.A1(_0389_),
    .A2(_0072_),
    .ZN(_0390_));
 NOR2_X1 _0994_ (.A1(_0144_),
    .A2(_0169_),
    .ZN(_0391_));
 MUX2_X1 _0995_ (.A(_0182_),
    .B(_0170_),
    .S(_0032_),
    .Z(_0392_));
 AOI221_X2 _0996_ (.A(_0391_),
    .B1(_0186_),
    .B2(_0039_),
    .C1(_0392_),
    .C2(net64),
    .ZN(_0393_));
 AOI21_X1 _0997_ (.A(_0390_),
    .B1(_0393_),
    .B2(_0074_),
    .ZN(_0394_));
 INV_X1 _0998_ (.A(_0210_),
    .ZN(_0395_));
 MUX2_X1 _0999_ (.A(_0216_),
    .B(_0218_),
    .S(net73),
    .Z(_0396_));
 OAI22_X2 _1000_ (.A1(_0128_),
    .A2(_0395_),
    .B1(_0396_),
    .B2(_0144_),
    .ZN(_0397_));
 OR3_X1 _1001_ (.A1(net80),
    .A2(_0562_),
    .A3(_0211_),
    .ZN(_0398_));
 OAI221_X1 _1002_ (.A(_0154_),
    .B1(_0562_),
    .B2(net80),
    .C1(_0113_),
    .C2(_0237_),
    .ZN(_0399_));
 AND3_X2 _1003_ (.A1(net62),
    .A2(_0398_),
    .A3(_0399_),
    .ZN(_0400_));
 NOR3_X2 _1004_ (.A1(net89),
    .A2(_0397_),
    .A3(_0400_),
    .ZN(_0401_));
 OAI21_X1 _1005_ (.A(_0110_),
    .B1(_0231_),
    .B2(_0041_),
    .ZN(_0402_));
 MUX2_X1 _1006_ (.A(_0179_),
    .B(_0402_),
    .S(_0173_),
    .Z(_0403_));
 AOI222_X2 _1007_ (.A1(_0228_),
    .A2(_0039_),
    .B1(_0185_),
    .B2(_0100_),
    .C1(_0403_),
    .C2(net64),
    .ZN(_0404_));
 AOI211_X2 _1008_ (.A(net59),
    .B(_0401_),
    .C1(net84),
    .C2(net79),
    .ZN(_0405_));
 MUX2_X1 _1009_ (.A(_0394_),
    .B(_0405_),
    .S(_0277_),
    .Z(net30));
 MUX2_X1 _1010_ (.A(_0102_),
    .B(net4),
    .S(_0000_),
    .Z(_0406_));
 AND2_X1 _1011_ (.A1(_0027_),
    .A2(_0406_),
    .ZN(_0407_));
 MUX2_X1 _1012_ (.A(net4),
    .B(_0102_),
    .S(_0000_),
    .Z(_0408_));
 NOR4_X1 _1013_ (.A1(_0047_),
    .A2(net63),
    .A3(_0002_),
    .A4(_0005_),
    .ZN(_0409_));
 AOI22_X1 _1014_ (.A1(_0311_),
    .A2(_0407_),
    .B1(_0408_),
    .B2(_0409_),
    .ZN(_0410_));
 NOR3_X1 _1015_ (.A1(_0104_),
    .A2(_0116_),
    .A3(net73),
    .ZN(_0411_));
 OAI21_X1 _1016_ (.A(_0411_),
    .B1(_0563_),
    .B2(_0560_),
    .ZN(_0412_));
 NOR3_X1 _1017_ (.A1(_0104_),
    .A2(_0233_),
    .A3(net73),
    .ZN(_0413_));
 NAND3_X1 _1018_ (.A1(_0030_),
    .A2(_0031_),
    .A3(_0413_),
    .ZN(_0414_));
 NAND3_X1 _1019_ (.A1(_0410_),
    .A2(_0412_),
    .A3(_0414_),
    .ZN(_0415_));
 MUX2_X1 _1020_ (.A(_0086_),
    .B(net3),
    .S(_0032_),
    .Z(_0416_));
 INV_X1 _1021_ (.A(_0298_),
    .ZN(_0417_));
 NAND2_X1 _1022_ (.A1(_0371_),
    .A2(_0372_),
    .ZN(_0418_));
 AOI221_X2 _1023_ (.A(_0415_),
    .B1(_0416_),
    .B2(_0417_),
    .C1(_0245_),
    .C2(_0418_),
    .ZN(_0419_));
 NAND3_X1 _1024_ (.A1(_0123_),
    .A2(_0124_),
    .A3(_0255_),
    .ZN(_0420_));
 OAI211_X2 _1025_ (.A(_0550_),
    .B(_0420_),
    .C1(_0222_),
    .C2(_0190_),
    .ZN(_0421_));
 AOI22_X2 _1026_ (.A1(_0100_),
    .A2(net102),
    .B1(_0258_),
    .B2(_0039_),
    .ZN(_0422_));
 AND2_X1 _1027_ (.A1(_0421_),
    .A2(_0422_),
    .ZN(_0423_));
 MUX2_X1 _1028_ (.A(_0419_),
    .B(_0423_),
    .S(_0073_),
    .Z(_0424_));
 MUX2_X1 _1029_ (.A(net6),
    .B(net7),
    .S(_0108_),
    .Z(_0425_));
 AOI21_X1 _1030_ (.A(_0425_),
    .B1(_0015_),
    .B2(_0013_),
    .ZN(_0426_));
 MUX2_X1 _1031_ (.A(net5),
    .B(_0035_),
    .S(_0108_),
    .Z(_0427_));
 NOR3_X1 _1032_ (.A1(_0059_),
    .A2(_0060_),
    .A3(_0427_),
    .ZN(_0428_));
 OR2_X1 _1033_ (.A1(_0426_),
    .A2(_0428_),
    .ZN(_0429_));
 MUX2_X1 _1034_ (.A(_0295_),
    .B(_0429_),
    .S(_0190_),
    .Z(_0430_));
 AND3_X1 _1035_ (.A1(_0190_),
    .A2(_0287_),
    .A3(_0290_),
    .ZN(_0431_));
 OAI22_X1 _1036_ (.A1(_0560_),
    .A2(_0563_),
    .B1(_0253_),
    .B2(_0028_),
    .ZN(_0432_));
 OR2_X1 _1037_ (.A1(_0018_),
    .A2(_0205_),
    .ZN(_0433_));
 OAI21_X1 _1038_ (.A(_0433_),
    .B1(net73),
    .B2(net18),
    .ZN(_0434_));
 AOI21_X1 _1039_ (.A(_0432_),
    .B1(_0434_),
    .B2(_0178_),
    .ZN(_0435_));
 OAI21_X1 _1040_ (.A(_0162_),
    .B1(_0431_),
    .B2(_0435_),
    .ZN(_0436_));
 MUX2_X1 _1041_ (.A(_0430_),
    .B(_0436_),
    .S(net79),
    .Z(_0437_));
 OAI22_X1 _1042_ (.A1(_0332_),
    .A2(_0424_),
    .B1(_0437_),
    .B2(_0322_),
    .ZN(net31));
 OAI22_X1 _1043_ (.A1(_0075_),
    .A2(_0322_),
    .B1(_0159_),
    .B2(_0332_),
    .ZN(net32));
 OR3_X1 _1044_ (.A1(_0102_),
    .A2(_0559_),
    .A3(_0562_),
    .ZN(_0438_));
 OAI21_X1 _1045_ (.A(_0119_),
    .B1(net78),
    .B2(_0562_),
    .ZN(_0439_));
 AND3_X1 _1046_ (.A1(_0309_),
    .A2(_0438_),
    .A3(_0439_),
    .ZN(_0440_));
 NOR3_X2 _1047_ (.A1(net62),
    .A2(_0061_),
    .A3(_0308_),
    .ZN(_0441_));
 OAI22_X4 _1048_ (.A1(_0267_),
    .A2(_0091_),
    .B1(_0099_),
    .B2(_0269_),
    .ZN(_0442_));
 NOR3_X1 _1049_ (.A1(_0440_),
    .A2(_0441_),
    .A3(_0442_),
    .ZN(_0443_));
 NOR3_X1 _1050_ (.A1(_0231_),
    .A2(_0059_),
    .A3(_0060_),
    .ZN(_0444_));
 AOI21_X1 _1051_ (.A(_0233_),
    .B1(_0013_),
    .B2(_0015_),
    .ZN(_0445_));
 OAI33_X1 _1052_ (.A1(_0128_),
    .A2(_0238_),
    .A3(_0240_),
    .B1(_0444_),
    .B2(_0144_),
    .B3(_0445_),
    .ZN(_0446_));
 OAI22_X2 _1053_ (.A1(_0267_),
    .A2(_0335_),
    .B1(_0341_),
    .B2(_0269_),
    .ZN(_0447_));
 OR2_X1 _1054_ (.A1(_0446_),
    .A2(_0447_),
    .ZN(_0448_));
 MUX2_X1 _1055_ (.A(_0443_),
    .B(_0448_),
    .S(_0074_),
    .Z(_0449_));
 AOI22_X2 _1056_ (.A1(_0039_),
    .A2(_0349_),
    .B1(_0378_),
    .B2(_0100_),
    .ZN(_0450_));
 NOR3_X2 _1057_ (.A1(_0348_),
    .A2(_0563_),
    .A3(_0560_),
    .ZN(_0451_));
 AOI21_X2 _1058_ (.A(_0383_),
    .B1(_0031_),
    .B2(_0030_),
    .ZN(_0452_));
 OR3_X4 _1059_ (.A1(_0451_),
    .A2(_0178_),
    .A3(_0452_),
    .ZN(_0453_));
 AND2_X1 _1060_ (.A1(_0450_),
    .A2(_0453_),
    .ZN(_0454_));
 NOR3_X1 _1061_ (.A1(_0174_),
    .A2(_0345_),
    .A3(_0346_),
    .ZN(_0455_));
 NAND3_X1 _1062_ (.A1(net81),
    .A2(_0015_),
    .A3(_0425_),
    .ZN(_0456_));
 OAI21_X1 _1063_ (.A(_0456_),
    .B1(_0292_),
    .B2(_0061_),
    .ZN(_0457_));
 AOI21_X2 _1064_ (.A(_0455_),
    .B1(_0457_),
    .B2(_0190_),
    .ZN(_0458_));
 MUX2_X1 _1065_ (.A(_0454_),
    .B(_0458_),
    .S(_0074_),
    .Z(_0459_));
 OAI22_X1 _1066_ (.A1(_0332_),
    .A2(_0449_),
    .B1(_0459_),
    .B2(_0163_),
    .ZN(net33));
 OAI21_X1 _1067_ (.A(_0167_),
    .B1(_0175_),
    .B2(_0176_),
    .ZN(_0460_));
 NOR2_X1 _1068_ (.A1(_0191_),
    .A2(_0193_),
    .ZN(_0461_));
 MUX2_X1 _1069_ (.A(_0208_),
    .B(_0212_),
    .S(_0204_),
    .Z(_0462_));
 MUX2_X1 _1070_ (.A(_0461_),
    .B(_0462_),
    .S(_0033_),
    .Z(_0463_));
 AOI22_X1 _1071_ (.A1(_0074_),
    .A2(_0460_),
    .B1(_0463_),
    .B2(_0243_),
    .ZN(_0464_));
 NAND3_X1 _1072_ (.A1(_0274_),
    .A2(_0184_),
    .A3(_0187_),
    .ZN(_0465_));
 OAI211_X2 _1073_ (.A(_0162_),
    .B(_0465_),
    .C1(_0242_),
    .C2(_0166_),
    .ZN(_0466_));
 OAI22_X1 _1074_ (.A1(_0322_),
    .A2(_0464_),
    .B1(_0466_),
    .B2(_0332_),
    .ZN(net34));
 NOR4_X2 _1075_ (.A1(_0274_),
    .A2(_0268_),
    .A3(_0270_),
    .A4(_0272_),
    .ZN(_0467_));
 AOI21_X2 _1076_ (.A(_0467_),
    .B1(_0320_),
    .B2(_0166_),
    .ZN(_0468_));
 NAND3_X1 _1077_ (.A1(_0166_),
    .A2(_0257_),
    .A3(_0264_),
    .ZN(_0469_));
 OAI211_X2 _1078_ (.A(_0074_),
    .B(_0291_),
    .C1(net94),
    .C2(_0033_),
    .ZN(_0470_));
 NAND3_X1 _1079_ (.A1(_0162_),
    .A2(_0469_),
    .A3(_0470_),
    .ZN(_0471_));
 OAI22_X1 _1080_ (.A1(_0332_),
    .A2(_0468_),
    .B1(_0471_),
    .B2(_0322_),
    .ZN(net35));
 OAI22_X1 _1081_ (.A1(_0163_),
    .A2(_0449_),
    .B1(_0459_),
    .B2(_0082_),
    .ZN(net36));
 AOI221_X2 _1082_ (.A(_0333_),
    .B1(_0124_),
    .B2(_0123_),
    .C1(_0178_),
    .C2(_0135_),
    .ZN(_0472_));
 AOI22_X1 _1083_ (.A1(_0007_),
    .A2(_0029_),
    .B1(_0204_),
    .B2(_0472_),
    .ZN(_0473_));
 MUX2_X1 _1084_ (.A(_0327_),
    .B(_0473_),
    .S(_0274_),
    .Z(_0474_));
 MUX2_X1 _1085_ (.A(_0112_),
    .B(_0156_),
    .S(_0174_),
    .Z(_0475_));
 MUX2_X1 _1086_ (.A(_0091_),
    .B(_0143_),
    .S(_0174_),
    .Z(_0476_));
 MUX2_X1 _1087_ (.A(_0475_),
    .B(_0476_),
    .S(_0178_),
    .Z(_0477_));
 MUX2_X1 _1088_ (.A(_0329_),
    .B(_0477_),
    .S(net99),
    .Z(_0478_));
 OAI22_X1 _1089_ (.A1(_0322_),
    .A2(_0474_),
    .B1(_0478_),
    .B2(_0331_),
    .ZN(net37));
 OR2_X4 _1090_ (.A1(_0347_),
    .A2(_0351_),
    .ZN(_0479_));
 AOI21_X1 _1091_ (.A(_0252_),
    .B1(_0380_),
    .B2(_0384_),
    .ZN(_0480_));
 AOI21_X1 _1092_ (.A(_0550_),
    .B1(_0018_),
    .B2(net67),
    .ZN(_0481_));
 NOR2_X1 _1093_ (.A1(_0028_),
    .A2(_0383_),
    .ZN(_0482_));
 NOR2_X1 _1094_ (.A1(_0481_),
    .A2(_0482_),
    .ZN(_0483_));
 NAND3_X1 _1095_ (.A1(_0190_),
    .A2(_0252_),
    .A3(_0483_),
    .ZN(_0484_));
 NAND2_X1 _1096_ (.A1(_0274_),
    .A2(_0484_),
    .ZN(_0485_));
 OAI22_X4 _1097_ (.A1(_0479_),
    .A2(_0166_),
    .B1(_0480_),
    .B2(_0485_),
    .ZN(_0486_));
 AOI21_X1 _1098_ (.A(net99),
    .B1(_0364_),
    .B2(_0366_),
    .ZN(_0487_));
 NOR4_X1 _1099_ (.A1(net79),
    .A2(_0370_),
    .A3(_0373_),
    .A4(_0376_),
    .ZN(_0488_));
 OR2_X1 _1100_ (.A1(_0487_),
    .A2(_0488_),
    .ZN(_0489_));
 OAI22_X1 _1101_ (.A1(_0486_),
    .A2(_0163_),
    .B1(_0489_),
    .B2(_0331_),
    .ZN(net38));
 NOR4_X4 _1102_ (.A1(_0118_),
    .A2(_0000_),
    .A3(_0002_),
    .A4(_0567_),
    .ZN(_0490_));
 NAND3_X1 _1103_ (.A1(_0146_),
    .A2(_0016_),
    .A3(_0490_),
    .ZN(_0491_));
 MUX2_X1 _1104_ (.A(_0393_),
    .B(_0404_),
    .S(_0073_),
    .Z(_0492_));
 OR3_X2 _1105_ (.A1(net58),
    .A2(_0397_),
    .A3(_0400_),
    .ZN(_0493_));
 AOI22_X2 _1106_ (.A1(_0074_),
    .A2(_0389_),
    .B1(_0243_),
    .B2(_0493_),
    .ZN(_0494_));
 OAI221_X1 _1107_ (.A(_0491_),
    .B1(_0492_),
    .B2(_0331_),
    .C1(_0322_),
    .C2(_0494_),
    .ZN(net39));
 NOR2_X1 _1108_ (.A1(_0176_),
    .A2(_0277_),
    .ZN(_0495_));
 OR3_X1 _1109_ (.A1(net79),
    .A2(_0431_),
    .A3(_0435_),
    .ZN(_0496_));
 AND2_X1 _1110_ (.A1(_0022_),
    .A2(_0245_),
    .ZN(_0497_));
 NAND2_X1 _1111_ (.A1(_0252_),
    .A2(_0497_),
    .ZN(_0498_));
 OAI21_X2 _1112_ (.A(_0274_),
    .B1(_0277_),
    .B2(_0498_),
    .ZN(_0499_));
 AOI21_X2 _1113_ (.A(_0252_),
    .B1(_0421_),
    .B2(_0422_),
    .ZN(_0500_));
 OAI211_X2 _1114_ (.A(_0495_),
    .B(_0496_),
    .C1(_0499_),
    .C2(_0500_),
    .ZN(_0501_));
 MUX2_X1 _1115_ (.A(_0419_),
    .B(_0430_),
    .S(_0165_),
    .Z(_0502_));
 NAND2_X1 _1116_ (.A1(_0016_),
    .A2(_0490_),
    .ZN(_0503_));
 OAI221_X1 _1117_ (.A(_0501_),
    .B1(_0502_),
    .B2(_0331_),
    .C1(_0503_),
    .C2(_0381_),
    .ZN(net40));
 MUX2_X1 _1118_ (.A(_0063_),
    .B(_0127_),
    .S(net99),
    .Z(_0504_));
 INV_X1 _1119_ (.A(_0146_),
    .ZN(_0505_));
 MUX2_X1 _1120_ (.A(_0505_),
    .B(_0237_),
    .S(_0016_),
    .Z(_0506_));
 OAI21_X1 _1121_ (.A(_0162_),
    .B1(_0157_),
    .B2(_0145_),
    .ZN(_0507_));
 MUX2_X1 _1122_ (.A(_0034_),
    .B(_0507_),
    .S(_0165_),
    .Z(_0508_));
 OAI222_X2 _1123_ (.A1(_0332_),
    .A2(_0504_),
    .B1(_0506_),
    .B2(_0283_),
    .C1(_0322_),
    .C2(_0508_),
    .ZN(net41));
 AOI22_X2 _1124_ (.A1(_0007_),
    .A2(_0350_),
    .B1(_0483_),
    .B2(_0033_),
    .ZN(_0509_));
 NOR4_X1 _1125_ (.A1(_0176_),
    .A2(_0277_),
    .A3(_0204_),
    .A4(_0509_),
    .ZN(_0510_));
 NOR2_X1 _1126_ (.A1(_0276_),
    .A2(net58),
    .ZN(_0511_));
 OAI21_X1 _1127_ (.A(_0164_),
    .B1(_0446_),
    .B2(_0447_),
    .ZN(_0512_));
 NAND3_X2 _1128_ (.A1(_0072_),
    .A2(_0450_),
    .A3(_0453_),
    .ZN(_0513_));
 AND3_X2 _1129_ (.A1(_0511_),
    .A2(_0512_),
    .A3(_0513_),
    .ZN(_0514_));
 NOR2_X1 _1130_ (.A1(_0135_),
    .A2(_0283_),
    .ZN(_0515_));
 NOR4_X4 _1131_ (.A1(net89),
    .A2(_0440_),
    .A3(_0441_),
    .A4(_0442_),
    .ZN(_0516_));
 AOI211_X2 _1132_ (.A(_0331_),
    .B(_0516_),
    .C1(_0458_),
    .C2(_0164_),
    .ZN(_0517_));
 OR4_X1 _1133_ (.A1(_0510_),
    .A2(_0514_),
    .A3(_0515_),
    .A4(_0517_),
    .ZN(net42));
 NOR2_X1 _1134_ (.A1(_0081_),
    .A2(_0252_),
    .ZN(_0518_));
 NAND3_X1 _1135_ (.A1(_0166_),
    .A2(_0167_),
    .A3(_0175_),
    .ZN(_0519_));
 OAI211_X2 _1136_ (.A(_0518_),
    .B(_0519_),
    .C1(_0166_),
    .C2(_0188_),
    .ZN(_0520_));
 OAI221_X1 _1137_ (.A(_0520_),
    .B1(_0283_),
    .B2(_0241_),
    .C1(_0322_),
    .C2(_0244_),
    .ZN(net43));
 NOR3_X2 _1138_ (.A1(_0176_),
    .A2(_0276_),
    .A3(_0204_),
    .ZN(_0521_));
 NAND2_X1 _1139_ (.A1(_0278_),
    .A2(_0281_),
    .ZN(_0522_));
 AOI22_X2 _1140_ (.A1(_0222_),
    .A2(_0490_),
    .B1(_0521_),
    .B2(_0522_),
    .ZN(_0523_));
 NOR3_X1 _1141_ (.A1(_0074_),
    .A2(_0176_),
    .A3(_0276_),
    .ZN(_0524_));
 AOI22_X2 _1142_ (.A1(_0265_),
    .A2(_0511_),
    .B1(_0524_),
    .B2(_0273_),
    .ZN(_0525_));
 OAI211_X2 _1143_ (.A(_0523_),
    .B(_0525_),
    .C1(_0321_),
    .C2(_0332_),
    .ZN(net44));
 AOI22_X1 _1144_ (.A1(net102),
    .A2(_0490_),
    .B1(_0521_),
    .B2(_0029_),
    .ZN(_0526_));
 NAND2_X2 _1145_ (.A1(_0081_),
    .A2(_0204_),
    .ZN(_0527_));
 OAI221_X1 _1146_ (.A(_0526_),
    .B1(_0527_),
    .B2(_0344_),
    .C1(_0330_),
    .C2(_0332_),
    .ZN(net45));
 OAI33_X1 _1147_ (.A1(_0352_),
    .A2(_0331_),
    .A3(_0367_),
    .B1(_0377_),
    .B2(_0385_),
    .B3(_0527_),
    .ZN(_0528_));
 NAND4_X1 _1148_ (.A1(_0162_),
    .A2(_0081_),
    .A3(_0252_),
    .A4(_0483_),
    .ZN(_0529_));
 OAI21_X1 _1149_ (.A(_0529_),
    .B1(_0283_),
    .B2(_0143_),
    .ZN(_0530_));
 OR2_X1 _1150_ (.A1(_0528_),
    .A2(_0530_),
    .ZN(net46));
 AOI221_X2 _1151_ (.A(_0081_),
    .B1(_0463_),
    .B2(_0243_),
    .C1(_0460_),
    .C2(net99),
    .ZN(_0531_));
 AOI21_X1 _1152_ (.A(_0531_),
    .B1(_0466_),
    .B2(_0082_),
    .ZN(net47));
 AOI211_X2 _1153_ (.A(_0401_),
    .B(_0527_),
    .C1(_0404_),
    .C2(net89),
    .ZN(_0532_));
 AND2_X1 _1154_ (.A1(_0208_),
    .A2(_0521_),
    .ZN(_0533_));
 NOR2_X1 _1155_ (.A1(_0236_),
    .A2(_0283_),
    .ZN(_0534_));
 AOI211_X2 _1156_ (.A(_0331_),
    .B(_0390_),
    .C1(_0393_),
    .C2(_0072_),
    .ZN(_0535_));
 OR4_X2 _1157_ (.A1(_0532_),
    .A2(_0533_),
    .A3(_0534_),
    .A4(_0535_),
    .ZN(net48));
 AOI22_X1 _1158_ (.A1(_0228_),
    .A2(_0490_),
    .B1(_0497_),
    .B2(_0521_),
    .ZN(_0536_));
 OAI221_X1 _1159_ (.A(_0536_),
    .B1(_0527_),
    .B2(_0424_),
    .C1(_0332_),
    .C2(_0437_),
    .ZN(net49));
 OAI22_X1 _1160_ (.A1(_0163_),
    .A2(_0468_),
    .B1(_0471_),
    .B2(_0082_),
    .ZN(net50));
 OAI22_X1 _1161_ (.A1(_0082_),
    .A2(_0474_),
    .B1(_0478_),
    .B2(_0163_),
    .ZN(net51));
 OAI22_X2 _1162_ (.A1(_0486_),
    .A2(_0082_),
    .B1(_0489_),
    .B2(_0163_),
    .ZN(net52));
 OAI22_X1 _1163_ (.A1(_0082_),
    .A2(_0494_),
    .B1(_0492_),
    .B2(_0163_),
    .ZN(net53));
 NAND2_X1 _1164_ (.A1(_0277_),
    .A2(_0496_),
    .ZN(_0537_));
 NOR2_X1 _1165_ (.A1(_0500_),
    .A2(_0499_),
    .ZN(_0538_));
 OAI22_X1 _1166_ (.A1(_0163_),
    .A2(_0502_),
    .B1(_0537_),
    .B2(_0538_),
    .ZN(net54));
 INV_X1 _1167_ (.A(_0243_),
    .ZN(_0539_));
 MUX2_X1 _1168_ (.A(_0063_),
    .B(_0158_),
    .S(_0277_),
    .Z(_0540_));
 MUX2_X1 _1169_ (.A(_0034_),
    .B(_0127_),
    .S(_0081_),
    .Z(_0541_));
 OAI22_X1 _1170_ (.A1(_0539_),
    .A2(_0540_),
    .B1(_0541_),
    .B2(_0166_),
    .ZN(net55));
 MUX2_X1 _1171_ (.A(_0443_),
    .B(_0458_),
    .S(_0274_),
    .Z(_0542_));
 AOI21_X1 _1172_ (.A(_0252_),
    .B1(_0512_),
    .B2(_0513_),
    .ZN(_0543_));
 OAI221_X1 _1173_ (.A(_0252_),
    .B1(_0283_),
    .B2(_0135_),
    .C1(_0509_),
    .C2(_0274_),
    .ZN(_0544_));
 NAND2_X1 _1174_ (.A1(_0277_),
    .A2(_0544_),
    .ZN(_0545_));
 OAI22_X1 _1175_ (.A1(_0163_),
    .A2(_0542_),
    .B1(_0543_),
    .B2(_0545_),
    .ZN(net56));
 HA_X1 _1176_ (.A(_0570_),
    .B(_0550_),
    .CO(_0571_),
    .S(_0572_));
 BUF_X4 clone1 (.A(_0547_),
    .Z(net1));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_59 ();
 BUF_X1 input1 (.A(data_in[12]),
    .Z(net2));
 BUF_X1 input2 (.A(data_in[13]),
    .Z(net3));
 BUF_X1 input3 (.A(data_in[14]),
    .Z(net4));
 BUF_X1 input4 (.A(data_in[15]),
    .Z(net5));
 BUF_X1 input5 (.A(data_in[17]),
    .Z(net6));
 BUF_X1 input6 (.A(data_in[18]),
    .Z(net7));
 BUF_X1 input7 (.A(data_in[19]),
    .Z(net8));
 BUF_X1 input8 (.A(data_in[1]),
    .Z(net9));
 BUF_X1 input9 (.A(data_in[20]),
    .Z(net10));
 BUF_X1 input10 (.A(data_in[21]),
    .Z(net11));
 BUF_X1 input11 (.A(data_in[22]),
    .Z(net12));
 BUF_X1 input12 (.A(data_in[23]),
    .Z(net13));
 BUF_X1 input13 (.A(data_in[24]),
    .Z(net14));
 BUF_X1 input14 (.A(data_in[25]),
    .Z(net15));
 BUF_X1 input15 (.A(data_in[26]),
    .Z(net16));
 BUF_X1 input16 (.A(data_in[27]),
    .Z(net17));
 CLKBUF_X2 input17 (.A(data_in[28]),
    .Z(net18));
 BUF_X1 input18 (.A(data_in[29]),
    .Z(net19));
 BUF_X1 input19 (.A(data_in[2]),
    .Z(net20));
 BUF_X1 input20 (.A(data_in[3]),
    .Z(net21));
 BUF_X1 input21 (.A(data_in[6]),
    .Z(net22));
 BUF_X1 input22 (.A(data_in[7]),
    .Z(net23));
 BUF_X1 input23 (.A(data_in[8]),
    .Z(net24));
 BUF_X1 output24 (.A(net25),
    .Z(data_out[0]));
 BUF_X1 output25 (.A(net26),
    .Z(data_out[10]));
 BUF_X1 output26 (.A(net27),
    .Z(data_out[11]));
 BUF_X1 output27 (.A(net28),
    .Z(data_out[12]));
 BUF_X1 output28 (.A(net29),
    .Z(data_out[13]));
 BUF_X1 output29 (.A(net30),
    .Z(data_out[14]));
 BUF_X1 output30 (.A(net31),
    .Z(data_out[15]));
 BUF_X1 output31 (.A(net32),
    .Z(data_out[16]));
 BUF_X1 output32 (.A(net33),
    .Z(data_out[17]));
 BUF_X1 output33 (.A(net34),
    .Z(data_out[18]));
 BUF_X1 output34 (.A(net35),
    .Z(data_out[19]));
 BUF_X1 output35 (.A(net36),
    .Z(data_out[1]));
 BUF_X1 output36 (.A(net37),
    .Z(data_out[20]));
 BUF_X1 output37 (.A(net38),
    .Z(data_out[21]));
 BUF_X1 output38 (.A(net39),
    .Z(data_out[22]));
 BUF_X1 output39 (.A(net40),
    .Z(data_out[23]));
 BUF_X1 output40 (.A(net41),
    .Z(data_out[24]));
 BUF_X1 output41 (.A(net42),
    .Z(data_out[25]));
 BUF_X1 output42 (.A(net43),
    .Z(data_out[26]));
 BUF_X1 output43 (.A(net44),
    .Z(data_out[27]));
 BUF_X1 output44 (.A(net45),
    .Z(data_out[28]));
 BUF_X1 output45 (.A(net46),
    .Z(data_out[29]));
 BUF_X1 output46 (.A(net47),
    .Z(data_out[2]));
 BUF_X1 output47 (.A(net48),
    .Z(data_out[30]));
 BUF_X1 output48 (.A(net49),
    .Z(data_out[31]));
 BUF_X1 output49 (.A(net50),
    .Z(data_out[3]));
 BUF_X1 output50 (.A(net51),
    .Z(data_out[4]));
 BUF_X1 output51 (.A(net52),
    .Z(data_out[5]));
 BUF_X1 output52 (.A(net53),
    .Z(data_out[6]));
 BUF_X1 output53 (.A(net54),
    .Z(data_out[7]));
 BUF_X1 output54 (.A(net55),
    .Z(data_out[8]));
 BUF_X1 output55 (.A(net56),
    .Z(data_out[9]));
 BUF_X1 rebuffer1 (.A(_0251_),
    .Z(net57));
 BUF_X1 rebuffer2 (.A(_0251_),
    .Z(net58));
 BUF_X1 rebuffer3 (.A(net58),
    .Z(net59));
 BUF_X1 rebuffer4 (.A(_0099_),
    .Z(net60));
 BUF_X1 rebuffer5 (.A(net60),
    .Z(net61));
 BUF_X16 clone6 (.A(net63),
    .Z(net62));
 BUF_X16 clone7 (.A(_0548_),
    .Z(net63));
 BUF_X16 clone8 (.A(net65),
    .Z(net64));
 BUF_X1 rebuffer9 (.A(_0550_),
    .Z(net65));
 BUF_X8 clone35 (.A(_0003_),
    .Z(net101));
 BUF_X2 rebuffer17 (.A(_0023_),
    .Z(net73));
 BUF_X1 rebuffer18 (.A(_0236_),
    .Z(net74));
 BUF_X1 rebuffer19 (.A(_0072_),
    .Z(net75));
 BUF_X2 clone23 (.A(_0164_),
    .Z(net79));
 BUF_X2 rebuffer28 (.A(_0404_),
    .Z(net84));
 XNOR2_X1 clone33 (.A(_0565_),
    .B(_0071_),
    .ZN(net89));
 BUF_X8 clone43 (.A(net100),
    .Z(net99));
 BUF_X2 rebuffer44 (.A(_0072_),
    .Z(net100));
 BUF_X1 rebuffer6 (.A(_0205_),
    .Z(net66));
 BUF_X1 rebuffer7 (.A(net66),
    .Z(net67));
 BUF_X1 rebuffer16 (.A(_0559_),
    .Z(net80));
 BUF_X2 clone17 (.A(_0012_),
    .Z(net81));
 BUF_X8 clone26 (.A(_0003_),
    .Z(net91));
 BUF_X1 rebuffer29 (.A(_0295_),
    .Z(net94));
 BUF_X4 rebuffer36 (.A(_0266_),
    .Z(net102));
 BUF_X4 rebuffer37 (.A(net102),
    .Z(net103));
 FILLCELL_X16 FILLER_0_1 ();
 FILLCELL_X4 FILLER_0_17 ();
 FILLCELL_X2 FILLER_0_21 ();
 FILLCELL_X32 FILLER_0_26 ();
 FILLCELL_X16 FILLER_0_58 ();
 FILLCELL_X4 FILLER_0_74 ();
 FILLCELL_X2 FILLER_0_82 ();
 FILLCELL_X1 FILLER_0_84 ();
 FILLCELL_X8 FILLER_0_88 ();
 FILLCELL_X2 FILLER_0_99 ();
 FILLCELL_X1 FILLER_0_101 ();
 FILLCELL_X4 FILLER_0_115 ();
 FILLCELL_X2 FILLER_0_119 ();
 FILLCELL_X4 FILLER_0_124 ();
 FILLCELL_X2 FILLER_0_128 ();
 FILLCELL_X4 FILLER_0_148 ();
 FILLCELL_X1 FILLER_0_156 ();
 FILLCELL_X32 FILLER_0_170 ();
 FILLCELL_X16 FILLER_0_202 ();
 FILLCELL_X8 FILLER_0_218 ();
 FILLCELL_X2 FILLER_0_226 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X2 FILLER_1_33 ();
 FILLCELL_X1 FILLER_1_35 ();
 FILLCELL_X4 FILLER_1_85 ();
 FILLCELL_X1 FILLER_1_89 ();
 FILLCELL_X1 FILLER_1_97 ();
 FILLCELL_X2 FILLER_1_105 ();
 FILLCELL_X1 FILLER_1_114 ();
 FILLCELL_X4 FILLER_1_122 ();
 FILLCELL_X16 FILLER_1_184 ();
 FILLCELL_X8 FILLER_1_200 ();
 FILLCELL_X2 FILLER_1_208 ();
 FILLCELL_X1 FILLER_1_210 ();
 FILLCELL_X8 FILLER_1_214 ();
 FILLCELL_X4 FILLER_1_222 ();
 FILLCELL_X2 FILLER_1_226 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X16 FILLER_2_33 ();
 FILLCELL_X1 FILLER_2_112 ();
 FILLCELL_X2 FILLER_2_128 ();
 FILLCELL_X1 FILLER_2_166 ();
 FILLCELL_X4 FILLER_2_174 ();
 FILLCELL_X1 FILLER_2_178 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X16 FILLER_3_33 ();
 FILLCELL_X2 FILLER_3_49 ();
 FILLCELL_X8 FILLER_3_65 ();
 FILLCELL_X4 FILLER_3_80 ();
 FILLCELL_X2 FILLER_3_84 ();
 FILLCELL_X1 FILLER_3_86 ();
 FILLCELL_X1 FILLER_3_101 ();
 FILLCELL_X1 FILLER_3_111 ();
 FILLCELL_X1 FILLER_3_141 ();
 FILLCELL_X32 FILLER_3_176 ();
 FILLCELL_X16 FILLER_3_208 ();
 FILLCELL_X4 FILLER_3_224 ();
 FILLCELL_X16 FILLER_4_1 ();
 FILLCELL_X8 FILLER_4_17 ();
 FILLCELL_X4 FILLER_4_25 ();
 FILLCELL_X2 FILLER_4_29 ();
 FILLCELL_X1 FILLER_4_56 ();
 FILLCELL_X2 FILLER_4_70 ();
 FILLCELL_X1 FILLER_4_72 ();
 FILLCELL_X4 FILLER_4_80 ();
 FILLCELL_X1 FILLER_4_84 ();
 FILLCELL_X4 FILLER_4_112 ();
 FILLCELL_X1 FILLER_4_116 ();
 FILLCELL_X2 FILLER_4_140 ();
 FILLCELL_X2 FILLER_4_164 ();
 FILLCELL_X16 FILLER_4_210 ();
 FILLCELL_X2 FILLER_4_226 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X8 FILLER_5_33 ();
 FILLCELL_X4 FILLER_5_41 ();
 FILLCELL_X2 FILLER_5_45 ();
 FILLCELL_X1 FILLER_5_47 ();
 FILLCELL_X2 FILLER_5_74 ();
 FILLCELL_X1 FILLER_5_94 ();
 FILLCELL_X2 FILLER_5_115 ();
 FILLCELL_X1 FILLER_5_117 ();
 FILLCELL_X1 FILLER_5_122 ();
 FILLCELL_X1 FILLER_5_132 ();
 FILLCELL_X32 FILLER_5_178 ();
 FILLCELL_X16 FILLER_5_210 ();
 FILLCELL_X2 FILLER_5_226 ();
 FILLCELL_X8 FILLER_6_1 ();
 FILLCELL_X4 FILLER_6_9 ();
 FILLCELL_X2 FILLER_6_13 ();
 FILLCELL_X1 FILLER_6_64 ();
 FILLCELL_X1 FILLER_6_113 ();
 FILLCELL_X8 FILLER_6_128 ();
 FILLCELL_X2 FILLER_6_136 ();
 FILLCELL_X2 FILLER_6_141 ();
 FILLCELL_X2 FILLER_6_147 ();
 FILLCELL_X1 FILLER_6_165 ();
 FILLCELL_X1 FILLER_6_173 ();
 FILLCELL_X16 FILLER_6_202 ();
 FILLCELL_X2 FILLER_6_218 ();
 FILLCELL_X1 FILLER_6_223 ();
 FILLCELL_X1 FILLER_6_227 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X16 FILLER_7_33 ();
 FILLCELL_X2 FILLER_7_49 ();
 FILLCELL_X1 FILLER_7_51 ();
 FILLCELL_X1 FILLER_7_123 ();
 FILLCELL_X4 FILLER_7_132 ();
 FILLCELL_X1 FILLER_7_147 ();
 FILLCELL_X4 FILLER_7_157 ();
 FILLCELL_X1 FILLER_7_178 ();
 FILLCELL_X1 FILLER_7_210 ();
 FILLCELL_X8 FILLER_7_219 ();
 FILLCELL_X1 FILLER_7_227 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X4 FILLER_8_33 ();
 FILLCELL_X1 FILLER_8_37 ();
 FILLCELL_X1 FILLER_8_103 ();
 FILLCELL_X2 FILLER_8_142 ();
 FILLCELL_X2 FILLER_8_203 ();
 FILLCELL_X8 FILLER_8_214 ();
 FILLCELL_X4 FILLER_8_222 ();
 FILLCELL_X2 FILLER_8_226 ();
 FILLCELL_X1 FILLER_9_1 ();
 FILLCELL_X16 FILLER_9_6 ();
 FILLCELL_X2 FILLER_9_22 ();
 FILLCELL_X8 FILLER_9_27 ();
 FILLCELL_X2 FILLER_9_35 ();
 FILLCELL_X1 FILLER_9_37 ();
 FILLCELL_X16 FILLER_9_47 ();
 FILLCELL_X2 FILLER_9_63 ();
 FILLCELL_X1 FILLER_9_92 ();
 FILLCELL_X1 FILLER_9_127 ();
 FILLCELL_X1 FILLER_9_142 ();
 FILLCELL_X1 FILLER_9_147 ();
 FILLCELL_X1 FILLER_9_152 ();
 FILLCELL_X1 FILLER_9_158 ();
 FILLCELL_X2 FILLER_9_179 ();
 FILLCELL_X1 FILLER_9_207 ();
 FILLCELL_X1 FILLER_9_215 ();
 FILLCELL_X2 FILLER_9_220 ();
 FILLCELL_X2 FILLER_9_225 ();
 FILLCELL_X1 FILLER_9_227 ();
 FILLCELL_X8 FILLER_10_1 ();
 FILLCELL_X4 FILLER_10_9 ();
 FILLCELL_X1 FILLER_10_13 ();
 FILLCELL_X4 FILLER_10_18 ();
 FILLCELL_X4 FILLER_10_38 ();
 FILLCELL_X2 FILLER_10_42 ();
 FILLCELL_X1 FILLER_10_47 ();
 FILLCELL_X4 FILLER_10_52 ();
 FILLCELL_X2 FILLER_10_56 ();
 FILLCELL_X1 FILLER_10_132 ();
 FILLCELL_X2 FILLER_10_184 ();
 FILLCELL_X2 FILLER_10_222 ();
 FILLCELL_X1 FILLER_10_227 ();
 FILLCELL_X4 FILLER_11_1 ();
 FILLCELL_X2 FILLER_11_5 ();
 FILLCELL_X1 FILLER_11_7 ();
 FILLCELL_X2 FILLER_11_44 ();
 FILLCELL_X2 FILLER_11_103 ();
 FILLCELL_X2 FILLER_11_113 ();
 FILLCELL_X8 FILLER_11_126 ();
 FILLCELL_X2 FILLER_11_134 ();
 FILLCELL_X1 FILLER_11_165 ();
 FILLCELL_X4 FILLER_11_198 ();
 FILLCELL_X1 FILLER_11_202 ();
 FILLCELL_X1 FILLER_11_214 ();
 FILLCELL_X2 FILLER_11_222 ();
 FILLCELL_X1 FILLER_11_224 ();
 FILLCELL_X8 FILLER_12_1 ();
 FILLCELL_X4 FILLER_12_9 ();
 FILLCELL_X1 FILLER_12_16 ();
 FILLCELL_X1 FILLER_12_22 ();
 FILLCELL_X2 FILLER_12_50 ();
 FILLCELL_X2 FILLER_12_61 ();
 FILLCELL_X2 FILLER_12_176 ();
 FILLCELL_X2 FILLER_12_200 ();
 FILLCELL_X2 FILLER_12_213 ();
 FILLCELL_X4 FILLER_12_224 ();
 FILLCELL_X2 FILLER_13_1 ();
 FILLCELL_X1 FILLER_13_3 ();
 FILLCELL_X4 FILLER_13_31 ();
 FILLCELL_X1 FILLER_13_35 ();
 FILLCELL_X8 FILLER_13_53 ();
 FILLCELL_X1 FILLER_13_61 ();
 FILLCELL_X2 FILLER_13_73 ();
 FILLCELL_X1 FILLER_13_75 ();
 FILLCELL_X1 FILLER_13_90 ();
 FILLCELL_X1 FILLER_13_98 ();
 FILLCELL_X4 FILLER_13_112 ();
 FILLCELL_X1 FILLER_13_116 ();
 FILLCELL_X1 FILLER_13_124 ();
 FILLCELL_X1 FILLER_13_134 ();
 FILLCELL_X1 FILLER_13_148 ();
 FILLCELL_X2 FILLER_13_160 ();
 FILLCELL_X1 FILLER_13_162 ();
 FILLCELL_X1 FILLER_13_187 ();
 FILLCELL_X4 FILLER_13_214 ();
 FILLCELL_X4 FILLER_13_221 ();
 FILLCELL_X2 FILLER_13_225 ();
 FILLCELL_X1 FILLER_13_227 ();
 FILLCELL_X8 FILLER_14_1 ();
 FILLCELL_X1 FILLER_14_9 ();
 FILLCELL_X4 FILLER_14_19 ();
 FILLCELL_X2 FILLER_14_23 ();
 FILLCELL_X1 FILLER_14_30 ();
 FILLCELL_X2 FILLER_14_51 ();
 FILLCELL_X8 FILLER_14_94 ();
 FILLCELL_X1 FILLER_14_183 ();
 FILLCELL_X4 FILLER_14_195 ();
 FILLCELL_X2 FILLER_14_199 ();
 FILLCELL_X16 FILLER_14_203 ();
 FILLCELL_X8 FILLER_14_219 ();
 FILLCELL_X1 FILLER_14_227 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X4 FILLER_15_33 ();
 FILLCELL_X2 FILLER_15_37 ();
 FILLCELL_X4 FILLER_15_52 ();
 FILLCELL_X2 FILLER_15_94 ();
 FILLCELL_X1 FILLER_15_114 ();
 FILLCELL_X1 FILLER_15_159 ();
 FILLCELL_X4 FILLER_15_171 ();
 FILLCELL_X1 FILLER_15_175 ();
 FILLCELL_X4 FILLER_15_194 ();
 FILLCELL_X2 FILLER_15_198 ();
 FILLCELL_X4 FILLER_15_211 ();
 FILLCELL_X1 FILLER_15_215 ();
 FILLCELL_X4 FILLER_15_219 ();
 FILLCELL_X1 FILLER_15_223 ();
 FILLCELL_X16 FILLER_16_1 ();
 FILLCELL_X4 FILLER_16_17 ();
 FILLCELL_X8 FILLER_16_24 ();
 FILLCELL_X1 FILLER_16_32 ();
 FILLCELL_X4 FILLER_16_63 ();
 FILLCELL_X2 FILLER_16_67 ();
 FILLCELL_X1 FILLER_16_73 ();
 FILLCELL_X1 FILLER_16_78 ();
 FILLCELL_X1 FILLER_16_95 ();
 FILLCELL_X4 FILLER_16_107 ();
 FILLCELL_X1 FILLER_16_111 ();
 FILLCELL_X1 FILLER_16_121 ();
 FILLCELL_X1 FILLER_16_127 ();
 FILLCELL_X1 FILLER_16_149 ();
 FILLCELL_X2 FILLER_16_154 ();
 FILLCELL_X2 FILLER_16_163 ();
 FILLCELL_X2 FILLER_16_169 ();
 FILLCELL_X2 FILLER_16_182 ();
 FILLCELL_X1 FILLER_16_184 ();
 FILLCELL_X1 FILLER_16_188 ();
 FILLCELL_X1 FILLER_16_193 ();
 FILLCELL_X2 FILLER_16_207 ();
 FILLCELL_X1 FILLER_16_209 ();
 FILLCELL_X2 FILLER_16_219 ();
 FILLCELL_X1 FILLER_16_221 ();
 FILLCELL_X2 FILLER_16_225 ();
 FILLCELL_X1 FILLER_16_227 ();
 FILLCELL_X4 FILLER_17_1 ();
 FILLCELL_X2 FILLER_17_46 ();
 FILLCELL_X1 FILLER_17_57 ();
 FILLCELL_X4 FILLER_17_74 ();
 FILLCELL_X2 FILLER_17_82 ();
 FILLCELL_X1 FILLER_17_84 ();
 FILLCELL_X2 FILLER_17_98 ();
 FILLCELL_X1 FILLER_17_100 ();
 FILLCELL_X2 FILLER_17_105 ();
 FILLCELL_X1 FILLER_17_107 ();
 FILLCELL_X4 FILLER_17_117 ();
 FILLCELL_X2 FILLER_17_121 ();
 FILLCELL_X1 FILLER_17_123 ();
 FILLCELL_X8 FILLER_17_194 ();
 FILLCELL_X16 FILLER_17_211 ();
 FILLCELL_X1 FILLER_17_227 ();
 FILLCELL_X16 FILLER_18_4 ();
 FILLCELL_X2 FILLER_18_20 ();
 FILLCELL_X16 FILLER_18_53 ();
 FILLCELL_X1 FILLER_18_73 ();
 FILLCELL_X1 FILLER_18_77 ();
 FILLCELL_X2 FILLER_18_85 ();
 FILLCELL_X2 FILLER_18_91 ();
 FILLCELL_X1 FILLER_18_93 ();
 FILLCELL_X16 FILLER_18_115 ();
 FILLCELL_X1 FILLER_18_146 ();
 FILLCELL_X4 FILLER_18_158 ();
 FILLCELL_X2 FILLER_18_173 ();
 FILLCELL_X1 FILLER_18_183 ();
 FILLCELL_X4 FILLER_18_221 ();
 FILLCELL_X8 FILLER_19_1 ();
 FILLCELL_X4 FILLER_19_12 ();
 FILLCELL_X2 FILLER_19_16 ();
 FILLCELL_X1 FILLER_19_43 ();
 FILLCELL_X4 FILLER_19_66 ();
 FILLCELL_X4 FILLER_19_98 ();
 FILLCELL_X1 FILLER_19_102 ();
 FILLCELL_X2 FILLER_19_141 ();
 FILLCELL_X2 FILLER_19_149 ();
 FILLCELL_X1 FILLER_19_151 ();
 FILLCELL_X1 FILLER_19_155 ();
 FILLCELL_X2 FILLER_19_186 ();
 FILLCELL_X2 FILLER_19_214 ();
 FILLCELL_X4 FILLER_19_221 ();
 FILLCELL_X4 FILLER_20_1 ();
 FILLCELL_X2 FILLER_20_5 ();
 FILLCELL_X1 FILLER_20_7 ();
 FILLCELL_X8 FILLER_20_17 ();
 FILLCELL_X1 FILLER_20_25 ();
 FILLCELL_X2 FILLER_20_63 ();
 FILLCELL_X1 FILLER_20_65 ();
 FILLCELL_X2 FILLER_20_73 ();
 FILLCELL_X1 FILLER_20_75 ();
 FILLCELL_X1 FILLER_20_110 ();
 FILLCELL_X1 FILLER_20_119 ();
 FILLCELL_X1 FILLER_20_124 ();
 FILLCELL_X4 FILLER_20_132 ();
 FILLCELL_X2 FILLER_20_140 ();
 FILLCELL_X4 FILLER_20_149 ();
 FILLCELL_X2 FILLER_20_156 ();
 FILLCELL_X2 FILLER_20_167 ();
 FILLCELL_X1 FILLER_20_169 ();
 FILLCELL_X4 FILLER_20_177 ();
 FILLCELL_X1 FILLER_20_181 ();
 FILLCELL_X1 FILLER_20_227 ();
 FILLCELL_X16 FILLER_21_1 ();
 FILLCELL_X8 FILLER_21_17 ();
 FILLCELL_X2 FILLER_21_25 ();
 FILLCELL_X1 FILLER_21_27 ();
 FILLCELL_X16 FILLER_21_30 ();
 FILLCELL_X8 FILLER_21_46 ();
 FILLCELL_X2 FILLER_21_78 ();
 FILLCELL_X1 FILLER_21_80 ();
 FILLCELL_X1 FILLER_21_89 ();
 FILLCELL_X1 FILLER_21_99 ();
 FILLCELL_X2 FILLER_21_104 ();
 FILLCELL_X1 FILLER_21_115 ();
 FILLCELL_X2 FILLER_21_119 ();
 FILLCELL_X1 FILLER_21_130 ();
 FILLCELL_X2 FILLER_21_146 ();
 FILLCELL_X4 FILLER_21_153 ();
 FILLCELL_X2 FILLER_21_157 ();
 FILLCELL_X4 FILLER_21_181 ();
 FILLCELL_X1 FILLER_21_185 ();
 FILLCELL_X1 FILLER_21_227 ();
 FILLCELL_X1 FILLER_22_1 ();
 FILLCELL_X8 FILLER_22_18 ();
 FILLCELL_X1 FILLER_22_26 ();
 FILLCELL_X8 FILLER_22_39 ();
 FILLCELL_X1 FILLER_22_47 ();
 FILLCELL_X2 FILLER_22_53 ();
 FILLCELL_X2 FILLER_22_62 ();
 FILLCELL_X1 FILLER_22_64 ();
 FILLCELL_X1 FILLER_22_72 ();
 FILLCELL_X4 FILLER_22_78 ();
 FILLCELL_X1 FILLER_22_82 ();
 FILLCELL_X2 FILLER_22_90 ();
 FILLCELL_X4 FILLER_22_110 ();
 FILLCELL_X2 FILLER_22_114 ();
 FILLCELL_X1 FILLER_22_116 ();
 FILLCELL_X4 FILLER_22_120 ();
 FILLCELL_X1 FILLER_22_124 ();
 FILLCELL_X4 FILLER_22_130 ();
 FILLCELL_X4 FILLER_22_147 ();
 FILLCELL_X2 FILLER_22_151 ();
 FILLCELL_X1 FILLER_22_153 ();
 FILLCELL_X2 FILLER_23_42 ();
 FILLCELL_X1 FILLER_23_55 ();
 FILLCELL_X2 FILLER_23_63 ();
 FILLCELL_X1 FILLER_23_65 ();
 FILLCELL_X8 FILLER_23_69 ();
 FILLCELL_X4 FILLER_23_77 ();
 FILLCELL_X2 FILLER_23_81 ();
 FILLCELL_X1 FILLER_23_83 ();
 FILLCELL_X2 FILLER_23_101 ();
 FILLCELL_X1 FILLER_23_103 ();
 FILLCELL_X1 FILLER_23_115 ();
 FILLCELL_X2 FILLER_23_147 ();
 FILLCELL_X1 FILLER_23_149 ();
 FILLCELL_X8 FILLER_23_164 ();
 FILLCELL_X4 FILLER_23_172 ();
 FILLCELL_X2 FILLER_23_179 ();
 FILLCELL_X2 FILLER_23_188 ();
 FILLCELL_X2 FILLER_23_214 ();
 FILLCELL_X16 FILLER_24_1 ();
 FILLCELL_X8 FILLER_24_17 ();
 FILLCELL_X1 FILLER_24_46 ();
 FILLCELL_X1 FILLER_24_54 ();
 FILLCELL_X8 FILLER_24_68 ();
 FILLCELL_X1 FILLER_24_97 ();
 FILLCELL_X1 FILLER_24_102 ();
 FILLCELL_X1 FILLER_24_112 ();
 FILLCELL_X4 FILLER_24_120 ();
 FILLCELL_X2 FILLER_24_124 ();
 FILLCELL_X1 FILLER_24_126 ();
 FILLCELL_X4 FILLER_24_154 ();
 FILLCELL_X1 FILLER_24_158 ();
 FILLCELL_X2 FILLER_24_167 ();
 FILLCELL_X1 FILLER_24_169 ();
 FILLCELL_X4 FILLER_24_174 ();
 FILLCELL_X2 FILLER_24_194 ();
 FILLCELL_X1 FILLER_24_210 ();
 FILLCELL_X1 FILLER_24_218 ();
 FILLCELL_X2 FILLER_24_222 ();
 FILLCELL_X1 FILLER_24_224 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X8 FILLER_25_33 ();
 FILLCELL_X4 FILLER_25_41 ();
 FILLCELL_X2 FILLER_25_45 ();
 FILLCELL_X16 FILLER_25_71 ();
 FILLCELL_X8 FILLER_25_87 ();
 FILLCELL_X1 FILLER_25_95 ();
 FILLCELL_X1 FILLER_25_122 ();
 FILLCELL_X4 FILLER_25_156 ();
 FILLCELL_X2 FILLER_25_160 ();
 FILLCELL_X1 FILLER_25_162 ();
 FILLCELL_X2 FILLER_25_178 ();
 FILLCELL_X1 FILLER_25_180 ();
 FILLCELL_X1 FILLER_25_206 ();
 FILLCELL_X2 FILLER_25_209 ();
 FILLCELL_X1 FILLER_25_227 ();
 FILLCELL_X16 FILLER_26_1 ();
 FILLCELL_X8 FILLER_26_30 ();
 FILLCELL_X4 FILLER_26_38 ();
 FILLCELL_X1 FILLER_26_65 ();
 FILLCELL_X8 FILLER_26_80 ();
 FILLCELL_X2 FILLER_26_88 ();
 FILLCELL_X1 FILLER_26_103 ();
 FILLCELL_X1 FILLER_26_107 ();
 FILLCELL_X1 FILLER_26_115 ();
 FILLCELL_X2 FILLER_26_123 ();
 FILLCELL_X1 FILLER_26_125 ();
 FILLCELL_X1 FILLER_26_137 ();
 FILLCELL_X2 FILLER_26_145 ();
 FILLCELL_X2 FILLER_26_152 ();
 FILLCELL_X2 FILLER_26_172 ();
 FILLCELL_X1 FILLER_26_174 ();
 FILLCELL_X1 FILLER_26_185 ();
 FILLCELL_X1 FILLER_26_202 ();
 FILLCELL_X2 FILLER_26_215 ();
 FILLCELL_X2 FILLER_26_222 ();
 FILLCELL_X1 FILLER_26_224 ();
 FILLCELL_X16 FILLER_27_1 ();
 FILLCELL_X4 FILLER_27_17 ();
 FILLCELL_X2 FILLER_27_21 ();
 FILLCELL_X16 FILLER_27_74 ();
 FILLCELL_X4 FILLER_27_90 ();
 FILLCELL_X2 FILLER_27_94 ();
 FILLCELL_X1 FILLER_27_115 ();
 FILLCELL_X2 FILLER_27_130 ();
 FILLCELL_X2 FILLER_27_165 ();
 FILLCELL_X2 FILLER_27_180 ();
 FILLCELL_X4 FILLER_27_205 ();
 FILLCELL_X8 FILLER_27_214 ();
 FILLCELL_X2 FILLER_27_222 ();
 FILLCELL_X1 FILLER_27_224 ();
 FILLCELL_X2 FILLER_28_62 ();
 FILLCELL_X16 FILLER_28_74 ();
 FILLCELL_X4 FILLER_28_90 ();
 FILLCELL_X1 FILLER_28_94 ();
 FILLCELL_X4 FILLER_28_119 ();
 FILLCELL_X1 FILLER_28_129 ();
 FILLCELL_X1 FILLER_28_173 ();
 FILLCELL_X8 FILLER_28_190 ();
 FILLCELL_X4 FILLER_28_198 ();
 FILLCELL_X1 FILLER_28_202 ();
 FILLCELL_X4 FILLER_28_221 ();
 FILLCELL_X2 FILLER_28_225 ();
 FILLCELL_X1 FILLER_28_227 ();
 FILLCELL_X16 FILLER_29_1 ();
 FILLCELL_X2 FILLER_29_17 ();
 FILLCELL_X1 FILLER_29_19 ();
 FILLCELL_X2 FILLER_29_33 ();
 FILLCELL_X1 FILLER_29_35 ();
 FILLCELL_X16 FILLER_29_59 ();
 FILLCELL_X8 FILLER_29_75 ();
 FILLCELL_X2 FILLER_29_83 ();
 FILLCELL_X16 FILLER_29_89 ();
 FILLCELL_X1 FILLER_29_105 ();
 FILLCELL_X1 FILLER_29_114 ();
 FILLCELL_X8 FILLER_29_118 ();
 FILLCELL_X1 FILLER_29_126 ();
 FILLCELL_X2 FILLER_29_130 ();
 FILLCELL_X1 FILLER_29_132 ();
 FILLCELL_X1 FILLER_29_139 ();
 FILLCELL_X1 FILLER_29_143 ();
 FILLCELL_X2 FILLER_29_147 ();
 FILLCELL_X2 FILLER_29_170 ();
 FILLCELL_X4 FILLER_29_175 ();
 FILLCELL_X2 FILLER_29_185 ();
 FILLCELL_X1 FILLER_29_187 ();
 FILLCELL_X8 FILLER_29_191 ();
 FILLCELL_X2 FILLER_29_199 ();
 FILLCELL_X16 FILLER_29_204 ();
 FILLCELL_X8 FILLER_29_220 ();
endmodule
